/* Verilog module written by vlog2Verilog (qflow) */

module mips(
    output MemRead,
    output MemWrite,
    input clk,
    output [31:0] memoryAddress,
    input [31:0] memoryOutData,
    output [31:0] memoryWriteData,
    input rst
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf2  ;
wire _5488__bF$buf0 ;
wire _5488__bF$buf1 ;
wire _5488__bF$buf2 ;
wire _5488__bF$buf3 ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire [31:0] _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire IRWrite_bF$buf0 ;
wire IRWrite_bF$buf1 ;
wire _1486_ ;
wire IRWrite_bF$buf2 ;
wire _1066_ ;
wire IRWrite_bF$buf3 ;
wire IRWrite_bF$buf4 ;
wire IRWrite_bF$buf5 ;
wire IRWrite_bF$buf6 ;
wire IRWrite_bF$buf7 ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire [31:0] _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf1  ;
wire \datapath_1.mux_wd3.dout_11_bF$buf4  ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6410_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf0  ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf0  ;
wire _57_ ;
wire _6504_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf4  ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf2  ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _5436__bF$buf0 ;
wire _5436__bF$buf1 ;
wire _5436__bF$buf2 ;
wire _5436__bF$buf3 ;
wire _1924_ ;
wire _5436__bF$buf4 ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6542_ ;
wire _6122_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf3  ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf0  ;
wire _6771_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf7  ;
wire _6351_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf3  ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf7  ;
wire _6580_ ;
wire _6160_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf5  ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _3947__bF$buf0 ;
wire _3947__bF$buf1 ;
wire _3947__bF$buf2 ;
wire _3947__bF$buf3 ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf3  ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire [31:0] \datapath_1.regfile_1.regOut[13]  ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire \datapath_1.PCJump_27_bF$buf2  ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _4643_ ;
wire _4223_ ;
wire [31:0] \datapath_1.regfile_1.regOut[7]  ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf2  ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf1  ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf5  ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _5518__bF$buf0 ;
wire _5518__bF$buf1 ;
wire _5518__bF$buf2 ;
wire _5518__bF$buf3 ;
wire _5518__bF$buf4 ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf1  ;
wire _54_ ;
wire _6501_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf4  ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf1  ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf0  ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf0  ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire PCWrite ;
wire _4678_ ;
wire _4258_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf4  ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf2  ;
wire _3282_ ;
wire RegWrite_bF$buf0 ;
wire RegWrite_bF$buf1 ;
wire RegWrite_bF$buf2 ;
wire RegWrite_bF$buf3 ;
wire RegWrite_bF$buf4 ;
wire RegWrite_bF$buf5 ;
wire RegWrite_bF$buf6 ;
wire RegWrite_bF$buf7 ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6442_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf0  ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf3  ;
wire _5713_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _2591_ ;
wire _2171_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf7  ;
wire _3796_ ;
wire _3376_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf3  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire \datapath_1.PCJump_22_bF$buf3  ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf7  ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf3  ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf7  ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6574_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _5506__bF$buf0 ;
wire _5506__bF$buf1 ;
wire _5506__bF$buf2 ;
wire _5506__bF$buf3 ;
wire _5506__bF$buf4 ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf2  ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf2  ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf1  ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf5  ;
wire _1286_ ;
wire _197_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf1  ;
wire _3717_ ;
wire _6189_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf4  ;
wire _3902__bF$buf0 ;
wire _3902__bF$buf1 ;
wire _3902__bF$buf2 ;
wire _3902__bF$buf3 ;
wire _3902__bF$buf4 ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _6401_ ;
wire _2741_ ;
wire _2321_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf1  ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf4  ;
wire _7_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf0  ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf4  ;
wire _3793_ ;
wire _3373_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf0  ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire Branch ;
wire \datapath_1.PCJump_22_bF$buf0  ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3894__bF$buf0 ;
wire _3894__bF$buf1 ;
wire _3894__bF$buf2 ;
wire _3894__bF$buf3 ;
wire _3894__bF$buf4 ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf4  ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6533_ ;
wire _6113_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf3  ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf0  ;
wire _6762_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf4  ;
wire _5613_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf7  ;
wire [31:0] _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6571_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire rst_bF$buf110 ;
wire rst_bF$buf111 ;
wire rst_bF$buf112 ;
wire rst_bF$buf113 ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _3957__bF$buf0 ;
wire _3957__bF$buf1 ;
wire _3957__bF$buf2 ;
wire _3957__bF$buf3 ;
wire _3957__bF$buf4 ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire RegDst ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6474_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _5513__bF$buf0 ;
wire _156_ ;
wire _5513__bF$buf1 ;
wire _5513__bF$buf2 ;
wire _5513__bF$buf3 ;
wire _5513__bF$buf4 ;
wire _3811_ ;
wire _6283_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire clk_bF$buf80 ;
wire clk_bF$buf81 ;
wire clk_bF$buf82 ;
wire clk_bF$buf83 ;
wire clk_bF$buf84 ;
wire clk_bF$buf85 ;
wire clk_bF$buf86 ;
wire _3620_ ;
wire clk_bF$buf87 ;
wire _3200_ ;
wire clk_bF$buf88 ;
wire clk_bF$buf89 ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _5783_ ;
wire _5363_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf2  ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf1  ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf5  ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf1  ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf5  ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _45_ ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf1  ;
wire _3790_ ;
wire _3370_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf4  ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf5  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf1  ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf0  ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf1  ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf4  ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6433_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _5704_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _2582_ ;
wire _3022__bF$buf0 ;
wire _2162_ ;
wire _3022__bF$buf1 ;
wire _3022__bF$buf2 ;
wire _3022__bF$buf3 ;
wire _3022__bF$buf4 ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire _1853_ ;
wire [31:0] _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6471_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _4060__bF$buf0 ;
wire _4060__bF$buf1 ;
wire _4060__bF$buf2 ;
wire _4060__bF$buf3 ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf2  ;
wire [31:0] \datapath_1.regfile_1.regOut[2]  ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6565_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf2  ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire [31:0] \datapath_1.regfile_1.regOut[25]  ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire _5520__bF$buf0 ;
wire _5520__bF$buf1 ;
wire _5520__bF$buf2 ;
wire _5520__bF$buf3 ;
wire _5520__bF$buf4 ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf2  ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire [31:0] _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _5683_ ;
wire _5263_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf2  ;
wire _2388_ ;
wire _2354__bF$buf0 ;
wire _2354__bF$buf1 ;
wire _2354__bF$buf2 ;
wire _2354__bF$buf3 ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire rst_bF$buf0 ;
wire rst_bF$buf1 ;
wire rst_bF$buf2 ;
wire rst_bF$buf3 ;
wire rst_bF$buf4 ;
wire rst_bF$buf5 ;
wire _5968_ ;
wire rst_bF$buf6 ;
wire _5548_ ;
wire rst_bF$buf7 ;
wire _5128_ ;
wire rst_bF$buf8 ;
wire rst_bF$buf9 ;
wire _42_ ;
wire [31:0] _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf1  ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf2  ;
wire _4628_ ;
wire _4208_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf5  ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf1  ;
wire \datapath_1.mux_wd3.dout_27_bF$buf4  ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf5  ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf4  ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6430_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire rst_bF$buf90 ;
wire rst_bF$buf91 ;
wire rst_bF$buf92 ;
wire rst_bF$buf93 ;
wire rst_bF$buf94 ;
wire rst_bF$buf95 ;
wire rst_bF$buf96 ;
wire rst_bF$buf97 ;
wire rst_bF$buf98 ;
wire rst_bF$buf99 ;
wire _5701_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire IorD ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6524_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _5460__bF$buf0 ;
wire _5460__bF$buf1 ;
wire _5460__bF$buf2 ;
wire _5460__bF$buf3 ;
wire _5460__bF$buf4 ;
wire _6562_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf2  ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf5  ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire [31:0] \datapath_1.regfile_1.regOut[15]  ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf4  ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf2  ;
wire _5583_ ;
wire _5163_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf6  ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire [3:0] _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire [31:0] \datapath_1.regfile_1.regOut[9]  ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf1  ;
wire _1788_ ;
wire [31:0] _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf2  ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf1  ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf5  ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire rst_bF$buf60 ;
wire rst_bF$buf61 ;
wire rst_bF$buf62 ;
wire rst_bF$buf63 ;
wire rst_bF$buf64 ;
wire rst_bF$buf65 ;
wire rst_bF$buf66 ;
wire rst_bF$buf67 ;
wire rst_bF$buf68 ;
wire rst_bF$buf69 ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _3915__bF$buf0 ;
wire _3915__bF$buf1 ;
wire _3915__bF$buf2 ;
wire _3915__bF$buf3 ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf5  ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire RegWrite ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6521_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf3  ;
wire _5601_ ;
wire [31:0] \datapath_1.mux_pcsrc.dout  ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire [31:0] \datapath_1.regfile_1.regOut[30]  ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire [5:0] \control_1.op  ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf2  ;
wire _2629_ ;
wire _2209_ ;
wire _6462_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf1  ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf5  ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf2  ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf3  ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf4  ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _5674_ ;
wire _5254_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf2  ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_31_bF$buf2  ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire rst_bF$buf30 ;
wire rst_bF$buf31 ;
wire rst_bF$buf32 ;
wire rst_bF$buf33 ;
wire rst_bF$buf34 ;
wire rst_bF$buf35 ;
wire rst_bF$buf36 ;
wire rst_bF$buf37 ;
wire rst_bF$buf38 ;
wire rst_bF$buf39 ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire [31:0] _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf2  ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _3185__bF$buf0 ;
wire _3185__bF$buf1 ;
wire _3185__bF$buf2 ;
wire _3185__bF$buf3 ;
wire _3185__bF$buf4 ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf0  ;
wire _4657_ ;
wire _4237_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6421_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf3  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire [31:0] _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf2  ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire [31:0] _68_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf6  ;
wire [31:0] \datapath_1.Data  ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire [31:0] \datapath_1.regfile_1.regOut[20]  ;
wire _5466__bF$buf0 ;
wire _5466__bF$buf1 ;
wire _5466__bF$buf2 ;
wire _5466__bF$buf3 ;
wire _5466__bF$buf4 ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6553_ ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf2  ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf0  ;
wire _5633_ ;
wire _5213_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf1  ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _5918_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf5  ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6456_ ;
wire _6036_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf2  ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf5  ;
wire _5727_ ;
wire _5307_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf3  ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire [31:0] _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _2185_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _3906__bF$buf0 ;
wire _3906__bF$buf1 ;
wire _3906__bF$buf2 ;
wire _3906__bF$buf3 ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire MemRead ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire \datapath_1.PCJump_17_bF$buf4  ;
wire _4616_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf6  ;
wire _2699_ ;
wire _2279_ ;
wire _2367__bF$buf0 ;
wire _2367__bF$buf1 ;
wire _3640_ ;
wire _2367__bF$buf2 ;
wire _3220_ ;
wire _2367__bF$buf3 ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire clk_hier0_bF$buf8 ;
wire clk_hier0_bF$buf9 ;
wire _2088_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf4  ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf0  ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire clk_bF$buf110 ;
wire clk_bF$buf111 ;
wire clk_bF$buf112 ;
wire clk_bF$buf113 ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _6703_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6512_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf3  ;
wire _3637_ ;
wire _3217_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf3  ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6550_ ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf2  ;
wire _5821_ ;
wire _5401_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf6  ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire [31:0] \datapath_1.regfile_1.regOut[10]  ;
wire \datapath_1.regfile_1.regEn_18_bF$buf2  ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6453_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf2  ;
wire _5724_ ;
wire _5304_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf0  ;
wire _6509_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf7  ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire \datapath_1.PCJump_17_bF$buf1  ;
wire _4613_ ;
wire [31:0] \datapath_1.regfile_1.regOut[4]  ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf5  ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf3  ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire [31:0] _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf4  ;
wire _4707_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf1  ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire [31:0] \datapath_1.regfile_1.regOut[27]  ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _5492__bF$buf0 ;
wire _5492__bF$buf1 ;
wire _5492__bF$buf2 ;
wire _5492__bF$buf3 ;
wire _5492__bF$buf4 ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire [31:0] _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _5421__bF$buf0 ;
wire _5421__bF$buf1 ;
wire _5421__bF$buf2 ;
wire _5421__bF$buf3 ;
wire \datapath_1.mux_wd3.dout_3_bF$buf4  ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf0  ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf0  ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _5555__bF$buf0 ;
wire _5555__bF$buf1 ;
wire _5555__bF$buf2 ;
wire _5555__bF$buf3 ;
wire _6603_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf3  ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6412_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire MemToReg ;
wire _6641_ ;
wire _6221_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf2  ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6450_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf6  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf2  ;
wire _59_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf6  ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf4  ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire [31:0] \datapath_1.rd1  ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf2  ;
wire _6773_ ;
wire _6353_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf0  ;
wire _2693_ ;
wire _2273_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire [5:0] \aluControl_1.inst  ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf7  ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf1  ;
wire _4704_ ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf5  ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire PCEn_bF$buf0 ;
wire PCEn_bF$buf1 ;
wire PCEn_bF$buf2 ;
wire PCEn_bF$buf3 ;
wire PCEn_bF$buf4 ;
wire PCEn_bF$buf5 ;
wire PCEn_bF$buf6 ;
wire PCEn_bF$buf7 ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _3916__bF$buf0 ;
wire _3916__bF$buf1 ;
wire _3916__bF$buf2 ;
wire _3916__bF$buf3 ;
wire _3916__bF$buf4 ;
wire _5756_ ;
wire _5336_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf1  ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire [31:0] \datapath_1.regfile_1.regOut[17]  ;
wire \datapath_1.PCJump_27_bF$buf4  ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf4  ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_11_bF$buf3  ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf7  ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _5558__bF$buf0 ;
wire _5558__bF$buf1 ;
wire _5558__bF$buf2 ;
wire _2614_ ;
wire _5558__bF$buf3 ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _3935__bF$buf0 ;
wire _3935__bF$buf1 ;
wire _3935__bF$buf2 ;
wire _3935__bF$buf3 ;
wire _4777_ ;
wire _4357_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf3  ;
wire _56_ ;
wire _6503_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf3  ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf1  ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6541_ ;
wire _6121_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf2  ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire [31:0] \datapath_1.alu_1.ALUInB  ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf6  ;
wire _6350_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf2  ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire [31:0] _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_5_bF$buf4  ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire [3:0] \control_1.reg_state.dout  ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf2  ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire \datapath_1.PCJump_27_bF$buf1  ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire [31:0] _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf1  ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf0  ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3875__bF$buf0 ;
wire _3875__bF$buf1 ;
wire _3875__bF$buf2 ;
wire _3875__bF$buf3 ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf4  ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf4  ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _4774_ ;
wire _4354_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf0  ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6500_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf3  ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _4583_ ;
wire _4163_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf0  ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf7  ;
wire _1288_ ;
wire _199_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf3  ;
wire _3719_ ;
wire _5565__bF$buf0 ;
wire _5565__bF$buf1 ;
wire _5565__bF$buf2 ;
wire _5565__bF$buf3 ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _6403_ ;
wire _2743_ ;
wire _2323_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf3  ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf1  ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire [31:0] _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire ALUOp_0_bF$buf0 ;
wire ALUOp_0_bF$buf1 ;
wire ALUOp_0_bF$buf2 ;
wire ALUOp_0_bF$buf3 ;
wire ALUOp_0_bF$buf4 ;
wire _2608_ ;
wire ALUOp_0_bF$buf5 ;
wire _6441_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf2  ;
wire _5712_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _2590_ ;
wire _2170_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf6  ;
wire _3795_ ;
wire _3375_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf2  ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire \datapath_1.PCJump_22_bF$buf2  ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf6  ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf2  ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf6  ;
wire _5615_ ;
wire [31:0] \datapath_1.regfile_1.regOut[22]  ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6573_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _3961__bF$buf0 ;
wire _3961__bF$buf1 ;
wire _3961__bF$buf2 ;
wire _3961__bF$buf3 ;
wire _3961__bF$buf4 ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf1  ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf1  ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf0  ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf4  ;
wire _1285_ ;
wire _196_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6379_ ;
wire _1094_ ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf0  ;
wire _3716_ ;
wire _6188_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf3  ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf0  ;
wire \datapath_1.regfile_1.regEn_17_bF$buf7  ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf3  ;
wire _6_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf7  ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf3  ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf7  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf3  ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6532_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _5803_ ;
wire _1723_ ;
wire [31:0] _1303_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf2  ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf3  ;
wire _5612_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf6  ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6570_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire rst_bF$buf100 ;
wire rst_bF$buf101 ;
wire rst_bF$buf102 ;
wire rst_bF$buf103 ;
wire rst_bF$buf104 ;
wire rst_bF$buf105 ;
wire rst_bF$buf106 ;
wire rst_bF$buf107 ;
wire rst_bF$buf108 ;
wire rst_bF$buf109 ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire rst ;
wire _3866__bF$buf0 ;
wire _3866__bF$buf1 ;
wire _3866__bF$buf2 ;
wire _3866__bF$buf3 ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _5493__bF$buf0 ;
wire _5493__bF$buf1 ;
wire _5493__bF$buf2 ;
wire _5493__bF$buf3 ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire [31:0] \datapath_1.regfile_1.regOut[12]  ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _3870__bF$buf0 ;
wire _766_ ;
wire _3870__bF$buf1 ;
wire _346_ ;
wire _3870__bF$buf2 ;
wire _3870__bF$buf3 ;
wire _6473_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf4  ;
wire MemWrite ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire clk_bF$buf76 ;
wire clk_bF$buf77 ;
wire clk_bF$buf78 ;
wire clk_bF$buf79 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf1  ;
wire _6567_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf4  ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire [31:0] \datapath_1.regfile_1.regOut[6]  ;
wire _5838_ ;
wire _5418_ ;
wire [31:0] _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf0  ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf4  ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf0  ;
wire [31:0] _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [31:0] \datapath_1.regfile_1.regOut[29]  ;
wire _1185_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf4  ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _2199_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_24_bF$buf3  ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf4  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf0  ;
wire \datapath_1.regfile_1.regEn_24_bF$buf7  ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf0  ;
wire _4668_ ;
wire _4248_ ;
wire [4:0] \datapath_1.a3  ;
wire \datapath_1.regfile_1.regEn_29_bF$buf3  ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _3952__bF$buf0 ;
wire _3952__bF$buf1 ;
wire _3952__bF$buf2 ;
wire _3952__bF$buf3 ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf7  ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6432_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _5703_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6470_ ;
wire _6050_ ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf1  ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6564_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf1  ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6373_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf4  ;
wire _5644_ ;
wire _5224_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf1  ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf7  ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf1  ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire [31:0] _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf0  ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf1  ;
wire _4627_ ;
wire _4207_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf4  ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire [31:0] \datapath_1.regfile_1.regOut[19]  ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_27_bF$buf3  ;
wire _2731_ ;
wire _2311_ ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf4  ;
wire [31:0] _913_ ;
wire _5679_ ;
wire _5259_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf7  ;
wire _6620_ ;
wire _6200_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf3  ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf7  ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire rst_bF$buf80 ;
wire rst_bF$buf81 ;
wire rst_bF$buf82 ;
wire rst_bF$buf83 ;
wire rst_bF$buf84 ;
wire rst_bF$buf85 ;
wire rst_bF$buf86 ;
wire rst_bF$buf87 ;
wire rst_bF$buf88 ;
wire rst_bF$buf89 ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _6714_ ;
wire _760_ ;
wire _340_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf7  ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6523_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _5511__bF$buf0 ;
wire _2672_ ;
wire _5511__bF$buf1 ;
wire _2252_ ;
wire _5511__bF$buf2 ;
wire _5511__bF$buf3 ;
wire _5511__bF$buf4 ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6561_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf1  ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf4  ;
wire _6464_ ;
wire _6044_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _5428__bF$buf0 ;
wire _5428__bF$buf1 ;
wire _5428__bF$buf2 ;
wire _5428__bF$buf3 ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _2193_ ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf3  ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire _6558_ ;
wire _6138_ ;
wire [31:0] _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf7  ;
wire _4624_ ;
wire _4204_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf1  ;
wire _5829_ ;
wire _5409_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf4  ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf5  ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf0  ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf1  ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf0  ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _4280_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf4  ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire rst_bF$buf50 ;
wire rst_bF$buf51 ;
wire rst_bF$buf52 ;
wire rst_bF$buf53 ;
wire rst_bF$buf54 ;
wire rst_bF$buf55 ;
wire rst_bF$buf56 ;
wire rst_bF$buf57 ;
wire rst_bF$buf58 ;
wire rst_bF$buf59 ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire [31:0] _6711_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf4  ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf2  ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _3962__bF$buf0 ;
wire _3962__bF$buf1 ;
wire _3962__bF$buf2 ;
wire _3962__bF$buf3 ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6423_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _5514__bF$buf0 ;
wire _5514__bF$buf1 ;
wire _5514__bF$buf2 ;
wire _5514__bF$buf3 ;
wire _5514__bF$buf4 ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf1  ;
wire _2628_ ;
wire _2208_ ;
wire _6461_ ;
wire _6041_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf4  ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _2190_ ;
wire [31:0] \datapath_1.regfile_1.regOut[1]  ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf0  ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire [31:0] _848_ ;
wire _428_ ;
wire _3879__bF$buf0 ;
wire _3879__bF$buf1 ;
wire _3879__bF$buf2 ;
wire _3879__bF$buf3 ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf4  ;
wire _4621_ ;
wire _4201_ ;
wire _5826_ ;
wire _5406_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf1  ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf2  ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire [31:0] \datapath_1.regfile_1.regOut[24]  ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf3  ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf7  ;
wire _5673_ ;
wire _5253_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf1  ;
wire _6458_ ;
wire _6038_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf4  ;
wire _1593_ ;
wire _3910__bF$buf0 ;
wire [31:0] _1173_ ;
wire _3910__bF$buf1 ;
wire _3910__bF$buf2 ;
wire _3910__bF$buf3 ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf7  ;
wire _5729_ ;
wire _5309_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf5  ;
wire _1649_ ;
wire _1229_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf1  ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire rst_bF$buf20 ;
wire rst_bF$buf21 ;
wire rst_bF$buf22 ;
wire rst_bF$buf23 ;
wire rst_bF$buf24 ;
wire rst_bF$buf25 ;
wire rst_bF$buf26 ;
wire rst_bF$buf27 ;
wire rst_bF$buf28 ;
wire rst_bF$buf29 ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire [31:0] \datapath_1.mux_wd3.dout  ;
wire _1687_ ;
wire _1267_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf1  ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _3019__bF$buf0 ;
wire _3019__bF$buf1 ;
wire _3019__bF$buf2 ;
wire _3019__bF$buf3 ;
wire _3019__bF$buf4 ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf2  ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf1  ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf5  ;
wire _3639_ ;
wire _3219_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _5517__bF$buf0 ;
wire _5517__bF$buf1 ;
wire _5517__bF$buf2 ;
wire _5517__bF$buf3 ;
wire _5517__bF$buf4 ;
wire _6743_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _5521__bF$buf0 ;
wire _5521__bF$buf1 ;
wire _5521__bF$buf2 ;
wire _5521__bF$buf3 ;
wire _5521__bF$buf4 ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6552_ ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf1  ;
wire _3677_ ;
wire _3257_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf4  ;
wire _5823_ ;
wire _5403_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf0  ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf4  ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire [31:0] _328_ ;
wire _6455_ ;
wire _6035_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf1  ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _3886__bF$buf0 ;
wire _3886__bF$buf1 ;
wire _3886__bF$buf2 ;
wire _3886__bF$buf3 ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf4  ;
wire _5726_ ;
wire _5306_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf2  ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire [31:0] \datapath_1.regfile_1.regOut[14]  ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire [31:0] _3410_ ;
wire \datapath_1.PCJump_17_bF$buf3  ;
wire _4615_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf7  ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf5  ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire _4653_ ;
wire [31:0] memoryWriteData ;
wire _4233_ ;
wire [31:0] \datapath_1.regfile_1.regOut[8]  ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf3  ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire clk_bF$buf100 ;
wire clk_bF$buf101 ;
wire clk_bF$buf102 ;
wire clk_bF$buf103 ;
wire clk_bF$buf104 ;
wire clk_bF$buf105 ;
wire clk_bF$buf106 ;
wire clk_bF$buf107 ;
wire clk_bF$buf108 ;
wire clk_bF$buf109 ;
wire _3771_ ;
wire _3351_ ;
wire _5457__bF$buf0 ;
wire _5457__bF$buf1 ;
wire _5457__bF$buf2 ;
wire _5457__bF$buf3 ;
wire _5457__bF$buf4 ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6511_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf2  ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf2  ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _3674_ ;
wire _3254_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf1  ;
wire ALUSrcA ;
wire [1:0] ALUSrcB ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf5  ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6414_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf1  ;
wire _1834_ ;
wire _1414_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf4  ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6452_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf1  ;
wire _5723_ ;
wire _5303_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf4  ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf6  ;
wire PCSource_1_bF$buf0 ;
wire _1032_ ;
wire PCSource_1_bF$buf1 ;
wire PCSource_1_bF$buf2 ;
wire PCSource_1_bF$buf3 ;
wire PCSource_1_bF$buf4 ;
wire [31:0] _783_ ;
wire _363_ ;
wire _2362__bF$buf0 ;
wire _2657_ ;
wire _2362__bF$buf1 ;
wire _2237_ ;
wire _2362__bF$buf2 ;
wire _2362__bF$buf3 ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire \datapath_1.PCJump_17_bF$buf0  ;
wire _4612_ ;
wire _5817_ ;
wire _3889__bF$buf0 ;
wire _3889__bF$buf1 ;
wire _3889__bF$buf2 ;
wire _3889__bF$buf3 ;
wire _3889__bF$buf4 ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf4  ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf2  ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _3183__bF$buf0 ;
wire _3183__bF$buf1 ;
wire _5855_ ;
wire _3183__bF$buf2 ;
wire _5435_ ;
wire _3183__bF$buf3 ;
wire _5015_ ;
wire _3183__bF$buf4 ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf3  ;
wire _4706_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf0  ;
wire _3098_ ;
wire _5664_ ;
wire _5244_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf7  ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf3  ;
wire _1678_ ;
wire _1258_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire BranchNe ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf2  ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6411_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire ALUZero ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire [31:0] _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf1  ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf1  ;
wire _58_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf5  ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf3  ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6543_ ;
wire _6123_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf4  ;
wire _3904__bF$buf0 ;
wire _3904__bF$buf1 ;
wire _3904__bF$buf2 ;
wire _3904__bF$buf3 ;
wire _3904__bF$buf4 ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire [31:0] \datapath_1.a  ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf1  ;
wire _6772_ ;
wire _6352_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf4  ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf6  ;
wire _2081_ ;
wire _2365__bF$buf0 ;
wire _2365__bF$buf1 ;
wire _2365__bF$buf2 ;
wire _2365__bF$buf3 ;
wire _2365__bF$buf4 ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire [31:0] _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf0  ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf4  ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _3186__bF$buf0 ;
wire _3186__bF$buf1 ;
wire _3186__bF$buf2 ;
wire _3186__bF$buf3 ;
wire _3186__bF$buf4 ;
wire _6484_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _3017__bF$buf0 ;
wire _3017__bF$buf1 ;
wire _3017__bF$buf2 ;
wire _3017__bF$buf3 ;
wire _3017__bF$buf4 ;
wire \datapath_1.mux_wd3.dout_3_bF$buf0  ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _3021__bF$buf0 ;
wire _3021__bF$buf1 ;
wire _3021__bF$buf2 ;
wire _3021__bF$buf3 ;
wire _3021__bF$buf4 ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire \datapath_1.PCJump_27_bF$buf3  ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _3923__bF$buf0 ;
wire _3923__bF$buf1 ;
wire _3923__bF$buf2 ;
wire _3923__bF$buf3 ;
wire _3923__bF$buf4 ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf3  ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf2  ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf6  ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [31:0] ALUOut ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf2  ;
wire _55_ ;
wire _6502_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _5471__bF$buf0 ;
wire _5471__bF$buf1 ;
wire _5471__bF$buf2 ;
wire _5471__bF$buf3 ;
wire _5471__bF$buf4 ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf2  ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf0  ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf1  ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire [31:0] \datapath_1.alu_1.ALUInA  ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf1  ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf5  ;
wire \datapath_1.regfile_1.regEn_5_bF$buf3  ;
wire ALUSrcB_1_bF$buf0 ;
wire ALUSrcB_1_bF$buf1 ;
wire ALUSrcB_1_bF$buf2 ;
wire ALUSrcB_1_bF$buf3 ;
wire ALUSrcB_1_bF$buf4 ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6443_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf1  ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf4  ;
wire _5714_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf4  ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _2368__bF$buf0 ;
wire _2368__bF$buf1 ;
wire _2368__bF$buf2 ;
wire _2368__bF$buf3 ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire [31:0] \datapath_1.regfile_1.regOut[3]  ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire \datapath_1.PCJump_27_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_1_bF$buf4  ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire [1:0] PCSource ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _3899__bF$buf0 ;
wire _3899__bF$buf1 ;
wire _3899__bF$buf2 ;
wire _3899__bF$buf3 ;
wire _3899__bF$buf4 ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf0  ;
wire _3089_ ;
wire _5455__bF$buf0 ;
wire _5455__bF$buf1 ;
wire _5455__bF$buf2 ;
wire _5455__bF$buf3 ;
wire _5455__bF$buf4 ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire [3:0] ALUControl ;
wire _5655_ ;
wire _5235_ ;
wire [31:0] \datapath_1.regfile_1.regOut[26]  ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf3  ;
wire _14_ ;
wire _4062__bF$buf0 ;
wire _4062__bF$buf1 ;
wire _4062__bF$buf2 ;
wire _4062__bF$buf3 ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf3  ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf2  ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf6  ;
wire _1287_ ;
wire [31:0] _198_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf2  ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6402_ ;
wire _2742_ ;
wire _2322_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf2  ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf0  ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6440_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf1  ;
wire _5711_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf5  ;
wire _3794_ ;
wire _3374_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf1  ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire \datapath_1.PCJump_22_bF$buf1  ;
wire MemToReg_bF$buf0 ;
wire MemToReg_bF$buf1 ;
wire MemToReg_bF$buf2 ;
wire MemToReg_bF$buf3 ;
wire MemToReg_bF$buf4 ;
wire MemToReg_bF$buf5 ;
wire MemToReg_bF$buf6 ;
wire MemToReg_bF$buf7 ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf5  ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _3181__bF$buf0 ;
wire _3181__bF$buf1 ;
wire _3181__bF$buf2 ;
wire _3181__bF$buf3 ;
wire _3181__bF$buf4 ;
wire _87_ ;
wire _6534_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf4  ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf1  ;
wire _6763_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf5  ;
wire _5614_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6572_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _5708_ ;
wire [31:0] _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf0  ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf0  ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _4770_ ;
wire _4350_ ;
wire _3929__bF$buf0 ;
wire _3929__bF$buf1 ;
wire _3929__bF$buf2 ;
wire _3929__bF$buf3 ;
wire _3929__bF$buf4 ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire [31:0] \datapath_1.regfile_1.regOut[16]  ;
wire _5462__bF$buf0 ;
wire _5462__bF$buf1 ;
wire _5462__bF$buf2 ;
wire _5462__bF$buf3 ;
wire _5462__bF$buf4 ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire clk_bF$buf90 ;
wire clk_bF$buf91 ;
wire clk_bF$buf92 ;
wire clk_bF$buf93 ;
wire clk_bF$buf94 ;
wire clk_bF$buf95 ;
wire clk_bF$buf96 ;
wire _3621_ ;
wire clk_bF$buf97 ;
wire _3201_ ;
wire clk_bF$buf98 ;
wire clk_bF$buf99 ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _5784_ ;
wire _5364_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf3  ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _5560__bF$buf0 ;
wire _5560__bF$buf1 ;
wire _5560__bF$buf2 ;
wire _5560__bF$buf3 ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf2  ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf6  ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf2  ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf6  ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf2  ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf2  ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6531_ ;
wire _6111_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf1  ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf2  ;
wire _5611_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf5  ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6434_ ;
wire _6014_ ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5705_ ;
wire [31:0] \datapath_1.regfile_1.regOut[31]  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6472_ ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf3  ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire [31:0] _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf0  ;
wire _859_ ;
wire _439_ ;
wire _6566_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf3  ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire IRWrite ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _5465__bF$buf0 ;
wire _5465__bF$buf1 ;
wire _5465__bF$buf2 ;
wire _5465__bF$buf3 ;
wire _5465__bF$buf4 ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf3  ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire [31:0] _2_ ;
wire _5563__bF$buf0 ;
wire _5563__bF$buf1 ;
wire _5563__bF$buf2 ;
wire _4726_ ;
wire _5563__bF$buf3 ;
wire _4306_ ;
wire _4068__bF$buf0 ;
wire _4068__bF$buf1 ;
wire _4068__bF$buf2 ;
wire _4068__bF$buf3 ;
wire _5684_ ;
wire _5264_ ;
wire _3940__bF$buf0 ;
wire _3940__bF$buf1 ;
wire _3940__bF$buf2 ;
wire _3940__bF$buf3 ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf3  ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire rst_hier0_bF$buf0 ;
wire rst_hier0_bF$buf1 ;
wire rst_hier0_bF$buf2 ;
wire rst_hier0_bF$buf3 ;
wire rst_hier0_bF$buf4 ;
wire rst_hier0_bF$buf5 ;
wire rst_hier0_bF$buf6 ;
wire rst_hier0_bF$buf7 ;
wire rst_hier0_bF$buf8 ;
wire rst_hier0_bF$buf9 ;
wire \datapath_1.mux_wd3.dout_24_bF$buf2  ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf3  ;
wire _4629_ ;
wire _4209_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf6  ;
wire ALUSrcB_0_bF$buf0 ;
wire ALUSrcB_0_bF$buf1 ;
wire ALUSrcB_0_bF$buf2 ;
wire ALUSrcB_0_bF$buf3 ;
wire ALUSrcB_0_bF$buf4 ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf2  ;
wire _2733_ ;
wire _2313_ ;
wire _5484__bF$buf0 ;
wire _5484__bF$buf1 ;
wire _5484__bF$buf2 ;
wire _5484__bF$buf3 ;
wire _5484__bF$buf4 ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf6  ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire [3:0] \control_1.next  ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6431_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire ALUSrcA_bF$buf0 ;
wire _533_ ;
wire ALUSrcA_bF$buf1 ;
wire _113_ ;
wire ALUSrcA_bF$buf2 ;
wire ALUSrcA_bF$buf3 ;
wire ALUSrcA_bF$buf4 ;
wire ALUSrcA_bF$buf5 ;
wire ALUSrcA_bF$buf6 ;
wire _2827_ ;
wire ALUSrcA_bF$buf7 ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf0  ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _3924__bF$buf0 ;
wire _3924__bF$buf1 ;
wire _3924__bF$buf2 ;
wire _3924__bF$buf3 ;
wire _5605_ ;
wire [31:0] \datapath_1.regfile_1.regOut[21]  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6563_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf0  ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf3  ;
wire _5643_ ;
wire _5223_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire [31:0] _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf0  ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf6  ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf0  ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _3939__bF$buf0 ;
wire _3939__bF$buf1 ;
wire _3939__bF$buf2 ;
wire _3939__bF$buf3 ;
wire _3939__bF$buf4 ;
wire _5472__bF$buf0 ;
wire _5472__bF$buf1 ;
wire _5472__bF$buf2 ;
wire _5472__bF$buf3 ;
wire _5472__bF$buf4 ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf0  ;
wire _4626_ ;
wire _4206_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf3  ;
wire _5584_ ;
wire _5164_ ;
wire _6369_ ;
wire _1084_ ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf7  ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf2  ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf3  ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf6  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf2  ;
wire _1598_ ;
wire _1178_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf6  ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire rst_bF$buf70 ;
wire rst_bF$buf71 ;
wire rst_bF$buf72 ;
wire rst_bF$buf73 ;
wire rst_bF$buf74 ;
wire rst_bF$buf75 ;
wire rst_bF$buf76 ;
wire rst_bF$buf77 ;
wire rst_bF$buf78 ;
wire rst_bF$buf79 ;
wire [31:0] \datapath_1.regfile_1.regEn  ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf6  ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6522_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6751_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf4  ;
wire _5602_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6560_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _3494_ ;
wire _3074_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf0  ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire [31:0] _718_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire [31:0] \datapath_1.regfile_1.regOut[11]  ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf3  ;
wire _6463_ ;
wire _6043_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire [31:0] _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf2  ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf6  ;
wire _4623_ ;
wire _4203_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf0  ;
wire [31:0] \datapath_1.regfile_1.regOut[5]  ;
wire _5828_ ;
wire _5408_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf3  ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf4  ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire [31:0] \datapath_1.ALUResult  ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf0  ;
wire _5675_ ;
wire _5255_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf3  ;
wire [31:0] \datapath_1.regfile_1.regOut[28]  ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _3950__bF$buf0 ;
wire _3950__bF$buf1 ;
wire _3950__bF$buf2 ;
wire _3950__bF$buf3 ;
wire \datapath_1.regfile_1.regEn_4_bF$buf7  ;
wire \datapath_1.regfile_1.regEn_31_bF$buf3  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire rst_bF$buf40 ;
wire rst_bF$buf41 ;
wire rst_bF$buf42 ;
wire rst_bF$buf43 ;
wire rst_bF$buf44 ;
wire rst_bF$buf45 ;
wire rst_bF$buf46 ;
wire rst_bF$buf47 ;
wire rst_bF$buf48 ;
wire rst_bF$buf49 ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _1689_ ;
wire _1269_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf3  ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire [31:0] _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [31:0] memoryAddress ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf1  ;
wire _4658_ ;
wire _4238_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire PCEn ;
wire _906_ ;
wire _6613_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6422_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _5423__bF$buf0 ;
wire _5423__bF$buf1 ;
wire _5423__bF$buf2 ;
wire _5423__bF$buf3 ;
wire \datapath_1.mux_wd3.dout_5_bF$buf4  ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf0  ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6460_ ;
wire _6040_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf3  ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf7  ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire [31:0] \datapath_1.PCJump  ;
wire _6554_ ;
wire _6134_ ;
wire _3934__bF$buf0 ;
wire _3934__bF$buf1 ;
wire _3934__bF$buf2 ;
wire _3934__bF$buf3 ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf3  ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5561__bF$buf0 ;
wire _5561__bF$buf1 ;
wire _5561__bF$buf2 ;
wire _5561__bF$buf3 ;
wire _5825_ ;
wire _5405_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf0  ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6363_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf1  ;
wire _5634_ ;
wire _5214_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf2  ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf6  ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf0  ;
wire _6457_ ;
wire _6037_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf3  ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf6  ;
wire _5728_ ;
wire _5308_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf4  ;
wire _1648_ ;
wire _1228_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf0  ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire rst_bF$buf10 ;
wire rst_bF$buf11 ;
wire rst_bF$buf12 ;
wire rst_bF$buf13 ;
wire rst_bF$buf14 ;
wire rst_bF$buf15 ;
wire rst_bF$buf16 ;
wire rst_bF$buf17 ;
wire rst_bF$buf18 ;
wire rst_bF$buf19 ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _5478__bF$buf0 ;
wire _5478__bF$buf1 ;
wire _5478__bF$buf2 ;
wire _5478__bF$buf3 ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf0  ;
wire _597_ ;
wire _177_ ;
wire _5482__bF$buf0 ;
wire _3832_ ;
wire _5482__bF$buf1 ;
wire _3412_ ;
wire _5482__bF$buf2 ;
wire _5482__bF$buf3 ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire [31:0] \datapath_1.regfile_1.regOut[18]  ;
wire _1495_ ;
wire _1075_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf7  ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf1  ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire [31:0] \datapath_1.mux_iord.din0  ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _6704_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf0  ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6513_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf4  ;
wire _3638_ ;
wire _3218_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire _2477__bF$buf0 ;
wire _2477__bF$buf1 ;
wire _2477__bF$buf2 ;
wire _2477__bF$buf3 ;
wire \datapath_1.mux_wd3.dout_8_bF$buf4  ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6551_ ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf0  ;
wire _3676_ ;
wire _3256_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf3  ;
wire _5822_ ;
wire _5402_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire [31:0] _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6360_ ;
wire _2280_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf7  ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf3  ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6454_ ;
wire _6034_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf0  ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf3  ;
wire _5725_ ;
wire _5305_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf1  ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire \datapath_1.PCJump_17_bF$buf2  ;
wire _4614_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf6  ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf4  ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf2  ;
wire _5485__bF$buf0 ;
wire _5485__bF$buf1 ;
wire _5485__bF$buf2 ;
wire _5485__bF$buf3 ;
wire _5485__bF$buf4 ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _3956__bF$buf0 ;
wire _3956__bF$buf1 ;
wire _3956__bF$buf2 ;
wire _3956__bF$buf3 ;
wire _3956__bF$buf4 ;
wire _4937_ ;
wire _4517_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf1  ;
wire _3635_ ;
wire _3215_ ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf1  ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _3673_ ;
wire _3253_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf0  ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _6604_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf4  ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6413_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5433__bF$buf0 ;
wire _5433__bF$buf1 ;
wire _5433__bF$buf2 ;
wire _5433__bF$buf3 ;
wire _5433__bF$buf4 ;
wire _5913_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf0  ;
wire _1833_ ;
wire _1413_ ;
wire IorD_bF$buf0 ;
wire IorD_bF$buf1 ;
wire IorD_bF$buf2 ;
wire IorD_bF$buf3 ;
wire IorD_bF$buf4 ;
wire \datapath_1.mux_wd3.dout_16_bF$buf3  ;
wire IorD_bF$buf5 ;
wire IorD_bF$buf6 ;
wire IorD_bF$buf7 ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6451_ ;
wire _6031_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf0  ;
wire _5722_ ;
wire _5302_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf7  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf3  ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire [31:0] _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _2180_ ;
wire [31:0] \datapath_1.regfile_1.regOut[0]  ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf7  ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf5  ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire [31:0] \datapath_1.rd2  ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _3944__bF$buf0 ;
wire _3944__bF$buf1 ;
wire _3944__bF$buf2 ;
wire _3944__bF$buf3 ;
wire _647_ ;
wire _227_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf3  ;
wire _6774_ ;
wire _6354_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf1  ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire [31:0] \datapath_1.regfile_1.regOut[23]  ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire [31:0] memoryOutData ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire [1:0] ALUOp ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf2  ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf6  ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;

BUFX2 BUFX2_insert1100 (
    .A(rst),
    .Y(rst_hier0_bF$buf0)
);

BUFX2 BUFX2_insert1099 (
    .A(rst),
    .Y(rst_hier0_bF$buf1)
);

BUFX2 BUFX2_insert1098 (
    .A(rst),
    .Y(rst_hier0_bF$buf2)
);

BUFX2 BUFX2_insert1097 (
    .A(rst),
    .Y(rst_hier0_bF$buf3)
);

BUFX2 BUFX2_insert1096 (
    .A(rst),
    .Y(rst_hier0_bF$buf4)
);

BUFX2 BUFX2_insert1095 (
    .A(rst),
    .Y(rst_hier0_bF$buf5)
);

BUFX2 BUFX2_insert1094 (
    .A(rst),
    .Y(rst_hier0_bF$buf6)
);

BUFX2 BUFX2_insert1093 (
    .A(rst),
    .Y(rst_hier0_bF$buf7)
);

BUFX2 BUFX2_insert1092 (
    .A(rst),
    .Y(rst_hier0_bF$buf8)
);

BUFX2 BUFX2_insert1091 (
    .A(rst),
    .Y(rst_hier0_bF$buf9)
);

CLKBUF1 CLKBUF1_insert1090 (
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert1089 (
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert1088 (
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1087 (
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1086 (
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1085 (
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1084 (
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1083 (
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

CLKBUF1 CLKBUF1_insert1082 (
    .A(clk),
    .Y(clk_hier0_bF$buf8)
);

CLKBUF1 CLKBUF1_insert1081 (
    .A(clk),
    .Y(clk_hier0_bF$buf9)
);

BUFX2 BUFX2_insert1080 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf0 )
);

BUFX2 BUFX2_insert1079 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf1 )
);

BUFX2 BUFX2_insert1078 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf2 )
);

BUFX2 BUFX2_insert1077 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf3 )
);

BUFX2 BUFX2_insert1076 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf4 )
);

BUFX2 BUFX2_insert1075 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf5 )
);

BUFX2 BUFX2_insert1074 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf6 )
);

BUFX2 BUFX2_insert1073 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf7 )
);

BUFX2 BUFX2_insert1072 (
    .A(_5472_),
    .Y(_5472__bF$buf0)
);

BUFX2 BUFX2_insert1071 (
    .A(_5472_),
    .Y(_5472__bF$buf1)
);

BUFX2 BUFX2_insert1070 (
    .A(_5472_),
    .Y(_5472__bF$buf2)
);

BUFX2 BUFX2_insert1069 (
    .A(_5472_),
    .Y(_5472__bF$buf3)
);

BUFX2 BUFX2_insert1068 (
    .A(_5472_),
    .Y(_5472__bF$buf4)
);

BUFX2 BUFX2_insert1067 (
    .A(_2368_),
    .Y(_2368__bF$buf0)
);

BUFX2 BUFX2_insert1066 (
    .A(_2368_),
    .Y(_2368__bF$buf1)
);

BUFX2 BUFX2_insert1065 (
    .A(_2368_),
    .Y(_2368__bF$buf2)
);

BUFX2 BUFX2_insert1064 (
    .A(_2368_),
    .Y(_2368__bF$buf3)
);

BUFX2 BUFX2_insert1063 (
    .A(_3899_),
    .Y(_3899__bF$buf0)
);

BUFX2 BUFX2_insert1062 (
    .A(_3899_),
    .Y(_3899__bF$buf1)
);

BUFX2 BUFX2_insert1061 (
    .A(_3899_),
    .Y(_3899__bF$buf2)
);

BUFX2 BUFX2_insert1060 (
    .A(_3899_),
    .Y(_3899__bF$buf3)
);

BUFX2 BUFX2_insert1059 (
    .A(_3899_),
    .Y(_3899__bF$buf4)
);

BUFX2 BUFX2_insert1058 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf0 )
);

BUFX2 BUFX2_insert1057 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf1 )
);

BUFX2 BUFX2_insert1056 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf2 )
);

BUFX2 BUFX2_insert1055 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf3 )
);

BUFX2 BUFX2_insert1054 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf4 )
);

BUFX2 BUFX2_insert1053 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf0 )
);

BUFX2 BUFX2_insert1052 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf1 )
);

BUFX2 BUFX2_insert1051 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf2 )
);

BUFX2 BUFX2_insert1050 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf3 )
);

BUFX2 BUFX2_insert1049 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf4 )
);

BUFX2 BUFX2_insert1048 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf5 )
);

BUFX2 BUFX2_insert1047 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf6 )
);

BUFX2 BUFX2_insert1046 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf7 )
);

BUFX2 BUFX2_insert1045 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf0 )
);

BUFX2 BUFX2_insert1044 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf1 )
);

BUFX2 BUFX2_insert1043 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf2 )
);

BUFX2 BUFX2_insert1042 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf3 )
);

BUFX2 BUFX2_insert1041 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf4 )
);

BUFX2 BUFX2_insert1040 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf0 )
);

BUFX2 BUFX2_insert1039 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf1 )
);

BUFX2 BUFX2_insert1038 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf2 )
);

BUFX2 BUFX2_insert1037 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf3 )
);

BUFX2 BUFX2_insert1036 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf4 )
);

BUFX2 BUFX2_insert1035 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf5 )
);

BUFX2 BUFX2_insert1034 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf6 )
);

BUFX2 BUFX2_insert1033 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf7 )
);

BUFX2 BUFX2_insert1032 (
    .A(_3961_),
    .Y(_3961__bF$buf0)
);

BUFX2 BUFX2_insert1031 (
    .A(_3961_),
    .Y(_3961__bF$buf1)
);

BUFX2 BUFX2_insert1030 (
    .A(_3961_),
    .Y(_3961__bF$buf2)
);

BUFX2 BUFX2_insert1029 (
    .A(_3961_),
    .Y(_3961__bF$buf3)
);

BUFX2 BUFX2_insert1028 (
    .A(_3961_),
    .Y(_3961__bF$buf4)
);

BUFX2 BUFX2_insert1027 (
    .A(_3923_),
    .Y(_3923__bF$buf0)
);

BUFX2 BUFX2_insert1026 (
    .A(_3923_),
    .Y(_3923__bF$buf1)
);

BUFX2 BUFX2_insert1025 (
    .A(_3923_),
    .Y(_3923__bF$buf2)
);

BUFX2 BUFX2_insert1024 (
    .A(_3923_),
    .Y(_3923__bF$buf3)
);

BUFX2 BUFX2_insert1023 (
    .A(_3923_),
    .Y(_3923__bF$buf4)
);

BUFX2 BUFX2_insert1022 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf0 )
);

BUFX2 BUFX2_insert1021 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf1 )
);

BUFX2 BUFX2_insert1020 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf2 )
);

BUFX2 BUFX2_insert1019 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf3 )
);

BUFX2 BUFX2_insert1018 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf4 )
);

BUFX2 BUFX2_insert1017 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf5 )
);

BUFX2 BUFX2_insert1016 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf6 )
);

BUFX2 BUFX2_insert1015 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf7 )
);

BUFX2 BUFX2_insert1014 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf0)
);

BUFX2 BUFX2_insert1013 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf1)
);

BUFX2 BUFX2_insert1012 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf2)
);

BUFX2 BUFX2_insert1011 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf3)
);

BUFX2 BUFX2_insert1010 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf4)
);

BUFX2 BUFX2_insert1009 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf0 )
);

BUFX2 BUFX2_insert1008 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf1 )
);

BUFX2 BUFX2_insert1007 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf2 )
);

BUFX2 BUFX2_insert1006 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf3 )
);

BUFX2 BUFX2_insert1005 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf4 )
);

BUFX2 BUFX2_insert1004 (
    .A(_5478_),
    .Y(_5478__bF$buf0)
);

BUFX2 BUFX2_insert1003 (
    .A(_5478_),
    .Y(_5478__bF$buf1)
);

BUFX2 BUFX2_insert1002 (
    .A(_5478_),
    .Y(_5478__bF$buf2)
);

BUFX2 BUFX2_insert1001 (
    .A(_5478_),
    .Y(_5478__bF$buf3)
);

BUFX2 BUFX2_insert1000 (
    .A(_3870_),
    .Y(_3870__bF$buf0)
);

BUFX2 BUFX2_insert999 (
    .A(_3870_),
    .Y(_3870__bF$buf1)
);

BUFX2 BUFX2_insert998 (
    .A(_3870_),
    .Y(_3870__bF$buf2)
);

BUFX2 BUFX2_insert997 (
    .A(_3870_),
    .Y(_3870__bF$buf3)
);

BUFX2 BUFX2_insert996 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf0 )
);

BUFX2 BUFX2_insert995 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf1 )
);

BUFX2 BUFX2_insert994 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf2 )
);

BUFX2 BUFX2_insert993 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf3 )
);

BUFX2 BUFX2_insert992 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf4 )
);

BUFX2 BUFX2_insert991 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf0 )
);

BUFX2 BUFX2_insert990 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf1 )
);

BUFX2 BUFX2_insert989 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf2 )
);

BUFX2 BUFX2_insert988 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf3 )
);

BUFX2 BUFX2_insert987 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf4 )
);

BUFX2 BUFX2_insert986 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf5 )
);

BUFX2 BUFX2_insert985 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf6 )
);

BUFX2 BUFX2_insert984 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf7 )
);

BUFX2 BUFX2_insert983 (
    .A(PCEn),
    .Y(PCEn_bF$buf0)
);

BUFX2 BUFX2_insert982 (
    .A(PCEn),
    .Y(PCEn_bF$buf1)
);

BUFX2 BUFX2_insert981 (
    .A(PCEn),
    .Y(PCEn_bF$buf2)
);

BUFX2 BUFX2_insert980 (
    .A(PCEn),
    .Y(PCEn_bF$buf3)
);

BUFX2 BUFX2_insert979 (
    .A(PCEn),
    .Y(PCEn_bF$buf4)
);

BUFX2 BUFX2_insert978 (
    .A(PCEn),
    .Y(PCEn_bF$buf5)
);

BUFX2 BUFX2_insert977 (
    .A(PCEn),
    .Y(PCEn_bF$buf6)
);

BUFX2 BUFX2_insert976 (
    .A(PCEn),
    .Y(PCEn_bF$buf7)
);

BUFX2 BUFX2_insert975 (
    .A(_3929_),
    .Y(_3929__bF$buf0)
);

BUFX2 BUFX2_insert974 (
    .A(_3929_),
    .Y(_3929__bF$buf1)
);

BUFX2 BUFX2_insert973 (
    .A(_3929_),
    .Y(_3929__bF$buf2)
);

BUFX2 BUFX2_insert972 (
    .A(_3929_),
    .Y(_3929__bF$buf3)
);

BUFX2 BUFX2_insert971 (
    .A(_3929_),
    .Y(_3929__bF$buf4)
);

BUFX2 BUFX2_insert970 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf0 )
);

BUFX2 BUFX2_insert969 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf1 )
);

BUFX2 BUFX2_insert968 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf2 )
);

BUFX2 BUFX2_insert967 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf3 )
);

BUFX2 BUFX2_insert966 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf4 )
);

BUFX2 BUFX2_insert965 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf0 )
);

BUFX2 BUFX2_insert964 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf1 )
);

BUFX2 BUFX2_insert963 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf2 )
);

BUFX2 BUFX2_insert962 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf3 )
);

BUFX2 BUFX2_insert961 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf4 )
);

BUFX2 BUFX2_insert960 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf5 )
);

BUFX2 BUFX2_insert959 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf6 )
);

BUFX2 BUFX2_insert958 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf7 )
);

BUFX2 BUFX2_insert957 (
    .A(_5484_),
    .Y(_5484__bF$buf0)
);

BUFX2 BUFX2_insert956 (
    .A(_5484_),
    .Y(_5484__bF$buf1)
);

BUFX2 BUFX2_insert955 (
    .A(_5484_),
    .Y(_5484__bF$buf2)
);

BUFX2 BUFX2_insert954 (
    .A(_5484_),
    .Y(_5484__bF$buf3)
);

BUFX2 BUFX2_insert953 (
    .A(_5484_),
    .Y(_5484__bF$buf4)
);

BUFX2 BUFX2_insert952 (
    .A(_2477_),
    .Y(_2477__bF$buf0)
);

BUFX2 BUFX2_insert951 (
    .A(_2477_),
    .Y(_2477__bF$buf1)
);

BUFX2 BUFX2_insert950 (
    .A(_2477_),
    .Y(_2477__bF$buf2)
);

BUFX2 BUFX2_insert949 (
    .A(_2477_),
    .Y(_2477__bF$buf3)
);

BUFX2 BUFX2_insert948 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf0 )
);

BUFX2 BUFX2_insert947 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf1 )
);

BUFX2 BUFX2_insert946 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf2 )
);

BUFX2 BUFX2_insert945 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf3 )
);

BUFX2 BUFX2_insert944 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf4 )
);

BUFX2 BUFX2_insert943 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf5 )
);

BUFX2 BUFX2_insert942 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf6 )
);

BUFX2 BUFX2_insert941 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf7 )
);

BUFX2 BUFX2_insert940 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf0 )
);

BUFX2 BUFX2_insert939 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf1 )
);

BUFX2 BUFX2_insert938 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf2 )
);

BUFX2 BUFX2_insert937 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf3 )
);

BUFX2 BUFX2_insert936 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf4 )
);

BUFX2 BUFX2_insert935 (
    .A(_3935_),
    .Y(_3935__bF$buf0)
);

BUFX2 BUFX2_insert934 (
    .A(_3935_),
    .Y(_3935__bF$buf1)
);

BUFX2 BUFX2_insert933 (
    .A(_3935_),
    .Y(_3935__bF$buf2)
);

BUFX2 BUFX2_insert932 (
    .A(_3935_),
    .Y(_3935__bF$buf3)
);

BUFX2 BUFX2_insert931 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf0 )
);

BUFX2 BUFX2_insert930 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf1 )
);

BUFX2 BUFX2_insert929 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf2 )
);

BUFX2 BUFX2_insert928 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf3 )
);

BUFX2 BUFX2_insert927 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf4 )
);

BUFX2 BUFX2_insert926 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf0 )
);

BUFX2 BUFX2_insert925 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf1 )
);

BUFX2 BUFX2_insert924 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf2 )
);

BUFX2 BUFX2_insert923 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf3 )
);

BUFX2 BUFX2_insert922 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf4 )
);

BUFX2 BUFX2_insert921 (
    .A(_3879_),
    .Y(_3879__bF$buf0)
);

BUFX2 BUFX2_insert920 (
    .A(_3879_),
    .Y(_3879__bF$buf1)
);

BUFX2 BUFX2_insert919 (
    .A(_3879_),
    .Y(_3879__bF$buf2)
);

BUFX2 BUFX2_insert918 (
    .A(_3879_),
    .Y(_3879__bF$buf3)
);

BUFX2 BUFX2_insert917 (
    .A(_5511_),
    .Y(_5511__bF$buf0)
);

BUFX2 BUFX2_insert916 (
    .A(_5511_),
    .Y(_5511__bF$buf1)
);

BUFX2 BUFX2_insert915 (
    .A(_5511_),
    .Y(_5511__bF$buf2)
);

BUFX2 BUFX2_insert914 (
    .A(_5511_),
    .Y(_5511__bF$buf3)
);

BUFX2 BUFX2_insert913 (
    .A(_5511_),
    .Y(_5511__bF$buf4)
);

BUFX2 BUFX2_insert912 (
    .A(_5493_),
    .Y(_5493__bF$buf0)
);

BUFX2 BUFX2_insert911 (
    .A(_5493_),
    .Y(_5493__bF$buf1)
);

BUFX2 BUFX2_insert910 (
    .A(_5493_),
    .Y(_5493__bF$buf2)
);

BUFX2 BUFX2_insert909 (
    .A(_5493_),
    .Y(_5493__bF$buf3)
);

BUFX2 BUFX2_insert908 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf0 )
);

BUFX2 BUFX2_insert907 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf1 )
);

BUFX2 BUFX2_insert906 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf2 )
);

BUFX2 BUFX2_insert905 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf3 )
);

BUFX2 BUFX2_insert904 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf4 )
);

BUFX2 BUFX2_insert903 (
    .A(_5455_),
    .Y(_5455__bF$buf0)
);

BUFX2 BUFX2_insert902 (
    .A(_5455_),
    .Y(_5455__bF$buf1)
);

BUFX2 BUFX2_insert901 (
    .A(_5455_),
    .Y(_5455__bF$buf2)
);

BUFX2 BUFX2_insert900 (
    .A(_5455_),
    .Y(_5455__bF$buf3)
);

BUFX2 BUFX2_insert899 (
    .A(_5455_),
    .Y(_5455__bF$buf4)
);

BUFX2 BUFX2_insert898 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf0)
);

BUFX2 BUFX2_insert897 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf1)
);

BUFX2 BUFX2_insert896 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf2)
);

BUFX2 BUFX2_insert895 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf3)
);

BUFX2 BUFX2_insert894 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf4)
);

BUFX2 BUFX2_insert893 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf5)
);

BUFX2 BUFX2_insert892 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf6)
);

BUFX2 BUFX2_insert891 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf7)
);

BUFX2 BUFX2_insert890 (
    .A(_5514_),
    .Y(_5514__bF$buf0)
);

BUFX2 BUFX2_insert889 (
    .A(_5514_),
    .Y(_5514__bF$buf1)
);

BUFX2 BUFX2_insert888 (
    .A(_5514_),
    .Y(_5514__bF$buf2)
);

BUFX2 BUFX2_insert887 (
    .A(_5514_),
    .Y(_5514__bF$buf3)
);

BUFX2 BUFX2_insert886 (
    .A(_5514_),
    .Y(_5514__bF$buf4)
);

BUFX2 BUFX2_insert885 (
    .A(_2354_),
    .Y(_2354__bF$buf0)
);

BUFX2 BUFX2_insert884 (
    .A(_2354_),
    .Y(_2354__bF$buf1)
);

BUFX2 BUFX2_insert883 (
    .A(_2354_),
    .Y(_2354__bF$buf2)
);

BUFX2 BUFX2_insert882 (
    .A(_2354_),
    .Y(_2354__bF$buf3)
);

BUFX2 BUFX2_insert881 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf0 )
);

BUFX2 BUFX2_insert880 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf1 )
);

BUFX2 BUFX2_insert879 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf2 )
);

BUFX2 BUFX2_insert878 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf3 )
);

BUFX2 BUFX2_insert877 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf4 )
);

BUFX2 BUFX2_insert876 (
    .A(_4062_),
    .Y(_4062__bF$buf0)
);

BUFX2 BUFX2_insert875 (
    .A(_4062_),
    .Y(_4062__bF$buf1)
);

BUFX2 BUFX2_insert874 (
    .A(_4062_),
    .Y(_4062__bF$buf2)
);

BUFX2 BUFX2_insert873 (
    .A(_4062_),
    .Y(_4062__bF$buf3)
);

BUFX2 BUFX2_insert872 (
    .A(_3944_),
    .Y(_3944__bF$buf0)
);

BUFX2 BUFX2_insert871 (
    .A(_3944_),
    .Y(_3944__bF$buf1)
);

BUFX2 BUFX2_insert870 (
    .A(_3944_),
    .Y(_3944__bF$buf2)
);

BUFX2 BUFX2_insert869 (
    .A(_3944_),
    .Y(_3944__bF$buf3)
);

BUFX2 BUFX2_insert868 (
    .A(_3906_),
    .Y(_3906__bF$buf0)
);

BUFX2 BUFX2_insert867 (
    .A(_3906_),
    .Y(_3906__bF$buf1)
);

BUFX2 BUFX2_insert866 (
    .A(_3906_),
    .Y(_3906__bF$buf2)
);

BUFX2 BUFX2_insert865 (
    .A(_3906_),
    .Y(_3906__bF$buf3)
);

BUFX2 BUFX2_insert864 (
    .A(_5555_),
    .Y(_5555__bF$buf0)
);

BUFX2 BUFX2_insert863 (
    .A(_5555_),
    .Y(_5555__bF$buf1)
);

BUFX2 BUFX2_insert862 (
    .A(_5555_),
    .Y(_5555__bF$buf2)
);

BUFX2 BUFX2_insert861 (
    .A(_5555_),
    .Y(_5555__bF$buf3)
);

BUFX2 BUFX2_insert860 (
    .A(_5517_),
    .Y(_5517__bF$buf0)
);

BUFX2 BUFX2_insert859 (
    .A(_5517_),
    .Y(_5517__bF$buf1)
);

BUFX2 BUFX2_insert858 (
    .A(_5517_),
    .Y(_5517__bF$buf2)
);

BUFX2 BUFX2_insert857 (
    .A(_5517_),
    .Y(_5517__bF$buf3)
);

BUFX2 BUFX2_insert856 (
    .A(_5517_),
    .Y(_5517__bF$buf4)
);

BUFX2 BUFX2_insert855 (
    .A(_5423_),
    .Y(_5423__bF$buf0)
);

BUFX2 BUFX2_insert854 (
    .A(_5423_),
    .Y(_5423__bF$buf1)
);

BUFX2 BUFX2_insert853 (
    .A(_5423_),
    .Y(_5423__bF$buf2)
);

BUFX2 BUFX2_insert852 (
    .A(_5423_),
    .Y(_5423__bF$buf3)
);

BUFX2 BUFX2_insert851 (
    .A(_3183_),
    .Y(_3183__bF$buf0)
);

BUFX2 BUFX2_insert850 (
    .A(_3183_),
    .Y(_3183__bF$buf1)
);

BUFX2 BUFX2_insert849 (
    .A(_3183_),
    .Y(_3183__bF$buf2)
);

BUFX2 BUFX2_insert848 (
    .A(_3183_),
    .Y(_3183__bF$buf3)
);

BUFX2 BUFX2_insert847 (
    .A(_3183_),
    .Y(_3183__bF$buf4)
);

BUFX2 BUFX2_insert846 (
    .A(_5520_),
    .Y(_5520__bF$buf0)
);

BUFX2 BUFX2_insert845 (
    .A(_5520_),
    .Y(_5520__bF$buf1)
);

BUFX2 BUFX2_insert844 (
    .A(_5520_),
    .Y(_5520__bF$buf2)
);

BUFX2 BUFX2_insert843 (
    .A(_5520_),
    .Y(_5520__bF$buf3)
);

BUFX2 BUFX2_insert842 (
    .A(_5520_),
    .Y(_5520__bF$buf4)
);

BUFX2 BUFX2_insert841 (
    .A(_3947_),
    .Y(_3947__bF$buf0)
);

BUFX2 BUFX2_insert840 (
    .A(_3947_),
    .Y(_3947__bF$buf1)
);

BUFX2 BUFX2_insert839 (
    .A(_3947_),
    .Y(_3947__bF$buf2)
);

BUFX2 BUFX2_insert838 (
    .A(_3947_),
    .Y(_3947__bF$buf3)
);

BUFX2 BUFX2_insert837 (
    .A(_5558_),
    .Y(_5558__bF$buf0)
);

BUFX2 BUFX2_insert836 (
    .A(_5558_),
    .Y(_5558__bF$buf1)
);

BUFX2 BUFX2_insert835 (
    .A(_5558_),
    .Y(_5558__bF$buf2)
);

BUFX2 BUFX2_insert834 (
    .A(_5558_),
    .Y(_5558__bF$buf3)
);

BUFX2 BUFX2_insert833 (
    .A(_3950_),
    .Y(_3950__bF$buf0)
);

BUFX2 BUFX2_insert832 (
    .A(_3950_),
    .Y(_3950__bF$buf1)
);

BUFX2 BUFX2_insert831 (
    .A(_3950_),
    .Y(_3950__bF$buf2)
);

BUFX2 BUFX2_insert830 (
    .A(_3950_),
    .Y(_3950__bF$buf3)
);

BUFX2 BUFX2_insert829 (
    .A(_5561_),
    .Y(_5561__bF$buf0)
);

BUFX2 BUFX2_insert828 (
    .A(_5561_),
    .Y(_5561__bF$buf1)
);

BUFX2 BUFX2_insert827 (
    .A(_5561_),
    .Y(_5561__bF$buf2)
);

BUFX2 BUFX2_insert826 (
    .A(_5561_),
    .Y(_5561__bF$buf3)
);

BUFX2 BUFX2_insert825 (
    .A(_3186_),
    .Y(_3186__bF$buf0)
);

BUFX2 BUFX2_insert824 (
    .A(_3186_),
    .Y(_3186__bF$buf1)
);

BUFX2 BUFX2_insert823 (
    .A(_3186_),
    .Y(_3186__bF$buf2)
);

BUFX2 BUFX2_insert822 (
    .A(_3186_),
    .Y(_3186__bF$buf3)
);

BUFX2 BUFX2_insert821 (
    .A(_3186_),
    .Y(_3186__bF$buf4)
);

BUFX2 BUFX2_insert820 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf0 )
);

BUFX2 BUFX2_insert819 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf1 )
);

BUFX2 BUFX2_insert818 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf2 )
);

BUFX2 BUFX2_insert817 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf3 )
);

BUFX2 BUFX2_insert816 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf4 )
);

BUFX2 BUFX2_insert815 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf5 )
);

BUFX2 BUFX2_insert814 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf6 )
);

BUFX2 BUFX2_insert813 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf7 )
);

BUFX2 BUFX2_insert812 (
    .A(_4068_),
    .Y(_4068__bF$buf0)
);

BUFX2 BUFX2_insert811 (
    .A(_4068_),
    .Y(_4068__bF$buf1)
);

BUFX2 BUFX2_insert810 (
    .A(_4068_),
    .Y(_4068__bF$buf2)
);

BUFX2 BUFX2_insert809 (
    .A(_4068_),
    .Y(_4068__bF$buf3)
);

BUFX2 BUFX2_insert808 (
    .A(_3894_),
    .Y(_3894__bF$buf0)
);

BUFX2 BUFX2_insert807 (
    .A(_3894_),
    .Y(_3894__bF$buf1)
);

BUFX2 BUFX2_insert806 (
    .A(_3894_),
    .Y(_3894__bF$buf2)
);

BUFX2 BUFX2_insert805 (
    .A(_3894_),
    .Y(_3894__bF$buf3)
);

BUFX2 BUFX2_insert804 (
    .A(_3894_),
    .Y(_3894__bF$buf4)
);

BUFX2 BUFX2_insert803 (
    .A(_3915_),
    .Y(_3915__bF$buf0)
);

BUFX2 BUFX2_insert802 (
    .A(_3915_),
    .Y(_3915__bF$buf1)
);

BUFX2 BUFX2_insert801 (
    .A(_3915_),
    .Y(_3915__bF$buf2)
);

BUFX2 BUFX2_insert800 (
    .A(_3915_),
    .Y(_3915__bF$buf3)
);

BUFX2 BUFX2_insert799 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf0 )
);

BUFX2 BUFX2_insert798 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf1 )
);

BUFX2 BUFX2_insert797 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf2 )
);

BUFX2 BUFX2_insert796 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf3 )
);

BUFX2 BUFX2_insert795 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf4 )
);

BUFX2 BUFX2_insert794 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf5 )
);

BUFX2 BUFX2_insert793 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf6 )
);

BUFX2 BUFX2_insert792 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf7 )
);

BUFX2 BUFX2_insert791 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf0 )
);

BUFX2 BUFX2_insert790 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf1 )
);

BUFX2 BUFX2_insert789 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf2 )
);

BUFX2 BUFX2_insert788 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf3 )
);

BUFX2 BUFX2_insert787 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf4 )
);

BUFX2 BUFX2_insert786 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf0 )
);

BUFX2 BUFX2_insert785 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf1 )
);

BUFX2 BUFX2_insert784 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf2 )
);

BUFX2 BUFX2_insert783 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf3 )
);

BUFX2 BUFX2_insert782 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf4 )
);

BUFX2 BUFX2_insert781 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf5 )
);

BUFX2 BUFX2_insert780 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf6 )
);

BUFX2 BUFX2_insert779 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf7 )
);

BUFX2 BUFX2_insert778 (
    .A(_3019_),
    .Y(_3019__bF$buf0)
);

BUFX2 BUFX2_insert777 (
    .A(_3019_),
    .Y(_3019__bF$buf1)
);

BUFX2 BUFX2_insert776 (
    .A(_3019_),
    .Y(_3019__bF$buf2)
);

BUFX2 BUFX2_insert775 (
    .A(_3019_),
    .Y(_3019__bF$buf3)
);

BUFX2 BUFX2_insert774 (
    .A(_3019_),
    .Y(_3019__bF$buf4)
);

BUFX2 BUFX2_insert773 (
    .A(_3956_),
    .Y(_3956__bF$buf0)
);

BUFX2 BUFX2_insert772 (
    .A(_3956_),
    .Y(_3956__bF$buf1)
);

BUFX2 BUFX2_insert771 (
    .A(_3956_),
    .Y(_3956__bF$buf2)
);

BUFX2 BUFX2_insert770 (
    .A(_3956_),
    .Y(_3956__bF$buf3)
);

BUFX2 BUFX2_insert769 (
    .A(_3956_),
    .Y(_3956__bF$buf4)
);

BUFX2 BUFX2_insert768 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf0 )
);

BUFX2 BUFX2_insert767 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf1 )
);

BUFX2 BUFX2_insert766 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf2 )
);

BUFX2 BUFX2_insert765 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf3 )
);

BUFX2 BUFX2_insert764 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf4 )
);

BUFX2 BUFX2_insert763 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf5 )
);

BUFX2 BUFX2_insert762 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf6 )
);

BUFX2 BUFX2_insert761 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf7 )
);

BUFX2 BUFX2_insert760 (
    .A(_3022_),
    .Y(_3022__bF$buf0)
);

BUFX2 BUFX2_insert759 (
    .A(_3022_),
    .Y(_3022__bF$buf1)
);

BUFX2 BUFX2_insert758 (
    .A(_3022_),
    .Y(_3022__bF$buf2)
);

BUFX2 BUFX2_insert757 (
    .A(_3022_),
    .Y(_3022__bF$buf3)
);

BUFX2 BUFX2_insert756 (
    .A(_3022_),
    .Y(_3022__bF$buf4)
);

BUFX2 BUFX2_insert755 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf0 )
);

BUFX2 BUFX2_insert754 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf1 )
);

BUFX2 BUFX2_insert753 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf2 )
);

BUFX2 BUFX2_insert752 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf3 )
);

BUFX2 BUFX2_insert751 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf4 )
);

BUFX2 BUFX2_insert750 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf0 )
);

BUFX2 BUFX2_insert749 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf1 )
);

BUFX2 BUFX2_insert748 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf2 )
);

BUFX2 BUFX2_insert747 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf3 )
);

BUFX2 BUFX2_insert746 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf4 )
);

BUFX2 BUFX2_insert745 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf5 )
);

BUFX2 BUFX2_insert744 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf6 )
);

BUFX2 BUFX2_insert743 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf7 )
);

BUFX2 BUFX2_insert742 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf0 )
);

BUFX2 BUFX2_insert741 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf1 )
);

BUFX2 BUFX2_insert740 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf2 )
);

BUFX2 BUFX2_insert739 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf3 )
);

BUFX2 BUFX2_insert738 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf4 )
);

BUFX2 BUFX2_insert737 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf5 )
);

BUFX2 BUFX2_insert736 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf6 )
);

BUFX2 BUFX2_insert735 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf7 )
);

BUFX2 BUFX2_insert734 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf0)
);

BUFX2 BUFX2_insert733 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf1)
);

BUFX2 BUFX2_insert732 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf2)
);

BUFX2 BUFX2_insert731 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf3)
);

BUFX2 BUFX2_insert730 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf4)
);

BUFX2 BUFX2_insert729 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf5)
);

BUFX2 BUFX2_insert728 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf6)
);

BUFX2 BUFX2_insert727 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf7)
);

BUFX2 BUFX2_insert726 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf0 )
);

BUFX2 BUFX2_insert725 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf1 )
);

BUFX2 BUFX2_insert724 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf2 )
);

BUFX2 BUFX2_insert723 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf3 )
);

BUFX2 BUFX2_insert722 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf4 )
);

BUFX2 BUFX2_insert721 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf5 )
);

BUFX2 BUFX2_insert720 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf6 )
);

BUFX2 BUFX2_insert719 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf7 )
);

BUFX2 BUFX2_insert718 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf0 )
);

BUFX2 BUFX2_insert717 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf1 )
);

BUFX2 BUFX2_insert716 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf2 )
);

BUFX2 BUFX2_insert715 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf3 )
);

BUFX2 BUFX2_insert714 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf4 )
);

BUFX2 BUFX2_insert713 (
    .A(_3962_),
    .Y(_3962__bF$buf0)
);

BUFX2 BUFX2_insert712 (
    .A(_3962_),
    .Y(_3962__bF$buf1)
);

BUFX2 BUFX2_insert711 (
    .A(_3962_),
    .Y(_3962__bF$buf2)
);

BUFX2 BUFX2_insert710 (
    .A(_3962_),
    .Y(_3962__bF$buf3)
);

BUFX2 BUFX2_insert709 (
    .A(_3924_),
    .Y(_3924__bF$buf0)
);

BUFX2 BUFX2_insert708 (
    .A(_3924_),
    .Y(_3924__bF$buf1)
);

BUFX2 BUFX2_insert707 (
    .A(_3924_),
    .Y(_3924__bF$buf2)
);

BUFX2 BUFX2_insert706 (
    .A(_3924_),
    .Y(_3924__bF$buf3)
);

BUFX2 BUFX2_insert705 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf0 )
);

BUFX2 BUFX2_insert704 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf1 )
);

BUFX2 BUFX2_insert703 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf2 )
);

BUFX2 BUFX2_insert702 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf3 )
);

BUFX2 BUFX2_insert701 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf4 )
);

BUFX2 BUFX2_insert700 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf5 )
);

BUFX2 BUFX2_insert699 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf6 )
);

BUFX2 BUFX2_insert698 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf7 )
);

BUFX2 BUFX2_insert697 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf0 )
);

BUFX2 BUFX2_insert696 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf1 )
);

BUFX2 BUFX2_insert695 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf2 )
);

BUFX2 BUFX2_insert694 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf3 )
);

BUFX2 BUFX2_insert693 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf4 )
);

BUFX2 BUFX2_insert692 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf0 )
);

BUFX2 BUFX2_insert691 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf1 )
);

BUFX2 BUFX2_insert690 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf2 )
);

BUFX2 BUFX2_insert689 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf3 )
);

BUFX2 BUFX2_insert688 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf4 )
);

BUFX2 BUFX2_insert687 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf0 )
);

BUFX2 BUFX2_insert686 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf1 )
);

BUFX2 BUFX2_insert685 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf2 )
);

BUFX2 BUFX2_insert684 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf3 )
);

BUFX2 BUFX2_insert683 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf4 )
);

BUFX2 BUFX2_insert682 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf5 )
);

BUFX2 BUFX2_insert681 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf6 )
);

BUFX2 BUFX2_insert680 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf7 )
);

BUFX2 BUFX2_insert679 (
    .A(_5482_),
    .Y(_5482__bF$buf0)
);

BUFX2 BUFX2_insert678 (
    .A(_5482_),
    .Y(_5482__bF$buf1)
);

BUFX2 BUFX2_insert677 (
    .A(_5482_),
    .Y(_5482__bF$buf2)
);

BUFX2 BUFX2_insert676 (
    .A(_5482_),
    .Y(_5482__bF$buf3)
);

BUFX2 BUFX2_insert675 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf0 )
);

BUFX2 BUFX2_insert674 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf1 )
);

BUFX2 BUFX2_insert673 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf2 )
);

BUFX2 BUFX2_insert672 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf3 )
);

BUFX2 BUFX2_insert671 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf4 )
);

BUFX2 BUFX2_insert670 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf0 )
);

BUFX2 BUFX2_insert669 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf1 )
);

BUFX2 BUFX2_insert668 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf2 )
);

BUFX2 BUFX2_insert667 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf3 )
);

BUFX2 BUFX2_insert666 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf4 )
);

BUFX2 BUFX2_insert665 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf0 )
);

BUFX2 BUFX2_insert664 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf1 )
);

BUFX2 BUFX2_insert663 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf2 )
);

BUFX2 BUFX2_insert662 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf3 )
);

BUFX2 BUFX2_insert661 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf4 )
);

BUFX2 BUFX2_insert660 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf5 )
);

BUFX2 BUFX2_insert659 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf6 )
);

BUFX2 BUFX2_insert658 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf7 )
);

BUFX2 BUFX2_insert657 (
    .A(_5485_),
    .Y(_5485__bF$buf0)
);

BUFX2 BUFX2_insert656 (
    .A(_5485_),
    .Y(_5485__bF$buf1)
);

BUFX2 BUFX2_insert655 (
    .A(_5485_),
    .Y(_5485__bF$buf2)
);

BUFX2 BUFX2_insert654 (
    .A(_5485_),
    .Y(_5485__bF$buf3)
);

BUFX2 BUFX2_insert653 (
    .A(_5485_),
    .Y(_5485__bF$buf4)
);

BUFX2 BUFX2_insert652 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf0 )
);

BUFX2 BUFX2_insert651 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf1 )
);

BUFX2 BUFX2_insert650 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf2 )
);

BUFX2 BUFX2_insert649 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf3 )
);

BUFX2 BUFX2_insert648 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf4 )
);

BUFX2 BUFX2_insert647 (
    .A(_5506_),
    .Y(_5506__bF$buf0)
);

BUFX2 BUFX2_insert646 (
    .A(_5506_),
    .Y(_5506__bF$buf1)
);

BUFX2 BUFX2_insert645 (
    .A(_5506_),
    .Y(_5506__bF$buf2)
);

BUFX2 BUFX2_insert644 (
    .A(_5506_),
    .Y(_5506__bF$buf3)
);

BUFX2 BUFX2_insert643 (
    .A(_5506_),
    .Y(_5506__bF$buf4)
);

BUFX2 BUFX2_insert642 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf0 )
);

BUFX2 BUFX2_insert641 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf1 )
);

BUFX2 BUFX2_insert640 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf2 )
);

BUFX2 BUFX2_insert639 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf3 )
);

BUFX2 BUFX2_insert638 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf4 )
);

BUFX2 BUFX2_insert637 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf0)
);

BUFX2 BUFX2_insert636 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf1)
);

BUFX2 BUFX2_insert635 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf2)
);

BUFX2 BUFX2_insert634 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf3)
);

BUFX2 BUFX2_insert633 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf4)
);

BUFX2 BUFX2_insert632 (
    .A(_5488_),
    .Y(_5488__bF$buf0)
);

BUFX2 BUFX2_insert631 (
    .A(_5488_),
    .Y(_5488__bF$buf1)
);

BUFX2 BUFX2_insert630 (
    .A(_5488_),
    .Y(_5488__bF$buf2)
);

BUFX2 BUFX2_insert629 (
    .A(_5488_),
    .Y(_5488__bF$buf3)
);

BUFX2 BUFX2_insert628 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf0 )
);

BUFX2 BUFX2_insert627 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf1 )
);

BUFX2 BUFX2_insert626 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf2 )
);

BUFX2 BUFX2_insert625 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf3 )
);

BUFX2 BUFX2_insert624 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf4 )
);

BUFX2 BUFX2_insert623 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf0 )
);

BUFX2 BUFX2_insert622 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf1 )
);

BUFX2 BUFX2_insert621 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf2 )
);

BUFX2 BUFX2_insert620 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf3 )
);

BUFX2 BUFX2_insert619 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf4 )
);

BUFX2 BUFX2_insert618 (
    .A(_3939_),
    .Y(_3939__bF$buf0)
);

BUFX2 BUFX2_insert617 (
    .A(_3939_),
    .Y(_3939__bF$buf1)
);

BUFX2 BUFX2_insert616 (
    .A(_3939_),
    .Y(_3939__bF$buf2)
);

BUFX2 BUFX2_insert615 (
    .A(_3939_),
    .Y(_3939__bF$buf3)
);

BUFX2 BUFX2_insert614 (
    .A(_3939_),
    .Y(_3939__bF$buf4)
);

BUFX2 BUFX2_insert613 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf0 )
);

BUFX2 BUFX2_insert612 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf1 )
);

BUFX2 BUFX2_insert611 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf2 )
);

BUFX2 BUFX2_insert610 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf3 )
);

BUFX2 BUFX2_insert609 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf4 )
);

BUFX2 BUFX2_insert608 (
    .A(_4060_),
    .Y(_4060__bF$buf0)
);

BUFX2 BUFX2_insert607 (
    .A(_4060_),
    .Y(_4060__bF$buf1)
);

BUFX2 BUFX2_insert606 (
    .A(_4060_),
    .Y(_4060__bF$buf2)
);

BUFX2 BUFX2_insert605 (
    .A(_4060_),
    .Y(_4060__bF$buf3)
);

BUFX2 BUFX2_insert604 (
    .A(_3904_),
    .Y(_3904__bF$buf0)
);

BUFX2 BUFX2_insert603 (
    .A(_3904_),
    .Y(_3904__bF$buf1)
);

BUFX2 BUFX2_insert602 (
    .A(_3904_),
    .Y(_3904__bF$buf2)
);

BUFX2 BUFX2_insert601 (
    .A(_3904_),
    .Y(_3904__bF$buf3)
);

BUFX2 BUFX2_insert600 (
    .A(_3904_),
    .Y(_3904__bF$buf4)
);

BUFX2 BUFX2_insert599 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf0)
);

BUFX2 BUFX2_insert598 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf1)
);

BUFX2 BUFX2_insert597 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf2)
);

BUFX2 BUFX2_insert596 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf3)
);

BUFX2 BUFX2_insert595 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf4)
);

BUFX2 BUFX2_insert594 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf5)
);

BUFX2 BUFX2_insert593 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf0)
);

BUFX2 BUFX2_insert592 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf1)
);

BUFX2 BUFX2_insert591 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf2)
);

BUFX2 BUFX2_insert590 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf3)
);

BUFX2 BUFX2_insert589 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf4)
);

BUFX2 BUFX2_insert588 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf5)
);

BUFX2 BUFX2_insert587 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf6)
);

BUFX2 BUFX2_insert586 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf7)
);

BUFX2 BUFX2_insert585 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf8)
);

BUFX2 BUFX2_insert584 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf9)
);

BUFX2 BUFX2_insert583 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf10)
);

BUFX2 BUFX2_insert582 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf11)
);

BUFX2 BUFX2_insert581 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf12)
);

BUFX2 BUFX2_insert580 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf13)
);

BUFX2 BUFX2_insert579 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf14)
);

BUFX2 BUFX2_insert578 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf15)
);

BUFX2 BUFX2_insert577 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf16)
);

BUFX2 BUFX2_insert576 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf17)
);

BUFX2 BUFX2_insert575 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf18)
);

BUFX2 BUFX2_insert574 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf19)
);

BUFX2 BUFX2_insert573 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf20)
);

BUFX2 BUFX2_insert572 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf21)
);

BUFX2 BUFX2_insert571 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf22)
);

BUFX2 BUFX2_insert570 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf23)
);

BUFX2 BUFX2_insert569 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf24)
);

BUFX2 BUFX2_insert568 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf25)
);

BUFX2 BUFX2_insert567 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf26)
);

BUFX2 BUFX2_insert566 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf27)
);

BUFX2 BUFX2_insert565 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf28)
);

BUFX2 BUFX2_insert564 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf29)
);

BUFX2 BUFX2_insert563 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf30)
);

BUFX2 BUFX2_insert562 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf31)
);

BUFX2 BUFX2_insert561 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf32)
);

BUFX2 BUFX2_insert560 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf33)
);

BUFX2 BUFX2_insert559 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf34)
);

BUFX2 BUFX2_insert558 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf35)
);

BUFX2 BUFX2_insert557 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf36)
);

BUFX2 BUFX2_insert556 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf37)
);

BUFX2 BUFX2_insert555 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf38)
);

BUFX2 BUFX2_insert554 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf39)
);

BUFX2 BUFX2_insert553 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf40)
);

BUFX2 BUFX2_insert552 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf41)
);

BUFX2 BUFX2_insert551 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf42)
);

BUFX2 BUFX2_insert550 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf43)
);

BUFX2 BUFX2_insert549 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf44)
);

BUFX2 BUFX2_insert548 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf45)
);

BUFX2 BUFX2_insert547 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf46)
);

BUFX2 BUFX2_insert546 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf47)
);

BUFX2 BUFX2_insert545 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf48)
);

BUFX2 BUFX2_insert544 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf49)
);

BUFX2 BUFX2_insert543 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf50)
);

BUFX2 BUFX2_insert542 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf51)
);

BUFX2 BUFX2_insert541 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf52)
);

BUFX2 BUFX2_insert540 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf53)
);

BUFX2 BUFX2_insert539 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf54)
);

BUFX2 BUFX2_insert538 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf55)
);

BUFX2 BUFX2_insert537 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf56)
);

BUFX2 BUFX2_insert536 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf57)
);

BUFX2 BUFX2_insert535 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf58)
);

BUFX2 BUFX2_insert534 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf59)
);

BUFX2 BUFX2_insert533 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf60)
);

BUFX2 BUFX2_insert532 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf61)
);

BUFX2 BUFX2_insert531 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf62)
);

BUFX2 BUFX2_insert530 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf63)
);

BUFX2 BUFX2_insert529 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf64)
);

BUFX2 BUFX2_insert528 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf65)
);

BUFX2 BUFX2_insert527 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf66)
);

BUFX2 BUFX2_insert526 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf67)
);

BUFX2 BUFX2_insert525 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf68)
);

BUFX2 BUFX2_insert524 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf69)
);

BUFX2 BUFX2_insert523 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf70)
);

BUFX2 BUFX2_insert522 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf71)
);

BUFX2 BUFX2_insert521 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf72)
);

BUFX2 BUFX2_insert520 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf73)
);

BUFX2 BUFX2_insert519 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf74)
);

BUFX2 BUFX2_insert518 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf75)
);

BUFX2 BUFX2_insert517 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf76)
);

BUFX2 BUFX2_insert516 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf77)
);

BUFX2 BUFX2_insert515 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf78)
);

BUFX2 BUFX2_insert514 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf79)
);

BUFX2 BUFX2_insert513 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf80)
);

BUFX2 BUFX2_insert512 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf81)
);

BUFX2 BUFX2_insert511 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf82)
);

BUFX2 BUFX2_insert510 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf83)
);

BUFX2 BUFX2_insert509 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf84)
);

BUFX2 BUFX2_insert508 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf85)
);

BUFX2 BUFX2_insert507 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf86)
);

BUFX2 BUFX2_insert506 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf87)
);

BUFX2 BUFX2_insert505 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf88)
);

BUFX2 BUFX2_insert504 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf89)
);

BUFX2 BUFX2_insert503 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf90)
);

BUFX2 BUFX2_insert502 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf91)
);

BUFX2 BUFX2_insert501 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf92)
);

BUFX2 BUFX2_insert500 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf93)
);

BUFX2 BUFX2_insert499 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf94)
);

BUFX2 BUFX2_insert498 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf95)
);

BUFX2 BUFX2_insert497 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf96)
);

BUFX2 BUFX2_insert496 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf97)
);

BUFX2 BUFX2_insert495 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf98)
);

BUFX2 BUFX2_insert494 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf99)
);

BUFX2 BUFX2_insert493 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf100)
);

BUFX2 BUFX2_insert492 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf101)
);

BUFX2 BUFX2_insert491 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf102)
);

BUFX2 BUFX2_insert490 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf103)
);

BUFX2 BUFX2_insert489 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf104)
);

BUFX2 BUFX2_insert488 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf105)
);

BUFX2 BUFX2_insert487 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf106)
);

BUFX2 BUFX2_insert486 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf107)
);

BUFX2 BUFX2_insert485 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf108)
);

BUFX2 BUFX2_insert484 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf109)
);

BUFX2 BUFX2_insert483 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf110)
);

BUFX2 BUFX2_insert482 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf111)
);

BUFX2 BUFX2_insert481 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf112)
);

BUFX2 BUFX2_insert480 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf113)
);

BUFX2 BUFX2_insert479 (
    .A(_5421_),
    .Y(_5421__bF$buf0)
);

BUFX2 BUFX2_insert478 (
    .A(_5421_),
    .Y(_5421__bF$buf1)
);

BUFX2 BUFX2_insert477 (
    .A(_5421_),
    .Y(_5421__bF$buf2)
);

BUFX2 BUFX2_insert476 (
    .A(_5421_),
    .Y(_5421__bF$buf3)
);

BUFX2 BUFX2_insert475 (
    .A(_3886_),
    .Y(_3886__bF$buf0)
);

BUFX2 BUFX2_insert474 (
    .A(_3886_),
    .Y(_3886__bF$buf1)
);

BUFX2 BUFX2_insert473 (
    .A(_3886_),
    .Y(_3886__bF$buf2)
);

BUFX2 BUFX2_insert472 (
    .A(_3886_),
    .Y(_3886__bF$buf3)
);

BUFX2 BUFX2_insert471 (
    .A(_3181_),
    .Y(_3181__bF$buf0)
);

BUFX2 BUFX2_insert470 (
    .A(_3181_),
    .Y(_3181__bF$buf1)
);

BUFX2 BUFX2_insert469 (
    .A(_3181_),
    .Y(_3181__bF$buf2)
);

BUFX2 BUFX2_insert468 (
    .A(_3181_),
    .Y(_3181__bF$buf3)
);

BUFX2 BUFX2_insert467 (
    .A(_3181_),
    .Y(_3181__bF$buf4)
);

BUFX2 BUFX2_insert466 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf0 )
);

BUFX2 BUFX2_insert465 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf1 )
);

BUFX2 BUFX2_insert464 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf2 )
);

BUFX2 BUFX2_insert463 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf3 )
);

BUFX2 BUFX2_insert462 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf4 )
);

BUFX2 BUFX2_insert461 (
    .A(_5518_),
    .Y(_5518__bF$buf0)
);

BUFX2 BUFX2_insert460 (
    .A(_5518_),
    .Y(_5518__bF$buf1)
);

BUFX2 BUFX2_insert459 (
    .A(_5518_),
    .Y(_5518__bF$buf2)
);

BUFX2 BUFX2_insert458 (
    .A(_5518_),
    .Y(_5518__bF$buf3)
);

BUFX2 BUFX2_insert457 (
    .A(_5518_),
    .Y(_5518__bF$buf4)
);

BUFX2 BUFX2_insert456 (
    .A(_5462_),
    .Y(_5462__bF$buf0)
);

BUFX2 BUFX2_insert455 (
    .A(_5462_),
    .Y(_5462__bF$buf1)
);

BUFX2 BUFX2_insert454 (
    .A(_5462_),
    .Y(_5462__bF$buf2)
);

BUFX2 BUFX2_insert453 (
    .A(_5462_),
    .Y(_5462__bF$buf3)
);

BUFX2 BUFX2_insert452 (
    .A(_5462_),
    .Y(_5462__bF$buf4)
);

BUFX2 BUFX2_insert451 (
    .A(_3910_),
    .Y(_3910__bF$buf0)
);

BUFX2 BUFX2_insert450 (
    .A(_3910_),
    .Y(_3910__bF$buf1)
);

BUFX2 BUFX2_insert449 (
    .A(_3910_),
    .Y(_3910__bF$buf2)
);

BUFX2 BUFX2_insert448 (
    .A(_3910_),
    .Y(_3910__bF$buf3)
);

BUFX2 BUFX2_insert447 (
    .A(_3889_),
    .Y(_3889__bF$buf0)
);

BUFX2 BUFX2_insert446 (
    .A(_3889_),
    .Y(_3889__bF$buf1)
);

BUFX2 BUFX2_insert445 (
    .A(_3889_),
    .Y(_3889__bF$buf2)
);

BUFX2 BUFX2_insert444 (
    .A(_3889_),
    .Y(_3889__bF$buf3)
);

BUFX2 BUFX2_insert443 (
    .A(_3889_),
    .Y(_3889__bF$buf4)
);

BUFX2 BUFX2_insert442 (
    .A(_5521_),
    .Y(_5521__bF$buf0)
);

BUFX2 BUFX2_insert441 (
    .A(_5521_),
    .Y(_5521__bF$buf1)
);

BUFX2 BUFX2_insert440 (
    .A(_5521_),
    .Y(_5521__bF$buf2)
);

BUFX2 BUFX2_insert439 (
    .A(_5521_),
    .Y(_5521__bF$buf3)
);

BUFX2 BUFX2_insert438 (
    .A(_5521_),
    .Y(_5521__bF$buf4)
);

BUFX2 BUFX2_insert437 (
    .A(_5465_),
    .Y(_5465__bF$buf0)
);

BUFX2 BUFX2_insert436 (
    .A(_5465_),
    .Y(_5465__bF$buf1)
);

BUFX2 BUFX2_insert435 (
    .A(_5465_),
    .Y(_5465__bF$buf2)
);

BUFX2 BUFX2_insert434 (
    .A(_5465_),
    .Y(_5465__bF$buf3)
);

BUFX2 BUFX2_insert433 (
    .A(_5465_),
    .Y(_5465__bF$buf4)
);

BUFX2 BUFX2_insert432 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf0 )
);

BUFX2 BUFX2_insert431 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf1 )
);

BUFX2 BUFX2_insert430 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf2 )
);

BUFX2 BUFX2_insert429 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf3 )
);

BUFX2 BUFX2_insert428 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf4 )
);

BUFX2 BUFX2_insert427 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf5 )
);

BUFX2 BUFX2_insert426 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf6 )
);

BUFX2 BUFX2_insert425 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf7 )
);

BUFX2 BUFX2_insert424 (
    .A(_3017_),
    .Y(_3017__bF$buf0)
);

BUFX2 BUFX2_insert423 (
    .A(_3017_),
    .Y(_3017__bF$buf1)
);

BUFX2 BUFX2_insert422 (
    .A(_3017_),
    .Y(_3017__bF$buf2)
);

BUFX2 BUFX2_insert421 (
    .A(_3017_),
    .Y(_3017__bF$buf3)
);

BUFX2 BUFX2_insert420 (
    .A(_3017_),
    .Y(_3017__bF$buf4)
);

BUFX2 BUFX2_insert419 (
    .A(_3916_),
    .Y(_3916__bF$buf0)
);

BUFX2 BUFX2_insert418 (
    .A(_3916_),
    .Y(_3916__bF$buf1)
);

BUFX2 BUFX2_insert417 (
    .A(_3916_),
    .Y(_3916__bF$buf2)
);

BUFX2 BUFX2_insert416 (
    .A(_3916_),
    .Y(_3916__bF$buf3)
);

BUFX2 BUFX2_insert415 (
    .A(_3916_),
    .Y(_3916__bF$buf4)
);

BUFX2 BUFX2_insert414 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf0 )
);

BUFX2 BUFX2_insert413 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf1 )
);

BUFX2 BUFX2_insert412 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf2 )
);

BUFX2 BUFX2_insert411 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf3 )
);

BUFX2 BUFX2_insert410 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf4 )
);

BUFX2 BUFX2_insert409 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf5 )
);

BUFX2 BUFX2_insert408 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf6 )
);

BUFX2 BUFX2_insert407 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf7 )
);

BUFX2 BUFX2_insert406 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf0 )
);

BUFX2 BUFX2_insert405 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf1 )
);

BUFX2 BUFX2_insert404 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf2 )
);

BUFX2 BUFX2_insert403 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf3 )
);

BUFX2 BUFX2_insert402 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf4 )
);

BUFX2 BUFX2_insert401 (
    .A(_5565_),
    .Y(_5565__bF$buf0)
);

BUFX2 BUFX2_insert400 (
    .A(_5565_),
    .Y(_5565__bF$buf1)
);

BUFX2 BUFX2_insert399 (
    .A(_5565_),
    .Y(_5565__bF$buf2)
);

BUFX2 BUFX2_insert398 (
    .A(_5565_),
    .Y(_5565__bF$buf3)
);

BUFX2 BUFX2_insert397 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf0 )
);

BUFX2 BUFX2_insert396 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf1 )
);

BUFX2 BUFX2_insert395 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf2 )
);

BUFX2 BUFX2_insert394 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf3 )
);

BUFX2 BUFX2_insert393 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf4 )
);

BUFX2 BUFX2_insert392 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf5 )
);

BUFX2 BUFX2_insert391 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf6 )
);

BUFX2 BUFX2_insert390 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf7 )
);

BUFX2 BUFX2_insert389 (
    .A(_5471_),
    .Y(_5471__bF$buf0)
);

BUFX2 BUFX2_insert388 (
    .A(_5471_),
    .Y(_5471__bF$buf1)
);

BUFX2 BUFX2_insert387 (
    .A(_5471_),
    .Y(_5471__bF$buf2)
);

BUFX2 BUFX2_insert386 (
    .A(_5471_),
    .Y(_5471__bF$buf3)
);

BUFX2 BUFX2_insert385 (
    .A(_5471_),
    .Y(_5471__bF$buf4)
);

BUFX2 BUFX2_insert384 (
    .A(_2367_),
    .Y(_2367__bF$buf0)
);

BUFX2 BUFX2_insert383 (
    .A(_2367_),
    .Y(_2367__bF$buf1)
);

BUFX2 BUFX2_insert382 (
    .A(_2367_),
    .Y(_2367__bF$buf2)
);

BUFX2 BUFX2_insert381 (
    .A(_2367_),
    .Y(_2367__bF$buf3)
);

BUFX2 BUFX2_insert380 (
    .A(_5433_),
    .Y(_5433__bF$buf0)
);

BUFX2 BUFX2_insert379 (
    .A(_5433_),
    .Y(_5433__bF$buf1)
);

BUFX2 BUFX2_insert378 (
    .A(_5433_),
    .Y(_5433__bF$buf2)
);

BUFX2 BUFX2_insert377 (
    .A(_5433_),
    .Y(_5433__bF$buf3)
);

BUFX2 BUFX2_insert376 (
    .A(_5433_),
    .Y(_5433__bF$buf4)
);

BUFX2 BUFX2_insert375 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf0)
);

BUFX2 BUFX2_insert374 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf1)
);

BUFX2 BUFX2_insert373 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf2)
);

BUFX2 BUFX2_insert372 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf3)
);

BUFX2 BUFX2_insert371 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf4)
);

BUFX2 BUFX2_insert370 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf5)
);

BUFX2 BUFX2_insert369 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf6)
);

BUFX2 BUFX2_insert368 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf7)
);

BUFX2 BUFX2_insert367 (
    .A(_3957_),
    .Y(_3957__bF$buf0)
);

BUFX2 BUFX2_insert366 (
    .A(_3957_),
    .Y(_3957__bF$buf1)
);

BUFX2 BUFX2_insert365 (
    .A(_3957_),
    .Y(_3957__bF$buf2)
);

BUFX2 BUFX2_insert364 (
    .A(_3957_),
    .Y(_3957__bF$buf3)
);

BUFX2 BUFX2_insert363 (
    .A(_3957_),
    .Y(_3957__bF$buf4)
);

BUFX2 BUFX2_insert362 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf0 )
);

BUFX2 BUFX2_insert361 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf1 )
);

BUFX2 BUFX2_insert360 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf2 )
);

BUFX2 BUFX2_insert359 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf3 )
);

BUFX2 BUFX2_insert358 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf4 )
);

BUFX2 BUFX2_insert357 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf5 )
);

BUFX2 BUFX2_insert356 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf6 )
);

BUFX2 BUFX2_insert355 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf7 )
);

BUFX2 BUFX2_insert354 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf0 )
);

BUFX2 BUFX2_insert353 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf1 )
);

BUFX2 BUFX2_insert352 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf2 )
);

BUFX2 BUFX2_insert351 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf3 )
);

BUFX2 BUFX2_insert350 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf4 )
);

BUFX2 BUFX2_insert349 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf0 )
);

BUFX2 BUFX2_insert348 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf1 )
);

BUFX2 BUFX2_insert347 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf2 )
);

BUFX2 BUFX2_insert346 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf3 )
);

BUFX2 BUFX2_insert345 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf4 )
);

BUFX2 BUFX2_insert344 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf5 )
);

BUFX2 BUFX2_insert343 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf6 )
);

BUFX2 BUFX2_insert342 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf7 )
);

BUFX2 BUFX2_insert341 (
    .A(_5436_),
    .Y(_5436__bF$buf0)
);

BUFX2 BUFX2_insert340 (
    .A(_5436_),
    .Y(_5436__bF$buf1)
);

BUFX2 BUFX2_insert339 (
    .A(_5436_),
    .Y(_5436__bF$buf2)
);

BUFX2 BUFX2_insert338 (
    .A(_5436_),
    .Y(_5436__bF$buf3)
);

BUFX2 BUFX2_insert337 (
    .A(_5436_),
    .Y(_5436__bF$buf4)
);

BUFX2 BUFX2_insert336 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf0 )
);

BUFX2 BUFX2_insert335 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf1 )
);

BUFX2 BUFX2_insert334 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf2 )
);

BUFX2 BUFX2_insert333 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf3 )
);

BUFX2 BUFX2_insert332 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf4 )
);

BUFX2 BUFX2_insert331 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf5 )
);

BUFX2 BUFX2_insert330 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf6 )
);

BUFX2 BUFX2_insert329 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf7 )
);

BUFX2 BUFX2_insert328 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf0 )
);

BUFX2 BUFX2_insert327 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf1 )
);

BUFX2 BUFX2_insert326 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf2 )
);

BUFX2 BUFX2_insert325 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf3 )
);

BUFX2 BUFX2_insert324 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf4 )
);

BUFX2 BUFX2_insert323 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf5 )
);

BUFX2 BUFX2_insert322 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf6 )
);

BUFX2 BUFX2_insert321 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf7 )
);

BUFX2 BUFX2_insert320 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf0)
);

BUFX2 BUFX2_insert319 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf1)
);

BUFX2 BUFX2_insert318 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf2)
);

BUFX2 BUFX2_insert317 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf3)
);

BUFX2 BUFX2_insert316 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf4)
);

BUFX2 BUFX2_insert315 (
    .A(_3866_),
    .Y(_3866__bF$buf0)
);

BUFX2 BUFX2_insert314 (
    .A(_3866_),
    .Y(_3866__bF$buf1)
);

BUFX2 BUFX2_insert313 (
    .A(_3866_),
    .Y(_3866__bF$buf2)
);

BUFX2 BUFX2_insert312 (
    .A(_3866_),
    .Y(_3866__bF$buf3)
);

BUFX2 BUFX2_insert311 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf0 )
);

BUFX2 BUFX2_insert310 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf1 )
);

BUFX2 BUFX2_insert309 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf2 )
);

BUFX2 BUFX2_insert308 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf3 )
);

BUFX2 BUFX2_insert307 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf4 )
);

BUFX2 BUFX2_insert306 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf0 )
);

BUFX2 BUFX2_insert305 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf1 )
);

BUFX2 BUFX2_insert304 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf2 )
);

BUFX2 BUFX2_insert303 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf3 )
);

BUFX2 BUFX2_insert302 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf0 )
);

BUFX2 BUFX2_insert301 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf1 )
);

BUFX2 BUFX2_insert300 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf2 )
);

BUFX2 BUFX2_insert299 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf3 )
);

BUFX2 BUFX2_insert298 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf4 )
);

BUFX2 BUFX2_insert297 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf0 )
);

BUFX2 BUFX2_insert296 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf1 )
);

BUFX2 BUFX2_insert295 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf2 )
);

BUFX2 BUFX2_insert294 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf3 )
);

BUFX2 BUFX2_insert293 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf4 )
);

BUFX2 BUFX2_insert292 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf5 )
);

BUFX2 BUFX2_insert291 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf6 )
);

BUFX2 BUFX2_insert290 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf7 )
);

BUFX2 BUFX2_insert289 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf0 )
);

BUFX2 BUFX2_insert288 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf1 )
);

BUFX2 BUFX2_insert287 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf2 )
);

BUFX2 BUFX2_insert286 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf3 )
);

BUFX2 BUFX2_insert285 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf4 )
);

BUFX2 BUFX2_insert284 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf0 )
);

BUFX2 BUFX2_insert283 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf1 )
);

BUFX2 BUFX2_insert282 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf2 )
);

BUFX2 BUFX2_insert281 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf3 )
);

BUFX2 BUFX2_insert280 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf4 )
);

BUFX2 BUFX2_insert279 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf5 )
);

BUFX2 BUFX2_insert278 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf6 )
);

BUFX2 BUFX2_insert277 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf7 )
);

BUFX2 BUFX2_insert276 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf0 )
);

BUFX2 BUFX2_insert275 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf1 )
);

BUFX2 BUFX2_insert274 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf2 )
);

BUFX2 BUFX2_insert273 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf3 )
);

BUFX2 BUFX2_insert272 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf4 )
);

BUFX2 BUFX2_insert271 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf5 )
);

BUFX2 BUFX2_insert270 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf6 )
);

BUFX2 BUFX2_insert269 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf7 )
);

BUFX2 BUFX2_insert268 (
    .A(_3875_),
    .Y(_3875__bF$buf0)
);

BUFX2 BUFX2_insert267 (
    .A(_3875_),
    .Y(_3875__bF$buf1)
);

BUFX2 BUFX2_insert266 (
    .A(_3875_),
    .Y(_3875__bF$buf2)
);

BUFX2 BUFX2_insert265 (
    .A(_3875_),
    .Y(_3875__bF$buf3)
);

BUFX2 BUFX2_insert264 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf0 )
);

BUFX2 BUFX2_insert263 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf1 )
);

BUFX2 BUFX2_insert262 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf2 )
);

BUFX2 BUFX2_insert261 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf3 )
);

BUFX2 BUFX2_insert260 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf4 )
);

BUFX2 BUFX2_insert259 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf0)
);

BUFX2 BUFX2_insert258 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf1)
);

BUFX2 BUFX2_insert257 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf2)
);

BUFX2 BUFX2_insert256 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf3)
);

BUFX2 BUFX2_insert255 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf4)
);

BUFX2 BUFX2_insert254 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf5)
);

BUFX2 BUFX2_insert253 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf6)
);

BUFX2 BUFX2_insert252 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf7)
);

BUFX2 BUFX2_insert251 (
    .A(_3934_),
    .Y(_3934__bF$buf0)
);

BUFX2 BUFX2_insert250 (
    .A(_3934_),
    .Y(_3934__bF$buf1)
);

BUFX2 BUFX2_insert249 (
    .A(_3934_),
    .Y(_3934__bF$buf2)
);

BUFX2 BUFX2_insert248 (
    .A(_3934_),
    .Y(_3934__bF$buf3)
);

BUFX2 BUFX2_insert247 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf0 )
);

BUFX2 BUFX2_insert246 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf1 )
);

BUFX2 BUFX2_insert245 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf2 )
);

BUFX2 BUFX2_insert244 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf3 )
);

BUFX2 BUFX2_insert243 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf4 )
);

BUFX2 BUFX2_insert242 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf0 )
);

BUFX2 BUFX2_insert241 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf1 )
);

BUFX2 BUFX2_insert240 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf2 )
);

BUFX2 BUFX2_insert239 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf3 )
);

BUFX2 BUFX2_insert238 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf4 )
);

CLKBUF1 CLKBUF1_insert237 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert236 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert235 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert234 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert233 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert232 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert231 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert230 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert229 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert228 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert227 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert226 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert225 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert224 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert223 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert222 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert221 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert220 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert219 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert218 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert217 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert216 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert215 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert214 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert213 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert212 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert211 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert210 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert209 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert208 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert207 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert206 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert205 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert204 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert203 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert202 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert201 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert200 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert199 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert198 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert197 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert196 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert195 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert194 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert193 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert192 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert191 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert190 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert189 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert188 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert187 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert186 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert185 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert184 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert183 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert182 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf55)
);

CLKBUF1 CLKBUF1_insert181 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert180 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert179 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf58)
);

CLKBUF1 CLKBUF1_insert178 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf59)
);

CLKBUF1 CLKBUF1_insert177 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf60)
);

CLKBUF1 CLKBUF1_insert176 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf61)
);

CLKBUF1 CLKBUF1_insert175 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf62)
);

CLKBUF1 CLKBUF1_insert174 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf63)
);

CLKBUF1 CLKBUF1_insert173 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf64)
);

CLKBUF1 CLKBUF1_insert172 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf65)
);

CLKBUF1 CLKBUF1_insert171 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert170 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf67)
);

CLKBUF1 CLKBUF1_insert169 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf68)
);

CLKBUF1 CLKBUF1_insert168 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert167 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf70)
);

CLKBUF1 CLKBUF1_insert166 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf71)
);

CLKBUF1 CLKBUF1_insert165 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf72)
);

CLKBUF1 CLKBUF1_insert164 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf73)
);

CLKBUF1 CLKBUF1_insert163 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf74)
);

CLKBUF1 CLKBUF1_insert162 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf75)
);

CLKBUF1 CLKBUF1_insert161 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf76)
);

CLKBUF1 CLKBUF1_insert160 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf77)
);

CLKBUF1 CLKBUF1_insert159 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf78)
);

CLKBUF1 CLKBUF1_insert158 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf79)
);

CLKBUF1 CLKBUF1_insert157 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf80)
);

CLKBUF1 CLKBUF1_insert156 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf81)
);

CLKBUF1 CLKBUF1_insert155 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf82)
);

CLKBUF1 CLKBUF1_insert154 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf83)
);

CLKBUF1 CLKBUF1_insert153 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf84)
);

CLKBUF1 CLKBUF1_insert152 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf85)
);

CLKBUF1 CLKBUF1_insert151 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf86)
);

CLKBUF1 CLKBUF1_insert150 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf87)
);

CLKBUF1 CLKBUF1_insert149 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf88)
);

CLKBUF1 CLKBUF1_insert148 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf89)
);

CLKBUF1 CLKBUF1_insert147 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf90)
);

CLKBUF1 CLKBUF1_insert146 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf91)
);

CLKBUF1 CLKBUF1_insert145 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf92)
);

CLKBUF1 CLKBUF1_insert144 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf93)
);

CLKBUF1 CLKBUF1_insert143 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf94)
);

CLKBUF1 CLKBUF1_insert142 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf95)
);

CLKBUF1 CLKBUF1_insert141 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf96)
);

CLKBUF1 CLKBUF1_insert140 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf97)
);

CLKBUF1 CLKBUF1_insert139 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf98)
);

CLKBUF1 CLKBUF1_insert138 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf99)
);

CLKBUF1 CLKBUF1_insert137 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf100)
);

CLKBUF1 CLKBUF1_insert136 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf101)
);

CLKBUF1 CLKBUF1_insert135 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf102)
);

CLKBUF1 CLKBUF1_insert134 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf103)
);

CLKBUF1 CLKBUF1_insert133 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf104)
);

CLKBUF1 CLKBUF1_insert132 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf105)
);

CLKBUF1 CLKBUF1_insert131 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf106)
);

CLKBUF1 CLKBUF1_insert130 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf107)
);

CLKBUF1 CLKBUF1_insert129 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf108)
);

CLKBUF1 CLKBUF1_insert128 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf109)
);

CLKBUF1 CLKBUF1_insert127 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf110)
);

CLKBUF1 CLKBUF1_insert126 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf111)
);

CLKBUF1 CLKBUF1_insert125 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf112)
);

CLKBUF1 CLKBUF1_insert124 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf113)
);

BUFX2 BUFX2_insert123 (
    .A(IorD),
    .Y(IorD_bF$buf0)
);

BUFX2 BUFX2_insert122 (
    .A(IorD),
    .Y(IorD_bF$buf1)
);

BUFX2 BUFX2_insert121 (
    .A(IorD),
    .Y(IorD_bF$buf2)
);

BUFX2 BUFX2_insert120 (
    .A(IorD),
    .Y(IorD_bF$buf3)
);

BUFX2 BUFX2_insert119 (
    .A(IorD),
    .Y(IorD_bF$buf4)
);

BUFX2 BUFX2_insert118 (
    .A(IorD),
    .Y(IorD_bF$buf5)
);

BUFX2 BUFX2_insert117 (
    .A(IorD),
    .Y(IorD_bF$buf6)
);

BUFX2 BUFX2_insert116 (
    .A(IorD),
    .Y(IorD_bF$buf7)
);

BUFX2 BUFX2_insert115 (
    .A(_5492_),
    .Y(_5492__bF$buf0)
);

BUFX2 BUFX2_insert114 (
    .A(_5492_),
    .Y(_5492__bF$buf1)
);

BUFX2 BUFX2_insert113 (
    .A(_5492_),
    .Y(_5492__bF$buf2)
);

BUFX2 BUFX2_insert112 (
    .A(_5492_),
    .Y(_5492__bF$buf3)
);

BUFX2 BUFX2_insert111 (
    .A(_5492_),
    .Y(_5492__bF$buf4)
);

BUFX2 BUFX2_insert110 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf0 )
);

BUFX2 BUFX2_insert109 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf1 )
);

BUFX2 BUFX2_insert108 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf2 )
);

BUFX2 BUFX2_insert107 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf3 )
);

BUFX2 BUFX2_insert106 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf4 )
);

BUFX2 BUFX2_insert105 (
    .A(_3940_),
    .Y(_3940__bF$buf0)
);

BUFX2 BUFX2_insert104 (
    .A(_3940_),
    .Y(_3940__bF$buf1)
);

BUFX2 BUFX2_insert103 (
    .A(_3940_),
    .Y(_3940__bF$buf2)
);

BUFX2 BUFX2_insert102 (
    .A(_3940_),
    .Y(_3940__bF$buf3)
);

BUFX2 BUFX2_insert101 (
    .A(_3902_),
    .Y(_3902__bF$buf0)
);

BUFX2 BUFX2_insert100 (
    .A(_3902_),
    .Y(_3902__bF$buf1)
);

BUFX2 BUFX2_insert99 (
    .A(_3902_),
    .Y(_3902__bF$buf2)
);

BUFX2 BUFX2_insert98 (
    .A(_3902_),
    .Y(_3902__bF$buf3)
);

BUFX2 BUFX2_insert97 (
    .A(_3902_),
    .Y(_3902__bF$buf4)
);

BUFX2 BUFX2_insert96 (
    .A(_5513_),
    .Y(_5513__bF$buf0)
);

BUFX2 BUFX2_insert95 (
    .A(_5513_),
    .Y(_5513__bF$buf1)
);

BUFX2 BUFX2_insert94 (
    .A(_5513_),
    .Y(_5513__bF$buf2)
);

BUFX2 BUFX2_insert93 (
    .A(_5513_),
    .Y(_5513__bF$buf3)
);

BUFX2 BUFX2_insert92 (
    .A(_5513_),
    .Y(_5513__bF$buf4)
);

BUFX2 BUFX2_insert91 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf0 )
);

BUFX2 BUFX2_insert90 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf1 )
);

BUFX2 BUFX2_insert89 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf2 )
);

BUFX2 BUFX2_insert88 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf3 )
);

BUFX2 BUFX2_insert87 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf4 )
);

BUFX2 BUFX2_insert86 (
    .A(_5457_),
    .Y(_5457__bF$buf0)
);

BUFX2 BUFX2_insert85 (
    .A(_5457_),
    .Y(_5457__bF$buf1)
);

BUFX2 BUFX2_insert84 (
    .A(_5457_),
    .Y(_5457__bF$buf2)
);

BUFX2 BUFX2_insert83 (
    .A(_5457_),
    .Y(_5457__bF$buf3)
);

BUFX2 BUFX2_insert82 (
    .A(_5457_),
    .Y(_5457__bF$buf4)
);

BUFX2 BUFX2_insert81 (
    .A(_5460_),
    .Y(_5460__bF$buf0)
);

BUFX2 BUFX2_insert80 (
    .A(_5460_),
    .Y(_5460__bF$buf1)
);

BUFX2 BUFX2_insert79 (
    .A(_5460_),
    .Y(_5460__bF$buf2)
);

BUFX2 BUFX2_insert78 (
    .A(_5460_),
    .Y(_5460__bF$buf3)
);

BUFX2 BUFX2_insert77 (
    .A(_5460_),
    .Y(_5460__bF$buf4)
);

BUFX2 BUFX2_insert76 (
    .A(_5560_),
    .Y(_5560__bF$buf0)
);

BUFX2 BUFX2_insert75 (
    .A(_5560_),
    .Y(_5560__bF$buf1)
);

BUFX2 BUFX2_insert74 (
    .A(_5560_),
    .Y(_5560__bF$buf2)
);

BUFX2 BUFX2_insert73 (
    .A(_5560_),
    .Y(_5560__bF$buf3)
);

BUFX2 BUFX2_insert72 (
    .A(_3185_),
    .Y(_3185__bF$buf0)
);

BUFX2 BUFX2_insert71 (
    .A(_3185_),
    .Y(_3185__bF$buf1)
);

BUFX2 BUFX2_insert70 (
    .A(_3185_),
    .Y(_3185__bF$buf2)
);

BUFX2 BUFX2_insert69 (
    .A(_3185_),
    .Y(_3185__bF$buf3)
);

BUFX2 BUFX2_insert68 (
    .A(_3185_),
    .Y(_3185__bF$buf4)
);

BUFX2 BUFX2_insert67 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf0 )
);

BUFX2 BUFX2_insert66 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf1 )
);

BUFX2 BUFX2_insert65 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf2 )
);

BUFX2 BUFX2_insert64 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf3 )
);

BUFX2 BUFX2_insert63 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf4 )
);

BUFX2 BUFX2_insert62 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf5 )
);

BUFX2 BUFX2_insert61 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf6 )
);

BUFX2 BUFX2_insert60 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf7 )
);

BUFX2 BUFX2_insert59 (
    .A(_2362_),
    .Y(_2362__bF$buf0)
);

BUFX2 BUFX2_insert58 (
    .A(_2362_),
    .Y(_2362__bF$buf1)
);

BUFX2 BUFX2_insert57 (
    .A(_2362_),
    .Y(_2362__bF$buf2)
);

BUFX2 BUFX2_insert56 (
    .A(_2362_),
    .Y(_2362__bF$buf3)
);

BUFX2 BUFX2_insert55 (
    .A(_3952_),
    .Y(_3952__bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .A(_3952_),
    .Y(_3952__bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .A(_3952_),
    .Y(_3952__bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .A(_3952_),
    .Y(_3952__bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .A(_5466_),
    .Y(_5466__bF$buf0)
);

BUFX2 BUFX2_insert50 (
    .A(_5466_),
    .Y(_5466__bF$buf1)
);

BUFX2 BUFX2_insert49 (
    .A(_5466_),
    .Y(_5466__bF$buf2)
);

BUFX2 BUFX2_insert48 (
    .A(_5466_),
    .Y(_5466__bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .A(_5466_),
    .Y(_5466__bF$buf4)
);

BUFX2 BUFX2_insert46 (
    .A(_5428_),
    .Y(_5428__bF$buf0)
);

BUFX2 BUFX2_insert45 (
    .A(_5428_),
    .Y(_5428__bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .A(_5428_),
    .Y(_5428__bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .A(_5428_),
    .Y(_5428__bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf0 )
);

BUFX2 BUFX2_insert41 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf1 )
);

BUFX2 BUFX2_insert40 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf2 )
);

BUFX2 BUFX2_insert39 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf3 )
);

BUFX2 BUFX2_insert38 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf4 )
);

BUFX2 BUFX2_insert37 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf5 )
);

BUFX2 BUFX2_insert36 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf6 )
);

BUFX2 BUFX2_insert35 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf7 )
);

BUFX2 BUFX2_insert34 (
    .A(_5563_),
    .Y(_5563__bF$buf0)
);

BUFX2 BUFX2_insert33 (
    .A(_5563_),
    .Y(_5563__bF$buf1)
);

BUFX2 BUFX2_insert32 (
    .A(_5563_),
    .Y(_5563__bF$buf2)
);

BUFX2 BUFX2_insert31 (
    .A(_5563_),
    .Y(_5563__bF$buf3)
);

BUFX2 BUFX2_insert30 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf0 )
);

BUFX2 BUFX2_insert29 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf1 )
);

BUFX2 BUFX2_insert28 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf2 )
);

BUFX2 BUFX2_insert27 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf3 )
);

BUFX2 BUFX2_insert26 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf4 )
);

BUFX2 BUFX2_insert25 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf5 )
);

BUFX2 BUFX2_insert24 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf6 )
);

BUFX2 BUFX2_insert23 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf7 )
);

BUFX2 BUFX2_insert22 (
    .A(_2365_),
    .Y(_2365__bF$buf0)
);

BUFX2 BUFX2_insert21 (
    .A(_2365_),
    .Y(_2365__bF$buf1)
);

BUFX2 BUFX2_insert20 (
    .A(_2365_),
    .Y(_2365__bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .A(_2365_),
    .Y(_2365__bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .A(_2365_),
    .Y(_2365__bF$buf4)
);

BUFX2 BUFX2_insert17 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf0 )
);

BUFX2 BUFX2_insert16 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf1 )
);

BUFX2 BUFX2_insert15 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf2 )
);

BUFX2 BUFX2_insert14 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf3 )
);

BUFX2 BUFX2_insert13 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf4 )
);

BUFX2 BUFX2_insert12 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf5 )
);

BUFX2 BUFX2_insert11 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf6 )
);

BUFX2 BUFX2_insert10 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf7 )
);

BUFX2 BUFX2_insert9 (
    .A(_3021_),
    .Y(_3021__bF$buf0)
);

BUFX2 BUFX2_insert8 (
    .A(_3021_),
    .Y(_3021__bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .A(_3021_),
    .Y(_3021__bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .A(_3021_),
    .Y(_3021__bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .A(_3021_),
    .Y(_3021__bF$buf4)
);

BUFX2 BUFX2_insert4 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf0 )
);

BUFX2 BUFX2_insert3 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf1 )
);

BUFX2 BUFX2_insert2 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf2 )
);

BUFX2 BUFX2_insert1 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf3 )
);

BUFX2 BUFX2_insert0 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf4 )
);

INVX1 _10000_ (
    .A(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_1618_)
);

NAND2X1 _10001_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1619_)
);

OAI21X1 _10002_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1618_),
    .C(_1619_),
    .Y(_1563_[28])
);

INVX1 _10003_ (
    .A(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_1620_)
);

NAND2X1 _10004_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1621_)
);

OAI21X1 _10005_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1620_),
    .C(_1621_),
    .Y(_1563_[29])
);

INVX1 _10006_ (
    .A(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_1622_)
);

NAND2X1 _10007_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1623_)
);

OAI21X1 _10008_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1622_),
    .C(_1623_),
    .Y(_1563_[30])
);

INVX1 _10009_ (
    .A(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_1624_)
);

NAND2X1 _10010_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1625_)
);

OAI21X1 _10011_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1624_),
    .C(_1625_),
    .Y(_1563_[31])
);

DFFSR _10012_ (
    .CLK(clk_bF$buf113),
    .D(_1563_[0]),
    .Q(\datapath_1.regfile_1.regOut[25] [0]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _10013_ (
    .CLK(clk_bF$buf112),
    .D(_1563_[1]),
    .Q(\datapath_1.regfile_1.regOut[25] [1]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _10014_ (
    .CLK(clk_bF$buf111),
    .D(_1563_[2]),
    .Q(\datapath_1.regfile_1.regOut[25] [2]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _10015_ (
    .CLK(clk_bF$buf110),
    .D(_1563_[3]),
    .Q(\datapath_1.regfile_1.regOut[25] [3]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _10016_ (
    .CLK(clk_bF$buf109),
    .D(_1563_[4]),
    .Q(\datapath_1.regfile_1.regOut[25] [4]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _10017_ (
    .CLK(clk_bF$buf108),
    .D(_1563_[5]),
    .Q(\datapath_1.regfile_1.regOut[25] [5]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _10018_ (
    .CLK(clk_bF$buf107),
    .D(_1563_[6]),
    .Q(\datapath_1.regfile_1.regOut[25] [6]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _10019_ (
    .CLK(clk_bF$buf106),
    .D(_1563_[7]),
    .Q(\datapath_1.regfile_1.regOut[25] [7]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _10020_ (
    .CLK(clk_bF$buf105),
    .D(_1563_[8]),
    .Q(\datapath_1.regfile_1.regOut[25] [8]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _10021_ (
    .CLK(clk_bF$buf104),
    .D(_1563_[9]),
    .Q(\datapath_1.regfile_1.regOut[25] [9]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _10022_ (
    .CLK(clk_bF$buf103),
    .D(_1563_[10]),
    .Q(\datapath_1.regfile_1.regOut[25] [10]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _10023_ (
    .CLK(clk_bF$buf102),
    .D(_1563_[11]),
    .Q(\datapath_1.regfile_1.regOut[25] [11]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _10024_ (
    .CLK(clk_bF$buf101),
    .D(_1563_[12]),
    .Q(\datapath_1.regfile_1.regOut[25] [12]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _10025_ (
    .CLK(clk_bF$buf100),
    .D(_1563_[13]),
    .Q(\datapath_1.regfile_1.regOut[25] [13]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _10026_ (
    .CLK(clk_bF$buf99),
    .D(_1563_[14]),
    .Q(\datapath_1.regfile_1.regOut[25] [14]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _10027_ (
    .CLK(clk_bF$buf98),
    .D(_1563_[15]),
    .Q(\datapath_1.regfile_1.regOut[25] [15]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _10028_ (
    .CLK(clk_bF$buf97),
    .D(_1563_[16]),
    .Q(\datapath_1.regfile_1.regOut[25] [16]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _10029_ (
    .CLK(clk_bF$buf96),
    .D(_1563_[17]),
    .Q(\datapath_1.regfile_1.regOut[25] [17]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _10030_ (
    .CLK(clk_bF$buf95),
    .D(_1563_[18]),
    .Q(\datapath_1.regfile_1.regOut[25] [18]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _10031_ (
    .CLK(clk_bF$buf94),
    .D(_1563_[19]),
    .Q(\datapath_1.regfile_1.regOut[25] [19]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _10032_ (
    .CLK(clk_bF$buf93),
    .D(_1563_[20]),
    .Q(\datapath_1.regfile_1.regOut[25] [20]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _10033_ (
    .CLK(clk_bF$buf92),
    .D(_1563_[21]),
    .Q(\datapath_1.regfile_1.regOut[25] [21]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _10034_ (
    .CLK(clk_bF$buf91),
    .D(_1563_[22]),
    .Q(\datapath_1.regfile_1.regOut[25] [22]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _10035_ (
    .CLK(clk_bF$buf90),
    .D(_1563_[23]),
    .Q(\datapath_1.regfile_1.regOut[25] [23]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _10036_ (
    .CLK(clk_bF$buf89),
    .D(_1563_[24]),
    .Q(\datapath_1.regfile_1.regOut[25] [24]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _10037_ (
    .CLK(clk_bF$buf88),
    .D(_1563_[25]),
    .Q(\datapath_1.regfile_1.regOut[25] [25]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _10038_ (
    .CLK(clk_bF$buf87),
    .D(_1563_[26]),
    .Q(\datapath_1.regfile_1.regOut[25] [26]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _10039_ (
    .CLK(clk_bF$buf86),
    .D(_1563_[27]),
    .Q(\datapath_1.regfile_1.regOut[25] [27]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _10040_ (
    .CLK(clk_bF$buf85),
    .D(_1563_[28]),
    .Q(\datapath_1.regfile_1.regOut[25] [28]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _10041_ (
    .CLK(clk_bF$buf84),
    .D(_1563_[29]),
    .Q(\datapath_1.regfile_1.regOut[25] [29]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _10042_ (
    .CLK(clk_bF$buf83),
    .D(_1563_[30]),
    .Q(\datapath_1.regfile_1.regOut[25] [30]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _10043_ (
    .CLK(clk_bF$buf82),
    .D(_1563_[31]),
    .Q(\datapath_1.regfile_1.regOut[25] [31]),
    .R(rst_bF$buf82),
    .S(vdd)
);

INVX1 _10044_ (
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_1691_)
);

NAND2X1 _10045_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .Y(_1692_)
);

OAI21X1 _10046_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1691_),
    .C(_1692_),
    .Y(_1628_[0])
);

INVX1 _10047_ (
    .A(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_1629_)
);

NAND2X1 _10048_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1630_)
);

OAI21X1 _10049_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1629_),
    .C(_1630_),
    .Y(_1628_[1])
);

INVX1 _10050_ (
    .A(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_1631_)
);

NAND2X1 _10051_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1632_)
);

OAI21X1 _10052_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1631_),
    .C(_1632_),
    .Y(_1628_[2])
);

INVX1 _10053_ (
    .A(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_1633_)
);

NAND2X1 _10054_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1634_)
);

OAI21X1 _10055_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1633_),
    .C(_1634_),
    .Y(_1628_[3])
);

INVX1 _10056_ (
    .A(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_1635_)
);

NAND2X1 _10057_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1636_)
);

OAI21X1 _10058_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1635_),
    .C(_1636_),
    .Y(_1628_[4])
);

INVX1 _10059_ (
    .A(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_1637_)
);

NAND2X1 _10060_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1638_)
);

OAI21X1 _10061_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1637_),
    .C(_1638_),
    .Y(_1628_[5])
);

INVX1 _10062_ (
    .A(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_1639_)
);

NAND2X1 _10063_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1640_)
);

OAI21X1 _10064_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1639_),
    .C(_1640_),
    .Y(_1628_[6])
);

INVX1 _10065_ (
    .A(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_1641_)
);

NAND2X1 _10066_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1642_)
);

OAI21X1 _10067_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1641_),
    .C(_1642_),
    .Y(_1628_[7])
);

INVX1 _10068_ (
    .A(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_1643_)
);

NAND2X1 _10069_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1644_)
);

OAI21X1 _10070_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1643_),
    .C(_1644_),
    .Y(_1628_[8])
);

INVX1 _10071_ (
    .A(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_1645_)
);

NAND2X1 _10072_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1646_)
);

OAI21X1 _10073_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1645_),
    .C(_1646_),
    .Y(_1628_[9])
);

INVX1 _10074_ (
    .A(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_1647_)
);

NAND2X1 _10075_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1648_)
);

OAI21X1 _10076_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1647_),
    .C(_1648_),
    .Y(_1628_[10])
);

INVX1 _10077_ (
    .A(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_1649_)
);

NAND2X1 _10078_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1650_)
);

OAI21X1 _10079_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1649_),
    .C(_1650_),
    .Y(_1628_[11])
);

INVX1 _10080_ (
    .A(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_1651_)
);

NAND2X1 _10081_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1652_)
);

OAI21X1 _10082_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1651_),
    .C(_1652_),
    .Y(_1628_[12])
);

INVX1 _10083_ (
    .A(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_1653_)
);

NAND2X1 _10084_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1654_)
);

OAI21X1 _10085_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1653_),
    .C(_1654_),
    .Y(_1628_[13])
);

INVX1 _10086_ (
    .A(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_1655_)
);

NAND2X1 _10087_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1656_)
);

OAI21X1 _10088_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1655_),
    .C(_1656_),
    .Y(_1628_[14])
);

INVX1 _10089_ (
    .A(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_1657_)
);

NAND2X1 _10090_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1658_)
);

OAI21X1 _10091_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1657_),
    .C(_1658_),
    .Y(_1628_[15])
);

INVX1 _10092_ (
    .A(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_1659_)
);

NAND2X1 _10093_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1660_)
);

OAI21X1 _10094_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1659_),
    .C(_1660_),
    .Y(_1628_[16])
);

INVX1 _10095_ (
    .A(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_1661_)
);

NAND2X1 _10096_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1662_)
);

OAI21X1 _10097_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1661_),
    .C(_1662_),
    .Y(_1628_[17])
);

INVX1 _10098_ (
    .A(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_1663_)
);

NAND2X1 _10099_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1664_)
);

OAI21X1 _10100_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1663_),
    .C(_1664_),
    .Y(_1628_[18])
);

INVX1 _10101_ (
    .A(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_1665_)
);

NAND2X1 _10102_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1666_)
);

OAI21X1 _10103_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1665_),
    .C(_1666_),
    .Y(_1628_[19])
);

INVX1 _10104_ (
    .A(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_1667_)
);

NAND2X1 _10105_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1668_)
);

OAI21X1 _10106_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1667_),
    .C(_1668_),
    .Y(_1628_[20])
);

INVX1 _10107_ (
    .A(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_1669_)
);

NAND2X1 _10108_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1670_)
);

OAI21X1 _10109_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1669_),
    .C(_1670_),
    .Y(_1628_[21])
);

INVX1 _10110_ (
    .A(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_1671_)
);

NAND2X1 _10111_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1672_)
);

OAI21X1 _10112_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1671_),
    .C(_1672_),
    .Y(_1628_[22])
);

INVX1 _10113_ (
    .A(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_1673_)
);

NAND2X1 _10114_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1674_)
);

OAI21X1 _10115_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1673_),
    .C(_1674_),
    .Y(_1628_[23])
);

INVX1 _10116_ (
    .A(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_1675_)
);

NAND2X1 _10117_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1676_)
);

OAI21X1 _10118_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1675_),
    .C(_1676_),
    .Y(_1628_[24])
);

INVX1 _10119_ (
    .A(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_1677_)
);

NAND2X1 _10120_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1678_)
);

OAI21X1 _10121_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1677_),
    .C(_1678_),
    .Y(_1628_[25])
);

INVX1 _10122_ (
    .A(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_1679_)
);

NAND2X1 _10123_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1680_)
);

OAI21X1 _10124_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1679_),
    .C(_1680_),
    .Y(_1628_[26])
);

INVX1 _10125_ (
    .A(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_1681_)
);

NAND2X1 _10126_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1682_)
);

OAI21X1 _10127_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1681_),
    .C(_1682_),
    .Y(_1628_[27])
);

INVX1 _10128_ (
    .A(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_1683_)
);

NAND2X1 _10129_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1684_)
);

OAI21X1 _10130_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(_1683_),
    .C(_1684_),
    .Y(_1628_[28])
);

INVX1 _10131_ (
    .A(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_1685_)
);

NAND2X1 _10132_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_1686_)
);

OAI21X1 _10133_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(_1685_),
    .C(_1686_),
    .Y(_1628_[29])
);

INVX1 _10134_ (
    .A(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_1687_)
);

NAND2X1 _10135_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1688_)
);

OAI21X1 _10136_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(_1687_),
    .C(_1688_),
    .Y(_1628_[30])
);

INVX1 _10137_ (
    .A(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_1689_)
);

NAND2X1 _10138_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_1690_)
);

OAI21X1 _10139_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(_1689_),
    .C(_1690_),
    .Y(_1628_[31])
);

DFFSR _10140_ (
    .CLK(clk_bF$buf81),
    .D(_1628_[0]),
    .Q(\datapath_1.regfile_1.regOut[26] [0]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _10141_ (
    .CLK(clk_bF$buf80),
    .D(_1628_[1]),
    .Q(\datapath_1.regfile_1.regOut[26] [1]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _10142_ (
    .CLK(clk_bF$buf79),
    .D(_1628_[2]),
    .Q(\datapath_1.regfile_1.regOut[26] [2]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _10143_ (
    .CLK(clk_bF$buf78),
    .D(_1628_[3]),
    .Q(\datapath_1.regfile_1.regOut[26] [3]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _10144_ (
    .CLK(clk_bF$buf77),
    .D(_1628_[4]),
    .Q(\datapath_1.regfile_1.regOut[26] [4]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _10145_ (
    .CLK(clk_bF$buf76),
    .D(_1628_[5]),
    .Q(\datapath_1.regfile_1.regOut[26] [5]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _10146_ (
    .CLK(clk_bF$buf75),
    .D(_1628_[6]),
    .Q(\datapath_1.regfile_1.regOut[26] [6]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _10147_ (
    .CLK(clk_bF$buf74),
    .D(_1628_[7]),
    .Q(\datapath_1.regfile_1.regOut[26] [7]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _10148_ (
    .CLK(clk_bF$buf73),
    .D(_1628_[8]),
    .Q(\datapath_1.regfile_1.regOut[26] [8]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _10149_ (
    .CLK(clk_bF$buf72),
    .D(_1628_[9]),
    .Q(\datapath_1.regfile_1.regOut[26] [9]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _10150_ (
    .CLK(clk_bF$buf71),
    .D(_1628_[10]),
    .Q(\datapath_1.regfile_1.regOut[26] [10]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _10151_ (
    .CLK(clk_bF$buf70),
    .D(_1628_[11]),
    .Q(\datapath_1.regfile_1.regOut[26] [11]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _10152_ (
    .CLK(clk_bF$buf69),
    .D(_1628_[12]),
    .Q(\datapath_1.regfile_1.regOut[26] [12]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _10153_ (
    .CLK(clk_bF$buf68),
    .D(_1628_[13]),
    .Q(\datapath_1.regfile_1.regOut[26] [13]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _10154_ (
    .CLK(clk_bF$buf67),
    .D(_1628_[14]),
    .Q(\datapath_1.regfile_1.regOut[26] [14]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _10155_ (
    .CLK(clk_bF$buf66),
    .D(_1628_[15]),
    .Q(\datapath_1.regfile_1.regOut[26] [15]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _10156_ (
    .CLK(clk_bF$buf65),
    .D(_1628_[16]),
    .Q(\datapath_1.regfile_1.regOut[26] [16]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _10157_ (
    .CLK(clk_bF$buf64),
    .D(_1628_[17]),
    .Q(\datapath_1.regfile_1.regOut[26] [17]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _10158_ (
    .CLK(clk_bF$buf63),
    .D(_1628_[18]),
    .Q(\datapath_1.regfile_1.regOut[26] [18]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _10159_ (
    .CLK(clk_bF$buf62),
    .D(_1628_[19]),
    .Q(\datapath_1.regfile_1.regOut[26] [19]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _10160_ (
    .CLK(clk_bF$buf61),
    .D(_1628_[20]),
    .Q(\datapath_1.regfile_1.regOut[26] [20]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _10161_ (
    .CLK(clk_bF$buf60),
    .D(_1628_[21]),
    .Q(\datapath_1.regfile_1.regOut[26] [21]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _10162_ (
    .CLK(clk_bF$buf59),
    .D(_1628_[22]),
    .Q(\datapath_1.regfile_1.regOut[26] [22]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _10163_ (
    .CLK(clk_bF$buf58),
    .D(_1628_[23]),
    .Q(\datapath_1.regfile_1.regOut[26] [23]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _10164_ (
    .CLK(clk_bF$buf57),
    .D(_1628_[24]),
    .Q(\datapath_1.regfile_1.regOut[26] [24]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _10165_ (
    .CLK(clk_bF$buf56),
    .D(_1628_[25]),
    .Q(\datapath_1.regfile_1.regOut[26] [25]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _10166_ (
    .CLK(clk_bF$buf55),
    .D(_1628_[26]),
    .Q(\datapath_1.regfile_1.regOut[26] [26]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _10167_ (
    .CLK(clk_bF$buf54),
    .D(_1628_[27]),
    .Q(\datapath_1.regfile_1.regOut[26] [27]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _10168_ (
    .CLK(clk_bF$buf53),
    .D(_1628_[28]),
    .Q(\datapath_1.regfile_1.regOut[26] [28]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _10169_ (
    .CLK(clk_bF$buf52),
    .D(_1628_[29]),
    .Q(\datapath_1.regfile_1.regOut[26] [29]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _10170_ (
    .CLK(clk_bF$buf51),
    .D(_1628_[30]),
    .Q(\datapath_1.regfile_1.regOut[26] [30]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _10171_ (
    .CLK(clk_bF$buf50),
    .D(_1628_[31]),
    .Q(\datapath_1.regfile_1.regOut[26] [31]),
    .R(rst_bF$buf50),
    .S(vdd)
);

INVX1 _10172_ (
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_1756_)
);

NAND2X1 _10173_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .Y(_1757_)
);

OAI21X1 _10174_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1756_),
    .C(_1757_),
    .Y(_1693_[0])
);

INVX1 _10175_ (
    .A(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_1694_)
);

NAND2X1 _10176_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1695_)
);

OAI21X1 _10177_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1694_),
    .C(_1695_),
    .Y(_1693_[1])
);

INVX1 _10178_ (
    .A(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_1696_)
);

NAND2X1 _10179_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1697_)
);

OAI21X1 _10180_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1696_),
    .C(_1697_),
    .Y(_1693_[2])
);

INVX1 _10181_ (
    .A(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_1698_)
);

NAND2X1 _10182_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_1699_)
);

OAI21X1 _10183_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1698_),
    .C(_1699_),
    .Y(_1693_[3])
);

INVX1 _10184_ (
    .A(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_1700_)
);

NAND2X1 _10185_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1701_)
);

OAI21X1 _10186_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1700_),
    .C(_1701_),
    .Y(_1693_[4])
);

INVX1 _10187_ (
    .A(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_1702_)
);

NAND2X1 _10188_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1703_)
);

OAI21X1 _10189_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1702_),
    .C(_1703_),
    .Y(_1693_[5])
);

INVX1 _10190_ (
    .A(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_1704_)
);

NAND2X1 _10191_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1705_)
);

OAI21X1 _10192_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1704_),
    .C(_1705_),
    .Y(_1693_[6])
);

INVX1 _10193_ (
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_1706_)
);

NAND2X1 _10194_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1707_)
);

OAI21X1 _10195_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1706_),
    .C(_1707_),
    .Y(_1693_[7])
);

INVX1 _10196_ (
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_1708_)
);

NAND2X1 _10197_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1709_)
);

OAI21X1 _10198_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1708_),
    .C(_1709_),
    .Y(_1693_[8])
);

INVX1 _10199_ (
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_1710_)
);

NAND2X1 _10200_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1711_)
);

OAI21X1 _10201_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1710_),
    .C(_1711_),
    .Y(_1693_[9])
);

INVX1 _10202_ (
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_1712_)
);

NAND2X1 _10203_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1713_)
);

OAI21X1 _10204_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1712_),
    .C(_1713_),
    .Y(_1693_[10])
);

INVX1 _10205_ (
    .A(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_1714_)
);

NAND2X1 _10206_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1715_)
);

OAI21X1 _10207_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1714_),
    .C(_1715_),
    .Y(_1693_[11])
);

INVX1 _10208_ (
    .A(\datapath_1.regfile_1.regOut[27] [12]),
    .Y(_1716_)
);

NAND2X1 _10209_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1717_)
);

OAI21X1 _10210_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1716_),
    .C(_1717_),
    .Y(_1693_[12])
);

INVX1 _10211_ (
    .A(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_1718_)
);

NAND2X1 _10212_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1719_)
);

OAI21X1 _10213_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1718_),
    .C(_1719_),
    .Y(_1693_[13])
);

INVX1 _10214_ (
    .A(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_1720_)
);

NAND2X1 _10215_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1721_)
);

OAI21X1 _10216_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1720_),
    .C(_1721_),
    .Y(_1693_[14])
);

INVX1 _10217_ (
    .A(\datapath_1.regfile_1.regOut[27] [15]),
    .Y(_1722_)
);

NAND2X1 _10218_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1723_)
);

OAI21X1 _10219_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1722_),
    .C(_1723_),
    .Y(_1693_[15])
);

INVX1 _10220_ (
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_1724_)
);

NAND2X1 _10221_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1725_)
);

OAI21X1 _10222_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1724_),
    .C(_1725_),
    .Y(_1693_[16])
);

INVX1 _10223_ (
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_1726_)
);

NAND2X1 _10224_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1727_)
);

OAI21X1 _10225_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1726_),
    .C(_1727_),
    .Y(_1693_[17])
);

INVX1 _10226_ (
    .A(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_1728_)
);

NAND2X1 _10227_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1729_)
);

OAI21X1 _10228_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1728_),
    .C(_1729_),
    .Y(_1693_[18])
);

INVX1 _10229_ (
    .A(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_1730_)
);

NAND2X1 _10230_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1731_)
);

OAI21X1 _10231_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1730_),
    .C(_1731_),
    .Y(_1693_[19])
);

INVX1 _10232_ (
    .A(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_1732_)
);

NAND2X1 _10233_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1733_)
);

OAI21X1 _10234_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1732_),
    .C(_1733_),
    .Y(_1693_[20])
);

INVX1 _10235_ (
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_1734_)
);

NAND2X1 _10236_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1735_)
);

OAI21X1 _10237_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1734_),
    .C(_1735_),
    .Y(_1693_[21])
);

INVX1 _10238_ (
    .A(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_1736_)
);

NAND2X1 _10239_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1737_)
);

OAI21X1 _10240_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1736_),
    .C(_1737_),
    .Y(_1693_[22])
);

INVX1 _10241_ (
    .A(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_1738_)
);

NAND2X1 _10242_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1739_)
);

OAI21X1 _10243_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1738_),
    .C(_1739_),
    .Y(_1693_[23])
);

INVX1 _10244_ (
    .A(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_1740_)
);

NAND2X1 _10245_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1741_)
);

OAI21X1 _10246_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1740_),
    .C(_1741_),
    .Y(_1693_[24])
);

INVX1 _10247_ (
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_1742_)
);

NAND2X1 _10248_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_1743_)
);

OAI21X1 _10249_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1742_),
    .C(_1743_),
    .Y(_1693_[25])
);

INVX1 _10250_ (
    .A(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_1744_)
);

NAND2X1 _10251_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1745_)
);

OAI21X1 _10252_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1744_),
    .C(_1745_),
    .Y(_1693_[26])
);

INVX1 _10253_ (
    .A(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_1746_)
);

NAND2X1 _10254_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1747_)
);

OAI21X1 _10255_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1746_),
    .C(_1747_),
    .Y(_1693_[27])
);

INVX1 _10256_ (
    .A(\datapath_1.regfile_1.regOut[27] [28]),
    .Y(_1748_)
);

NAND2X1 _10257_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1749_)
);

OAI21X1 _10258_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(_1748_),
    .C(_1749_),
    .Y(_1693_[28])
);

INVX1 _10259_ (
    .A(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_1750_)
);

NAND2X1 _10260_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1751_)
);

OAI21X1 _10261_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(_1750_),
    .C(_1751_),
    .Y(_1693_[29])
);

INVX1 _10262_ (
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_1752_)
);

NAND2X1 _10263_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1753_)
);

OAI21X1 _10264_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(_1752_),
    .C(_1753_),
    .Y(_1693_[30])
);

INVX1 _10265_ (
    .A(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_1754_)
);

NAND2X1 _10266_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1755_)
);

OAI21X1 _10267_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(_1754_),
    .C(_1755_),
    .Y(_1693_[31])
);

DFFSR _10268_ (
    .CLK(clk_bF$buf49),
    .D(_1693_[0]),
    .Q(\datapath_1.regfile_1.regOut[27] [0]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _10269_ (
    .CLK(clk_bF$buf48),
    .D(_1693_[1]),
    .Q(\datapath_1.regfile_1.regOut[27] [1]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _10270_ (
    .CLK(clk_bF$buf47),
    .D(_1693_[2]),
    .Q(\datapath_1.regfile_1.regOut[27] [2]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _10271_ (
    .CLK(clk_bF$buf46),
    .D(_1693_[3]),
    .Q(\datapath_1.regfile_1.regOut[27] [3]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _10272_ (
    .CLK(clk_bF$buf45),
    .D(_1693_[4]),
    .Q(\datapath_1.regfile_1.regOut[27] [4]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _10273_ (
    .CLK(clk_bF$buf44),
    .D(_1693_[5]),
    .Q(\datapath_1.regfile_1.regOut[27] [5]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _10274_ (
    .CLK(clk_bF$buf43),
    .D(_1693_[6]),
    .Q(\datapath_1.regfile_1.regOut[27] [6]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _10275_ (
    .CLK(clk_bF$buf42),
    .D(_1693_[7]),
    .Q(\datapath_1.regfile_1.regOut[27] [7]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _10276_ (
    .CLK(clk_bF$buf41),
    .D(_1693_[8]),
    .Q(\datapath_1.regfile_1.regOut[27] [8]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _10277_ (
    .CLK(clk_bF$buf40),
    .D(_1693_[9]),
    .Q(\datapath_1.regfile_1.regOut[27] [9]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _10278_ (
    .CLK(clk_bF$buf39),
    .D(_1693_[10]),
    .Q(\datapath_1.regfile_1.regOut[27] [10]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _10279_ (
    .CLK(clk_bF$buf38),
    .D(_1693_[11]),
    .Q(\datapath_1.regfile_1.regOut[27] [11]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _10280_ (
    .CLK(clk_bF$buf37),
    .D(_1693_[12]),
    .Q(\datapath_1.regfile_1.regOut[27] [12]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _10281_ (
    .CLK(clk_bF$buf36),
    .D(_1693_[13]),
    .Q(\datapath_1.regfile_1.regOut[27] [13]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _10282_ (
    .CLK(clk_bF$buf35),
    .D(_1693_[14]),
    .Q(\datapath_1.regfile_1.regOut[27] [14]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _10283_ (
    .CLK(clk_bF$buf34),
    .D(_1693_[15]),
    .Q(\datapath_1.regfile_1.regOut[27] [15]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _10284_ (
    .CLK(clk_bF$buf33),
    .D(_1693_[16]),
    .Q(\datapath_1.regfile_1.regOut[27] [16]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _10285_ (
    .CLK(clk_bF$buf32),
    .D(_1693_[17]),
    .Q(\datapath_1.regfile_1.regOut[27] [17]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _10286_ (
    .CLK(clk_bF$buf31),
    .D(_1693_[18]),
    .Q(\datapath_1.regfile_1.regOut[27] [18]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _10287_ (
    .CLK(clk_bF$buf30),
    .D(_1693_[19]),
    .Q(\datapath_1.regfile_1.regOut[27] [19]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _10288_ (
    .CLK(clk_bF$buf29),
    .D(_1693_[20]),
    .Q(\datapath_1.regfile_1.regOut[27] [20]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _10289_ (
    .CLK(clk_bF$buf28),
    .D(_1693_[21]),
    .Q(\datapath_1.regfile_1.regOut[27] [21]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _10290_ (
    .CLK(clk_bF$buf27),
    .D(_1693_[22]),
    .Q(\datapath_1.regfile_1.regOut[27] [22]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _10291_ (
    .CLK(clk_bF$buf26),
    .D(_1693_[23]),
    .Q(\datapath_1.regfile_1.regOut[27] [23]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _10292_ (
    .CLK(clk_bF$buf25),
    .D(_1693_[24]),
    .Q(\datapath_1.regfile_1.regOut[27] [24]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _10293_ (
    .CLK(clk_bF$buf24),
    .D(_1693_[25]),
    .Q(\datapath_1.regfile_1.regOut[27] [25]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _10294_ (
    .CLK(clk_bF$buf23),
    .D(_1693_[26]),
    .Q(\datapath_1.regfile_1.regOut[27] [26]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _10295_ (
    .CLK(clk_bF$buf22),
    .D(_1693_[27]),
    .Q(\datapath_1.regfile_1.regOut[27] [27]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _10296_ (
    .CLK(clk_bF$buf21),
    .D(_1693_[28]),
    .Q(\datapath_1.regfile_1.regOut[27] [28]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _10297_ (
    .CLK(clk_bF$buf20),
    .D(_1693_[29]),
    .Q(\datapath_1.regfile_1.regOut[27] [29]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _10298_ (
    .CLK(clk_bF$buf19),
    .D(_1693_[30]),
    .Q(\datapath_1.regfile_1.regOut[27] [30]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _10299_ (
    .CLK(clk_bF$buf18),
    .D(_1693_[31]),
    .Q(\datapath_1.regfile_1.regOut[27] [31]),
    .R(rst_bF$buf18),
    .S(vdd)
);

INVX1 _10300_ (
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_1821_)
);

NAND2X1 _10301_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .Y(_1822_)
);

OAI21X1 _10302_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1821_),
    .C(_1822_),
    .Y(_1758_[0])
);

INVX1 _10303_ (
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .Y(_1759_)
);

NAND2X1 _10304_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1760_)
);

OAI21X1 _10305_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1759_),
    .C(_1760_),
    .Y(_1758_[1])
);

INVX1 _10306_ (
    .A(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_1761_)
);

NAND2X1 _10307_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1762_)
);

OAI21X1 _10308_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1761_),
    .C(_1762_),
    .Y(_1758_[2])
);

INVX1 _10309_ (
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .Y(_1763_)
);

NAND2X1 _10310_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1764_)
);

OAI21X1 _10311_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1763_),
    .C(_1764_),
    .Y(_1758_[3])
);

INVX1 _10312_ (
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_1765_)
);

NAND2X1 _10313_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1766_)
);

OAI21X1 _10314_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1765_),
    .C(_1766_),
    .Y(_1758_[4])
);

INVX1 _10315_ (
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_1767_)
);

NAND2X1 _10316_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1768_)
);

OAI21X1 _10317_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1767_),
    .C(_1768_),
    .Y(_1758_[5])
);

INVX1 _10318_ (
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_1769_)
);

NAND2X1 _10319_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1770_)
);

OAI21X1 _10320_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1769_),
    .C(_1770_),
    .Y(_1758_[6])
);

INVX1 _10321_ (
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .Y(_1771_)
);

NAND2X1 _10322_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1772_)
);

OAI21X1 _10323_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1771_),
    .C(_1772_),
    .Y(_1758_[7])
);

INVX1 _10324_ (
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_1773_)
);

NAND2X1 _10325_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1774_)
);

OAI21X1 _10326_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1773_),
    .C(_1774_),
    .Y(_1758_[8])
);

INVX1 _10327_ (
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_1775_)
);

NAND2X1 _10328_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1776_)
);

OAI21X1 _10329_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1775_),
    .C(_1776_),
    .Y(_1758_[9])
);

INVX1 _10330_ (
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_1777_)
);

NAND2X1 _10331_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1778_)
);

OAI21X1 _10332_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1777_),
    .C(_1778_),
    .Y(_1758_[10])
);

INVX1 _10333_ (
    .A(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_1779_)
);

NAND2X1 _10334_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1780_)
);

OAI21X1 _10335_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1779_),
    .C(_1780_),
    .Y(_1758_[11])
);

INVX1 _10336_ (
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_1781_)
);

NAND2X1 _10337_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1782_)
);

OAI21X1 _10338_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1781_),
    .C(_1782_),
    .Y(_1758_[12])
);

INVX1 _10339_ (
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_1783_)
);

NAND2X1 _10340_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1784_)
);

OAI21X1 _10341_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1783_),
    .C(_1784_),
    .Y(_1758_[13])
);

INVX1 _10342_ (
    .A(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_1785_)
);

NAND2X1 _10343_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1786_)
);

OAI21X1 _10344_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1785_),
    .C(_1786_),
    .Y(_1758_[14])
);

INVX1 _10345_ (
    .A(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_1787_)
);

NAND2X1 _10346_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1788_)
);

OAI21X1 _10347_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1787_),
    .C(_1788_),
    .Y(_1758_[15])
);

INVX1 _10348_ (
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_1789_)
);

NAND2X1 _10349_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1790_)
);

OAI21X1 _10350_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1789_),
    .C(_1790_),
    .Y(_1758_[16])
);

INVX1 _10351_ (
    .A(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_1791_)
);

NAND2X1 _10352_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1792_)
);

OAI21X1 _10353_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1791_),
    .C(_1792_),
    .Y(_1758_[17])
);

INVX1 _10354_ (
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_1793_)
);

NAND2X1 _10355_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1794_)
);

OAI21X1 _10356_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1793_),
    .C(_1794_),
    .Y(_1758_[18])
);

INVX1 _10357_ (
    .A(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_1795_)
);

NAND2X1 _10358_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1796_)
);

OAI21X1 _10359_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1795_),
    .C(_1796_),
    .Y(_1758_[19])
);

INVX1 _10360_ (
    .A(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_1797_)
);

NAND2X1 _10361_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1798_)
);

OAI21X1 _10362_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1797_),
    .C(_1798_),
    .Y(_1758_[20])
);

INVX1 _10363_ (
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .Y(_1799_)
);

NAND2X1 _10364_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1800_)
);

OAI21X1 _10365_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1799_),
    .C(_1800_),
    .Y(_1758_[21])
);

INVX1 _10366_ (
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_1801_)
);

NAND2X1 _10367_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1802_)
);

OAI21X1 _10368_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1801_),
    .C(_1802_),
    .Y(_1758_[22])
);

INVX1 _10369_ (
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_1803_)
);

NAND2X1 _10370_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1804_)
);

OAI21X1 _10371_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1803_),
    .C(_1804_),
    .Y(_1758_[23])
);

INVX1 _10372_ (
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_1805_)
);

NAND2X1 _10373_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1806_)
);

OAI21X1 _10374_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1805_),
    .C(_1806_),
    .Y(_1758_[24])
);

INVX1 _10375_ (
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_1807_)
);

NAND2X1 _10376_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1808_)
);

OAI21X1 _10377_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1807_),
    .C(_1808_),
    .Y(_1758_[25])
);

INVX1 _10378_ (
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_1809_)
);

NAND2X1 _10379_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1810_)
);

OAI21X1 _10380_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1809_),
    .C(_1810_),
    .Y(_1758_[26])
);

INVX1 _10381_ (
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_1811_)
);

NAND2X1 _10382_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1812_)
);

OAI21X1 _10383_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1811_),
    .C(_1812_),
    .Y(_1758_[27])
);

INVX1 _10384_ (
    .A(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_1813_)
);

NAND2X1 _10385_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1814_)
);

OAI21X1 _10386_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(_1813_),
    .C(_1814_),
    .Y(_1758_[28])
);

INVX1 _10387_ (
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_1815_)
);

NAND2X1 _10388_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1816_)
);

OAI21X1 _10389_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(_1815_),
    .C(_1816_),
    .Y(_1758_[29])
);

INVX1 _10390_ (
    .A(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_1817_)
);

NAND2X1 _10391_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1818_)
);

OAI21X1 _10392_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(_1817_),
    .C(_1818_),
    .Y(_1758_[30])
);

INVX1 _10393_ (
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_1819_)
);

NAND2X1 _10394_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1820_)
);

OAI21X1 _10395_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(_1819_),
    .C(_1820_),
    .Y(_1758_[31])
);

DFFSR _10396_ (
    .CLK(clk_bF$buf17),
    .D(_1758_[0]),
    .Q(\datapath_1.regfile_1.regOut[28] [0]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _10397_ (
    .CLK(clk_bF$buf16),
    .D(_1758_[1]),
    .Q(\datapath_1.regfile_1.regOut[28] [1]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _10398_ (
    .CLK(clk_bF$buf15),
    .D(_1758_[2]),
    .Q(\datapath_1.regfile_1.regOut[28] [2]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _10399_ (
    .CLK(clk_bF$buf14),
    .D(_1758_[3]),
    .Q(\datapath_1.regfile_1.regOut[28] [3]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _10400_ (
    .CLK(clk_bF$buf13),
    .D(_1758_[4]),
    .Q(\datapath_1.regfile_1.regOut[28] [4]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _10401_ (
    .CLK(clk_bF$buf12),
    .D(_1758_[5]),
    .Q(\datapath_1.regfile_1.regOut[28] [5]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _10402_ (
    .CLK(clk_bF$buf11),
    .D(_1758_[6]),
    .Q(\datapath_1.regfile_1.regOut[28] [6]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _10403_ (
    .CLK(clk_bF$buf10),
    .D(_1758_[7]),
    .Q(\datapath_1.regfile_1.regOut[28] [7]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _10404_ (
    .CLK(clk_bF$buf9),
    .D(_1758_[8]),
    .Q(\datapath_1.regfile_1.regOut[28] [8]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _10405_ (
    .CLK(clk_bF$buf8),
    .D(_1758_[9]),
    .Q(\datapath_1.regfile_1.regOut[28] [9]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _10406_ (
    .CLK(clk_bF$buf7),
    .D(_1758_[10]),
    .Q(\datapath_1.regfile_1.regOut[28] [10]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _10407_ (
    .CLK(clk_bF$buf6),
    .D(_1758_[11]),
    .Q(\datapath_1.regfile_1.regOut[28] [11]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _10408_ (
    .CLK(clk_bF$buf5),
    .D(_1758_[12]),
    .Q(\datapath_1.regfile_1.regOut[28] [12]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _10409_ (
    .CLK(clk_bF$buf4),
    .D(_1758_[13]),
    .Q(\datapath_1.regfile_1.regOut[28] [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _10410_ (
    .CLK(clk_bF$buf3),
    .D(_1758_[14]),
    .Q(\datapath_1.regfile_1.regOut[28] [14]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _10411_ (
    .CLK(clk_bF$buf2),
    .D(_1758_[15]),
    .Q(\datapath_1.regfile_1.regOut[28] [15]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _10412_ (
    .CLK(clk_bF$buf1),
    .D(_1758_[16]),
    .Q(\datapath_1.regfile_1.regOut[28] [16]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _10413_ (
    .CLK(clk_bF$buf0),
    .D(_1758_[17]),
    .Q(\datapath_1.regfile_1.regOut[28] [17]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _10414_ (
    .CLK(clk_bF$buf113),
    .D(_1758_[18]),
    .Q(\datapath_1.regfile_1.regOut[28] [18]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _10415_ (
    .CLK(clk_bF$buf112),
    .D(_1758_[19]),
    .Q(\datapath_1.regfile_1.regOut[28] [19]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _10416_ (
    .CLK(clk_bF$buf111),
    .D(_1758_[20]),
    .Q(\datapath_1.regfile_1.regOut[28] [20]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _10417_ (
    .CLK(clk_bF$buf110),
    .D(_1758_[21]),
    .Q(\datapath_1.regfile_1.regOut[28] [21]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _10418_ (
    .CLK(clk_bF$buf109),
    .D(_1758_[22]),
    .Q(\datapath_1.regfile_1.regOut[28] [22]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _10419_ (
    .CLK(clk_bF$buf108),
    .D(_1758_[23]),
    .Q(\datapath_1.regfile_1.regOut[28] [23]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _10420_ (
    .CLK(clk_bF$buf107),
    .D(_1758_[24]),
    .Q(\datapath_1.regfile_1.regOut[28] [24]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _10421_ (
    .CLK(clk_bF$buf106),
    .D(_1758_[25]),
    .Q(\datapath_1.regfile_1.regOut[28] [25]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _10422_ (
    .CLK(clk_bF$buf105),
    .D(_1758_[26]),
    .Q(\datapath_1.regfile_1.regOut[28] [26]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _10423_ (
    .CLK(clk_bF$buf104),
    .D(_1758_[27]),
    .Q(\datapath_1.regfile_1.regOut[28] [27]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _10424_ (
    .CLK(clk_bF$buf103),
    .D(_1758_[28]),
    .Q(\datapath_1.regfile_1.regOut[28] [28]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _10425_ (
    .CLK(clk_bF$buf102),
    .D(_1758_[29]),
    .Q(\datapath_1.regfile_1.regOut[28] [29]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _10426_ (
    .CLK(clk_bF$buf101),
    .D(_1758_[30]),
    .Q(\datapath_1.regfile_1.regOut[28] [30]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _10427_ (
    .CLK(clk_bF$buf100),
    .D(_1758_[31]),
    .Q(\datapath_1.regfile_1.regOut[28] [31]),
    .R(rst_bF$buf100),
    .S(vdd)
);

INVX1 _10428_ (
    .A(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_1886_)
);

NAND2X1 _10429_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .Y(_1887_)
);

OAI21X1 _10430_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1886_),
    .C(_1887_),
    .Y(_1823_[0])
);

INVX1 _10431_ (
    .A(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_1824_)
);

NAND2X1 _10432_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1825_)
);

OAI21X1 _10433_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1824_),
    .C(_1825_),
    .Y(_1823_[1])
);

INVX1 _10434_ (
    .A(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_1826_)
);

NAND2X1 _10435_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1827_)
);

OAI21X1 _10436_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1826_),
    .C(_1827_),
    .Y(_1823_[2])
);

INVX1 _10437_ (
    .A(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_1828_)
);

NAND2X1 _10438_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1829_)
);

OAI21X1 _10439_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1828_),
    .C(_1829_),
    .Y(_1823_[3])
);

INVX1 _10440_ (
    .A(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_1830_)
);

NAND2X1 _10441_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1831_)
);

OAI21X1 _10442_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1830_),
    .C(_1831_),
    .Y(_1823_[4])
);

INVX1 _10443_ (
    .A(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_1832_)
);

NAND2X1 _10444_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1833_)
);

OAI21X1 _10445_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1832_),
    .C(_1833_),
    .Y(_1823_[5])
);

INVX1 _10446_ (
    .A(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_1834_)
);

NAND2X1 _10447_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1835_)
);

OAI21X1 _10448_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1834_),
    .C(_1835_),
    .Y(_1823_[6])
);

INVX1 _10449_ (
    .A(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_1836_)
);

NAND2X1 _10450_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1837_)
);

OAI21X1 _10451_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1836_),
    .C(_1837_),
    .Y(_1823_[7])
);

INVX1 _10452_ (
    .A(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_1838_)
);

NAND2X1 _10453_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1839_)
);

OAI21X1 _10454_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1838_),
    .C(_1839_),
    .Y(_1823_[8])
);

INVX1 _10455_ (
    .A(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_1840_)
);

NAND2X1 _10456_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1841_)
);

OAI21X1 _10457_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1840_),
    .C(_1841_),
    .Y(_1823_[9])
);

INVX1 _10458_ (
    .A(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_1842_)
);

NAND2X1 _10459_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1843_)
);

OAI21X1 _10460_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1842_),
    .C(_1843_),
    .Y(_1823_[10])
);

INVX1 _10461_ (
    .A(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_1844_)
);

NAND2X1 _10462_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1845_)
);

OAI21X1 _10463_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1844_),
    .C(_1845_),
    .Y(_1823_[11])
);

INVX1 _10464_ (
    .A(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_1846_)
);

NAND2X1 _10465_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1847_)
);

OAI21X1 _10466_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1846_),
    .C(_1847_),
    .Y(_1823_[12])
);

INVX1 _10467_ (
    .A(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_1848_)
);

NAND2X1 _10468_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1849_)
);

OAI21X1 _10469_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1848_),
    .C(_1849_),
    .Y(_1823_[13])
);

INVX1 _10470_ (
    .A(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_1850_)
);

NAND2X1 _10471_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1851_)
);

OAI21X1 _10472_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1850_),
    .C(_1851_),
    .Y(_1823_[14])
);

INVX1 _10473_ (
    .A(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_1852_)
);

NAND2X1 _10474_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1853_)
);

OAI21X1 _10475_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1852_),
    .C(_1853_),
    .Y(_1823_[15])
);

INVX1 _10476_ (
    .A(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_1854_)
);

NAND2X1 _10477_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1855_)
);

OAI21X1 _10478_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1854_),
    .C(_1855_),
    .Y(_1823_[16])
);

INVX1 _10479_ (
    .A(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_1856_)
);

NAND2X1 _10480_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1857_)
);

OAI21X1 _10481_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1856_),
    .C(_1857_),
    .Y(_1823_[17])
);

INVX1 _10482_ (
    .A(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_1858_)
);

NAND2X1 _10483_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1859_)
);

OAI21X1 _10484_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1858_),
    .C(_1859_),
    .Y(_1823_[18])
);

INVX1 _10485_ (
    .A(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_1860_)
);

NAND2X1 _10486_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1861_)
);

OAI21X1 _10487_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1860_),
    .C(_1861_),
    .Y(_1823_[19])
);

INVX1 _10488_ (
    .A(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_1862_)
);

NAND2X1 _10489_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1863_)
);

OAI21X1 _10490_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1862_),
    .C(_1863_),
    .Y(_1823_[20])
);

INVX1 _10491_ (
    .A(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_1864_)
);

NAND2X1 _10492_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1865_)
);

OAI21X1 _10493_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1864_),
    .C(_1865_),
    .Y(_1823_[21])
);

INVX1 _10494_ (
    .A(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_1866_)
);

NAND2X1 _10495_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_1867_)
);

OAI21X1 _10496_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1866_),
    .C(_1867_),
    .Y(_1823_[22])
);

INVX1 _10497_ (
    .A(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_1868_)
);

NAND2X1 _10498_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1869_)
);

OAI21X1 _10499_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1868_),
    .C(_1869_),
    .Y(_1823_[23])
);

INVX1 _10500_ (
    .A(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_1870_)
);

NAND2X1 _10501_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1871_)
);

OAI21X1 _10502_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1870_),
    .C(_1871_),
    .Y(_1823_[24])
);

INVX1 _10503_ (
    .A(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_1872_)
);

NAND2X1 _10504_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1873_)
);

OAI21X1 _10505_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1872_),
    .C(_1873_),
    .Y(_1823_[25])
);

INVX1 _10506_ (
    .A(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_1874_)
);

NAND2X1 _10507_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1875_)
);

OAI21X1 _10508_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1874_),
    .C(_1875_),
    .Y(_1823_[26])
);

INVX1 _10509_ (
    .A(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_1876_)
);

NAND2X1 _10510_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1877_)
);

OAI21X1 _10511_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1876_),
    .C(_1877_),
    .Y(_1823_[27])
);

INVX1 _10512_ (
    .A(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_1878_)
);

NAND2X1 _10513_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1879_)
);

OAI21X1 _10514_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(_1878_),
    .C(_1879_),
    .Y(_1823_[28])
);

INVX1 _10515_ (
    .A(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_1880_)
);

NAND2X1 _10516_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1881_)
);

OAI21X1 _10517_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(_1880_),
    .C(_1881_),
    .Y(_1823_[29])
);

INVX1 _10518_ (
    .A(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_1882_)
);

NAND2X1 _10519_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1883_)
);

OAI21X1 _10520_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(_1882_),
    .C(_1883_),
    .Y(_1823_[30])
);

INVX1 _10521_ (
    .A(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_1884_)
);

NAND2X1 _10522_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1885_)
);

OAI21X1 _10523_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(_1884_),
    .C(_1885_),
    .Y(_1823_[31])
);

DFFSR _10524_ (
    .CLK(clk_bF$buf99),
    .D(_1823_[0]),
    .Q(\datapath_1.regfile_1.regOut[29] [0]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _10525_ (
    .CLK(clk_bF$buf98),
    .D(_1823_[1]),
    .Q(\datapath_1.regfile_1.regOut[29] [1]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _10526_ (
    .CLK(clk_bF$buf97),
    .D(_1823_[2]),
    .Q(\datapath_1.regfile_1.regOut[29] [2]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _10527_ (
    .CLK(clk_bF$buf96),
    .D(_1823_[3]),
    .Q(\datapath_1.regfile_1.regOut[29] [3]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _10528_ (
    .CLK(clk_bF$buf95),
    .D(_1823_[4]),
    .Q(\datapath_1.regfile_1.regOut[29] [4]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _10529_ (
    .CLK(clk_bF$buf94),
    .D(_1823_[5]),
    .Q(\datapath_1.regfile_1.regOut[29] [5]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _10530_ (
    .CLK(clk_bF$buf93),
    .D(_1823_[6]),
    .Q(\datapath_1.regfile_1.regOut[29] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _10531_ (
    .CLK(clk_bF$buf92),
    .D(_1823_[7]),
    .Q(\datapath_1.regfile_1.regOut[29] [7]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _10532_ (
    .CLK(clk_bF$buf91),
    .D(_1823_[8]),
    .Q(\datapath_1.regfile_1.regOut[29] [8]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _10533_ (
    .CLK(clk_bF$buf90),
    .D(_1823_[9]),
    .Q(\datapath_1.regfile_1.regOut[29] [9]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _10534_ (
    .CLK(clk_bF$buf89),
    .D(_1823_[10]),
    .Q(\datapath_1.regfile_1.regOut[29] [10]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _10535_ (
    .CLK(clk_bF$buf88),
    .D(_1823_[11]),
    .Q(\datapath_1.regfile_1.regOut[29] [11]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _10536_ (
    .CLK(clk_bF$buf87),
    .D(_1823_[12]),
    .Q(\datapath_1.regfile_1.regOut[29] [12]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _10537_ (
    .CLK(clk_bF$buf86),
    .D(_1823_[13]),
    .Q(\datapath_1.regfile_1.regOut[29] [13]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _10538_ (
    .CLK(clk_bF$buf85),
    .D(_1823_[14]),
    .Q(\datapath_1.regfile_1.regOut[29] [14]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _10539_ (
    .CLK(clk_bF$buf84),
    .D(_1823_[15]),
    .Q(\datapath_1.regfile_1.regOut[29] [15]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _10540_ (
    .CLK(clk_bF$buf83),
    .D(_1823_[16]),
    .Q(\datapath_1.regfile_1.regOut[29] [16]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _10541_ (
    .CLK(clk_bF$buf82),
    .D(_1823_[17]),
    .Q(\datapath_1.regfile_1.regOut[29] [17]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _10542_ (
    .CLK(clk_bF$buf81),
    .D(_1823_[18]),
    .Q(\datapath_1.regfile_1.regOut[29] [18]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _10543_ (
    .CLK(clk_bF$buf80),
    .D(_1823_[19]),
    .Q(\datapath_1.regfile_1.regOut[29] [19]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _10544_ (
    .CLK(clk_bF$buf79),
    .D(_1823_[20]),
    .Q(\datapath_1.regfile_1.regOut[29] [20]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _10545_ (
    .CLK(clk_bF$buf78),
    .D(_1823_[21]),
    .Q(\datapath_1.regfile_1.regOut[29] [21]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _10546_ (
    .CLK(clk_bF$buf77),
    .D(_1823_[22]),
    .Q(\datapath_1.regfile_1.regOut[29] [22]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _10547_ (
    .CLK(clk_bF$buf76),
    .D(_1823_[23]),
    .Q(\datapath_1.regfile_1.regOut[29] [23]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _10548_ (
    .CLK(clk_bF$buf75),
    .D(_1823_[24]),
    .Q(\datapath_1.regfile_1.regOut[29] [24]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _10549_ (
    .CLK(clk_bF$buf74),
    .D(_1823_[25]),
    .Q(\datapath_1.regfile_1.regOut[29] [25]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _10550_ (
    .CLK(clk_bF$buf73),
    .D(_1823_[26]),
    .Q(\datapath_1.regfile_1.regOut[29] [26]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _10551_ (
    .CLK(clk_bF$buf72),
    .D(_1823_[27]),
    .Q(\datapath_1.regfile_1.regOut[29] [27]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _10552_ (
    .CLK(clk_bF$buf71),
    .D(_1823_[28]),
    .Q(\datapath_1.regfile_1.regOut[29] [28]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _10553_ (
    .CLK(clk_bF$buf70),
    .D(_1823_[29]),
    .Q(\datapath_1.regfile_1.regOut[29] [29]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _10554_ (
    .CLK(clk_bF$buf69),
    .D(_1823_[30]),
    .Q(\datapath_1.regfile_1.regOut[29] [30]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _10555_ (
    .CLK(clk_bF$buf68),
    .D(_1823_[31]),
    .Q(\datapath_1.regfile_1.regOut[29] [31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

INVX1 _10556_ (
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .Y(_1951_)
);

NAND2X1 _10557_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .Y(_1952_)
);

OAI21X1 _10558_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1951_),
    .C(_1952_),
    .Y(_1888_[0])
);

INVX1 _10559_ (
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_1889_)
);

NAND2X1 _10560_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1890_)
);

OAI21X1 _10561_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1889_),
    .C(_1890_),
    .Y(_1888_[1])
);

INVX1 _10562_ (
    .A(\datapath_1.regfile_1.regOut[30] [2]),
    .Y(_1891_)
);

NAND2X1 _10563_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1892_)
);

OAI21X1 _10564_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1891_),
    .C(_1892_),
    .Y(_1888_[2])
);

INVX1 _10565_ (
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_1893_)
);

NAND2X1 _10566_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1894_)
);

OAI21X1 _10567_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1893_),
    .C(_1894_),
    .Y(_1888_[3])
);

INVX1 _10568_ (
    .A(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_1895_)
);

NAND2X1 _10569_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1896_)
);

OAI21X1 _10570_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1895_),
    .C(_1896_),
    .Y(_1888_[4])
);

INVX1 _10571_ (
    .A(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_1897_)
);

NAND2X1 _10572_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1898_)
);

OAI21X1 _10573_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1897_),
    .C(_1898_),
    .Y(_1888_[5])
);

INVX1 _10574_ (
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_1899_)
);

NAND2X1 _10575_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1900_)
);

OAI21X1 _10576_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1899_),
    .C(_1900_),
    .Y(_1888_[6])
);

INVX1 _10577_ (
    .A(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_1901_)
);

NAND2X1 _10578_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1902_)
);

OAI21X1 _10579_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1901_),
    .C(_1902_),
    .Y(_1888_[7])
);

INVX1 _10580_ (
    .A(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_1903_)
);

NAND2X1 _10581_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1904_)
);

OAI21X1 _10582_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1903_),
    .C(_1904_),
    .Y(_1888_[8])
);

INVX1 _10583_ (
    .A(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_1905_)
);

NAND2X1 _10584_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1906_)
);

OAI21X1 _10585_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1905_),
    .C(_1906_),
    .Y(_1888_[9])
);

INVX1 _10586_ (
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_1907_)
);

NAND2X1 _10587_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1908_)
);

OAI21X1 _10588_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1907_),
    .C(_1908_),
    .Y(_1888_[10])
);

INVX1 _10589_ (
    .A(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_1909_)
);

NAND2X1 _10590_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1910_)
);

OAI21X1 _10591_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1909_),
    .C(_1910_),
    .Y(_1888_[11])
);

INVX1 _10592_ (
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_1911_)
);

NAND2X1 _10593_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1912_)
);

OAI21X1 _10594_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1911_),
    .C(_1912_),
    .Y(_1888_[12])
);

INVX1 _10595_ (
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_1913_)
);

NAND2X1 _10596_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1914_)
);

OAI21X1 _10597_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1913_),
    .C(_1914_),
    .Y(_1888_[13])
);

INVX1 _10598_ (
    .A(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_1915_)
);

NAND2X1 _10599_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1916_)
);

OAI21X1 _10600_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1915_),
    .C(_1916_),
    .Y(_1888_[14])
);

INVX1 _10601_ (
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_1917_)
);

NAND2X1 _10602_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1918_)
);

OAI21X1 _10603_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1917_),
    .C(_1918_),
    .Y(_1888_[15])
);

INVX1 _10604_ (
    .A(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_1919_)
);

NAND2X1 _10605_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1920_)
);

OAI21X1 _10606_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1919_),
    .C(_1920_),
    .Y(_1888_[16])
);

INVX1 _10607_ (
    .A(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_1921_)
);

NAND2X1 _10608_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1922_)
);

OAI21X1 _10609_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1921_),
    .C(_1922_),
    .Y(_1888_[17])
);

INVX1 _10610_ (
    .A(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_1923_)
);

NAND2X1 _10611_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1924_)
);

OAI21X1 _10612_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1923_),
    .C(_1924_),
    .Y(_1888_[18])
);

INVX1 _10613_ (
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_1925_)
);

NAND2X1 _10614_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1926_)
);

OAI21X1 _10615_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1925_),
    .C(_1926_),
    .Y(_1888_[19])
);

INVX1 _10616_ (
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_1927_)
);

NAND2X1 _10617_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1928_)
);

OAI21X1 _10618_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1927_),
    .C(_1928_),
    .Y(_1888_[20])
);

INVX1 _10619_ (
    .A(\datapath_1.regfile_1.regOut[30] [21]),
    .Y(_1929_)
);

NAND2X1 _10620_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1930_)
);

OAI21X1 _10621_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1929_),
    .C(_1930_),
    .Y(_1888_[21])
);

INVX1 _10622_ (
    .A(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_1931_)
);

NAND2X1 _10623_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1932_)
);

OAI21X1 _10624_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1931_),
    .C(_1932_),
    .Y(_1888_[22])
);

INVX1 _10625_ (
    .A(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_1933_)
);

NAND2X1 _10626_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1934_)
);

OAI21X1 _10627_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1933_),
    .C(_1934_),
    .Y(_1888_[23])
);

INVX1 _10628_ (
    .A(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_1935_)
);

NAND2X1 _10629_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1936_)
);

OAI21X1 _10630_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1935_),
    .C(_1936_),
    .Y(_1888_[24])
);

INVX1 _10631_ (
    .A(\datapath_1.regfile_1.regOut[30] [25]),
    .Y(_1937_)
);

NAND2X1 _10632_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1938_)
);

OAI21X1 _10633_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1937_),
    .C(_1938_),
    .Y(_1888_[25])
);

INVX1 _10634_ (
    .A(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_1939_)
);

NAND2X1 _10635_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1940_)
);

OAI21X1 _10636_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1939_),
    .C(_1940_),
    .Y(_1888_[26])
);

INVX1 _10637_ (
    .A(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_1941_)
);

NAND2X1 _10638_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1942_)
);

OAI21X1 _10639_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1941_),
    .C(_1942_),
    .Y(_1888_[27])
);

INVX1 _10640_ (
    .A(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_1943_)
);

NAND2X1 _10641_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1944_)
);

OAI21X1 _10642_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(_1943_),
    .C(_1944_),
    .Y(_1888_[28])
);

INVX1 _10643_ (
    .A(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_1945_)
);

NAND2X1 _10644_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1946_)
);

OAI21X1 _10645_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(_1945_),
    .C(_1946_),
    .Y(_1888_[29])
);

INVX1 _10646_ (
    .A(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_1947_)
);

NAND2X1 _10647_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1948_)
);

OAI21X1 _10648_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(_1947_),
    .C(_1948_),
    .Y(_1888_[30])
);

INVX1 _10649_ (
    .A(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_1949_)
);

NAND2X1 _10650_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1950_)
);

OAI21X1 _10651_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(_1949_),
    .C(_1950_),
    .Y(_1888_[31])
);

DFFSR _10652_ (
    .CLK(clk_bF$buf67),
    .D(_1888_[0]),
    .Q(\datapath_1.regfile_1.regOut[30] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _10653_ (
    .CLK(clk_bF$buf66),
    .D(_1888_[1]),
    .Q(\datapath_1.regfile_1.regOut[30] [1]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _10654_ (
    .CLK(clk_bF$buf65),
    .D(_1888_[2]),
    .Q(\datapath_1.regfile_1.regOut[30] [2]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _10655_ (
    .CLK(clk_bF$buf64),
    .D(_1888_[3]),
    .Q(\datapath_1.regfile_1.regOut[30] [3]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _10656_ (
    .CLK(clk_bF$buf63),
    .D(_1888_[4]),
    .Q(\datapath_1.regfile_1.regOut[30] [4]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _10657_ (
    .CLK(clk_bF$buf62),
    .D(_1888_[5]),
    .Q(\datapath_1.regfile_1.regOut[30] [5]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _10658_ (
    .CLK(clk_bF$buf61),
    .D(_1888_[6]),
    .Q(\datapath_1.regfile_1.regOut[30] [6]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _10659_ (
    .CLK(clk_bF$buf60),
    .D(_1888_[7]),
    .Q(\datapath_1.regfile_1.regOut[30] [7]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _10660_ (
    .CLK(clk_bF$buf59),
    .D(_1888_[8]),
    .Q(\datapath_1.regfile_1.regOut[30] [8]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _10661_ (
    .CLK(clk_bF$buf58),
    .D(_1888_[9]),
    .Q(\datapath_1.regfile_1.regOut[30] [9]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _10662_ (
    .CLK(clk_bF$buf57),
    .D(_1888_[10]),
    .Q(\datapath_1.regfile_1.regOut[30] [10]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _10663_ (
    .CLK(clk_bF$buf56),
    .D(_1888_[11]),
    .Q(\datapath_1.regfile_1.regOut[30] [11]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _10664_ (
    .CLK(clk_bF$buf55),
    .D(_1888_[12]),
    .Q(\datapath_1.regfile_1.regOut[30] [12]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _10665_ (
    .CLK(clk_bF$buf54),
    .D(_1888_[13]),
    .Q(\datapath_1.regfile_1.regOut[30] [13]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _10666_ (
    .CLK(clk_bF$buf53),
    .D(_1888_[14]),
    .Q(\datapath_1.regfile_1.regOut[30] [14]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _10667_ (
    .CLK(clk_bF$buf52),
    .D(_1888_[15]),
    .Q(\datapath_1.regfile_1.regOut[30] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _10668_ (
    .CLK(clk_bF$buf51),
    .D(_1888_[16]),
    .Q(\datapath_1.regfile_1.regOut[30] [16]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _10669_ (
    .CLK(clk_bF$buf50),
    .D(_1888_[17]),
    .Q(\datapath_1.regfile_1.regOut[30] [17]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _10670_ (
    .CLK(clk_bF$buf49),
    .D(_1888_[18]),
    .Q(\datapath_1.regfile_1.regOut[30] [18]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _10671_ (
    .CLK(clk_bF$buf48),
    .D(_1888_[19]),
    .Q(\datapath_1.regfile_1.regOut[30] [19]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _10672_ (
    .CLK(clk_bF$buf47),
    .D(_1888_[20]),
    .Q(\datapath_1.regfile_1.regOut[30] [20]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _10673_ (
    .CLK(clk_bF$buf46),
    .D(_1888_[21]),
    .Q(\datapath_1.regfile_1.regOut[30] [21]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _10674_ (
    .CLK(clk_bF$buf45),
    .D(_1888_[22]),
    .Q(\datapath_1.regfile_1.regOut[30] [22]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _10675_ (
    .CLK(clk_bF$buf44),
    .D(_1888_[23]),
    .Q(\datapath_1.regfile_1.regOut[30] [23]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _10676_ (
    .CLK(clk_bF$buf43),
    .D(_1888_[24]),
    .Q(\datapath_1.regfile_1.regOut[30] [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _10677_ (
    .CLK(clk_bF$buf42),
    .D(_1888_[25]),
    .Q(\datapath_1.regfile_1.regOut[30] [25]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _10678_ (
    .CLK(clk_bF$buf41),
    .D(_1888_[26]),
    .Q(\datapath_1.regfile_1.regOut[30] [26]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _10679_ (
    .CLK(clk_bF$buf40),
    .D(_1888_[27]),
    .Q(\datapath_1.regfile_1.regOut[30] [27]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _10680_ (
    .CLK(clk_bF$buf39),
    .D(_1888_[28]),
    .Q(\datapath_1.regfile_1.regOut[30] [28]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _10681_ (
    .CLK(clk_bF$buf38),
    .D(_1888_[29]),
    .Q(\datapath_1.regfile_1.regOut[30] [29]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _10682_ (
    .CLK(clk_bF$buf37),
    .D(_1888_[30]),
    .Q(\datapath_1.regfile_1.regOut[30] [30]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _10683_ (
    .CLK(clk_bF$buf36),
    .D(_1888_[31]),
    .Q(\datapath_1.regfile_1.regOut[30] [31]),
    .R(rst_bF$buf36),
    .S(vdd)
);

INVX1 _10684_ (
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_2016_)
);

NAND2X1 _10685_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .Y(_2017_)
);

OAI21X1 _10686_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_2016_),
    .C(_2017_),
    .Y(_1953_[0])
);

INVX1 _10687_ (
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_1954_)
);

NAND2X1 _10688_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1955_)
);

OAI21X1 _10689_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_1954_),
    .C(_1955_),
    .Y(_1953_[1])
);

INVX1 _10690_ (
    .A(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_1956_)
);

NAND2X1 _10691_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1957_)
);

OAI21X1 _10692_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_1956_),
    .C(_1957_),
    .Y(_1953_[2])
);

INVX1 _10693_ (
    .A(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_1958_)
);

NAND2X1 _10694_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1959_)
);

OAI21X1 _10695_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_1958_),
    .C(_1959_),
    .Y(_1953_[3])
);

INVX1 _10696_ (
    .A(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_1960_)
);

NAND2X1 _10697_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1961_)
);

OAI21X1 _10698_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_1960_),
    .C(_1961_),
    .Y(_1953_[4])
);

INVX1 _10699_ (
    .A(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_1962_)
);

NAND2X1 _10700_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1963_)
);

OAI21X1 _10701_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_1962_),
    .C(_1963_),
    .Y(_1953_[5])
);

INVX1 _10702_ (
    .A(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_1964_)
);

NAND2X1 _10703_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1965_)
);

OAI21X1 _10704_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_1964_),
    .C(_1965_),
    .Y(_1953_[6])
);

INVX1 _10705_ (
    .A(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_1966_)
);

NAND2X1 _10706_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1967_)
);

OAI21X1 _10707_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_1966_),
    .C(_1967_),
    .Y(_1953_[7])
);

INVX1 _10708_ (
    .A(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_1968_)
);

NAND2X1 _10709_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1969_)
);

OAI21X1 _10710_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_1968_),
    .C(_1969_),
    .Y(_1953_[8])
);

INVX1 _10711_ (
    .A(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_1970_)
);

NAND2X1 _10712_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1971_)
);

OAI21X1 _10713_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_1970_),
    .C(_1971_),
    .Y(_1953_[9])
);

INVX1 _10714_ (
    .A(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_1972_)
);

NAND2X1 _10715_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1973_)
);

OAI21X1 _10716_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_1972_),
    .C(_1973_),
    .Y(_1953_[10])
);

INVX1 _10717_ (
    .A(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_1974_)
);

NAND2X1 _10718_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1975_)
);

OAI21X1 _10719_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_1974_),
    .C(_1975_),
    .Y(_1953_[11])
);

INVX1 _10720_ (
    .A(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_1976_)
);

NAND2X1 _10721_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1977_)
);

OAI21X1 _10722_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_1976_),
    .C(_1977_),
    .Y(_1953_[12])
);

INVX1 _10723_ (
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_1978_)
);

NAND2X1 _10724_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1979_)
);

OAI21X1 _10725_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_1978_),
    .C(_1979_),
    .Y(_1953_[13])
);

INVX1 _10726_ (
    .A(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_1980_)
);

NAND2X1 _10727_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1981_)
);

OAI21X1 _10728_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_1980_),
    .C(_1981_),
    .Y(_1953_[14])
);

INVX1 _10729_ (
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_1982_)
);

NAND2X1 _10730_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1983_)
);

OAI21X1 _10731_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_1982_),
    .C(_1983_),
    .Y(_1953_[15])
);

INVX1 _10732_ (
    .A(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_1984_)
);

NAND2X1 _10733_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1985_)
);

OAI21X1 _10734_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_1984_),
    .C(_1985_),
    .Y(_1953_[16])
);

INVX1 _10735_ (
    .A(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_1986_)
);

NAND2X1 _10736_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1987_)
);

OAI21X1 _10737_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_1986_),
    .C(_1987_),
    .Y(_1953_[17])
);

INVX1 _10738_ (
    .A(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_1988_)
);

NAND2X1 _10739_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1989_)
);

OAI21X1 _10740_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_1988_),
    .C(_1989_),
    .Y(_1953_[18])
);

INVX1 _10741_ (
    .A(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_1990_)
);

NAND2X1 _10742_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1991_)
);

OAI21X1 _10743_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_1990_),
    .C(_1991_),
    .Y(_1953_[19])
);

INVX1 _10744_ (
    .A(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_1992_)
);

NAND2X1 _10745_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1993_)
);

OAI21X1 _10746_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_1992_),
    .C(_1993_),
    .Y(_1953_[20])
);

INVX1 _10747_ (
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_1994_)
);

NAND2X1 _10748_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1995_)
);

OAI21X1 _10749_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_1994_),
    .C(_1995_),
    .Y(_1953_[21])
);

INVX1 _10750_ (
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_1996_)
);

NAND2X1 _10751_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1997_)
);

OAI21X1 _10752_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_1996_),
    .C(_1997_),
    .Y(_1953_[22])
);

INVX1 _10753_ (
    .A(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_1998_)
);

NAND2X1 _10754_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1999_)
);

OAI21X1 _10755_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_1998_),
    .C(_1999_),
    .Y(_1953_[23])
);

INVX1 _10756_ (
    .A(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_2000_)
);

NAND2X1 _10757_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_2001_)
);

OAI21X1 _10758_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_2000_),
    .C(_2001_),
    .Y(_1953_[24])
);

INVX1 _10759_ (
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_2002_)
);

NAND2X1 _10760_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_2003_)
);

OAI21X1 _10761_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_2002_),
    .C(_2003_),
    .Y(_1953_[25])
);

INVX1 _10762_ (
    .A(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_2004_)
);

NAND2X1 _10763_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_2005_)
);

OAI21X1 _10764_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_2004_),
    .C(_2005_),
    .Y(_1953_[26])
);

INVX1 _10765_ (
    .A(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_2006_)
);

NAND2X1 _10766_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_2007_)
);

OAI21X1 _10767_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_2006_),
    .C(_2007_),
    .Y(_1953_[27])
);

INVX1 _10768_ (
    .A(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_2008_)
);

NAND2X1 _10769_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_2009_)
);

OAI21X1 _10770_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(_2008_),
    .C(_2009_),
    .Y(_1953_[28])
);

INVX1 _10771_ (
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_2010_)
);

NAND2X1 _10772_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_2011_)
);

OAI21X1 _10773_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(_2010_),
    .C(_2011_),
    .Y(_1953_[29])
);

INVX1 _10774_ (
    .A(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_2012_)
);

NAND2X1 _10775_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_2013_)
);

OAI21X1 _10776_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(_2012_),
    .C(_2013_),
    .Y(_1953_[30])
);

INVX1 _10777_ (
    .A(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_2014_)
);

NAND2X1 _10778_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_2015_)
);

OAI21X1 _10779_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(_2014_),
    .C(_2015_),
    .Y(_1953_[31])
);

DFFSR _10780_ (
    .CLK(clk_bF$buf35),
    .D(_1953_[0]),
    .Q(\datapath_1.regfile_1.regOut[31] [0]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _10781_ (
    .CLK(clk_bF$buf34),
    .D(_1953_[1]),
    .Q(\datapath_1.regfile_1.regOut[31] [1]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _10782_ (
    .CLK(clk_bF$buf33),
    .D(_1953_[2]),
    .Q(\datapath_1.regfile_1.regOut[31] [2]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _10783_ (
    .CLK(clk_bF$buf32),
    .D(_1953_[3]),
    .Q(\datapath_1.regfile_1.regOut[31] [3]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _10784_ (
    .CLK(clk_bF$buf31),
    .D(_1953_[4]),
    .Q(\datapath_1.regfile_1.regOut[31] [4]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _10785_ (
    .CLK(clk_bF$buf30),
    .D(_1953_[5]),
    .Q(\datapath_1.regfile_1.regOut[31] [5]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _10786_ (
    .CLK(clk_bF$buf29),
    .D(_1953_[6]),
    .Q(\datapath_1.regfile_1.regOut[31] [6]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _10787_ (
    .CLK(clk_bF$buf28),
    .D(_1953_[7]),
    .Q(\datapath_1.regfile_1.regOut[31] [7]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _10788_ (
    .CLK(clk_bF$buf27),
    .D(_1953_[8]),
    .Q(\datapath_1.regfile_1.regOut[31] [8]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _10789_ (
    .CLK(clk_bF$buf26),
    .D(_1953_[9]),
    .Q(\datapath_1.regfile_1.regOut[31] [9]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _10790_ (
    .CLK(clk_bF$buf25),
    .D(_1953_[10]),
    .Q(\datapath_1.regfile_1.regOut[31] [10]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _10791_ (
    .CLK(clk_bF$buf24),
    .D(_1953_[11]),
    .Q(\datapath_1.regfile_1.regOut[31] [11]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _10792_ (
    .CLK(clk_bF$buf23),
    .D(_1953_[12]),
    .Q(\datapath_1.regfile_1.regOut[31] [12]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _10793_ (
    .CLK(clk_bF$buf22),
    .D(_1953_[13]),
    .Q(\datapath_1.regfile_1.regOut[31] [13]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _10794_ (
    .CLK(clk_bF$buf21),
    .D(_1953_[14]),
    .Q(\datapath_1.regfile_1.regOut[31] [14]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _10795_ (
    .CLK(clk_bF$buf20),
    .D(_1953_[15]),
    .Q(\datapath_1.regfile_1.regOut[31] [15]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _10796_ (
    .CLK(clk_bF$buf19),
    .D(_1953_[16]),
    .Q(\datapath_1.regfile_1.regOut[31] [16]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _10797_ (
    .CLK(clk_bF$buf18),
    .D(_1953_[17]),
    .Q(\datapath_1.regfile_1.regOut[31] [17]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _10798_ (
    .CLK(clk_bF$buf17),
    .D(_1953_[18]),
    .Q(\datapath_1.regfile_1.regOut[31] [18]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _10799_ (
    .CLK(clk_bF$buf16),
    .D(_1953_[19]),
    .Q(\datapath_1.regfile_1.regOut[31] [19]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _10800_ (
    .CLK(clk_bF$buf15),
    .D(_1953_[20]),
    .Q(\datapath_1.regfile_1.regOut[31] [20]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _10801_ (
    .CLK(clk_bF$buf14),
    .D(_1953_[21]),
    .Q(\datapath_1.regfile_1.regOut[31] [21]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _10802_ (
    .CLK(clk_bF$buf13),
    .D(_1953_[22]),
    .Q(\datapath_1.regfile_1.regOut[31] [22]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _10803_ (
    .CLK(clk_bF$buf12),
    .D(_1953_[23]),
    .Q(\datapath_1.regfile_1.regOut[31] [23]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _10804_ (
    .CLK(clk_bF$buf11),
    .D(_1953_[24]),
    .Q(\datapath_1.regfile_1.regOut[31] [24]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _10805_ (
    .CLK(clk_bF$buf10),
    .D(_1953_[25]),
    .Q(\datapath_1.regfile_1.regOut[31] [25]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _10806_ (
    .CLK(clk_bF$buf9),
    .D(_1953_[26]),
    .Q(\datapath_1.regfile_1.regOut[31] [26]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _10807_ (
    .CLK(clk_bF$buf8),
    .D(_1953_[27]),
    .Q(\datapath_1.regfile_1.regOut[31] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _10808_ (
    .CLK(clk_bF$buf7),
    .D(_1953_[28]),
    .Q(\datapath_1.regfile_1.regOut[31] [28]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _10809_ (
    .CLK(clk_bF$buf6),
    .D(_1953_[29]),
    .Q(\datapath_1.regfile_1.regOut[31] [29]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _10810_ (
    .CLK(clk_bF$buf5),
    .D(_1953_[30]),
    .Q(\datapath_1.regfile_1.regOut[31] [30]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _10811_ (
    .CLK(clk_bF$buf4),
    .D(_1953_[31]),
    .Q(\datapath_1.regfile_1.regOut[31] [31]),
    .R(rst_bF$buf4),
    .S(vdd)
);

INVX1 _10812_ (
    .A(\aluControl_1.inst [4]),
    .Y(_2018_)
);

NAND2X1 _10813_ (
    .A(\aluControl_1.inst [5]),
    .B(_2018_),
    .Y(_2019_)
);

INVX1 _10814_ (
    .A(\aluControl_1.inst [3]),
    .Y(_2020_)
);

NAND2X1 _10815_ (
    .A(\aluControl_1.inst [2]),
    .B(_2020_),
    .Y(_2021_)
);

NOR2X1 _10816_ (
    .A(_2021_),
    .B(_2019_),
    .Y(_2022_)
);

INVX1 _10817_ (
    .A(ALUOp[1]),
    .Y(_2023_)
);

NOR2X1 _10818_ (
    .A(ALUOp_0_bF$buf5),
    .B(_2023_),
    .Y(_2024_)
);

OAI21X1 _10819_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .C(_2024_),
    .Y(_2025_)
);

AOI21X1 _10820_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .C(_2025_),
    .Y(_2026_)
);

AND2X2 _10821_ (
    .A(_2026_),
    .B(_2022_),
    .Y(ALUControl[0])
);

NOR2X1 _10822_ (
    .A(\aluControl_1.inst [1]),
    .B(\aluControl_1.inst [0]),
    .Y(_2027_)
);

OR2X2 _10823_ (
    .A(\aluControl_1.inst [2]),
    .B(\aluControl_1.inst [3]),
    .Y(_2028_)
);

NOR2X1 _10824_ (
    .A(_2028_),
    .B(_2019_),
    .Y(_2029_)
);

NAND2X1 _10825_ (
    .A(_2027_),
    .B(_2029_),
    .Y(_2030_)
);

INVX1 _10826_ (
    .A(\aluControl_1.inst [1]),
    .Y(_2031_)
);

NOR2X1 _10827_ (
    .A(\aluControl_1.inst [0]),
    .B(_2031_),
    .Y(_2032_)
);

OAI21X1 _10828_ (
    .A(_2029_),
    .B(_2022_),
    .C(_2032_),
    .Y(_2033_)
);

NAND3X1 _10829_ (
    .A(_2030_),
    .B(_2024_),
    .C(_2033_),
    .Y(ALUControl[1])
);

INVX1 _10830_ (
    .A(ALUOp_0_bF$buf4),
    .Y(_2034_)
);

INVX1 _10831_ (
    .A(_2019_),
    .Y(_2035_)
);

INVX1 _10832_ (
    .A(\aluControl_1.inst [2]),
    .Y(_2036_)
);

NAND2X1 _10833_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2037_)
);

NOR3X1 _10834_ (
    .A(\aluControl_1.inst [3]),
    .B(_2036_),
    .C(_2037_),
    .Y(_2038_)
);

AOI22X1 _10835_ (
    .A(_2035_),
    .B(_2038_),
    .C(_2032_),
    .D(_2029_),
    .Y(_2039_)
);

OAI21X1 _10836_ (
    .A(_2023_),
    .B(_2039_),
    .C(_2034_),
    .Y(ALUControl[2])
);

INVX1 _10837_ (
    .A(\control_1.reg_state.dout [3]),
    .Y(_2042_)
);

NOR2X1 _10838_ (
    .A(\control_1.reg_state.dout [2]),
    .B(_2042_),
    .Y(_2043_)
);

INVX2 _10839_ (
    .A(_2043_),
    .Y(_2044_)
);

INVX1 _10840_ (
    .A(\control_1.reg_state.dout [1]),
    .Y(_2045_)
);

NAND2X1 _10841_ (
    .A(\control_1.reg_state.dout [0]),
    .B(_2045_),
    .Y(_2046_)
);

NOR2X1 _10842_ (
    .A(_2046_),
    .B(_2044_),
    .Y(BranchNe)
);

INVX1 _10843_ (
    .A(\control_1.reg_state.dout [0]),
    .Y(_2047_)
);

NAND2X1 _10844_ (
    .A(_2045_),
    .B(_2047_),
    .Y(_2048_)
);

NOR2X1 _10845_ (
    .A(_2048_),
    .B(_2044_),
    .Y(Branch)
);

NAND2X1 _10846_ (
    .A(\control_1.reg_state.dout [2]),
    .B(_2042_),
    .Y(_2049_)
);

NAND2X1 _10847_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2047_),
    .Y(_2050_)
);

NOR2X1 _10848_ (
    .A(_2050_),
    .B(_2049_),
    .Y(ALUOp[1])
);

INVX1 _10849_ (
    .A(\control_1.reg_state.dout [2]),
    .Y(_2051_)
);

NOR2X1 _10850_ (
    .A(_2051_),
    .B(_2042_),
    .Y(_2052_)
);

OAI22X1 _10851_ (
    .A(_2052_),
    .B(_2050_),
    .C(\control_1.reg_state.dout [1]),
    .D(_2044_),
    .Y(ALUSrcA)
);

NOR2X1 _10852_ (
    .A(\control_1.reg_state.dout [2]),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2053_)
);

INVX2 _10853_ (
    .A(_2053_),
    .Y(_2054_)
);

NOR2X1 _10854_ (
    .A(_2048_),
    .B(_2054_),
    .Y(IRWrite)
);

INVX1 _10855_ (
    .A(_2052_),
    .Y(_2055_)
);

NOR2X1 _10856_ (
    .A(_2048_),
    .B(_2055_),
    .Y(PCSource[1])
);

NOR2X1 _10857_ (
    .A(_2053_),
    .B(_2052_),
    .Y(_2056_)
);

NOR2X1 _10858_ (
    .A(_2048_),
    .B(_2056_),
    .Y(PCWrite)
);

NAND2X1 _10859_ (
    .A(\control_1.reg_state.dout [1]),
    .B(\control_1.reg_state.dout [0]),
    .Y(_2057_)
);

NOR2X1 _10860_ (
    .A(_2057_),
    .B(_2049_),
    .Y(RegDst)
);

NOR2X1 _10861_ (
    .A(_2049_),
    .B(_2048_),
    .Y(MemToReg)
);

NAND3X1 _10862_ (
    .A(\control_1.reg_state.dout [0]),
    .B(\control_1.reg_state.dout [1]),
    .C(_2056_),
    .Y(_2058_)
);

OAI21X1 _10863_ (
    .A(_2048_),
    .B(_2049_),
    .C(_2058_),
    .Y(RegWrite)
);

NOR2X1 _10864_ (
    .A(_2049_),
    .B(_2046_),
    .Y(_0_)
);

NOR2X1 _10865_ (
    .A(_2057_),
    .B(_2054_),
    .Y(_2059_)
);

OR2X2 _10866_ (
    .A(_2059_),
    .B(_0_),
    .Y(IorD)
);

NOR2X1 _10867_ (
    .A(\control_1.op [5]),
    .B(\control_1.op [4]),
    .Y(_2060_)
);

INVX1 _10868_ (
    .A(_2060_),
    .Y(_2061_)
);

INVX1 _10869_ (
    .A(\control_1.op [1]),
    .Y(_2062_)
);

INVX1 _10870_ (
    .A(\control_1.op [3]),
    .Y(_2063_)
);

NAND3X1 _10871_ (
    .A(\control_1.op [2]),
    .B(_2062_),
    .C(_2063_),
    .Y(_2064_)
);

NOR2X1 _10872_ (
    .A(_2064_),
    .B(_2061_),
    .Y(_2065_)
);

NOR2X1 _10873_ (
    .A(_2046_),
    .B(_2054_),
    .Y(_2066_)
);

NAND3X1 _10874_ (
    .A(\control_1.op [0]),
    .B(_2066_),
    .C(_2065_),
    .Y(_2067_)
);

INVX1 _10875_ (
    .A(\control_1.op [2]),
    .Y(_2068_)
);

NOR2X1 _10876_ (
    .A(_2050_),
    .B(_2054_),
    .Y(_2069_)
);

INVX1 _10877_ (
    .A(\control_1.op [4]),
    .Y(_2070_)
);

NAND2X1 _10878_ (
    .A(\control_1.op [5]),
    .B(_2070_),
    .Y(_2071_)
);

NAND2X1 _10879_ (
    .A(\control_1.op [0]),
    .B(\control_1.op [1]),
    .Y(_2072_)
);

NOR2X1 _10880_ (
    .A(_2072_),
    .B(_2071_),
    .Y(_2073_)
);

NAND3X1 _10881_ (
    .A(_2068_),
    .B(_2073_),
    .C(_2069_),
    .Y(_2074_)
);

INVX1 _10882_ (
    .A(_2050_),
    .Y(_2075_)
);

AOI21X1 _10883_ (
    .A(_2056_),
    .B(_2075_),
    .C(IRWrite_bF$buf7),
    .Y(_2076_)
);

NAND3X1 _10884_ (
    .A(_2074_),
    .B(_2067_),
    .C(_2076_),
    .Y(\control_1.next [0])
);

NAND2X1 _10885_ (
    .A(_2075_),
    .B(_2056_),
    .Y(_2077_)
);

INVX1 _10886_ (
    .A(\control_1.op [0]),
    .Y(_2078_)
);

NAND3X1 _10887_ (
    .A(_2062_),
    .B(_2078_),
    .C(_2060_),
    .Y(_2079_)
);

OAI21X1 _10888_ (
    .A(_2071_),
    .B(_2072_),
    .C(_2079_),
    .Y(_2080_)
);

NAND3X1 _10889_ (
    .A(_2068_),
    .B(_2066_),
    .C(_2080_),
    .Y(_2081_)
);

INVX1 _10890_ (
    .A(_2071_),
    .Y(_2082_)
);

NOR2X1 _10891_ (
    .A(\control_1.op [3]),
    .B(\control_1.op [2]),
    .Y(_2083_)
);

INVX1 _10892_ (
    .A(_2083_),
    .Y(_2084_)
);

NOR2X1 _10893_ (
    .A(_2072_),
    .B(_2084_),
    .Y(_2085_)
);

NAND3X1 _10894_ (
    .A(_2082_),
    .B(_2085_),
    .C(_2069_),
    .Y(_2086_)
);

NAND3X1 _10895_ (
    .A(_2077_),
    .B(_2086_),
    .C(_2081_),
    .Y(\control_1.next [1])
);

NAND2X1 _10896_ (
    .A(\control_1.op [3]),
    .B(_2068_),
    .Y(_2087_)
);

NOR2X1 _10897_ (
    .A(_2072_),
    .B(_2087_),
    .Y(_2088_)
);

NAND3X1 _10898_ (
    .A(_2082_),
    .B(_2088_),
    .C(_2069_),
    .Y(_2089_)
);

NAND2X1 _10899_ (
    .A(_2060_),
    .B(_2083_),
    .Y(_2090_)
);

INVX1 _10900_ (
    .A(_2090_),
    .Y(_2091_)
);

NAND3X1 _10901_ (
    .A(_2078_),
    .B(_2091_),
    .C(_2066_),
    .Y(_2092_)
);

NOR2X1 _10902_ (
    .A(ALUOp[1]),
    .B(_2059_),
    .Y(_2093_)
);

NAND3X1 _10903_ (
    .A(_2089_),
    .B(_2093_),
    .C(_2092_),
    .Y(\control_1.next [2])
);

NAND2X1 _10904_ (
    .A(_2043_),
    .B(_2075_),
    .Y(_2094_)
);

NOR2X1 _10905_ (
    .A(_2087_),
    .B(_2079_),
    .Y(_2095_)
);

NAND2X1 _10906_ (
    .A(\control_1.op [1]),
    .B(_2078_),
    .Y(_2096_)
);

OAI22X1 _10907_ (
    .A(_2064_),
    .B(_2061_),
    .C(_2096_),
    .D(_2090_),
    .Y(_2040_)
);

OAI21X1 _10908_ (
    .A(_2095_),
    .B(_2040_),
    .C(_2066_),
    .Y(_2041_)
);

NAND2X1 _10909_ (
    .A(_2094_),
    .B(_2041_),
    .Y(\control_1.next [3])
);

NOR2X1 _10910_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2044_),
    .Y(ALUOp[0])
);

NOR2X1 _10911_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2054_),
    .Y(ALUSrcB[0])
);

OAI22X1 _10912_ (
    .A(\control_1.reg_state.dout [2]),
    .B(_2050_),
    .C(_2046_),
    .D(_2054_),
    .Y(ALUSrcB[1])
);

INVX1 _10913_ (
    .A(\control_1.reg_state.dout [0]),
    .Y(_2098_)
);

NAND2X1 _10914_ (
    .A(\control_1.next [0]),
    .B(vdd),
    .Y(_2099_)
);

OAI21X1 _10915_ (
    .A(vdd),
    .B(_2098_),
    .C(_2099_),
    .Y(_2097_[0])
);

INVX1 _10916_ (
    .A(\control_1.reg_state.dout [1]),
    .Y(_2100_)
);

NAND2X1 _10917_ (
    .A(vdd),
    .B(\control_1.next [1]),
    .Y(_2101_)
);

OAI21X1 _10918_ (
    .A(vdd),
    .B(_2100_),
    .C(_2101_),
    .Y(_2097_[1])
);

INVX1 _10919_ (
    .A(\control_1.reg_state.dout [2]),
    .Y(_2102_)
);

NAND2X1 _10920_ (
    .A(vdd),
    .B(\control_1.next [2]),
    .Y(_2103_)
);

OAI21X1 _10921_ (
    .A(vdd),
    .B(_2102_),
    .C(_2103_),
    .Y(_2097_[2])
);

INVX1 _10922_ (
    .A(\control_1.reg_state.dout [3]),
    .Y(_2104_)
);

NAND2X1 _10923_ (
    .A(vdd),
    .B(\control_1.next [3]),
    .Y(_2105_)
);

OAI21X1 _10924_ (
    .A(vdd),
    .B(_2104_),
    .C(_2105_),
    .Y(_2097_[3])
);

DFFSR _10925_ (
    .CLK(clk_bF$buf3),
    .D(_2097_[0]),
    .Q(\control_1.reg_state.dout [0]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _10926_ (
    .CLK(clk_bF$buf2),
    .D(_2097_[1]),
    .Q(\control_1.reg_state.dout [1]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _10927_ (
    .CLK(clk_bF$buf1),
    .D(_2097_[2]),
    .Q(\control_1.reg_state.dout [2]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _10928_ (
    .CLK(clk_bF$buf0),
    .D(_2097_[3]),
    .Q(\control_1.reg_state.dout [3]),
    .R(rst_bF$buf0),
    .S(vdd)
);

NOR2X1 _10929_ (
    .A(\datapath_1.alu_1.ALUInB [31]),
    .B(\datapath_1.alu_1.ALUInA [31]),
    .Y(_2106_)
);

NAND2X1 _10930_ (
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2107_)
);

INVX1 _10931_ (
    .A(_2107_),
    .Y(_2108_)
);

NOR2X1 _10932_ (
    .A(_2106_),
    .B(_2108_),
    .Y(_2109_)
);

INVX1 _10933_ (
    .A(\datapath_1.alu_1.ALUInA [30]),
    .Y(_2110_)
);

NOR2X1 _10934_ (
    .A(\datapath_1.alu_1.ALUInB [30]),
    .B(_2110_),
    .Y(_2111_)
);

INVX1 _10935_ (
    .A(_2111_),
    .Y(_2112_)
);

INVX1 _10936_ (
    .A(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2113_)
);

NOR2X1 _10937_ (
    .A(_2113_),
    .B(_2110_),
    .Y(_2114_)
);

NOR2X1 _10938_ (
    .A(\datapath_1.alu_1.ALUInB [30]),
    .B(\datapath_1.alu_1.ALUInA [30]),
    .Y(_2115_)
);

INVX1 _10939_ (
    .A(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2116_)
);

INVX1 _10940_ (
    .A(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2117_)
);

NOR2X1 _10941_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(_2117_),
    .Y(_2118_)
);

AND2X2 _10942_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2119_)
);

NOR2X1 _10943_ (
    .A(\datapath_1.alu_1.ALUInA [3]),
    .B(\datapath_1.alu_1.ALUInB [3]),
    .Y(_2120_)
);

OAI21X1 _10944_ (
    .A(_2119_),
    .B(_2120_),
    .C(_2118_),
    .Y(_2121_)
);

OAI21X1 _10945_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2116_),
    .C(_2121_),
    .Y(_2122_)
);

INVX1 _10946_ (
    .A(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2123_)
);

NOR2X1 _10947_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(_2123_),
    .Y(_2124_)
);

INVX1 _10948_ (
    .A(_2124_),
    .Y(_2125_)
);

INVX2 _10949_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .Y(_2126_)
);

AND2X2 _10950_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2127_)
);

NOR2X1 _10951_ (
    .A(\datapath_1.alu_1.ALUInA [1]),
    .B(\datapath_1.alu_1.ALUInB [1]),
    .Y(_2128_)
);

OAI22X1 _10952_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .B(_2126_),
    .C(_2128_),
    .D(_2127_),
    .Y(_2129_)
);

AND2X2 _10953_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2130_)
);

NOR2X1 _10954_ (
    .A(\datapath_1.alu_1.ALUInA [2]),
    .B(\datapath_1.alu_1.ALUInB [2]),
    .Y(_2131_)
);

OAI22X1 _10955_ (
    .A(_2131_),
    .B(_2130_),
    .C(_2120_),
    .D(_2119_),
    .Y(_2132_)
);

AOI21X1 _10956_ (
    .A(_2125_),
    .B(_2129_),
    .C(_2132_),
    .Y(_2133_)
);

AND2X2 _10957_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2134_)
);

NOR2X1 _10958_ (
    .A(\datapath_1.alu_1.ALUInA [7]),
    .B(\datapath_1.alu_1.ALUInB [7]),
    .Y(_2135_)
);

AND2X2 _10959_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2136_)
);

NOR2X1 _10960_ (
    .A(\datapath_1.alu_1.ALUInA [6]),
    .B(\datapath_1.alu_1.ALUInB [6]),
    .Y(_2137_)
);

OAI22X1 _10961_ (
    .A(_2135_),
    .B(_2134_),
    .C(_2137_),
    .D(_2136_),
    .Y(_2138_)
);

AND2X2 _10962_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2139_)
);

NOR2X1 _10963_ (
    .A(\datapath_1.alu_1.ALUInA [5]),
    .B(\datapath_1.alu_1.ALUInB [5]),
    .Y(_2140_)
);

AND2X2 _10964_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2141_)
);

NOR2X1 _10965_ (
    .A(\datapath_1.alu_1.ALUInA [4]),
    .B(\datapath_1.alu_1.ALUInB [4]),
    .Y(_2142_)
);

OAI22X1 _10966_ (
    .A(_2140_),
    .B(_2139_),
    .C(_2142_),
    .D(_2141_),
    .Y(_2143_)
);

NOR2X1 _10967_ (
    .A(_2143_),
    .B(_2138_),
    .Y(_2144_)
);

OAI21X1 _10968_ (
    .A(_2122_),
    .B(_2133_),
    .C(_2144_),
    .Y(_2145_)
);

INVX1 _10969_ (
    .A(_2138_),
    .Y(_2146_)
);

NOR2X1 _10970_ (
    .A(_2140_),
    .B(_2139_),
    .Y(_2147_)
);

INVX1 _10971_ (
    .A(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2148_)
);

NOR2X1 _10972_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(_2148_),
    .Y(_2149_)
);

INVX1 _10973_ (
    .A(_2149_),
    .Y(_2150_)
);

INVX1 _10974_ (
    .A(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2151_)
);

OR2X2 _10975_ (
    .A(_2151_),
    .B(\datapath_1.alu_1.ALUInB [4]),
    .Y(_2152_)
);

OAI21X1 _10976_ (
    .A(_2152_),
    .B(_2147_),
    .C(_2150_),
    .Y(_2153_)
);

INVX1 _10977_ (
    .A(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2154_)
);

INVX1 _10978_ (
    .A(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2155_)
);

NOR2X1 _10979_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(_2155_),
    .Y(_2156_)
);

OAI21X1 _10980_ (
    .A(_2134_),
    .B(_2135_),
    .C(_2156_),
    .Y(_2157_)
);

OAI21X1 _10981_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2154_),
    .C(_2157_),
    .Y(_2158_)
);

AOI21X1 _10982_ (
    .A(_2153_),
    .B(_2146_),
    .C(_2158_),
    .Y(_2159_)
);

NAND2X1 _10983_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2160_)
);

INVX1 _10984_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .Y(_2161_)
);

INVX1 _10985_ (
    .A(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2162_)
);

NAND2X1 _10986_ (
    .A(_2161_),
    .B(_2162_),
    .Y(_2163_)
);

NAND2X1 _10987_ (
    .A(_2160_),
    .B(_2163_),
    .Y(_2164_)
);

AND2X2 _10988_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2165_)
);

NOR2X1 _10989_ (
    .A(\datapath_1.alu_1.ALUInA [14]),
    .B(\datapath_1.alu_1.ALUInB [14]),
    .Y(_2166_)
);

OAI21X1 _10990_ (
    .A(_2165_),
    .B(_2166_),
    .C(_2164_),
    .Y(_2167_)
);

NAND2X1 _10991_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2168_)
);

OR2X2 _10992_ (
    .A(\datapath_1.alu_1.ALUInA [13]),
    .B(\datapath_1.alu_1.ALUInB [13]),
    .Y(_2169_)
);

NAND2X1 _10993_ (
    .A(_2168_),
    .B(_2169_),
    .Y(_2170_)
);

AND2X2 _10994_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2171_)
);

NOR2X1 _10995_ (
    .A(\datapath_1.alu_1.ALUInA [12]),
    .B(\datapath_1.alu_1.ALUInB [12]),
    .Y(_2172_)
);

OAI21X1 _10996_ (
    .A(_2171_),
    .B(_2172_),
    .C(_2170_),
    .Y(_2173_)
);

NOR2X1 _10997_ (
    .A(_2173_),
    .B(_2167_),
    .Y(_2174_)
);

NAND2X1 _10998_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2175_)
);

OR2X2 _10999_ (
    .A(\datapath_1.alu_1.ALUInA [9]),
    .B(\datapath_1.alu_1.ALUInB [9]),
    .Y(_2176_)
);

NAND2X1 _11000_ (
    .A(_2175_),
    .B(_2176_),
    .Y(_2177_)
);

AND2X2 _11001_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2178_)
);

NOR2X1 _11002_ (
    .A(\datapath_1.alu_1.ALUInA [8]),
    .B(\datapath_1.alu_1.ALUInB [8]),
    .Y(_2179_)
);

OAI21X1 _11003_ (
    .A(_2178_),
    .B(_2179_),
    .C(_2177_),
    .Y(_2180_)
);

NAND2X1 _11004_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2181_)
);

OR2X2 _11005_ (
    .A(\datapath_1.alu_1.ALUInA [11]),
    .B(\datapath_1.alu_1.ALUInB [11]),
    .Y(_2182_)
);

NAND2X1 _11006_ (
    .A(_2181_),
    .B(_2182_),
    .Y(_2183_)
);

AND2X2 _11007_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2184_)
);

NOR2X1 _11008_ (
    .A(\datapath_1.alu_1.ALUInA [10]),
    .B(\datapath_1.alu_1.ALUInB [10]),
    .Y(_2185_)
);

OAI21X1 _11009_ (
    .A(_2184_),
    .B(_2185_),
    .C(_2183_),
    .Y(_2186_)
);

NOR2X1 _11010_ (
    .A(_2180_),
    .B(_2186_),
    .Y(_2187_)
);

NAND2X1 _11011_ (
    .A(_2187_),
    .B(_2174_),
    .Y(_2188_)
);

AOI21X1 _11012_ (
    .A(_2145_),
    .B(_2159_),
    .C(_2188_),
    .Y(_2189_)
);

AND2X2 _11013_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2190_)
);

NOR2X1 _11014_ (
    .A(\datapath_1.alu_1.ALUInA [15]),
    .B(\datapath_1.alu_1.ALUInB [15]),
    .Y(_2191_)
);

NOR2X1 _11015_ (
    .A(_2191_),
    .B(_2190_),
    .Y(_2192_)
);

NOR2X1 _11016_ (
    .A(_2166_),
    .B(_2165_),
    .Y(_2193_)
);

NOR2X1 _11017_ (
    .A(_2193_),
    .B(_2192_),
    .Y(_2194_)
);

NAND2X1 _11018_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2195_)
);

INVX1 _11019_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .Y(_2196_)
);

INVX1 _11020_ (
    .A(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2197_)
);

NAND2X1 _11021_ (
    .A(_2196_),
    .B(_2197_),
    .Y(_2198_)
);

NAND2X1 _11022_ (
    .A(_2195_),
    .B(_2198_),
    .Y(_2199_)
);

NAND3X1 _11023_ (
    .A(_2170_),
    .B(_2199_),
    .C(_2194_),
    .Y(_2200_)
);

AND2X2 _11024_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2201_)
);

NOR2X1 _11025_ (
    .A(\datapath_1.alu_1.ALUInA [11]),
    .B(\datapath_1.alu_1.ALUInB [11]),
    .Y(_2202_)
);

NOR2X1 _11026_ (
    .A(_2202_),
    .B(_2201_),
    .Y(_2203_)
);

NOR2X1 _11027_ (
    .A(_2185_),
    .B(_2184_),
    .Y(_2204_)
);

NOR2X1 _11028_ (
    .A(_2204_),
    .B(_2203_),
    .Y(_2205_)
);

AND2X2 _11029_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2206_)
);

NOR2X1 _11030_ (
    .A(\datapath_1.alu_1.ALUInA [9]),
    .B(\datapath_1.alu_1.ALUInB [9]),
    .Y(_2207_)
);

NOR2X1 _11031_ (
    .A(_2207_),
    .B(_2206_),
    .Y(_2208_)
);

INVX1 _11032_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .Y(_2209_)
);

NAND2X1 _11033_ (
    .A(\datapath_1.alu_1.ALUInA [9]),
    .B(_2209_),
    .Y(_2210_)
);

INVX1 _11034_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .Y(_2211_)
);

NAND2X1 _11035_ (
    .A(\datapath_1.alu_1.ALUInA [8]),
    .B(_2211_),
    .Y(_2212_)
);

OAI21X1 _11036_ (
    .A(_2212_),
    .B(_2208_),
    .C(_2210_),
    .Y(_2213_)
);

INVX1 _11037_ (
    .A(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2214_)
);

INVX1 _11038_ (
    .A(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2215_)
);

NOR2X1 _11039_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2215_),
    .Y(_2216_)
);

OAI21X1 _11040_ (
    .A(_2201_),
    .B(_2202_),
    .C(_2216_),
    .Y(_2217_)
);

OAI21X1 _11041_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(_2214_),
    .C(_2217_),
    .Y(_2218_)
);

AOI21X1 _11042_ (
    .A(_2213_),
    .B(_2205_),
    .C(_2218_),
    .Y(_2219_)
);

AND2X2 _11043_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2220_)
);

NOR2X1 _11044_ (
    .A(\datapath_1.alu_1.ALUInA [13]),
    .B(\datapath_1.alu_1.ALUInB [13]),
    .Y(_2221_)
);

NOR2X1 _11045_ (
    .A(_2221_),
    .B(_2220_),
    .Y(_2222_)
);

INVX1 _11046_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .Y(_2223_)
);

NAND2X1 _11047_ (
    .A(\datapath_1.alu_1.ALUInA [13]),
    .B(_2223_),
    .Y(_2224_)
);

NAND2X1 _11048_ (
    .A(\datapath_1.alu_1.ALUInA [12]),
    .B(_2196_),
    .Y(_2225_)
);

OAI21X1 _11049_ (
    .A(_2225_),
    .B(_2222_),
    .C(_2224_),
    .Y(_2226_)
);

INVX1 _11050_ (
    .A(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2227_)
);

NOR2X1 _11051_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(_2227_),
    .Y(_2228_)
);

OAI21X1 _11052_ (
    .A(_2190_),
    .B(_2191_),
    .C(_2228_),
    .Y(_2229_)
);

OAI21X1 _11053_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(_2162_),
    .C(_2229_),
    .Y(_2230_)
);

AOI21X1 _11054_ (
    .A(_2226_),
    .B(_2194_),
    .C(_2230_),
    .Y(_2231_)
);

OAI21X1 _11055_ (
    .A(_2200_),
    .B(_2219_),
    .C(_2231_),
    .Y(_2232_)
);

NOR2X1 _11056_ (
    .A(\datapath_1.alu_1.ALUInB [22]),
    .B(\datapath_1.alu_1.ALUInA [22]),
    .Y(_2233_)
);

NAND2X1 _11057_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2234_)
);

INVX2 _11058_ (
    .A(_2234_),
    .Y(_2235_)
);

NOR2X1 _11059_ (
    .A(_2233_),
    .B(_2235_),
    .Y(_2236_)
);

INVX1 _11060_ (
    .A(\datapath_1.alu_1.ALUInA [23]),
    .Y(_2237_)
);

INVX1 _11061_ (
    .A(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2238_)
);

NOR2X1 _11062_ (
    .A(_2238_),
    .B(_2237_),
    .Y(_2239_)
);

NOR2X1 _11063_ (
    .A(\datapath_1.alu_1.ALUInB [23]),
    .B(\datapath_1.alu_1.ALUInA [23]),
    .Y(_2240_)
);

NOR2X1 _11064_ (
    .A(_2240_),
    .B(_2239_),
    .Y(_2241_)
);

NOR2X1 _11065_ (
    .A(_2236_),
    .B(_2241_),
    .Y(_2242_)
);

INVX1 _11066_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .Y(_2243_)
);

INVX1 _11067_ (
    .A(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2244_)
);

NOR2X1 _11068_ (
    .A(_2244_),
    .B(_2243_),
    .Y(_2245_)
);

NOR2X1 _11069_ (
    .A(\datapath_1.alu_1.ALUInB [21]),
    .B(\datapath_1.alu_1.ALUInA [21]),
    .Y(_2246_)
);

NOR2X1 _11070_ (
    .A(_2246_),
    .B(_2245_),
    .Y(_2247_)
);

NAND2X1 _11071_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .B(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2248_)
);

INVX1 _11072_ (
    .A(_2248_),
    .Y(_2249_)
);

NOR2X1 _11073_ (
    .A(\datapath_1.alu_1.ALUInB [20]),
    .B(\datapath_1.alu_1.ALUInA [20]),
    .Y(_2250_)
);

NOR2X1 _11074_ (
    .A(_2250_),
    .B(_2249_),
    .Y(_2251_)
);

NOR2X1 _11075_ (
    .A(_2251_),
    .B(_2247_),
    .Y(_2252_)
);

NAND2X1 _11076_ (
    .A(_2242_),
    .B(_2252_),
    .Y(_2253_)
);

NOR2X1 _11077_ (
    .A(\datapath_1.alu_1.ALUInB [18]),
    .B(\datapath_1.alu_1.ALUInA [18]),
    .Y(_2254_)
);

NAND2X1 _11078_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2255_)
);

INVX1 _11079_ (
    .A(_2255_),
    .Y(_2256_)
);

NOR2X1 _11080_ (
    .A(_2254_),
    .B(_2256_),
    .Y(_2257_)
);

INVX1 _11081_ (
    .A(\datapath_1.alu_1.ALUInA [19]),
    .Y(_2258_)
);

INVX1 _11082_ (
    .A(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2259_)
);

NOR2X1 _11083_ (
    .A(_2259_),
    .B(_2258_),
    .Y(_2260_)
);

NOR2X1 _11084_ (
    .A(\datapath_1.alu_1.ALUInB [19]),
    .B(\datapath_1.alu_1.ALUInA [19]),
    .Y(_2261_)
);

NOR2X1 _11085_ (
    .A(_2261_),
    .B(_2260_),
    .Y(_2262_)
);

NOR2X1 _11086_ (
    .A(_2257_),
    .B(_2262_),
    .Y(_2263_)
);

INVX1 _11087_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .Y(_2264_)
);

INVX1 _11088_ (
    .A(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2265_)
);

NOR2X1 _11089_ (
    .A(_2265_),
    .B(_2264_),
    .Y(_2266_)
);

NOR2X1 _11090_ (
    .A(\datapath_1.alu_1.ALUInB [17]),
    .B(\datapath_1.alu_1.ALUInA [17]),
    .Y(_2267_)
);

NAND2X1 _11091_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2268_)
);

INVX2 _11092_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .Y(_2269_)
);

INVX1 _11093_ (
    .A(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2270_)
);

NAND2X1 _11094_ (
    .A(_2269_),
    .B(_2270_),
    .Y(_2271_)
);

NAND2X1 _11095_ (
    .A(_2268_),
    .B(_2271_),
    .Y(_2272_)
);

OAI21X1 _11096_ (
    .A(_2266_),
    .B(_2267_),
    .C(_2272_),
    .Y(_2273_)
);

INVX1 _11097_ (
    .A(_2273_),
    .Y(_2274_)
);

NAND2X1 _11098_ (
    .A(_2263_),
    .B(_2274_),
    .Y(_2275_)
);

NOR2X1 _11099_ (
    .A(_2253_),
    .B(_2275_),
    .Y(_2276_)
);

OAI21X1 _11100_ (
    .A(_2232_),
    .B(_2189_),
    .C(_2276_),
    .Y(_2277_)
);

NOR2X1 _11101_ (
    .A(\datapath_1.alu_1.ALUInB [16]),
    .B(_2269_),
    .Y(_2278_)
);

OAI21X1 _11102_ (
    .A(_2267_),
    .B(_2266_),
    .C(_2278_),
    .Y(_2279_)
);

OAI21X1 _11103_ (
    .A(_2264_),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .C(_2279_),
    .Y(_2280_)
);

INVX1 _11104_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .Y(_2281_)
);

NOR2X1 _11105_ (
    .A(\datapath_1.alu_1.ALUInB [18]),
    .B(_2281_),
    .Y(_2282_)
);

OAI21X1 _11106_ (
    .A(_2261_),
    .B(_2260_),
    .C(_2282_),
    .Y(_2283_)
);

OAI21X1 _11107_ (
    .A(_2258_),
    .B(\datapath_1.alu_1.ALUInB [19]),
    .C(_2283_),
    .Y(_2284_)
);

AOI21X1 _11108_ (
    .A(_2280_),
    .B(_2263_),
    .C(_2284_),
    .Y(_2285_)
);

INVX1 _11109_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .Y(_2286_)
);

NOR2X1 _11110_ (
    .A(\datapath_1.alu_1.ALUInB [20]),
    .B(_2286_),
    .Y(_2287_)
);

OAI21X1 _11111_ (
    .A(_2246_),
    .B(_2245_),
    .C(_2287_),
    .Y(_2288_)
);

OAI21X1 _11112_ (
    .A(_2243_),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .C(_2288_),
    .Y(_2289_)
);

INVX1 _11113_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .Y(_2290_)
);

NOR2X1 _11114_ (
    .A(\datapath_1.alu_1.ALUInB [22]),
    .B(_2290_),
    .Y(_2291_)
);

OAI21X1 _11115_ (
    .A(_2240_),
    .B(_2239_),
    .C(_2291_),
    .Y(_2292_)
);

OAI21X1 _11116_ (
    .A(_2237_),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .C(_2292_),
    .Y(_2293_)
);

AOI21X1 _11117_ (
    .A(_2289_),
    .B(_2242_),
    .C(_2293_),
    .Y(_2294_)
);

OAI21X1 _11118_ (
    .A(_2253_),
    .B(_2285_),
    .C(_2294_),
    .Y(_2295_)
);

INVX1 _11119_ (
    .A(_2295_),
    .Y(_2296_)
);

NOR2X1 _11120_ (
    .A(\datapath_1.alu_1.ALUInB [26]),
    .B(\datapath_1.alu_1.ALUInA [26]),
    .Y(_2297_)
);

INVX1 _11121_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .Y(_2298_)
);

INVX1 _11122_ (
    .A(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2299_)
);

NOR2X1 _11123_ (
    .A(_2299_),
    .B(_2298_),
    .Y(_2300_)
);

NOR2X1 _11124_ (
    .A(_2297_),
    .B(_2300_),
    .Y(_2301_)
);

INVX1 _11125_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .Y(_2302_)
);

INVX1 _11126_ (
    .A(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2303_)
);

NOR2X1 _11127_ (
    .A(_2303_),
    .B(_2302_),
    .Y(_2304_)
);

NOR2X1 _11128_ (
    .A(\datapath_1.alu_1.ALUInB [27]),
    .B(\datapath_1.alu_1.ALUInA [27]),
    .Y(_2305_)
);

NOR2X1 _11129_ (
    .A(_2305_),
    .B(_2304_),
    .Y(_2306_)
);

NOR2X1 _11130_ (
    .A(_2306_),
    .B(_2301_),
    .Y(_2307_)
);

NAND2X1 _11131_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2308_)
);

NOR2X1 _11132_ (
    .A(\datapath_1.alu_1.ALUInB [25]),
    .B(\datapath_1.alu_1.ALUInA [25]),
    .Y(_2309_)
);

INVX1 _11133_ (
    .A(_2309_),
    .Y(_2310_)
);

NAND2X1 _11134_ (
    .A(_2308_),
    .B(_2310_),
    .Y(_2311_)
);

INVX1 _11135_ (
    .A(\datapath_1.alu_1.ALUInA [24]),
    .Y(_2312_)
);

INVX1 _11136_ (
    .A(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2313_)
);

NOR2X1 _11137_ (
    .A(_2313_),
    .B(_2312_),
    .Y(_2314_)
);

NOR2X1 _11138_ (
    .A(\datapath_1.alu_1.ALUInB [24]),
    .B(\datapath_1.alu_1.ALUInA [24]),
    .Y(_2315_)
);

OAI21X1 _11139_ (
    .A(_2314_),
    .B(_2315_),
    .C(_2311_),
    .Y(_2316_)
);

INVX1 _11140_ (
    .A(_2316_),
    .Y(_2317_)
);

NAND2X1 _11141_ (
    .A(_2307_),
    .B(_2317_),
    .Y(_2318_)
);

AOI21X1 _11142_ (
    .A(_2277_),
    .B(_2296_),
    .C(_2318_),
    .Y(_2319_)
);

INVX1 _11143_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .Y(_2320_)
);

INVX1 _11144_ (
    .A(_2308_),
    .Y(_2321_)
);

NOR2X1 _11145_ (
    .A(\datapath_1.alu_1.ALUInB [24]),
    .B(_2312_),
    .Y(_2322_)
);

OAI21X1 _11146_ (
    .A(_2309_),
    .B(_2321_),
    .C(_2322_),
    .Y(_2323_)
);

OAI21X1 _11147_ (
    .A(_2320_),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .C(_2323_),
    .Y(_2324_)
);

AND2X2 _11148_ (
    .A(_2307_),
    .B(_2324_),
    .Y(_2325_)
);

NOR2X1 _11149_ (
    .A(\datapath_1.alu_1.ALUInB [26]),
    .B(_2298_),
    .Y(_2326_)
);

OAI21X1 _11150_ (
    .A(_2305_),
    .B(_2304_),
    .C(_2326_),
    .Y(_2327_)
);

OAI21X1 _11151_ (
    .A(_2302_),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .C(_2327_),
    .Y(_2328_)
);

NOR2X1 _11152_ (
    .A(_2328_),
    .B(_2325_),
    .Y(_2329_)
);

INVX1 _11153_ (
    .A(_2329_),
    .Y(_2330_)
);

INVX1 _11154_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .Y(_2331_)
);

INVX1 _11155_ (
    .A(\datapath_1.alu_1.ALUInB [29]),
    .Y(_2332_)
);

NOR2X1 _11156_ (
    .A(_2332_),
    .B(_2331_),
    .Y(_2333_)
);

NOR2X1 _11157_ (
    .A(\datapath_1.alu_1.ALUInB [29]),
    .B(\datapath_1.alu_1.ALUInA [29]),
    .Y(_2334_)
);

AND2X2 _11158_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2335_)
);

NOR2X1 _11159_ (
    .A(\datapath_1.alu_1.ALUInB [28]),
    .B(\datapath_1.alu_1.ALUInA [28]),
    .Y(_2336_)
);

NOR2X1 _11160_ (
    .A(_2336_),
    .B(_2335_),
    .Y(_2337_)
);

INVX2 _11161_ (
    .A(_2337_),
    .Y(_2338_)
);

OAI21X1 _11162_ (
    .A(_2333_),
    .B(_2334_),
    .C(_2338_),
    .Y(_2339_)
);

INVX1 _11163_ (
    .A(_2339_),
    .Y(_2340_)
);

OAI21X1 _11164_ (
    .A(_2330_),
    .B(_2319_),
    .C(_2340_),
    .Y(_2341_)
);

INVX1 _11165_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .Y(_2342_)
);

NOR2X1 _11166_ (
    .A(\datapath_1.alu_1.ALUInB [28]),
    .B(_2342_),
    .Y(_2343_)
);

OAI21X1 _11167_ (
    .A(_2334_),
    .B(_2333_),
    .C(_2343_),
    .Y(_2344_)
);

NAND2X1 _11168_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(_2332_),
    .Y(_2345_)
);

NAND3X1 _11169_ (
    .A(_2344_),
    .B(_2345_),
    .C(_2341_),
    .Y(_2346_)
);

OAI21X1 _11170_ (
    .A(_2114_),
    .B(_2115_),
    .C(_2346_),
    .Y(_2347_)
);

NAND3X1 _11171_ (
    .A(_2112_),
    .B(_2109_),
    .C(_2347_),
    .Y(_2348_)
);

INVX1 _11172_ (
    .A(ALUControl[1]),
    .Y(_2349_)
);

NOR2X1 _11173_ (
    .A(ALUControl[0]),
    .B(_2349_),
    .Y(_2350_)
);

INVX1 _11174_ (
    .A(ALUControl[2]),
    .Y(_2351_)
);

NOR2X1 _11175_ (
    .A(gnd),
    .B(_2351_),
    .Y(_2352_)
);

NAND2X1 _11176_ (
    .A(_2350_),
    .B(_2352_),
    .Y(_2353_)
);

INVX8 _11177_ (
    .A(_2353_),
    .Y(_2354_)
);

INVX1 _11178_ (
    .A(_2109_),
    .Y(_2355_)
);

NOR2X1 _11179_ (
    .A(_2115_),
    .B(_2114_),
    .Y(_2356_)
);

INVX2 _11180_ (
    .A(_2356_),
    .Y(_2357_)
);

AND2X2 _11181_ (
    .A(_2346_),
    .B(_2357_),
    .Y(_2358_)
);

OAI21X1 _11182_ (
    .A(_2111_),
    .B(_2358_),
    .C(_2355_),
    .Y(_2359_)
);

NAND3X1 _11183_ (
    .A(_2354__bF$buf3),
    .B(_2348_),
    .C(_2359_),
    .Y(_2360_)
);

NOR2X1 _11184_ (
    .A(ALUControl[0]),
    .B(ALUControl[1]),
    .Y(_2361_)
);

AND2X2 _11185_ (
    .A(_2352_),
    .B(_2361_),
    .Y(_2362_)
);

NAND2X1 _11186_ (
    .A(_2106_),
    .B(_2362__bF$buf3),
    .Y(_2363_)
);

NOR2X1 _11187_ (
    .A(ALUControl[2]),
    .B(gnd),
    .Y(_2364_)
);

NAND3X1 _11188_ (
    .A(ALUControl[0]),
    .B(ALUControl[1]),
    .C(_2364_),
    .Y(_2365_)
);

OAI21X1 _11189_ (
    .A(_2365__bF$buf4),
    .B(_2355_),
    .C(_2363_),
    .Y(_2366_)
);

NAND2X1 _11190_ (
    .A(_2361_),
    .B(_2364_),
    .Y(_2367_)
);

NAND3X1 _11191_ (
    .A(ALUControl[0]),
    .B(_2349_),
    .C(_2364_),
    .Y(_2368_)
);

OAI22X1 _11192_ (
    .A(_2367__bF$buf3),
    .B(_2107_),
    .C(_2106_),
    .D(_2368__bF$buf3),
    .Y(_2369_)
);

NOR2X1 _11193_ (
    .A(_2369_),
    .B(_2366_),
    .Y(_2370_)
);

INVX1 _11194_ (
    .A(_2114_),
    .Y(_2371_)
);

NOR2X1 _11195_ (
    .A(_2131_),
    .B(_2130_),
    .Y(_2372_)
);

NOR2X1 _11196_ (
    .A(_2120_),
    .B(_2119_),
    .Y(_2373_)
);

NAND2X1 _11197_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2374_)
);

NAND2X1 _11198_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2375_)
);

OAI21X1 _11199_ (
    .A(_2375_),
    .B(_2128_),
    .C(_2374_),
    .Y(_2376_)
);

NAND3X1 _11200_ (
    .A(_2372_),
    .B(_2376_),
    .C(_2373_),
    .Y(_2377_)
);

OR2X2 _11201_ (
    .A(\datapath_1.alu_1.ALUInA [3]),
    .B(\datapath_1.alu_1.ALUInB [3]),
    .Y(_2378_)
);

AOI21X1 _11202_ (
    .A(_2378_),
    .B(_2130_),
    .C(_2119_),
    .Y(_2379_)
);

NAND2X1 _11203_ (
    .A(_2379_),
    .B(_2377_),
    .Y(_2380_)
);

NOR2X1 _11204_ (
    .A(_2135_),
    .B(_2134_),
    .Y(_2381_)
);

NOR2X1 _11205_ (
    .A(_2137_),
    .B(_2136_),
    .Y(_2382_)
);

NAND2X1 _11206_ (
    .A(_2381_),
    .B(_2382_),
    .Y(_2383_)
);

NOR2X1 _11207_ (
    .A(_2142_),
    .B(_2141_),
    .Y(_2384_)
);

NAND2X1 _11208_ (
    .A(_2147_),
    .B(_2384_),
    .Y(_2385_)
);

NOR2X1 _11209_ (
    .A(_2385_),
    .B(_2383_),
    .Y(_2386_)
);

NAND2X1 _11210_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2387_)
);

NAND2X1 _11211_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2388_)
);

OAI21X1 _11212_ (
    .A(_2388_),
    .B(_2140_),
    .C(_2387_),
    .Y(_2389_)
);

INVX1 _11213_ (
    .A(_2389_),
    .Y(_2390_)
);

OR2X2 _11214_ (
    .A(\datapath_1.alu_1.ALUInA [7]),
    .B(\datapath_1.alu_1.ALUInB [7]),
    .Y(_2391_)
);

AOI21X1 _11215_ (
    .A(_2391_),
    .B(_2136_),
    .C(_2134_),
    .Y(_2392_)
);

OAI21X1 _11216_ (
    .A(_2390_),
    .B(_2383_),
    .C(_2392_),
    .Y(_2393_)
);

AOI21X1 _11217_ (
    .A(_2386_),
    .B(_2380_),
    .C(_2393_),
    .Y(_2394_)
);

NAND2X1 _11218_ (
    .A(_2192_),
    .B(_2193_),
    .Y(_2395_)
);

NOR2X1 _11219_ (
    .A(_2172_),
    .B(_2171_),
    .Y(_2396_)
);

NAND2X1 _11220_ (
    .A(_2222_),
    .B(_2396_),
    .Y(_2397_)
);

NOR2X1 _11221_ (
    .A(_2397_),
    .B(_2395_),
    .Y(_2398_)
);

NAND2X1 _11222_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2399_)
);

OR2X2 _11223_ (
    .A(\datapath_1.alu_1.ALUInA [8]),
    .B(\datapath_1.alu_1.ALUInB [8]),
    .Y(_2400_)
);

NAND2X1 _11224_ (
    .A(_2399_),
    .B(_2400_),
    .Y(_2401_)
);

NOR2X1 _11225_ (
    .A(_2177_),
    .B(_2401_),
    .Y(_2402_)
);

NAND2X1 _11226_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2403_)
);

INVX1 _11227_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .Y(_2404_)
);

NAND2X1 _11228_ (
    .A(_2404_),
    .B(_2215_),
    .Y(_2405_)
);

NAND2X1 _11229_ (
    .A(_2403_),
    .B(_2405_),
    .Y(_2406_)
);

NOR2X1 _11230_ (
    .A(_2183_),
    .B(_2406_),
    .Y(_2407_)
);

NAND3X1 _11231_ (
    .A(_2402_),
    .B(_2407_),
    .C(_2398_),
    .Y(_2408_)
);

NAND2X1 _11232_ (
    .A(_2203_),
    .B(_2204_),
    .Y(_2409_)
);

OAI21X1 _11233_ (
    .A(_2399_),
    .B(_2207_),
    .C(_2175_),
    .Y(_2410_)
);

INVX1 _11234_ (
    .A(_2410_),
    .Y(_2411_)
);

OAI21X1 _11235_ (
    .A(_2403_),
    .B(_2202_),
    .C(_2181_),
    .Y(_2412_)
);

INVX1 _11236_ (
    .A(_2412_),
    .Y(_2413_)
);

OAI21X1 _11237_ (
    .A(_2411_),
    .B(_2409_),
    .C(_2413_),
    .Y(_2414_)
);

OAI21X1 _11238_ (
    .A(_2195_),
    .B(_2221_),
    .C(_2168_),
    .Y(_2415_)
);

INVX1 _11239_ (
    .A(_2415_),
    .Y(_2416_)
);

AOI21X1 _11240_ (
    .A(_2163_),
    .B(_2165_),
    .C(_2190_),
    .Y(_2417_)
);

OAI21X1 _11241_ (
    .A(_2416_),
    .B(_2395_),
    .C(_2417_),
    .Y(_2418_)
);

AOI21X1 _11242_ (
    .A(_2414_),
    .B(_2398_),
    .C(_2418_),
    .Y(_2419_)
);

OAI21X1 _11243_ (
    .A(_2408_),
    .B(_2394_),
    .C(_2419_),
    .Y(_2420_)
);

NAND2X1 _11244_ (
    .A(_2236_),
    .B(_2241_),
    .Y(_2421_)
);

NAND2X1 _11245_ (
    .A(_2251_),
    .B(_2247_),
    .Y(_2422_)
);

NOR2X1 _11246_ (
    .A(_2422_),
    .B(_2421_),
    .Y(_2423_)
);

NAND2X1 _11247_ (
    .A(_2257_),
    .B(_2262_),
    .Y(_2424_)
);

NOR2X1 _11248_ (
    .A(_2267_),
    .B(_2266_),
    .Y(_2425_)
);

INVX2 _11249_ (
    .A(_2272_),
    .Y(_2426_)
);

NAND2X1 _11250_ (
    .A(_2425_),
    .B(_2426_),
    .Y(_2427_)
);

NOR2X1 _11251_ (
    .A(_2424_),
    .B(_2427_),
    .Y(_2428_)
);

NAND2X1 _11252_ (
    .A(_2423_),
    .B(_2428_),
    .Y(_2429_)
);

INVX1 _11253_ (
    .A(_2429_),
    .Y(_2430_)
);

OAI21X1 _11254_ (
    .A(_2264_),
    .B(_2265_),
    .C(_2268_),
    .Y(_2431_)
);

OAI21X1 _11255_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .C(_2431_),
    .Y(_2432_)
);

INVX1 _11256_ (
    .A(_2261_),
    .Y(_2433_)
);

AOI21X1 _11257_ (
    .A(_2433_),
    .B(_2256_),
    .C(_2260_),
    .Y(_2434_)
);

OAI21X1 _11258_ (
    .A(_2432_),
    .B(_2424_),
    .C(_2434_),
    .Y(_2435_)
);

NAND2X1 _11259_ (
    .A(_2423_),
    .B(_2435_),
    .Y(_2436_)
);

INVX1 _11260_ (
    .A(_2245_),
    .Y(_2437_)
);

OAI21X1 _11261_ (
    .A(_2248_),
    .B(_2246_),
    .C(_2437_),
    .Y(_2438_)
);

INVX2 _11262_ (
    .A(_2438_),
    .Y(_2439_)
);

OR2X2 _11263_ (
    .A(_2439_),
    .B(_2421_),
    .Y(_2440_)
);

INVX1 _11264_ (
    .A(_2240_),
    .Y(_2441_)
);

AOI21X1 _11265_ (
    .A(_2441_),
    .B(_2235_),
    .C(_2239_),
    .Y(_2442_)
);

NAND3X1 _11266_ (
    .A(_2440_),
    .B(_2442_),
    .C(_2436_),
    .Y(_2443_)
);

AOI21X1 _11267_ (
    .A(_2420_),
    .B(_2430_),
    .C(_2443_),
    .Y(_2444_)
);

NAND2X1 _11268_ (
    .A(_2301_),
    .B(_2306_),
    .Y(_2445_)
);

NOR2X1 _11269_ (
    .A(_2315_),
    .B(_2314_),
    .Y(_2446_)
);

INVX2 _11270_ (
    .A(_2446_),
    .Y(_2447_)
);

NOR2X1 _11271_ (
    .A(_2311_),
    .B(_2447_),
    .Y(_2448_)
);

INVX1 _11272_ (
    .A(_2448_),
    .Y(_2449_)
);

NOR2X1 _11273_ (
    .A(_2445_),
    .B(_2449_),
    .Y(_2450_)
);

INVX1 _11274_ (
    .A(_2450_),
    .Y(_2451_)
);

INVX1 _11275_ (
    .A(_2445_),
    .Y(_2452_)
);

INVX1 _11276_ (
    .A(_2314_),
    .Y(_2453_)
);

OAI21X1 _11277_ (
    .A(_2309_),
    .B(_2453_),
    .C(_2308_),
    .Y(_2454_)
);

INVX1 _11278_ (
    .A(_2300_),
    .Y(_2455_)
);

INVX1 _11279_ (
    .A(_2304_),
    .Y(_2456_)
);

OAI21X1 _11280_ (
    .A(_2305_),
    .B(_2455_),
    .C(_2456_),
    .Y(_2457_)
);

AOI21X1 _11281_ (
    .A(_2452_),
    .B(_2454_),
    .C(_2457_),
    .Y(_2458_)
);

OAI21X1 _11282_ (
    .A(_2451_),
    .B(_2444_),
    .C(_2458_),
    .Y(_2459_)
);

NOR2X1 _11283_ (
    .A(_2334_),
    .B(_2333_),
    .Y(_2460_)
);

INVX1 _11284_ (
    .A(_2460_),
    .Y(_2461_)
);

NOR2X1 _11285_ (
    .A(_2338_),
    .B(_2461_),
    .Y(_2462_)
);

OAI21X1 _11286_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .C(_2335_),
    .Y(_2463_)
);

OAI21X1 _11287_ (
    .A(_2331_),
    .B(_2332_),
    .C(_2463_),
    .Y(_2464_)
);

AOI21X1 _11288_ (
    .A(_2459_),
    .B(_2462_),
    .C(_2464_),
    .Y(_2465_)
);

OAI21X1 _11289_ (
    .A(_2115_),
    .B(_2465_),
    .C(_2371_),
    .Y(_2466_)
);

NAND2X1 _11290_ (
    .A(_2364_),
    .B(_2350_),
    .Y(_2467_)
);

AOI21X1 _11291_ (
    .A(_2466_),
    .B(_2109_),
    .C(_2467_),
    .Y(_2468_)
);

OAI21X1 _11292_ (
    .A(_2109_),
    .B(_2466_),
    .C(_2468_),
    .Y(_2469_)
);

NAND3X1 _11293_ (
    .A(_2370_),
    .B(_2469_),
    .C(_2360_),
    .Y(\datapath_1.ALUResult [31])
);

OR2X2 _11294_ (
    .A(_2346_),
    .B(_2357_),
    .Y(_2470_)
);

NOR2X1 _11295_ (
    .A(_2353_),
    .B(_2358_),
    .Y(_2471_)
);

NAND2X1 _11296_ (
    .A(_2115_),
    .B(_2362__bF$buf2),
    .Y(_2472_)
);

OAI21X1 _11297_ (
    .A(_2365__bF$buf3),
    .B(_2357_),
    .C(_2472_),
    .Y(_2473_)
);

OAI22X1 _11298_ (
    .A(_2115_),
    .B(_2368__bF$buf2),
    .C(_2367__bF$buf2),
    .D(_2371_),
    .Y(_2474_)
);

NOR2X1 _11299_ (
    .A(_2474_),
    .B(_2473_),
    .Y(_2475_)
);

AND2X2 _11300_ (
    .A(_2465_),
    .B(_2357_),
    .Y(_2476_)
);

INVX8 _11301_ (
    .A(_2467_),
    .Y(_2477_)
);

OAI21X1 _11302_ (
    .A(_2357_),
    .B(_2465_),
    .C(_2477__bF$buf3),
    .Y(_2478_)
);

OAI21X1 _11303_ (
    .A(_2476_),
    .B(_2478_),
    .C(_2475_),
    .Y(_2479_)
);

AOI21X1 _11304_ (
    .A(_2471_),
    .B(_2470_),
    .C(_2479_),
    .Y(_2480_)
);

INVX1 _11305_ (
    .A(_2480_),
    .Y(\datapath_1.ALUResult [30])
);

AOI21X1 _11306_ (
    .A(_2459_),
    .B(_2337_),
    .C(_2335_),
    .Y(_2481_)
);

AND2X2 _11307_ (
    .A(_2481_),
    .B(_2461_),
    .Y(_2482_)
);

OAI21X1 _11308_ (
    .A(_2461_),
    .B(_2481_),
    .C(_2477__bF$buf2),
    .Y(_2483_)
);

INVX2 _11309_ (
    .A(_2365__bF$buf2),
    .Y(_2484_)
);

INVX1 _11310_ (
    .A(_2334_),
    .Y(_2485_)
);

NAND2X1 _11311_ (
    .A(_2361_),
    .B(_2352_),
    .Y(_2486_)
);

INVX8 _11312_ (
    .A(_2367__bF$buf1),
    .Y(_2487_)
);

NAND2X1 _11313_ (
    .A(_2333_),
    .B(_2487_),
    .Y(_2488_)
);

OAI21X1 _11314_ (
    .A(_2485_),
    .B(_2486_),
    .C(_2488_),
    .Y(_2489_)
);

AOI21X1 _11315_ (
    .A(_2460_),
    .B(_2484_),
    .C(_2489_),
    .Y(_2490_)
);

OAI21X1 _11316_ (
    .A(_2334_),
    .B(_2368__bF$buf1),
    .C(_2490_),
    .Y(_2491_)
);

INVX1 _11317_ (
    .A(_2343_),
    .Y(_2492_)
);

OAI21X1 _11318_ (
    .A(_2330_),
    .B(_2319_),
    .C(_2338_),
    .Y(_2493_)
);

NAND3X1 _11319_ (
    .A(_2492_),
    .B(_2460_),
    .C(_2493_),
    .Y(_2494_)
);

NOR2X1 _11320_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2116_),
    .Y(_2495_)
);

NAND2X1 _11321_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2496_)
);

NAND2X1 _11322_ (
    .A(_2496_),
    .B(_2378_),
    .Y(_2497_)
);

AOI21X1 _11323_ (
    .A(_2497_),
    .B(_2118_),
    .C(_2495_),
    .Y(_2498_)
);

INVX2 _11324_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2499_)
);

OR2X2 _11325_ (
    .A(\datapath_1.alu_1.ALUInA [1]),
    .B(\datapath_1.alu_1.ALUInB [1]),
    .Y(_2500_)
);

AOI22X1 _11326_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(_2499_),
    .C(_2374_),
    .D(_2500_),
    .Y(_2501_)
);

NAND2X1 _11327_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2502_)
);

INVX1 _11328_ (
    .A(_2131_),
    .Y(_2503_)
);

AOI22X1 _11329_ (
    .A(_2496_),
    .B(_2378_),
    .C(_2502_),
    .D(_2503_),
    .Y(_2504_)
);

OAI21X1 _11330_ (
    .A(_2124_),
    .B(_2501_),
    .C(_2504_),
    .Y(_2505_)
);

NAND2X1 _11331_ (
    .A(_2498_),
    .B(_2505_),
    .Y(_2506_)
);

INVX1 _11332_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .Y(_2507_)
);

NAND2X1 _11333_ (
    .A(_2507_),
    .B(_2148_),
    .Y(_2508_)
);

NAND2X1 _11334_ (
    .A(_2387_),
    .B(_2508_),
    .Y(_2509_)
);

NOR2X1 _11335_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(_2151_),
    .Y(_2510_)
);

AOI21X1 _11336_ (
    .A(_2509_),
    .B(_2510_),
    .C(_2149_),
    .Y(_2511_)
);

NAND2X1 _11337_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2512_)
);

NAND2X1 _11338_ (
    .A(_2512_),
    .B(_2391_),
    .Y(_2513_)
);

NOR2X1 _11339_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2154_),
    .Y(_2514_)
);

AOI21X1 _11340_ (
    .A(_2513_),
    .B(_2156_),
    .C(_2514_),
    .Y(_2515_)
);

OAI21X1 _11341_ (
    .A(_2138_),
    .B(_2511_),
    .C(_2515_),
    .Y(_2516_)
);

AOI21X1 _11342_ (
    .A(_2506_),
    .B(_2144_),
    .C(_2516_),
    .Y(_2517_)
);

INVX1 _11343_ (
    .A(_2210_),
    .Y(_2518_)
);

INVX1 _11344_ (
    .A(_2212_),
    .Y(_2519_)
);

AOI21X1 _11345_ (
    .A(_2177_),
    .B(_2519_),
    .C(_2518_),
    .Y(_2520_)
);

NOR2X1 _11346_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(_2214_),
    .Y(_2521_)
);

AOI21X1 _11347_ (
    .A(_2183_),
    .B(_2216_),
    .C(_2521_),
    .Y(_2522_)
);

OAI21X1 _11348_ (
    .A(_2186_),
    .B(_2520_),
    .C(_2522_),
    .Y(_2523_)
);

NAND2X1 _11349_ (
    .A(_2194_),
    .B(_2226_),
    .Y(_2524_)
);

NAND2X1 _11350_ (
    .A(\datapath_1.alu_1.ALUInA [15]),
    .B(_2161_),
    .Y(_2525_)
);

NAND3X1 _11351_ (
    .A(_2229_),
    .B(_2525_),
    .C(_2524_),
    .Y(_2526_)
);

AOI21X1 _11352_ (
    .A(_2174_),
    .B(_2523_),
    .C(_2526_),
    .Y(_2527_)
);

OAI21X1 _11353_ (
    .A(_2517_),
    .B(_2188_),
    .C(_2527_),
    .Y(_2528_)
);

AOI21X1 _11354_ (
    .A(_2528_),
    .B(_2276_),
    .C(_2295_),
    .Y(_2529_)
);

OAI21X1 _11355_ (
    .A(_2318_),
    .B(_2529_),
    .C(_2329_),
    .Y(_2530_)
);

OAI21X1 _11356_ (
    .A(_2492_),
    .B(_2460_),
    .C(_2354__bF$buf2),
    .Y(_2531_)
);

AOI21X1 _11357_ (
    .A(_2530_),
    .B(_2340_),
    .C(_2531_),
    .Y(_2532_)
);

AOI21X1 _11358_ (
    .A(_2532_),
    .B(_2494_),
    .C(_2491_),
    .Y(_2533_)
);

OAI21X1 _11359_ (
    .A(_2482_),
    .B(_2483_),
    .C(_2533_),
    .Y(\datapath_1.ALUResult [29])
);

OR2X2 _11360_ (
    .A(_2143_),
    .B(_2138_),
    .Y(_2534_)
);

AOI21X1 _11361_ (
    .A(_2505_),
    .B(_2498_),
    .C(_2534_),
    .Y(_2535_)
);

AND2X2 _11362_ (
    .A(_2174_),
    .B(_2187_),
    .Y(_2536_)
);

OAI21X1 _11363_ (
    .A(_2516_),
    .B(_2535_),
    .C(_2536_),
    .Y(_2537_)
);

INVX1 _11364_ (
    .A(_2276_),
    .Y(_2538_)
);

AOI21X1 _11365_ (
    .A(_2537_),
    .B(_2527_),
    .C(_2538_),
    .Y(_2539_)
);

INVX1 _11366_ (
    .A(_2318_),
    .Y(_2540_)
);

OAI21X1 _11367_ (
    .A(_2295_),
    .B(_2539_),
    .C(_2540_),
    .Y(_2541_)
);

NAND3X1 _11368_ (
    .A(_2329_),
    .B(_2337_),
    .C(_2541_),
    .Y(_2542_)
);

NAND3X1 _11369_ (
    .A(_2354__bF$buf1),
    .B(_2493_),
    .C(_2542_),
    .Y(_2543_)
);

NAND2X1 _11370_ (
    .A(_2336_),
    .B(_2362__bF$buf1),
    .Y(_2544_)
);

OAI21X1 _11371_ (
    .A(_2365__bF$buf1),
    .B(_2338_),
    .C(_2544_),
    .Y(_2545_)
);

NAND2X1 _11372_ (
    .A(_2335_),
    .B(_2487_),
    .Y(_2546_)
);

OAI21X1 _11373_ (
    .A(_2336_),
    .B(_2368__bF$buf0),
    .C(_2546_),
    .Y(_2547_)
);

NOR2X1 _11374_ (
    .A(_2547_),
    .B(_2545_),
    .Y(_2548_)
);

NAND2X1 _11375_ (
    .A(_2337_),
    .B(_2459_),
    .Y(_2549_)
);

NAND2X1 _11376_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2550_)
);

OR2X2 _11377_ (
    .A(\datapath_1.alu_1.ALUInA [6]),
    .B(\datapath_1.alu_1.ALUInB [6]),
    .Y(_2551_)
);

NAND2X1 _11378_ (
    .A(_2550_),
    .B(_2551_),
    .Y(_2552_)
);

NOR2X1 _11379_ (
    .A(_2552_),
    .B(_2513_),
    .Y(_2553_)
);

OR2X2 _11380_ (
    .A(\datapath_1.alu_1.ALUInA [4]),
    .B(\datapath_1.alu_1.ALUInB [4]),
    .Y(_2554_)
);

NAND2X1 _11381_ (
    .A(_2388_),
    .B(_2554_),
    .Y(_2555_)
);

NOR2X1 _11382_ (
    .A(_2555_),
    .B(_2509_),
    .Y(_2556_)
);

NAND2X1 _11383_ (
    .A(_2553_),
    .B(_2556_),
    .Y(_2557_)
);

AOI21X1 _11384_ (
    .A(_2377_),
    .B(_2379_),
    .C(_2557_),
    .Y(_2558_)
);

NOR2X1 _11385_ (
    .A(_2170_),
    .B(_2199_),
    .Y(_2559_)
);

NAND3X1 _11386_ (
    .A(_2193_),
    .B(_2192_),
    .C(_2559_),
    .Y(_2560_)
);

NAND2X1 _11387_ (
    .A(_2402_),
    .B(_2407_),
    .Y(_2561_)
);

NOR2X1 _11388_ (
    .A(_2561_),
    .B(_2560_),
    .Y(_2562_)
);

OAI21X1 _11389_ (
    .A(_2393_),
    .B(_2558_),
    .C(_2562_),
    .Y(_2563_)
);

AOI21X1 _11390_ (
    .A(_2563_),
    .B(_2419_),
    .C(_2429_),
    .Y(_2564_)
);

OAI21X1 _11391_ (
    .A(_2443_),
    .B(_2564_),
    .C(_2450_),
    .Y(_2565_)
);

NAND3X1 _11392_ (
    .A(_2338_),
    .B(_2458_),
    .C(_2565_),
    .Y(_2566_)
);

NAND3X1 _11393_ (
    .A(_2477__bF$buf1),
    .B(_2566_),
    .C(_2549_),
    .Y(_2567_)
);

NAND3X1 _11394_ (
    .A(_2548_),
    .B(_2543_),
    .C(_2567_),
    .Y(\datapath_1.ALUResult [28])
);

INVX1 _11395_ (
    .A(_2326_),
    .Y(_2568_)
);

INVX2 _11396_ (
    .A(_2301_),
    .Y(_2569_)
);

AOI21X1 _11397_ (
    .A(_2277_),
    .B(_2296_),
    .C(_2316_),
    .Y(_2570_)
);

OAI21X1 _11398_ (
    .A(_2324_),
    .B(_2570_),
    .C(_2569_),
    .Y(_2571_)
);

NAND3X1 _11399_ (
    .A(_2568_),
    .B(_2306_),
    .C(_2571_),
    .Y(_2572_)
);

INVX1 _11400_ (
    .A(_2306_),
    .Y(_2573_)
);

INVX1 _11401_ (
    .A(_2324_),
    .Y(_2574_)
);

OAI21X1 _11402_ (
    .A(_2295_),
    .B(_2539_),
    .C(_2317_),
    .Y(_2575_)
);

AOI21X1 _11403_ (
    .A(_2575_),
    .B(_2574_),
    .C(_2301_),
    .Y(_2576_)
);

OAI21X1 _11404_ (
    .A(_2326_),
    .B(_2576_),
    .C(_2573_),
    .Y(_2577_)
);

NAND3X1 _11405_ (
    .A(_2572_),
    .B(_2354__bF$buf0),
    .C(_2577_),
    .Y(_2578_)
);

INVX1 _11406_ (
    .A(_2305_),
    .Y(_2579_)
);

OAI22X1 _11407_ (
    .A(_2367__bF$buf0),
    .B(_2456_),
    .C(_2579_),
    .D(_2486_),
    .Y(_2580_)
);

OAI21X1 _11408_ (
    .A(_2304_),
    .B(_2365__bF$buf0),
    .C(_2368__bF$buf3),
    .Y(_2581_)
);

AOI21X1 _11409_ (
    .A(_2581_),
    .B(_2579_),
    .C(_2580_),
    .Y(_2582_)
);

INVX1 _11410_ (
    .A(_2454_),
    .Y(_2583_)
);

OAI21X1 _11411_ (
    .A(_2449_),
    .B(_2444_),
    .C(_2583_),
    .Y(_2584_)
);

NAND2X1 _11412_ (
    .A(_2301_),
    .B(_2584_),
    .Y(_2585_)
);

NAND3X1 _11413_ (
    .A(_2573_),
    .B(_2455_),
    .C(_2585_),
    .Y(_2586_)
);

OAI21X1 _11414_ (
    .A(_2443_),
    .B(_2564_),
    .C(_2448_),
    .Y(_2587_)
);

AOI21X1 _11415_ (
    .A(_2587_),
    .B(_2583_),
    .C(_2569_),
    .Y(_2588_)
);

OAI21X1 _11416_ (
    .A(_2300_),
    .B(_2588_),
    .C(_2306_),
    .Y(_2589_)
);

NAND3X1 _11417_ (
    .A(_2586_),
    .B(_2477__bF$buf0),
    .C(_2589_),
    .Y(_2590_)
);

NAND3X1 _11418_ (
    .A(_2582_),
    .B(_2578_),
    .C(_2590_),
    .Y(\datapath_1.ALUResult [27])
);

NAND3X1 _11419_ (
    .A(_2574_),
    .B(_2301_),
    .C(_2575_),
    .Y(_2591_)
);

NAND3X1 _11420_ (
    .A(_2354__bF$buf3),
    .B(_2571_),
    .C(_2591_),
    .Y(_2592_)
);

NAND2X1 _11421_ (
    .A(_2297_),
    .B(_2362__bF$buf0),
    .Y(_2593_)
);

OAI21X1 _11422_ (
    .A(_2365__bF$buf4),
    .B(_2569_),
    .C(_2593_),
    .Y(_2594_)
);

OAI22X1 _11423_ (
    .A(_2297_),
    .B(_2368__bF$buf2),
    .C(_2367__bF$buf3),
    .D(_2455_),
    .Y(_2595_)
);

NOR2X1 _11424_ (
    .A(_2595_),
    .B(_2594_),
    .Y(_2596_)
);

NAND3X1 _11425_ (
    .A(_2583_),
    .B(_2569_),
    .C(_2587_),
    .Y(_2597_)
);

NAND3X1 _11426_ (
    .A(_2477__bF$buf3),
    .B(_2597_),
    .C(_2585_),
    .Y(_2598_)
);

NAND3X1 _11427_ (
    .A(_2596_),
    .B(_2592_),
    .C(_2598_),
    .Y(\datapath_1.ALUResult [26])
);

INVX1 _11428_ (
    .A(_2311_),
    .Y(_2599_)
);

OAI21X1 _11429_ (
    .A(_2447_),
    .B(_2444_),
    .C(_2453_),
    .Y(_2600_)
);

XNOR2X1 _11430_ (
    .A(_2600_),
    .B(_2599_),
    .Y(_2601_)
);

OAI22X1 _11431_ (
    .A(_2367__bF$buf2),
    .B(_2308_),
    .C(_2310_),
    .D(_2486_),
    .Y(_2602_)
);

AOI21X1 _11432_ (
    .A(_2599_),
    .B(_2484_),
    .C(_2602_),
    .Y(_2603_)
);

OAI21X1 _11433_ (
    .A(_2309_),
    .B(_2368__bF$buf1),
    .C(_2603_),
    .Y(_2604_)
);

NOR2X1 _11434_ (
    .A(_2322_),
    .B(_2311_),
    .Y(_2605_)
);

OAI21X1 _11435_ (
    .A(_2446_),
    .B(_2529_),
    .C(_2605_),
    .Y(_2606_)
);

NAND2X1 _11436_ (
    .A(_2354__bF$buf2),
    .B(_2323_),
    .Y(_2607_)
);

NOR2X1 _11437_ (
    .A(_2607_),
    .B(_2570_),
    .Y(_2608_)
);

AOI21X1 _11438_ (
    .A(_2608_),
    .B(_2606_),
    .C(_2604_),
    .Y(_2609_)
);

OAI21X1 _11439_ (
    .A(_2467_),
    .B(_2601_),
    .C(_2609_),
    .Y(\datapath_1.ALUResult [25])
);

NAND2X1 _11440_ (
    .A(_2296_),
    .B(_2277_),
    .Y(_2610_)
);

AOI21X1 _11441_ (
    .A(_2610_),
    .B(_2447_),
    .C(_2353_),
    .Y(_2611_)
);

OAI21X1 _11442_ (
    .A(_2610_),
    .B(_2447_),
    .C(_2611_),
    .Y(_2612_)
);

NAND2X1 _11443_ (
    .A(_2315_),
    .B(_2362__bF$buf3),
    .Y(_2613_)
);

OAI21X1 _11444_ (
    .A(_2365__bF$buf3),
    .B(_2447_),
    .C(_2613_),
    .Y(_2614_)
);

OAI22X1 _11445_ (
    .A(_2315_),
    .B(_2368__bF$buf0),
    .C(_2367__bF$buf1),
    .D(_2453_),
    .Y(_2615_)
);

NOR2X1 _11446_ (
    .A(_2615_),
    .B(_2614_),
    .Y(_2616_)
);

INVX1 _11447_ (
    .A(_2616_),
    .Y(_2617_)
);

XNOR2X1 _11448_ (
    .A(_2444_),
    .B(_2446_),
    .Y(_2618_)
);

AOI21X1 _11449_ (
    .A(_2618_),
    .B(_2477__bF$buf2),
    .C(_2617_),
    .Y(_2619_)
);

NAND2X1 _11450_ (
    .A(_2612_),
    .B(_2619_),
    .Y(\datapath_1.ALUResult [24])
);

INVX1 _11451_ (
    .A(_2291_),
    .Y(_2620_)
);

INVX2 _11452_ (
    .A(_2236_),
    .Y(_2621_)
);

INVX1 _11453_ (
    .A(_2252_),
    .Y(_2622_)
);

INVX1 _11454_ (
    .A(_2275_),
    .Y(_2623_)
);

OAI21X1 _11455_ (
    .A(_2232_),
    .B(_2189_),
    .C(_2623_),
    .Y(_2624_)
);

AOI21X1 _11456_ (
    .A(_2624_),
    .B(_2285_),
    .C(_2622_),
    .Y(_2625_)
);

OAI21X1 _11457_ (
    .A(_2289_),
    .B(_2625_),
    .C(_2621_),
    .Y(_2626_)
);

NAND3X1 _11458_ (
    .A(_2620_),
    .B(_2241_),
    .C(_2626_),
    .Y(_2627_)
);

INVX1 _11459_ (
    .A(_2241_),
    .Y(_2628_)
);

INVX1 _11460_ (
    .A(_2233_),
    .Y(_2629_)
);

INVX1 _11461_ (
    .A(_2289_),
    .Y(_2630_)
);

INVX1 _11462_ (
    .A(_2285_),
    .Y(_2631_)
);

AOI21X1 _11463_ (
    .A(_2537_),
    .B(_2527_),
    .C(_2275_),
    .Y(_2632_)
);

OAI21X1 _11464_ (
    .A(_2631_),
    .B(_2632_),
    .C(_2252_),
    .Y(_2633_)
);

AOI22X1 _11465_ (
    .A(_2629_),
    .B(_2234_),
    .C(_2630_),
    .D(_2633_),
    .Y(_2634_)
);

OAI21X1 _11466_ (
    .A(_2291_),
    .B(_2634_),
    .C(_2628_),
    .Y(_2635_)
);

NAND3X1 _11467_ (
    .A(_2627_),
    .B(_2354__bF$buf1),
    .C(_2635_),
    .Y(_2636_)
);

INVX4 _11468_ (
    .A(_2368__bF$buf3),
    .Y(_2637_)
);

AOI22X1 _11469_ (
    .A(_2239_),
    .B(_2487_),
    .C(_2240_),
    .D(_2362__bF$buf2),
    .Y(_2638_)
);

OAI21X1 _11470_ (
    .A(_2628_),
    .B(_2365__bF$buf2),
    .C(_2638_),
    .Y(_2639_)
);

AOI21X1 _11471_ (
    .A(_2441_),
    .B(_2637_),
    .C(_2639_),
    .Y(_2640_)
);

AOI21X1 _11472_ (
    .A(_2420_),
    .B(_2428_),
    .C(_2435_),
    .Y(_2641_)
);

OAI21X1 _11473_ (
    .A(_2422_),
    .B(_2641_),
    .C(_2439_),
    .Y(_2642_)
);

NAND2X1 _11474_ (
    .A(_2236_),
    .B(_2642_),
    .Y(_2643_)
);

NAND3X1 _11475_ (
    .A(_2628_),
    .B(_2234_),
    .C(_2643_),
    .Y(_2644_)
);

INVX1 _11476_ (
    .A(_2422_),
    .Y(_2645_)
);

INVX1 _11477_ (
    .A(_2428_),
    .Y(_2646_)
);

AOI21X1 _11478_ (
    .A(_2563_),
    .B(_2419_),
    .C(_2646_),
    .Y(_2647_)
);

OAI21X1 _11479_ (
    .A(_2435_),
    .B(_2647_),
    .C(_2645_),
    .Y(_2648_)
);

AOI21X1 _11480_ (
    .A(_2648_),
    .B(_2439_),
    .C(_2621_),
    .Y(_2649_)
);

OAI21X1 _11481_ (
    .A(_2235_),
    .B(_2649_),
    .C(_2241_),
    .Y(_2650_)
);

NAND3X1 _11482_ (
    .A(_2644_),
    .B(_2477__bF$buf1),
    .C(_2650_),
    .Y(_2651_)
);

NAND3X1 _11483_ (
    .A(_2640_),
    .B(_2636_),
    .C(_2651_),
    .Y(\datapath_1.ALUResult [23])
);

NAND3X1 _11484_ (
    .A(_2630_),
    .B(_2236_),
    .C(_2633_),
    .Y(_2652_)
);

NAND3X1 _11485_ (
    .A(_2354__bF$buf0),
    .B(_2626_),
    .C(_2652_),
    .Y(_2653_)
);

AOI22X1 _11486_ (
    .A(_2487_),
    .B(_2235_),
    .C(_2233_),
    .D(_2362__bF$buf1),
    .Y(_2654_)
);

OAI21X1 _11487_ (
    .A(_2621_),
    .B(_2365__bF$buf1),
    .C(_2654_),
    .Y(_2655_)
);

AOI21X1 _11488_ (
    .A(_2629_),
    .B(_2637_),
    .C(_2655_),
    .Y(_2656_)
);

NAND3X1 _11489_ (
    .A(_2439_),
    .B(_2621_),
    .C(_2648_),
    .Y(_2657_)
);

NAND3X1 _11490_ (
    .A(_2477__bF$buf0),
    .B(_2657_),
    .C(_2643_),
    .Y(_2658_)
);

NAND3X1 _11491_ (
    .A(_2656_),
    .B(_2653_),
    .C(_2658_),
    .Y(\datapath_1.ALUResult [22])
);

INVX2 _11492_ (
    .A(_2251_),
    .Y(_2659_)
);

OAI21X1 _11493_ (
    .A(_2659_),
    .B(_2641_),
    .C(_2248_),
    .Y(_2660_)
);

NAND2X1 _11494_ (
    .A(_2247_),
    .B(_2660_),
    .Y(_2661_)
);

OR2X2 _11495_ (
    .A(_2660_),
    .B(_2247_),
    .Y(_2662_)
);

NAND3X1 _11496_ (
    .A(_2477__bF$buf3),
    .B(_2661_),
    .C(_2662_),
    .Y(_2663_)
);

INVX1 _11497_ (
    .A(_2246_),
    .Y(_2664_)
);

INVX1 _11498_ (
    .A(_2247_),
    .Y(_2665_)
);

AOI22X1 _11499_ (
    .A(_2245_),
    .B(_2487_),
    .C(_2246_),
    .D(_2362__bF$buf0),
    .Y(_2666_)
);

OAI21X1 _11500_ (
    .A(_2665_),
    .B(_2365__bF$buf0),
    .C(_2666_),
    .Y(_2667_)
);

AOI21X1 _11501_ (
    .A(_2664_),
    .B(_2637_),
    .C(_2667_),
    .Y(_2668_)
);

INVX1 _11502_ (
    .A(_2668_),
    .Y(_2669_)
);

INVX1 _11503_ (
    .A(_2287_),
    .Y(_2670_)
);

OAI21X1 _11504_ (
    .A(_2631_),
    .B(_2632_),
    .C(_2659_),
    .Y(_2671_)
);

NAND3X1 _11505_ (
    .A(_2670_),
    .B(_2247_),
    .C(_2671_),
    .Y(_2672_)
);

OAI21X1 _11506_ (
    .A(_2670_),
    .B(_2247_),
    .C(_2354__bF$buf3),
    .Y(_2673_)
);

NOR2X1 _11507_ (
    .A(_2673_),
    .B(_2625_),
    .Y(_2674_)
);

AOI21X1 _11508_ (
    .A(_2672_),
    .B(_2674_),
    .C(_2669_),
    .Y(_2675_)
);

NAND2X1 _11509_ (
    .A(_2675_),
    .B(_2663_),
    .Y(\datapath_1.ALUResult [21])
);

NAND3X1 _11510_ (
    .A(_2285_),
    .B(_2251_),
    .C(_2624_),
    .Y(_2676_)
);

AND2X2 _11511_ (
    .A(_2671_),
    .B(_2354__bF$buf2),
    .Y(_2677_)
);

NAND2X1 _11512_ (
    .A(_2250_),
    .B(_2362__bF$buf3),
    .Y(_2678_)
);

OAI21X1 _11513_ (
    .A(_2659_),
    .B(_2365__bF$buf4),
    .C(_2678_),
    .Y(_2679_)
);

OAI22X1 _11514_ (
    .A(_2367__bF$buf0),
    .B(_2248_),
    .C(_2250_),
    .D(_2368__bF$buf2),
    .Y(_2680_)
);

NOR2X1 _11515_ (
    .A(_2680_),
    .B(_2679_),
    .Y(_2681_)
);

AND2X2 _11516_ (
    .A(_2641_),
    .B(_2659_),
    .Y(_2682_)
);

OAI21X1 _11517_ (
    .A(_2659_),
    .B(_2641_),
    .C(_2477__bF$buf2),
    .Y(_2683_)
);

OAI21X1 _11518_ (
    .A(_2682_),
    .B(_2683_),
    .C(_2681_),
    .Y(_2684_)
);

AOI21X1 _11519_ (
    .A(_2677_),
    .B(_2676_),
    .C(_2684_),
    .Y(_2685_)
);

INVX1 _11520_ (
    .A(_2685_),
    .Y(\datapath_1.ALUResult [20])
);

INVX1 _11521_ (
    .A(_2262_),
    .Y(_2686_)
);

INVX1 _11522_ (
    .A(_2254_),
    .Y(_2687_)
);

INVX1 _11523_ (
    .A(_2280_),
    .Y(_2688_)
);

OAI21X1 _11524_ (
    .A(_2232_),
    .B(_2189_),
    .C(_2274_),
    .Y(_2689_)
);

AOI22X1 _11525_ (
    .A(_2687_),
    .B(_2255_),
    .C(_2688_),
    .D(_2689_),
    .Y(_2690_)
);

OAI21X1 _11526_ (
    .A(_2282_),
    .B(_2690_),
    .C(_2686_),
    .Y(_2691_)
);

INVX1 _11527_ (
    .A(_2282_),
    .Y(_2692_)
);

INVX2 _11528_ (
    .A(_2257_),
    .Y(_2693_)
);

AOI21X1 _11529_ (
    .A(_2537_),
    .B(_2527_),
    .C(_2273_),
    .Y(_2694_)
);

OAI21X1 _11530_ (
    .A(_2280_),
    .B(_2694_),
    .C(_2693_),
    .Y(_2695_)
);

NAND3X1 _11531_ (
    .A(_2692_),
    .B(_2262_),
    .C(_2695_),
    .Y(_2696_)
);

NAND3X1 _11532_ (
    .A(_2354__bF$buf1),
    .B(_2691_),
    .C(_2696_),
    .Y(_2697_)
);

OAI22X1 _11533_ (
    .A(_2486_),
    .B(_2433_),
    .C(_2365__bF$buf3),
    .D(_2686_),
    .Y(_2698_)
);

NAND2X1 _11534_ (
    .A(_2260_),
    .B(_2487_),
    .Y(_2699_)
);

OAI21X1 _11535_ (
    .A(_2261_),
    .B(_2368__bF$buf1),
    .C(_2699_),
    .Y(_2700_)
);

NOR2X1 _11536_ (
    .A(_2700_),
    .B(_2698_),
    .Y(_2701_)
);

INVX1 _11537_ (
    .A(_2432_),
    .Y(_2702_)
);

AOI21X1 _11538_ (
    .A(_2563_),
    .B(_2419_),
    .C(_2427_),
    .Y(_2703_)
);

OAI21X1 _11539_ (
    .A(_2702_),
    .B(_2703_),
    .C(_2257_),
    .Y(_2704_)
);

NAND3X1 _11540_ (
    .A(_2686_),
    .B(_2255_),
    .C(_2704_),
    .Y(_2705_)
);

INVX1 _11541_ (
    .A(_2267_),
    .Y(_2706_)
);

INVX1 _11542_ (
    .A(_2427_),
    .Y(_2707_)
);

AOI22X1 _11543_ (
    .A(_2431_),
    .B(_2706_),
    .C(_2707_),
    .D(_2420_),
    .Y(_2708_)
);

OAI21X1 _11544_ (
    .A(_2693_),
    .B(_2708_),
    .C(_2255_),
    .Y(_2709_)
);

NAND2X1 _11545_ (
    .A(_2262_),
    .B(_2709_),
    .Y(_2710_)
);

NAND3X1 _11546_ (
    .A(_2477__bF$buf1),
    .B(_2710_),
    .C(_2705_),
    .Y(_2711_)
);

NAND3X1 _11547_ (
    .A(_2701_),
    .B(_2697_),
    .C(_2711_),
    .Y(\datapath_1.ALUResult [19])
);

NAND3X1 _11548_ (
    .A(_2688_),
    .B(_2257_),
    .C(_2689_),
    .Y(_2712_)
);

NOR2X1 _11549_ (
    .A(_2353_),
    .B(_2690_),
    .Y(_2713_)
);

AOI22X1 _11550_ (
    .A(_2487_),
    .B(_2256_),
    .C(_2254_),
    .D(_2362__bF$buf2),
    .Y(_2714_)
);

OAI21X1 _11551_ (
    .A(_2693_),
    .B(_2365__bF$buf2),
    .C(_2714_),
    .Y(_2715_)
);

AOI21X1 _11552_ (
    .A(_2687_),
    .B(_2637_),
    .C(_2715_),
    .Y(_2716_)
);

AND2X2 _11553_ (
    .A(_2708_),
    .B(_2693_),
    .Y(_2717_)
);

OAI21X1 _11554_ (
    .A(_2693_),
    .B(_2708_),
    .C(_2477__bF$buf0),
    .Y(_2718_)
);

OAI21X1 _11555_ (
    .A(_2717_),
    .B(_2718_),
    .C(_2716_),
    .Y(_2719_)
);

AOI21X1 _11556_ (
    .A(_2712_),
    .B(_2713_),
    .C(_2719_),
    .Y(_2720_)
);

INVX1 _11557_ (
    .A(_2720_),
    .Y(\datapath_1.ALUResult [18])
);

NAND2X1 _11558_ (
    .A(_2426_),
    .B(_2420_),
    .Y(_2721_)
);

OAI21X1 _11559_ (
    .A(_2269_),
    .B(_2270_),
    .C(_2721_),
    .Y(_2722_)
);

OR2X2 _11560_ (
    .A(_2722_),
    .B(_2425_),
    .Y(_2723_)
);

AOI21X1 _11561_ (
    .A(_2722_),
    .B(_2425_),
    .C(_2467_),
    .Y(_2724_)
);

AOI22X1 _11562_ (
    .A(_2425_),
    .B(_2484_),
    .C(_2362__bF$buf1),
    .D(_2267_),
    .Y(_2725_)
);

AOI22X1 _11563_ (
    .A(_2487_),
    .B(_2266_),
    .C(_2637_),
    .D(_2706_),
    .Y(_2726_)
);

AND2X2 _11564_ (
    .A(_2725_),
    .B(_2726_),
    .Y(_2727_)
);

OAI21X1 _11565_ (
    .A(_2269_),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .C(_2425_),
    .Y(_2728_)
);

AOI21X1 _11566_ (
    .A(_2528_),
    .B(_2272_),
    .C(_2728_),
    .Y(_2729_)
);

NAND3X1 _11567_ (
    .A(_2354__bF$buf0),
    .B(_2279_),
    .C(_2689_),
    .Y(_2730_)
);

OAI21X1 _11568_ (
    .A(_2730_),
    .B(_2729_),
    .C(_2727_),
    .Y(_2731_)
);

AOI21X1 _11569_ (
    .A(_2723_),
    .B(_2724_),
    .C(_2731_),
    .Y(_2732_)
);

INVX1 _11570_ (
    .A(_2732_),
    .Y(\datapath_1.ALUResult [17])
);

OAI21X1 _11571_ (
    .A(_2232_),
    .B(_2189_),
    .C(_2272_),
    .Y(_2733_)
);

NAND3X1 _11572_ (
    .A(_2426_),
    .B(_2527_),
    .C(_2537_),
    .Y(_2734_)
);

NAND3X1 _11573_ (
    .A(_2354__bF$buf3),
    .B(_2733_),
    .C(_2734_),
    .Y(_2735_)
);

OAI22X1 _11574_ (
    .A(_2272_),
    .B(_2365__bF$buf1),
    .C(_2271_),
    .D(_2486_),
    .Y(_2736_)
);

OAI21X1 _11575_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .C(_2637_),
    .Y(_2737_)
);

OAI21X1 _11576_ (
    .A(_2268_),
    .B(_2367__bF$buf3),
    .C(_2737_),
    .Y(_2738_)
);

NOR2X1 _11577_ (
    .A(_2736_),
    .B(_2738_),
    .Y(_2739_)
);

AOI21X1 _11578_ (
    .A(_2420_),
    .B(_2426_),
    .C(_2467_),
    .Y(_2740_)
);

OAI21X1 _11579_ (
    .A(_2426_),
    .B(_2420_),
    .C(_2740_),
    .Y(_2741_)
);

NAND3X1 _11580_ (
    .A(_2739_),
    .B(_2735_),
    .C(_2741_),
    .Y(\datapath_1.ALUResult [16])
);

INVX1 _11581_ (
    .A(_2226_),
    .Y(_2742_)
);

NAND2X1 _11582_ (
    .A(_2159_),
    .B(_2145_),
    .Y(_2743_)
);

AOI21X1 _11583_ (
    .A(_2743_),
    .B(_2187_),
    .C(_2523_),
    .Y(_2744_)
);

OAI21X1 _11584_ (
    .A(_2173_),
    .B(_2744_),
    .C(_2742_),
    .Y(_2745_)
);

OAI21X1 _11585_ (
    .A(_2165_),
    .B(_2166_),
    .C(_2745_),
    .Y(_2746_)
);

OAI21X1 _11586_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(_2227_),
    .C(_2746_),
    .Y(_2747_)
);

OAI21X1 _11587_ (
    .A(_2190_),
    .B(_2191_),
    .C(_2747_),
    .Y(_2748_)
);

INVX1 _11588_ (
    .A(_2228_),
    .Y(_2749_)
);

NAND3X1 _11589_ (
    .A(_2749_),
    .B(_2192_),
    .C(_2746_),
    .Y(_2750_)
);

NAND3X1 _11590_ (
    .A(_2354__bF$buf2),
    .B(_2750_),
    .C(_2748_),
    .Y(_2751_)
);

OAI22X1 _11591_ (
    .A(_2367__bF$buf2),
    .B(_2160_),
    .C(_2163_),
    .D(_2486_),
    .Y(_2752_)
);

OAI21X1 _11592_ (
    .A(_2190_),
    .B(_2365__bF$buf0),
    .C(_2368__bF$buf0),
    .Y(_2753_)
);

AOI21X1 _11593_ (
    .A(_2753_),
    .B(_2163_),
    .C(_2752_),
    .Y(_2754_)
);

INVX1 _11594_ (
    .A(_2165_),
    .Y(_2755_)
);

INVX2 _11595_ (
    .A(_2193_),
    .Y(_2756_)
);

INVX1 _11596_ (
    .A(_2414_),
    .Y(_2757_)
);

OAI21X1 _11597_ (
    .A(_2561_),
    .B(_2394_),
    .C(_2757_),
    .Y(_2758_)
);

AOI21X1 _11598_ (
    .A(_2758_),
    .B(_2559_),
    .C(_2415_),
    .Y(_2759_)
);

NOR2X1 _11599_ (
    .A(_2756_),
    .B(_2759_),
    .Y(_2760_)
);

INVX1 _11600_ (
    .A(_2760_),
    .Y(_2761_)
);

NAND3X1 _11601_ (
    .A(_2755_),
    .B(_2164_),
    .C(_2761_),
    .Y(_2762_)
);

OAI21X1 _11602_ (
    .A(_2165_),
    .B(_2760_),
    .C(_2192_),
    .Y(_2763_)
);

NAND3X1 _11603_ (
    .A(_2477__bF$buf3),
    .B(_2763_),
    .C(_2762_),
    .Y(_2764_)
);

NAND3X1 _11604_ (
    .A(_2754_),
    .B(_2764_),
    .C(_2751_),
    .Y(\datapath_1.ALUResult [15])
);

OR2X2 _11605_ (
    .A(_2745_),
    .B(_2756_),
    .Y(_2765_)
);

AOI21X1 _11606_ (
    .A(_2745_),
    .B(_2756_),
    .C(_2353_),
    .Y(_2766_)
);

NAND2X1 _11607_ (
    .A(_2166_),
    .B(_2362__bF$buf0),
    .Y(_2767_)
);

OAI21X1 _11608_ (
    .A(_2756_),
    .B(_2365__bF$buf4),
    .C(_2767_),
    .Y(_2768_)
);

OAI22X1 _11609_ (
    .A(_2367__bF$buf1),
    .B(_2755_),
    .C(_2166_),
    .D(_2368__bF$buf3),
    .Y(_2769_)
);

NOR2X1 _11610_ (
    .A(_2769_),
    .B(_2768_),
    .Y(_2770_)
);

AND2X2 _11611_ (
    .A(_2759_),
    .B(_2756_),
    .Y(_2771_)
);

OAI21X1 _11612_ (
    .A(_2756_),
    .B(_2759_),
    .C(_2477__bF$buf2),
    .Y(_2772_)
);

OAI21X1 _11613_ (
    .A(_2771_),
    .B(_2772_),
    .C(_2770_),
    .Y(_2773_)
);

AOI21X1 _11614_ (
    .A(_2765_),
    .B(_2766_),
    .C(_2773_),
    .Y(_2774_)
);

INVX1 _11615_ (
    .A(_2774_),
    .Y(\datapath_1.ALUResult [14])
);

NAND2X1 _11616_ (
    .A(_2396_),
    .B(_2758_),
    .Y(_2775_)
);

OAI21X1 _11617_ (
    .A(_2196_),
    .B(_2197_),
    .C(_2775_),
    .Y(_2776_)
);

OR2X2 _11618_ (
    .A(_2776_),
    .B(_2222_),
    .Y(_2777_)
);

AOI21X1 _11619_ (
    .A(_2776_),
    .B(_2222_),
    .C(_2467_),
    .Y(_2778_)
);

OAI22X1 _11620_ (
    .A(_2170_),
    .B(_2365__bF$buf3),
    .C(_2169_),
    .D(_2486_),
    .Y(_2779_)
);

OAI22X1 _11621_ (
    .A(_2367__bF$buf0),
    .B(_2168_),
    .C(_2221_),
    .D(_2368__bF$buf2),
    .Y(_2780_)
);

NOR2X1 _11622_ (
    .A(_2780_),
    .B(_2779_),
    .Y(_2781_)
);

OAI21X1 _11623_ (
    .A(_2396_),
    .B(_2744_),
    .C(_2225_),
    .Y(_2782_)
);

NOR2X1 _11624_ (
    .A(_2170_),
    .B(_2782_),
    .Y(_2783_)
);

INVX1 _11625_ (
    .A(_2225_),
    .Y(_2784_)
);

AOI21X1 _11626_ (
    .A(_2170_),
    .B(_2784_),
    .C(_2353_),
    .Y(_2785_)
);

OAI21X1 _11627_ (
    .A(_2173_),
    .B(_2744_),
    .C(_2785_),
    .Y(_2786_)
);

OAI21X1 _11628_ (
    .A(_2786_),
    .B(_2783_),
    .C(_2781_),
    .Y(_2787_)
);

AOI21X1 _11629_ (
    .A(_2777_),
    .B(_2778_),
    .C(_2787_),
    .Y(_2788_)
);

INVX1 _11630_ (
    .A(_2788_),
    .Y(\datapath_1.ALUResult [13])
);

AND2X2 _11631_ (
    .A(_2744_),
    .B(_2396_),
    .Y(_2789_)
);

OAI21X1 _11632_ (
    .A(_2396_),
    .B(_2744_),
    .C(_2354__bF$buf1),
    .Y(_2790_)
);

OR2X2 _11633_ (
    .A(_2790_),
    .B(_2789_),
    .Y(_2791_)
);

OAI22X1 _11634_ (
    .A(_2199_),
    .B(_2365__bF$buf2),
    .C(_2198_),
    .D(_2486_),
    .Y(_2792_)
);

OAI22X1 _11635_ (
    .A(_2367__bF$buf3),
    .B(_2195_),
    .C(_2172_),
    .D(_2368__bF$buf1),
    .Y(_2793_)
);

NOR2X1 _11636_ (
    .A(_2793_),
    .B(_2792_),
    .Y(_2794_)
);

AOI21X1 _11637_ (
    .A(_2758_),
    .B(_2396_),
    .C(_2467_),
    .Y(_2795_)
);

OAI21X1 _11638_ (
    .A(_2396_),
    .B(_2758_),
    .C(_2795_),
    .Y(_2796_)
);

NAND3X1 _11639_ (
    .A(_2794_),
    .B(_2796_),
    .C(_2791_),
    .Y(\datapath_1.ALUResult [12])
);

AOI21X1 _11640_ (
    .A(_2145_),
    .B(_2159_),
    .C(_2180_),
    .Y(_2797_)
);

OAI21X1 _11641_ (
    .A(_2213_),
    .B(_2797_),
    .C(_2406_),
    .Y(_2798_)
);

OAI21X1 _11642_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2215_),
    .C(_2798_),
    .Y(_2799_)
);

OAI21X1 _11643_ (
    .A(_2201_),
    .B(_2202_),
    .C(_2799_),
    .Y(_2800_)
);

NOR2X1 _11644_ (
    .A(_2183_),
    .B(_2799_),
    .Y(_2801_)
);

NOR2X1 _11645_ (
    .A(_2353_),
    .B(_2801_),
    .Y(_2802_)
);

OAI22X1 _11646_ (
    .A(_2183_),
    .B(_2365__bF$buf1),
    .C(_2182_),
    .D(_2486_),
    .Y(_2803_)
);

OAI22X1 _11647_ (
    .A(_2367__bF$buf2),
    .B(_2181_),
    .C(_2202_),
    .D(_2368__bF$buf0),
    .Y(_2804_)
);

NOR2X1 _11648_ (
    .A(_2804_),
    .B(_2803_),
    .Y(_2805_)
);

INVX1 _11649_ (
    .A(_2402_),
    .Y(_2806_)
);

OAI21X1 _11650_ (
    .A(_2806_),
    .B(_2394_),
    .C(_2411_),
    .Y(_2807_)
);

AOI21X1 _11651_ (
    .A(_2807_),
    .B(_2204_),
    .C(_2184_),
    .Y(_2808_)
);

AND2X2 _11652_ (
    .A(_2808_),
    .B(_2183_),
    .Y(_2809_)
);

OAI21X1 _11653_ (
    .A(_2183_),
    .B(_2808_),
    .C(_2477__bF$buf1),
    .Y(_2810_)
);

OAI21X1 _11654_ (
    .A(_2809_),
    .B(_2810_),
    .C(_2805_),
    .Y(_2811_)
);

AOI21X1 _11655_ (
    .A(_2802_),
    .B(_2800_),
    .C(_2811_),
    .Y(_2812_)
);

INVX1 _11656_ (
    .A(_2812_),
    .Y(\datapath_1.ALUResult [11])
);

NOR2X1 _11657_ (
    .A(_2213_),
    .B(_2797_),
    .Y(_2813_)
);

NAND2X1 _11658_ (
    .A(_2204_),
    .B(_2813_),
    .Y(_2814_)
);

NAND3X1 _11659_ (
    .A(_2798_),
    .B(_2354__bF$buf0),
    .C(_2814_),
    .Y(_2815_)
);

AOI22X1 _11660_ (
    .A(_2184_),
    .B(_2487_),
    .C(_2185_),
    .D(_2362__bF$buf3),
    .Y(_2816_)
);

OAI21X1 _11661_ (
    .A(_2406_),
    .B(_2365__bF$buf0),
    .C(_2816_),
    .Y(_2817_)
);

AOI21X1 _11662_ (
    .A(_2405_),
    .B(_2637_),
    .C(_2817_),
    .Y(_2818_)
);

AOI21X1 _11663_ (
    .A(_2807_),
    .B(_2204_),
    .C(_2467_),
    .Y(_2819_)
);

OAI21X1 _11664_ (
    .A(_2204_),
    .B(_2807_),
    .C(_2819_),
    .Y(_2820_)
);

NAND3X1 _11665_ (
    .A(_2818_),
    .B(_2820_),
    .C(_2815_),
    .Y(\datapath_1.ALUResult [10])
);

OAI21X1 _11666_ (
    .A(_2179_),
    .B(_2394_),
    .C(_2399_),
    .Y(_2821_)
);

AND2X2 _11667_ (
    .A(_2821_),
    .B(_2208_),
    .Y(_2822_)
);

OAI21X1 _11668_ (
    .A(_2208_),
    .B(_2821_),
    .C(_2477__bF$buf0),
    .Y(_2823_)
);

OAI22X1 _11669_ (
    .A(_2367__bF$buf1),
    .B(_2175_),
    .C(_2176_),
    .D(_2486_),
    .Y(_2824_)
);

AOI21X1 _11670_ (
    .A(_2208_),
    .B(_2484_),
    .C(_2824_),
    .Y(_2825_)
);

OAI21X1 _11671_ (
    .A(_2207_),
    .B(_2368__bF$buf3),
    .C(_2825_),
    .Y(_2826_)
);

NOR2X1 _11672_ (
    .A(_2179_),
    .B(_2178_),
    .Y(_2827_)
);

NOR2X1 _11673_ (
    .A(_2519_),
    .B(_2177_),
    .Y(_2828_)
);

OAI21X1 _11674_ (
    .A(_2827_),
    .B(_2517_),
    .C(_2828_),
    .Y(_2829_)
);

OAI21X1 _11675_ (
    .A(_2208_),
    .B(_2212_),
    .C(_2354__bF$buf3),
    .Y(_2830_)
);

NOR2X1 _11676_ (
    .A(_2830_),
    .B(_2797_),
    .Y(_2831_)
);

AOI21X1 _11677_ (
    .A(_2829_),
    .B(_2831_),
    .C(_2826_),
    .Y(_2832_)
);

OAI21X1 _11678_ (
    .A(_2822_),
    .B(_2823_),
    .C(_2832_),
    .Y(\datapath_1.ALUResult [9])
);

OAI21X1 _11679_ (
    .A(_2827_),
    .B(_2517_),
    .C(_2354__bF$buf2),
    .Y(_2833_)
);

AOI21X1 _11680_ (
    .A(_2517_),
    .B(_2827_),
    .C(_2833_),
    .Y(_2834_)
);

OAI22X1 _11681_ (
    .A(_2367__bF$buf0),
    .B(_2399_),
    .C(_2400_),
    .D(_2486_),
    .Y(_2835_)
);

OAI21X1 _11682_ (
    .A(_2178_),
    .B(_2365__bF$buf4),
    .C(_2368__bF$buf2),
    .Y(_2836_)
);

AOI21X1 _11683_ (
    .A(_2836_),
    .B(_2400_),
    .C(_2835_),
    .Y(_2837_)
);

AND2X2 _11684_ (
    .A(_2394_),
    .B(_2401_),
    .Y(_2838_)
);

OAI21X1 _11685_ (
    .A(_2401_),
    .B(_2394_),
    .C(_2477__bF$buf3),
    .Y(_2839_)
);

OAI21X1 _11686_ (
    .A(_2838_),
    .B(_2839_),
    .C(_2837_),
    .Y(_2840_)
);

NOR2X1 _11687_ (
    .A(_2840_),
    .B(_2834_),
    .Y(_2841_)
);

INVX1 _11688_ (
    .A(_2841_),
    .Y(\datapath_1.ALUResult [8])
);

AOI21X1 _11689_ (
    .A(_2505_),
    .B(_2498_),
    .C(_2143_),
    .Y(_2842_)
);

OAI21X1 _11690_ (
    .A(_2153_),
    .B(_2842_),
    .C(_2552_),
    .Y(_2843_)
);

OAI21X1 _11691_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(_2155_),
    .C(_2843_),
    .Y(_2844_)
);

AOI21X1 _11692_ (
    .A(_2844_),
    .B(_2513_),
    .C(_2353_),
    .Y(_2845_)
);

OAI21X1 _11693_ (
    .A(_2513_),
    .B(_2844_),
    .C(_2845_),
    .Y(_2846_)
);

AOI22X1 _11694_ (
    .A(_2134_),
    .B(_2487_),
    .C(_2135_),
    .D(_2362__bF$buf2),
    .Y(_2847_)
);

OAI21X1 _11695_ (
    .A(_2513_),
    .B(_2365__bF$buf3),
    .C(_2847_),
    .Y(_2848_)
);

AOI21X1 _11696_ (
    .A(_2391_),
    .B(_2637_),
    .C(_2848_),
    .Y(_2849_)
);

AOI21X1 _11697_ (
    .A(_2380_),
    .B(_2556_),
    .C(_2389_),
    .Y(_2850_)
);

OAI21X1 _11698_ (
    .A(_2137_),
    .B(_2850_),
    .C(_2550_),
    .Y(_2851_)
);

AOI21X1 _11699_ (
    .A(_2851_),
    .B(_2381_),
    .C(_2467_),
    .Y(_2852_)
);

OAI21X1 _11700_ (
    .A(_2381_),
    .B(_2851_),
    .C(_2852_),
    .Y(_2853_)
);

NAND3X1 _11701_ (
    .A(_2849_),
    .B(_2853_),
    .C(_2846_),
    .Y(\datapath_1.ALUResult [7])
);

AOI21X1 _11702_ (
    .A(_2505_),
    .B(_2498_),
    .C(_2384_),
    .Y(_2854_)
);

OAI21X1 _11703_ (
    .A(_2510_),
    .B(_2854_),
    .C(_2509_),
    .Y(_2855_)
);

NAND3X1 _11704_ (
    .A(_2150_),
    .B(_2382_),
    .C(_2855_),
    .Y(_2856_)
);

NAND3X1 _11705_ (
    .A(_2843_),
    .B(_2354__bF$buf1),
    .C(_2856_),
    .Y(_2857_)
);

AOI22X1 _11706_ (
    .A(_2362__bF$buf1),
    .B(_2137_),
    .C(_2136_),
    .D(_2487_),
    .Y(_2858_)
);

OAI21X1 _11707_ (
    .A(_2552_),
    .B(_2365__bF$buf2),
    .C(_2858_),
    .Y(_2859_)
);

AOI21X1 _11708_ (
    .A(_2551_),
    .B(_2637_),
    .C(_2859_),
    .Y(_2860_)
);

AND2X2 _11709_ (
    .A(_2850_),
    .B(_2552_),
    .Y(_2861_)
);

OAI21X1 _11710_ (
    .A(_2552_),
    .B(_2850_),
    .C(_2477__bF$buf2),
    .Y(_2862_)
);

OR2X2 _11711_ (
    .A(_2862_),
    .B(_2861_),
    .Y(_2863_)
);

NAND3X1 _11712_ (
    .A(_2860_),
    .B(_2863_),
    .C(_2857_),
    .Y(\datapath_1.ALUResult [6])
);

OAI21X1 _11713_ (
    .A(_2122_),
    .B(_2133_),
    .C(_2555_),
    .Y(_2864_)
);

NAND3X1 _11714_ (
    .A(_2152_),
    .B(_2147_),
    .C(_2864_),
    .Y(_2865_)
);

NAND3X1 _11715_ (
    .A(_2354__bF$buf0),
    .B(_2865_),
    .C(_2855_),
    .Y(_2866_)
);

AOI22X1 _11716_ (
    .A(_2139_),
    .B(_2487_),
    .C(_2140_),
    .D(_2362__bF$buf0),
    .Y(_2867_)
);

OAI21X1 _11717_ (
    .A(_2509_),
    .B(_2365__bF$buf1),
    .C(_2867_),
    .Y(_2868_)
);

AOI21X1 _11718_ (
    .A(_2508_),
    .B(_2637_),
    .C(_2868_),
    .Y(_2869_)
);

AOI21X1 _11719_ (
    .A(_2377_),
    .B(_2379_),
    .C(_2555_),
    .Y(_2870_)
);

INVX1 _11720_ (
    .A(_2870_),
    .Y(_2871_)
);

NAND3X1 _11721_ (
    .A(_2388_),
    .B(_2509_),
    .C(_2871_),
    .Y(_2872_)
);

OAI21X1 _11722_ (
    .A(_2141_),
    .B(_2870_),
    .C(_2147_),
    .Y(_2873_)
);

NAND3X1 _11723_ (
    .A(_2477__bF$buf1),
    .B(_2873_),
    .C(_2872_),
    .Y(_2874_)
);

NAND3X1 _11724_ (
    .A(_2869_),
    .B(_2866_),
    .C(_2874_),
    .Y(\datapath_1.ALUResult [5])
);

NAND3X1 _11725_ (
    .A(_2498_),
    .B(_2384_),
    .C(_2505_),
    .Y(_2875_)
);

NAND3X1 _11726_ (
    .A(_2354__bF$buf3),
    .B(_2864_),
    .C(_2875_),
    .Y(_2876_)
);

AOI22X1 _11727_ (
    .A(_2141_),
    .B(_2487_),
    .C(_2142_),
    .D(_2362__bF$buf3),
    .Y(_2877_)
);

OAI21X1 _11728_ (
    .A(_2555_),
    .B(_2365__bF$buf0),
    .C(_2877_),
    .Y(_2878_)
);

AOI21X1 _11729_ (
    .A(_2554_),
    .B(_2637_),
    .C(_2878_),
    .Y(_2879_)
);

NOR2X1 _11730_ (
    .A(_2467_),
    .B(_2870_),
    .Y(_2880_)
);

OAI21X1 _11731_ (
    .A(_2384_),
    .B(_2380_),
    .C(_2880_),
    .Y(_2881_)
);

NAND3X1 _11732_ (
    .A(_2879_),
    .B(_2876_),
    .C(_2881_),
    .Y(\datapath_1.ALUResult [4])
);

AOI21X1 _11733_ (
    .A(_2125_),
    .B(_2129_),
    .C(_2372_),
    .Y(_2882_)
);

NOR2X1 _11734_ (
    .A(_2118_),
    .B(_2882_),
    .Y(_2883_)
);

NAND2X1 _11735_ (
    .A(_2373_),
    .B(_2883_),
    .Y(_2884_)
);

OAI21X1 _11736_ (
    .A(_2118_),
    .B(_2882_),
    .C(_2497_),
    .Y(_2885_)
);

NAND3X1 _11737_ (
    .A(_2354__bF$buf2),
    .B(_2885_),
    .C(_2884_),
    .Y(_2886_)
);

AOI22X1 _11738_ (
    .A(_2119_),
    .B(_2487_),
    .C(_2120_),
    .D(_2362__bF$buf2),
    .Y(_2887_)
);

OAI21X1 _11739_ (
    .A(_2497_),
    .B(_2365__bF$buf4),
    .C(_2887_),
    .Y(_2888_)
);

AOI21X1 _11740_ (
    .A(_2378_),
    .B(_2637_),
    .C(_2888_),
    .Y(_2889_)
);

NAND2X1 _11741_ (
    .A(_2372_),
    .B(_2376_),
    .Y(_2890_)
);

AOI21X1 _11742_ (
    .A(_2890_),
    .B(_2502_),
    .C(_2497_),
    .Y(_2891_)
);

NAND2X1 _11743_ (
    .A(_2502_),
    .B(_2890_),
    .Y(_2892_)
);

OAI21X1 _11744_ (
    .A(_2373_),
    .B(_2892_),
    .C(_2477__bF$buf0),
    .Y(_2893_)
);

OR2X2 _11745_ (
    .A(_2893_),
    .B(_2891_),
    .Y(_2894_)
);

NAND3X1 _11746_ (
    .A(_2889_),
    .B(_2894_),
    .C(_2886_),
    .Y(\datapath_1.ALUResult [3])
);

INVX1 _11747_ (
    .A(_2882_),
    .Y(_2895_)
);

NAND3X1 _11748_ (
    .A(_2372_),
    .B(_2129_),
    .C(_2125_),
    .Y(_2896_)
);

NAND3X1 _11749_ (
    .A(_2354__bF$buf1),
    .B(_2896_),
    .C(_2895_),
    .Y(_2897_)
);

AOI22X1 _11750_ (
    .A(_2484_),
    .B(_2372_),
    .C(_2131_),
    .D(_2362__bF$buf1),
    .Y(_2898_)
);

AOI22X1 _11751_ (
    .A(_2487_),
    .B(_2130_),
    .C(_2637_),
    .D(_2503_),
    .Y(_2899_)
);

AND2X2 _11752_ (
    .A(_2898_),
    .B(_2899_),
    .Y(_2900_)
);

AOI21X1 _11753_ (
    .A(_2372_),
    .B(_2376_),
    .C(_2467_),
    .Y(_2901_)
);

OAI21X1 _11754_ (
    .A(_2372_),
    .B(_2376_),
    .C(_2901_),
    .Y(_2902_)
);

NAND3X1 _11755_ (
    .A(_2902_),
    .B(_2900_),
    .C(_2897_),
    .Y(\datapath_1.ALUResult [2])
);

NOR2X1 _11756_ (
    .A(_2128_),
    .B(_2127_),
    .Y(_2903_)
);

AOI22X1 _11757_ (
    .A(_2484_),
    .B(_2903_),
    .C(_2128_),
    .D(_2362__bF$buf0),
    .Y(_2904_)
);

AOI22X1 _11758_ (
    .A(_2487_),
    .B(_2127_),
    .C(_2637_),
    .D(_2500_),
    .Y(_2905_)
);

AND2X2 _11759_ (
    .A(_2904_),
    .B(_2905_),
    .Y(_2906_)
);

XNOR2X1 _11760_ (
    .A(_2903_),
    .B(_2375_),
    .Y(_2907_)
);

NOR2X1 _11761_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .B(_2126_),
    .Y(_2908_)
);

AOI21X1 _11762_ (
    .A(_2903_),
    .B(_2908_),
    .C(_2353_),
    .Y(_2909_)
);

AOI22X1 _11763_ (
    .A(_2129_),
    .B(_2909_),
    .C(_2477__bF$buf3),
    .D(_2907_),
    .Y(_2910_)
);

NAND2X1 _11764_ (
    .A(_2910_),
    .B(_2906_),
    .Y(\datapath_1.ALUResult [1])
);

INVX1 _11765_ (
    .A(gnd),
    .Y(_2911_)
);

NAND2X1 _11766_ (
    .A(_2911_),
    .B(_2350_),
    .Y(_2912_)
);

NOR2X1 _11767_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(_2499_),
    .Y(_2913_)
);

NOR2X1 _11768_ (
    .A(_2913_),
    .B(_2908_),
    .Y(_2914_)
);

AOI21X1 _11769_ (
    .A(_2912_),
    .B(_2365__bF$buf3),
    .C(_2914_),
    .Y(_2915_)
);

AOI21X1 _11770_ (
    .A(_2126_),
    .B(_2499_),
    .C(_2368__bF$buf1),
    .Y(_2916_)
);

NAND2X1 _11771_ (
    .A(_2126_),
    .B(_2499_),
    .Y(_2917_)
);

OAI22X1 _11772_ (
    .A(_2375_),
    .B(_2367__bF$buf3),
    .C(_2917_),
    .D(_2486_),
    .Y(_2918_)
);

NOR3X1 _11773_ (
    .A(_2916_),
    .B(_2918_),
    .C(_2915_),
    .Y(_2919_)
);

INVX1 _11774_ (
    .A(_2919_),
    .Y(\datapath_1.ALUResult [0])
);

INVX1 _11775_ (
    .A(\datapath_1.ALUResult [12]),
    .Y(_2920_)
);

INVX1 _11776_ (
    .A(\datapath_1.ALUResult [5]),
    .Y(_2921_)
);

NAND3X1 _11777_ (
    .A(_2910_),
    .B(_2906_),
    .C(_2919_),
    .Y(_2922_)
);

OR2X2 _11778_ (
    .A(_2922_),
    .B(\datapath_1.ALUResult [2]),
    .Y(_2923_)
);

NOR3X1 _11779_ (
    .A(\datapath_1.ALUResult [3]),
    .B(\datapath_1.ALUResult [4]),
    .C(_2923_),
    .Y(_2924_)
);

NAND3X1 _11780_ (
    .A(_2921_),
    .B(_2841_),
    .C(_2924_),
    .Y(_2925_)
);

NOR2X1 _11781_ (
    .A(\datapath_1.ALUResult [9]),
    .B(_2925_),
    .Y(_2926_)
);

NAND3X1 _11782_ (
    .A(_2732_),
    .B(_2920_),
    .C(_2926_),
    .Y(_2927_)
);

NAND3X1 _11783_ (
    .A(_2675_),
    .B(_2774_),
    .C(_2663_),
    .Y(_2928_)
);

NOR3X1 _11784_ (
    .A(\datapath_1.ALUResult [25]),
    .B(_2927_),
    .C(_2928_),
    .Y(_2929_)
);

INVX1 _11785_ (
    .A(\datapath_1.ALUResult [7]),
    .Y(_2930_)
);

NAND3X1 _11786_ (
    .A(_2930_),
    .B(_2788_),
    .C(_2812_),
    .Y(_2931_)
);

NAND2X1 _11787_ (
    .A(_2720_),
    .B(_2685_),
    .Y(_2932_)
);

NOR3X1 _11788_ (
    .A(\datapath_1.ALUResult [6]),
    .B(\datapath_1.ALUResult [16]),
    .C(\datapath_1.ALUResult [10]),
    .Y(_2933_)
);

NAND3X1 _11789_ (
    .A(_2612_),
    .B(_2619_),
    .C(_2933_),
    .Y(_2934_)
);

NOR3X1 _11790_ (
    .A(_2932_),
    .B(_2934_),
    .C(_2931_),
    .Y(_2935_)
);

NOR2X1 _11791_ (
    .A(\datapath_1.ALUResult [15]),
    .B(\datapath_1.ALUResult [29]),
    .Y(_2936_)
);

NAND3X1 _11792_ (
    .A(_2929_),
    .B(_2935_),
    .C(_2936_),
    .Y(_2937_)
);

NOR2X1 _11793_ (
    .A(\datapath_1.ALUResult [26]),
    .B(\datapath_1.ALUResult [28]),
    .Y(_2938_)
);

NOR2X1 _11794_ (
    .A(\datapath_1.ALUResult [19]),
    .B(\datapath_1.ALUResult [22]),
    .Y(_2939_)
);

AND2X2 _11795_ (
    .A(_2938_),
    .B(_2939_),
    .Y(_2940_)
);

NOR2X1 _11796_ (
    .A(\datapath_1.ALUResult [23]),
    .B(\datapath_1.ALUResult [27]),
    .Y(_2941_)
);

NAND3X1 _11797_ (
    .A(_2480_),
    .B(_2940_),
    .C(_2941_),
    .Y(_2942_)
);

NOR3X1 _11798_ (
    .A(_2937_),
    .B(\datapath_1.ALUResult [31]),
    .C(_2942_),
    .Y(ALUZero)
);

INVX1 _11799_ (
    .A(\datapath_1.PCJump [18]),
    .Y(_2943_)
);

NAND2X1 _11800_ (
    .A(\datapath_1.PCJump [13]),
    .B(RegDst),
    .Y(_2944_)
);

OAI21X1 _11801_ (
    .A(RegDst),
    .B(_2943_),
    .C(_2944_),
    .Y(\datapath_1.a3 [0])
);

INVX1 _11802_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_2945_)
);

NAND2X1 _11803_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [14]),
    .Y(_2946_)
);

OAI21X1 _11804_ (
    .A(RegDst),
    .B(_2945_),
    .C(_2946_),
    .Y(\datapath_1.a3 [1])
);

INVX1 _11805_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_2947_)
);

NAND2X1 _11806_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [15]),
    .Y(_2948_)
);

OAI21X1 _11807_ (
    .A(RegDst),
    .B(_2947_),
    .C(_2948_),
    .Y(\datapath_1.a3 [2])
);

INVX1 _11808_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_2949_)
);

NAND2X1 _11809_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [16]),
    .Y(_2950_)
);

OAI21X1 _11810_ (
    .A(RegDst),
    .B(_2949_),
    .C(_2950_),
    .Y(\datapath_1.a3 [3])
);

INVX1 _11811_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_2951_)
);

NAND2X1 _11812_ (
    .A(RegDst),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_2952_)
);

OAI21X1 _11813_ (
    .A(RegDst),
    .B(_2951_),
    .C(_2952_),
    .Y(\datapath_1.a3 [4])
);

INVX1 _11814_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3015_)
);

NAND2X1 _11815_ (
    .A(ALUOut[0]),
    .B(IorD_bF$buf7),
    .Y(_3016_)
);

OAI21X1 _11816_ (
    .A(IorD_bF$buf6),
    .B(_3015_),
    .C(_3016_),
    .Y(_1_[0])
);

INVX1 _11817_ (
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_2953_)
);

NAND2X1 _11818_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[1]),
    .Y(_2954_)
);

OAI21X1 _11819_ (
    .A(IorD_bF$buf4),
    .B(_2953_),
    .C(_2954_),
    .Y(_1_[1])
);

INVX1 _11820_ (
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_2955_)
);

NAND2X1 _11821_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[2]),
    .Y(_2956_)
);

OAI21X1 _11822_ (
    .A(IorD_bF$buf2),
    .B(_2955_),
    .C(_2956_),
    .Y(_1_[2])
);

INVX1 _11823_ (
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_2957_)
);

NAND2X1 _11824_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[3]),
    .Y(_2958_)
);

OAI21X1 _11825_ (
    .A(IorD_bF$buf0),
    .B(_2957_),
    .C(_2958_),
    .Y(_1_[3])
);

INVX1 _11826_ (
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_2959_)
);

NAND2X1 _11827_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[4]),
    .Y(_2960_)
);

OAI21X1 _11828_ (
    .A(IorD_bF$buf6),
    .B(_2959_),
    .C(_2960_),
    .Y(_1_[4])
);

INVX1 _11829_ (
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_2961_)
);

NAND2X1 _11830_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[5]),
    .Y(_2962_)
);

OAI21X1 _11831_ (
    .A(IorD_bF$buf4),
    .B(_2961_),
    .C(_2962_),
    .Y(_1_[5])
);

INVX1 _11832_ (
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_2963_)
);

NAND2X1 _11833_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[6]),
    .Y(_2964_)
);

OAI21X1 _11834_ (
    .A(IorD_bF$buf2),
    .B(_2963_),
    .C(_2964_),
    .Y(_1_[6])
);

INVX1 _11835_ (
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_2965_)
);

NAND2X1 _11836_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[7]),
    .Y(_2966_)
);

OAI21X1 _11837_ (
    .A(IorD_bF$buf0),
    .B(_2965_),
    .C(_2966_),
    .Y(_1_[7])
);

INVX1 _11838_ (
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_2967_)
);

NAND2X1 _11839_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[8]),
    .Y(_2968_)
);

OAI21X1 _11840_ (
    .A(IorD_bF$buf6),
    .B(_2967_),
    .C(_2968_),
    .Y(_1_[8])
);

INVX1 _11841_ (
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_2969_)
);

NAND2X1 _11842_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[9]),
    .Y(_2970_)
);

OAI21X1 _11843_ (
    .A(IorD_bF$buf4),
    .B(_2969_),
    .C(_2970_),
    .Y(_1_[9])
);

INVX1 _11844_ (
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_2971_)
);

NAND2X1 _11845_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[10]),
    .Y(_2972_)
);

OAI21X1 _11846_ (
    .A(IorD_bF$buf2),
    .B(_2971_),
    .C(_2972_),
    .Y(_1_[10])
);

INVX1 _11847_ (
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_2973_)
);

NAND2X1 _11848_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[11]),
    .Y(_2974_)
);

OAI21X1 _11849_ (
    .A(IorD_bF$buf0),
    .B(_2973_),
    .C(_2974_),
    .Y(_1_[11])
);

INVX1 _11850_ (
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_2975_)
);

NAND2X1 _11851_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[12]),
    .Y(_2976_)
);

OAI21X1 _11852_ (
    .A(IorD_bF$buf6),
    .B(_2975_),
    .C(_2976_),
    .Y(_1_[12])
);

INVX1 _11853_ (
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_2977_)
);

NAND2X1 _11854_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[13]),
    .Y(_2978_)
);

OAI21X1 _11855_ (
    .A(IorD_bF$buf4),
    .B(_2977_),
    .C(_2978_),
    .Y(_1_[13])
);

INVX1 _11856_ (
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_2979_)
);

NAND2X1 _11857_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[14]),
    .Y(_2980_)
);

OAI21X1 _11858_ (
    .A(IorD_bF$buf2),
    .B(_2979_),
    .C(_2980_),
    .Y(_1_[14])
);

INVX1 _11859_ (
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_2981_)
);

NAND2X1 _11860_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[15]),
    .Y(_2982_)
);

OAI21X1 _11861_ (
    .A(IorD_bF$buf0),
    .B(_2981_),
    .C(_2982_),
    .Y(_1_[15])
);

INVX1 _11862_ (
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_2983_)
);

NAND2X1 _11863_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[16]),
    .Y(_2984_)
);

OAI21X1 _11864_ (
    .A(IorD_bF$buf6),
    .B(_2983_),
    .C(_2984_),
    .Y(_1_[16])
);

INVX1 _11865_ (
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_2985_)
);

NAND2X1 _11866_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[17]),
    .Y(_2986_)
);

OAI21X1 _11867_ (
    .A(IorD_bF$buf4),
    .B(_2985_),
    .C(_2986_),
    .Y(_1_[17])
);

INVX1 _11868_ (
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_2987_)
);

NAND2X1 _11869_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[18]),
    .Y(_2988_)
);

OAI21X1 _11870_ (
    .A(IorD_bF$buf2),
    .B(_2987_),
    .C(_2988_),
    .Y(_1_[18])
);

INVX1 _11871_ (
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_2989_)
);

NAND2X1 _11872_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[19]),
    .Y(_2990_)
);

OAI21X1 _11873_ (
    .A(IorD_bF$buf0),
    .B(_2989_),
    .C(_2990_),
    .Y(_1_[19])
);

INVX1 _11874_ (
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_2991_)
);

NAND2X1 _11875_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[20]),
    .Y(_2992_)
);

OAI21X1 _11876_ (
    .A(IorD_bF$buf6),
    .B(_2991_),
    .C(_2992_),
    .Y(_1_[20])
);

INVX1 _11877_ (
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_2993_)
);

NAND2X1 _11878_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[21]),
    .Y(_2994_)
);

OAI21X1 _11879_ (
    .A(IorD_bF$buf4),
    .B(_2993_),
    .C(_2994_),
    .Y(_1_[21])
);

INVX1 _11880_ (
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_2995_)
);

NAND2X1 _11881_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[22]),
    .Y(_2996_)
);

OAI21X1 _11882_ (
    .A(IorD_bF$buf2),
    .B(_2995_),
    .C(_2996_),
    .Y(_1_[22])
);

INVX1 _11883_ (
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_2997_)
);

NAND2X1 _11884_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[23]),
    .Y(_2998_)
);

OAI21X1 _11885_ (
    .A(IorD_bF$buf0),
    .B(_2997_),
    .C(_2998_),
    .Y(_1_[23])
);

INVX1 _11886_ (
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_2999_)
);

NAND2X1 _11887_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[24]),
    .Y(_3000_)
);

OAI21X1 _11888_ (
    .A(IorD_bF$buf6),
    .B(_2999_),
    .C(_3000_),
    .Y(_1_[24])
);

INVX1 _11889_ (
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3001_)
);

NAND2X1 _11890_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[25]),
    .Y(_3002_)
);

OAI21X1 _11891_ (
    .A(IorD_bF$buf4),
    .B(_3001_),
    .C(_3002_),
    .Y(_1_[25])
);

INVX1 _11892_ (
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3003_)
);

NAND2X1 _11893_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[26]),
    .Y(_3004_)
);

OAI21X1 _11894_ (
    .A(IorD_bF$buf2),
    .B(_3003_),
    .C(_3004_),
    .Y(_1_[26])
);

INVX1 _11895_ (
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3005_)
);

NAND2X1 _11896_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[27]),
    .Y(_3006_)
);

OAI21X1 _11897_ (
    .A(IorD_bF$buf0),
    .B(_3005_),
    .C(_3006_),
    .Y(_1_[27])
);

INVX1 _11898_ (
    .A(\datapath_1.PCJump [28]),
    .Y(_3007_)
);

NAND2X1 _11899_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[28]),
    .Y(_3008_)
);

OAI21X1 _11900_ (
    .A(IorD_bF$buf6),
    .B(_3007_),
    .C(_3008_),
    .Y(_1_[28])
);

INVX1 _11901_ (
    .A(\datapath_1.PCJump [29]),
    .Y(_3009_)
);

NAND2X1 _11902_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[29]),
    .Y(_3010_)
);

OAI21X1 _11903_ (
    .A(IorD_bF$buf4),
    .B(_3009_),
    .C(_3010_),
    .Y(_1_[29])
);

INVX1 _11904_ (
    .A(\datapath_1.PCJump [30]),
    .Y(_3011_)
);

NAND2X1 _11905_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[30]),
    .Y(_3012_)
);

OAI21X1 _11906_ (
    .A(IorD_bF$buf2),
    .B(_3011_),
    .C(_3012_),
    .Y(_1_[30])
);

INVX1 _11907_ (
    .A(\datapath_1.PCJump [31]),
    .Y(_3013_)
);

NAND2X1 _11908_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[31]),
    .Y(_3014_)
);

OAI21X1 _11909_ (
    .A(IorD_bF$buf0),
    .B(_3013_),
    .C(_3014_),
    .Y(_1_[31])
);

INVX8 _11910_ (
    .A(PCSource_1_bF$buf4),
    .Y(_3017_)
);

NAND3X1 _11911_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[0]),
    .C(_3017__bF$buf4),
    .Y(_3018_)
);

INVX8 _11912_ (
    .A(ALUOp_0_bF$buf2),
    .Y(_3019_)
);

NAND3X1 _11913_ (
    .A(PCSource_1_bF$buf3),
    .B(gnd),
    .C(_3019__bF$buf4),
    .Y(_3020_)
);

NOR2X1 _11914_ (
    .A(ALUOp_0_bF$buf1),
    .B(PCSource_1_bF$buf2),
    .Y(_3021_)
);

AND2X2 _11915_ (
    .A(PCSource_1_bF$buf1),
    .B(ALUOp_0_bF$buf0),
    .Y(_3022_)
);

AOI22X1 _11916_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [0]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3023_)
);

NAND3X1 _11917_ (
    .A(_3020_),
    .B(_3018_),
    .C(_3023_),
    .Y(\datapath_1.mux_pcsrc.dout [0])
);

NAND3X1 _11918_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[1]),
    .C(_3017__bF$buf3),
    .Y(_3024_)
);

NAND3X1 _11919_ (
    .A(PCSource_1_bF$buf0),
    .B(gnd),
    .C(_3019__bF$buf3),
    .Y(_3025_)
);

AOI22X1 _11920_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [1]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3026_)
);

NAND3X1 _11921_ (
    .A(_3025_),
    .B(_3024_),
    .C(_3026_),
    .Y(\datapath_1.mux_pcsrc.dout [1])
);

NAND3X1 _11922_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[2]),
    .C(_3017__bF$buf2),
    .Y(_3027_)
);

NAND3X1 _11923_ (
    .A(PCSource_1_bF$buf4),
    .B(\aluControl_1.inst [0]),
    .C(_3019__bF$buf2),
    .Y(_3028_)
);

AOI22X1 _11924_ (
    .A(_3021__bF$buf2),
    .B(\datapath_1.ALUResult [2]),
    .C(gnd),
    .D(_3022__bF$buf2),
    .Y(_3029_)
);

NAND3X1 _11925_ (
    .A(_3028_),
    .B(_3027_),
    .C(_3029_),
    .Y(\datapath_1.mux_pcsrc.dout [2])
);

NAND3X1 _11926_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[3]),
    .C(_3017__bF$buf1),
    .Y(_3030_)
);

NAND3X1 _11927_ (
    .A(PCSource_1_bF$buf3),
    .B(\aluControl_1.inst [1]),
    .C(_3019__bF$buf1),
    .Y(_3031_)
);

AOI22X1 _11928_ (
    .A(_3021__bF$buf1),
    .B(\datapath_1.ALUResult [3]),
    .C(gnd),
    .D(_3022__bF$buf1),
    .Y(_3032_)
);

NAND3X1 _11929_ (
    .A(_3031_),
    .B(_3030_),
    .C(_3032_),
    .Y(\datapath_1.mux_pcsrc.dout [3])
);

NAND3X1 _11930_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[4]),
    .C(_3017__bF$buf0),
    .Y(_3033_)
);

NAND3X1 _11931_ (
    .A(PCSource_1_bF$buf2),
    .B(\aluControl_1.inst [2]),
    .C(_3019__bF$buf0),
    .Y(_3034_)
);

AOI22X1 _11932_ (
    .A(_3021__bF$buf0),
    .B(\datapath_1.ALUResult [4]),
    .C(gnd),
    .D(_3022__bF$buf0),
    .Y(_3035_)
);

NAND3X1 _11933_ (
    .A(_3034_),
    .B(_3033_),
    .C(_3035_),
    .Y(\datapath_1.mux_pcsrc.dout [4])
);

NAND3X1 _11934_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[5]),
    .C(_3017__bF$buf4),
    .Y(_3036_)
);

NAND3X1 _11935_ (
    .A(PCSource_1_bF$buf1),
    .B(\aluControl_1.inst [3]),
    .C(_3019__bF$buf4),
    .Y(_3037_)
);

AOI22X1 _11936_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [5]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3038_)
);

NAND3X1 _11937_ (
    .A(_3037_),
    .B(_3036_),
    .C(_3038_),
    .Y(\datapath_1.mux_pcsrc.dout [5])
);

NAND3X1 _11938_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[6]),
    .C(_3017__bF$buf3),
    .Y(_3039_)
);

NAND3X1 _11939_ (
    .A(PCSource_1_bF$buf0),
    .B(\aluControl_1.inst [4]),
    .C(_3019__bF$buf3),
    .Y(_3040_)
);

AOI22X1 _11940_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [6]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3041_)
);

NAND3X1 _11941_ (
    .A(_3040_),
    .B(_3039_),
    .C(_3041_),
    .Y(\datapath_1.mux_pcsrc.dout [6])
);

NAND3X1 _11942_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[7]),
    .C(_3017__bF$buf2),
    .Y(_3042_)
);

NAND3X1 _11943_ (
    .A(PCSource_1_bF$buf4),
    .B(\aluControl_1.inst [5]),
    .C(_3019__bF$buf2),
    .Y(_3043_)
);

AOI22X1 _11944_ (
    .A(_3021__bF$buf2),
    .B(\datapath_1.ALUResult [7]),
    .C(gnd),
    .D(_3022__bF$buf2),
    .Y(_3044_)
);

NAND3X1 _11945_ (
    .A(_3043_),
    .B(_3042_),
    .C(_3044_),
    .Y(\datapath_1.mux_pcsrc.dout [7])
);

NAND3X1 _11946_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[8]),
    .C(_3017__bF$buf1),
    .Y(_3045_)
);

NAND3X1 _11947_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [8]),
    .C(_3019__bF$buf1),
    .Y(_3046_)
);

AOI22X1 _11948_ (
    .A(_3021__bF$buf1),
    .B(\datapath_1.ALUResult [8]),
    .C(gnd),
    .D(_3022__bF$buf1),
    .Y(_3047_)
);

NAND3X1 _11949_ (
    .A(_3046_),
    .B(_3045_),
    .C(_3047_),
    .Y(\datapath_1.mux_pcsrc.dout [8])
);

NAND3X1 _11950_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[9]),
    .C(_3017__bF$buf0),
    .Y(_3048_)
);

NAND3X1 _11951_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [9]),
    .C(_3019__bF$buf0),
    .Y(_3049_)
);

AOI22X1 _11952_ (
    .A(_3021__bF$buf0),
    .B(\datapath_1.ALUResult [9]),
    .C(gnd),
    .D(_3022__bF$buf0),
    .Y(_3050_)
);

NAND3X1 _11953_ (
    .A(_3049_),
    .B(_3048_),
    .C(_3050_),
    .Y(\datapath_1.mux_pcsrc.dout [9])
);

NAND3X1 _11954_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[10]),
    .C(_3017__bF$buf4),
    .Y(_3051_)
);

NAND3X1 _11955_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [10]),
    .C(_3019__bF$buf4),
    .Y(_3052_)
);

AOI22X1 _11956_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [10]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3053_)
);

NAND3X1 _11957_ (
    .A(_3052_),
    .B(_3051_),
    .C(_3053_),
    .Y(\datapath_1.mux_pcsrc.dout [10])
);

NAND3X1 _11958_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[11]),
    .C(_3017__bF$buf3),
    .Y(_3054_)
);

NAND3X1 _11959_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [11]),
    .C(_3019__bF$buf3),
    .Y(_3055_)
);

AOI22X1 _11960_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [11]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3056_)
);

NAND3X1 _11961_ (
    .A(_3055_),
    .B(_3054_),
    .C(_3056_),
    .Y(\datapath_1.mux_pcsrc.dout [11])
);

NAND3X1 _11962_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[12]),
    .C(_3017__bF$buf2),
    .Y(_3057_)
);

NAND3X1 _11963_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump [12]),
    .C(_3019__bF$buf2),
    .Y(_3058_)
);

AOI22X1 _11964_ (
    .A(_3021__bF$buf2),
    .B(\datapath_1.ALUResult [12]),
    .C(gnd),
    .D(_3022__bF$buf2),
    .Y(_3059_)
);

NAND3X1 _11965_ (
    .A(_3058_),
    .B(_3057_),
    .C(_3059_),
    .Y(\datapath_1.mux_pcsrc.dout [12])
);

NAND3X1 _11966_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[13]),
    .C(_3017__bF$buf1),
    .Y(_3060_)
);

NAND3X1 _11967_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [13]),
    .C(_3019__bF$buf1),
    .Y(_3061_)
);

AOI22X1 _11968_ (
    .A(_3021__bF$buf1),
    .B(\datapath_1.ALUResult [13]),
    .C(gnd),
    .D(_3022__bF$buf1),
    .Y(_3062_)
);

NAND3X1 _11969_ (
    .A(_3061_),
    .B(_3060_),
    .C(_3062_),
    .Y(\datapath_1.mux_pcsrc.dout [13])
);

NAND3X1 _11970_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[14]),
    .C(_3017__bF$buf0),
    .Y(_3063_)
);

NAND3X1 _11971_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [14]),
    .C(_3019__bF$buf0),
    .Y(_3064_)
);

AOI22X1 _11972_ (
    .A(_3021__bF$buf0),
    .B(\datapath_1.ALUResult [14]),
    .C(gnd),
    .D(_3022__bF$buf0),
    .Y(_3065_)
);

NAND3X1 _11973_ (
    .A(_3064_),
    .B(_3063_),
    .C(_3065_),
    .Y(\datapath_1.mux_pcsrc.dout [14])
);

NAND3X1 _11974_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[15]),
    .C(_3017__bF$buf4),
    .Y(_3066_)
);

NAND3X1 _11975_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [15]),
    .C(_3019__bF$buf4),
    .Y(_3067_)
);

AOI22X1 _11976_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [15]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3068_)
);

NAND3X1 _11977_ (
    .A(_3067_),
    .B(_3066_),
    .C(_3068_),
    .Y(\datapath_1.mux_pcsrc.dout [15])
);

NAND3X1 _11978_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[16]),
    .C(_3017__bF$buf3),
    .Y(_3069_)
);

NAND3X1 _11979_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [16]),
    .C(_3019__bF$buf3),
    .Y(_3070_)
);

AOI22X1 _11980_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [16]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3071_)
);

NAND3X1 _11981_ (
    .A(_3070_),
    .B(_3069_),
    .C(_3071_),
    .Y(\datapath_1.mux_pcsrc.dout [16])
);

NAND3X1 _11982_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[17]),
    .C(_3017__bF$buf2),
    .Y(_3072_)
);

NAND3X1 _11983_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3019__bF$buf2),
    .Y(_3073_)
);

AOI22X1 _11984_ (
    .A(_3021__bF$buf2),
    .B(\datapath_1.ALUResult [17]),
    .C(gnd),
    .D(_3022__bF$buf2),
    .Y(_3074_)
);

NAND3X1 _11985_ (
    .A(_3073_),
    .B(_3072_),
    .C(_3074_),
    .Y(\datapath_1.mux_pcsrc.dout [17])
);

NAND3X1 _11986_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[18]),
    .C(_3017__bF$buf1),
    .Y(_3075_)
);

NAND3X1 _11987_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [18]),
    .C(_3019__bF$buf1),
    .Y(_3076_)
);

AOI22X1 _11988_ (
    .A(_3021__bF$buf1),
    .B(\datapath_1.ALUResult [18]),
    .C(gnd),
    .D(_3022__bF$buf1),
    .Y(_3077_)
);

NAND3X1 _11989_ (
    .A(_3076_),
    .B(_3075_),
    .C(_3077_),
    .Y(\datapath_1.mux_pcsrc.dout [18])
);

NAND3X1 _11990_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[19]),
    .C(_3017__bF$buf0),
    .Y(_3078_)
);

NAND3X1 _11991_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [19]),
    .C(_3019__bF$buf0),
    .Y(_3079_)
);

AOI22X1 _11992_ (
    .A(_3021__bF$buf0),
    .B(\datapath_1.ALUResult [19]),
    .C(gnd),
    .D(_3022__bF$buf0),
    .Y(_3080_)
);

NAND3X1 _11993_ (
    .A(_3079_),
    .B(_3078_),
    .C(_3080_),
    .Y(\datapath_1.mux_pcsrc.dout [19])
);

NAND3X1 _11994_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[20]),
    .C(_3017__bF$buf4),
    .Y(_3081_)
);

NAND3X1 _11995_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [20]),
    .C(_3019__bF$buf4),
    .Y(_3082_)
);

AOI22X1 _11996_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [20]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3083_)
);

NAND3X1 _11997_ (
    .A(_3082_),
    .B(_3081_),
    .C(_3083_),
    .Y(\datapath_1.mux_pcsrc.dout [20])
);

NAND3X1 _11998_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[21]),
    .C(_3017__bF$buf3),
    .Y(_3084_)
);

NAND3X1 _11999_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [21]),
    .C(_3019__bF$buf3),
    .Y(_3085_)
);

AOI22X1 _12000_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [21]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3086_)
);

NAND3X1 _12001_ (
    .A(_3085_),
    .B(_3084_),
    .C(_3086_),
    .Y(\datapath_1.mux_pcsrc.dout [21])
);

NAND3X1 _12002_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[22]),
    .C(_3017__bF$buf2),
    .Y(_3087_)
);

NAND3X1 _12003_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .C(_3019__bF$buf2),
    .Y(_3088_)
);

AOI22X1 _12004_ (
    .A(_3021__bF$buf2),
    .B(\datapath_1.ALUResult [22]),
    .C(gnd),
    .D(_3022__bF$buf2),
    .Y(_3089_)
);

NAND3X1 _12005_ (
    .A(_3088_),
    .B(_3087_),
    .C(_3089_),
    .Y(\datapath_1.mux_pcsrc.dout [22])
);

NAND3X1 _12006_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[23]),
    .C(_3017__bF$buf1),
    .Y(_3090_)
);

NAND3X1 _12007_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [23]),
    .C(_3019__bF$buf1),
    .Y(_3091_)
);

AOI22X1 _12008_ (
    .A(_3021__bF$buf1),
    .B(\datapath_1.ALUResult [23]),
    .C(gnd),
    .D(_3022__bF$buf1),
    .Y(_3092_)
);

NAND3X1 _12009_ (
    .A(_3091_),
    .B(_3090_),
    .C(_3092_),
    .Y(\datapath_1.mux_pcsrc.dout [23])
);

NAND3X1 _12010_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[24]),
    .C(_3017__bF$buf0),
    .Y(_3093_)
);

NAND3X1 _12011_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [24]),
    .C(_3019__bF$buf0),
    .Y(_3094_)
);

AOI22X1 _12012_ (
    .A(_3021__bF$buf0),
    .B(\datapath_1.ALUResult [24]),
    .C(gnd),
    .D(_3022__bF$buf0),
    .Y(_3095_)
);

NAND3X1 _12013_ (
    .A(_3094_),
    .B(_3093_),
    .C(_3095_),
    .Y(\datapath_1.mux_pcsrc.dout [24])
);

NAND3X1 _12014_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[25]),
    .C(_3017__bF$buf4),
    .Y(_3096_)
);

NAND3X1 _12015_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [25]),
    .C(_3019__bF$buf4),
    .Y(_3097_)
);

AOI22X1 _12016_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [25]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3098_)
);

NAND3X1 _12017_ (
    .A(_3097_),
    .B(_3096_),
    .C(_3098_),
    .Y(\datapath_1.mux_pcsrc.dout [25])
);

NAND3X1 _12018_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[26]),
    .C(_3017__bF$buf3),
    .Y(_3099_)
);

NAND3X1 _12019_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [26]),
    .C(_3019__bF$buf3),
    .Y(_3100_)
);

AOI22X1 _12020_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [26]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3101_)
);

NAND3X1 _12021_ (
    .A(_3100_),
    .B(_3099_),
    .C(_3101_),
    .Y(\datapath_1.mux_pcsrc.dout [26])
);

NAND3X1 _12022_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[27]),
    .C(_3017__bF$buf2),
    .Y(_3102_)
);

NAND3X1 _12023_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_27_bF$buf4 ),
    .C(_3019__bF$buf2),
    .Y(_3103_)
);

AOI22X1 _12024_ (
    .A(_3021__bF$buf2),
    .B(\datapath_1.ALUResult [27]),
    .C(gnd),
    .D(_3022__bF$buf2),
    .Y(_3104_)
);

NAND3X1 _12025_ (
    .A(_3103_),
    .B(_3102_),
    .C(_3104_),
    .Y(\datapath_1.mux_pcsrc.dout [27])
);

NAND3X1 _12026_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[28]),
    .C(_3017__bF$buf1),
    .Y(_3105_)
);

NAND3X1 _12027_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [28]),
    .C(_3019__bF$buf1),
    .Y(_3106_)
);

AOI22X1 _12028_ (
    .A(_3021__bF$buf1),
    .B(\datapath_1.ALUResult [28]),
    .C(gnd),
    .D(_3022__bF$buf1),
    .Y(_3107_)
);

NAND3X1 _12029_ (
    .A(_3106_),
    .B(_3105_),
    .C(_3107_),
    .Y(\datapath_1.mux_pcsrc.dout [28])
);

NAND3X1 _12030_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[29]),
    .C(_3017__bF$buf0),
    .Y(_3108_)
);

NAND3X1 _12031_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [29]),
    .C(_3019__bF$buf0),
    .Y(_3109_)
);

AOI22X1 _12032_ (
    .A(_3021__bF$buf0),
    .B(\datapath_1.ALUResult [29]),
    .C(gnd),
    .D(_3022__bF$buf0),
    .Y(_3110_)
);

NAND3X1 _12033_ (
    .A(_3109_),
    .B(_3108_),
    .C(_3110_),
    .Y(\datapath_1.mux_pcsrc.dout [29])
);

NAND3X1 _12034_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[30]),
    .C(_3017__bF$buf4),
    .Y(_3111_)
);

NAND3X1 _12035_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [30]),
    .C(_3019__bF$buf4),
    .Y(_3112_)
);

AOI22X1 _12036_ (
    .A(_3021__bF$buf4),
    .B(\datapath_1.ALUResult [30]),
    .C(gnd),
    .D(_3022__bF$buf4),
    .Y(_3113_)
);

NAND3X1 _12037_ (
    .A(_3112_),
    .B(_3111_),
    .C(_3113_),
    .Y(\datapath_1.mux_pcsrc.dout [30])
);

NAND3X1 _12038_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[31]),
    .C(_3017__bF$buf3),
    .Y(_3114_)
);

NAND3X1 _12039_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [31]),
    .C(_3019__bF$buf3),
    .Y(_3115_)
);

AOI22X1 _12040_ (
    .A(_3021__bF$buf3),
    .B(\datapath_1.ALUResult [31]),
    .C(gnd),
    .D(_3022__bF$buf3),
    .Y(_3116_)
);

NAND3X1 _12041_ (
    .A(_3115_),
    .B(_3114_),
    .C(_3116_),
    .Y(\datapath_1.mux_pcsrc.dout [31])
);

INVX1 _12042_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3179_)
);

NAND2X1 _12043_ (
    .A(\datapath_1.a [0]),
    .B(ALUSrcA_bF$buf7),
    .Y(_3180_)
);

OAI21X1 _12044_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3179_),
    .C(_3180_),
    .Y(\datapath_1.alu_1.ALUInA [0])
);

INVX1 _12045_ (
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_3117_)
);

NAND2X1 _12046_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [1]),
    .Y(_3118_)
);

OAI21X1 _12047_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3117_),
    .C(_3118_),
    .Y(\datapath_1.alu_1.ALUInA [1])
);

INVX1 _12048_ (
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_3119_)
);

NAND2X1 _12049_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [2]),
    .Y(_3120_)
);

OAI21X1 _12050_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3119_),
    .C(_3120_),
    .Y(\datapath_1.alu_1.ALUInA [2])
);

INVX1 _12051_ (
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_3121_)
);

NAND2X1 _12052_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [3]),
    .Y(_3122_)
);

OAI21X1 _12053_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3121_),
    .C(_3122_),
    .Y(\datapath_1.alu_1.ALUInA [3])
);

INVX1 _12054_ (
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_3123_)
);

NAND2X1 _12055_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [4]),
    .Y(_3124_)
);

OAI21X1 _12056_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3123_),
    .C(_3124_),
    .Y(\datapath_1.alu_1.ALUInA [4])
);

INVX1 _12057_ (
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_3125_)
);

NAND2X1 _12058_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [5]),
    .Y(_3126_)
);

OAI21X1 _12059_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3125_),
    .C(_3126_),
    .Y(\datapath_1.alu_1.ALUInA [5])
);

INVX1 _12060_ (
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_3127_)
);

NAND2X1 _12061_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [6]),
    .Y(_3128_)
);

OAI21X1 _12062_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3127_),
    .C(_3128_),
    .Y(\datapath_1.alu_1.ALUInA [6])
);

INVX1 _12063_ (
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_3129_)
);

NAND2X1 _12064_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [7]),
    .Y(_3130_)
);

OAI21X1 _12065_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3129_),
    .C(_3130_),
    .Y(\datapath_1.alu_1.ALUInA [7])
);

INVX1 _12066_ (
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_3131_)
);

NAND2X1 _12067_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [8]),
    .Y(_3132_)
);

OAI21X1 _12068_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3131_),
    .C(_3132_),
    .Y(\datapath_1.alu_1.ALUInA [8])
);

INVX1 _12069_ (
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_3133_)
);

NAND2X1 _12070_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [9]),
    .Y(_3134_)
);

OAI21X1 _12071_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3133_),
    .C(_3134_),
    .Y(\datapath_1.alu_1.ALUInA [9])
);

INVX1 _12072_ (
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_3135_)
);

NAND2X1 _12073_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [10]),
    .Y(_3136_)
);

OAI21X1 _12074_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3135_),
    .C(_3136_),
    .Y(\datapath_1.alu_1.ALUInA [10])
);

INVX1 _12075_ (
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_3137_)
);

NAND2X1 _12076_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [11]),
    .Y(_3138_)
);

OAI21X1 _12077_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3137_),
    .C(_3138_),
    .Y(\datapath_1.alu_1.ALUInA [11])
);

INVX1 _12078_ (
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_3139_)
);

NAND2X1 _12079_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [12]),
    .Y(_3140_)
);

OAI21X1 _12080_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3139_),
    .C(_3140_),
    .Y(\datapath_1.alu_1.ALUInA [12])
);

INVX1 _12081_ (
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_3141_)
);

NAND2X1 _12082_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [13]),
    .Y(_3142_)
);

OAI21X1 _12083_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3141_),
    .C(_3142_),
    .Y(\datapath_1.alu_1.ALUInA [13])
);

INVX1 _12084_ (
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_3143_)
);

NAND2X1 _12085_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [14]),
    .Y(_3144_)
);

OAI21X1 _12086_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3143_),
    .C(_3144_),
    .Y(\datapath_1.alu_1.ALUInA [14])
);

INVX1 _12087_ (
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_3145_)
);

NAND2X1 _12088_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [15]),
    .Y(_3146_)
);

OAI21X1 _12089_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3145_),
    .C(_3146_),
    .Y(\datapath_1.alu_1.ALUInA [15])
);

INVX1 _12090_ (
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_3147_)
);

NAND2X1 _12091_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [16]),
    .Y(_3148_)
);

OAI21X1 _12092_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3147_),
    .C(_3148_),
    .Y(\datapath_1.alu_1.ALUInA [16])
);

INVX1 _12093_ (
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3149_)
);

NAND2X1 _12094_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [17]),
    .Y(_3150_)
);

OAI21X1 _12095_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3149_),
    .C(_3150_),
    .Y(\datapath_1.alu_1.ALUInA [17])
);

INVX1 _12096_ (
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3151_)
);

NAND2X1 _12097_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [18]),
    .Y(_3152_)
);

OAI21X1 _12098_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3151_),
    .C(_3152_),
    .Y(\datapath_1.alu_1.ALUInA [18])
);

INVX1 _12099_ (
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3153_)
);

NAND2X1 _12100_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [19]),
    .Y(_3154_)
);

OAI21X1 _12101_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3153_),
    .C(_3154_),
    .Y(\datapath_1.alu_1.ALUInA [19])
);

INVX1 _12102_ (
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3155_)
);

NAND2X1 _12103_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [20]),
    .Y(_3156_)
);

OAI21X1 _12104_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3155_),
    .C(_3156_),
    .Y(\datapath_1.alu_1.ALUInA [20])
);

INVX1 _12105_ (
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3157_)
);

NAND2X1 _12106_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [21]),
    .Y(_3158_)
);

OAI21X1 _12107_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3157_),
    .C(_3158_),
    .Y(\datapath_1.alu_1.ALUInA [21])
);

INVX1 _12108_ (
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3159_)
);

NAND2X1 _12109_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [22]),
    .Y(_3160_)
);

OAI21X1 _12110_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3159_),
    .C(_3160_),
    .Y(\datapath_1.alu_1.ALUInA [22])
);

INVX1 _12111_ (
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3161_)
);

NAND2X1 _12112_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [23]),
    .Y(_3162_)
);

OAI21X1 _12113_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3161_),
    .C(_3162_),
    .Y(\datapath_1.alu_1.ALUInA [23])
);

INVX1 _12114_ (
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3163_)
);

NAND2X1 _12115_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [24]),
    .Y(_3164_)
);

OAI21X1 _12116_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3163_),
    .C(_3164_),
    .Y(\datapath_1.alu_1.ALUInA [24])
);

INVX1 _12117_ (
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3165_)
);

NAND2X1 _12118_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [25]),
    .Y(_3166_)
);

OAI21X1 _12119_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3165_),
    .C(_3166_),
    .Y(\datapath_1.alu_1.ALUInA [25])
);

INVX1 _12120_ (
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3167_)
);

NAND2X1 _12121_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [26]),
    .Y(_3168_)
);

OAI21X1 _12122_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3167_),
    .C(_3168_),
    .Y(\datapath_1.alu_1.ALUInA [26])
);

INVX1 _12123_ (
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3169_)
);

NAND2X1 _12124_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [27]),
    .Y(_3170_)
);

OAI21X1 _12125_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3169_),
    .C(_3170_),
    .Y(\datapath_1.alu_1.ALUInA [27])
);

INVX1 _12126_ (
    .A(\datapath_1.PCJump [28]),
    .Y(_3171_)
);

NAND2X1 _12127_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [28]),
    .Y(_3172_)
);

OAI21X1 _12128_ (
    .A(ALUSrcA_bF$buf6),
    .B(_3171_),
    .C(_3172_),
    .Y(\datapath_1.alu_1.ALUInA [28])
);

INVX1 _12129_ (
    .A(\datapath_1.PCJump [29]),
    .Y(_3173_)
);

NAND2X1 _12130_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [29]),
    .Y(_3174_)
);

OAI21X1 _12131_ (
    .A(ALUSrcA_bF$buf4),
    .B(_3173_),
    .C(_3174_),
    .Y(\datapath_1.alu_1.ALUInA [29])
);

INVX1 _12132_ (
    .A(\datapath_1.PCJump [30]),
    .Y(_3175_)
);

NAND2X1 _12133_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [30]),
    .Y(_3176_)
);

OAI21X1 _12134_ (
    .A(ALUSrcA_bF$buf2),
    .B(_3175_),
    .C(_3176_),
    .Y(\datapath_1.alu_1.ALUInA [30])
);

INVX1 _12135_ (
    .A(\datapath_1.PCJump [31]),
    .Y(_3177_)
);

NAND2X1 _12136_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [31]),
    .Y(_3178_)
);

OAI21X1 _12137_ (
    .A(ALUSrcA_bF$buf0),
    .B(_3177_),
    .C(_3178_),
    .Y(\datapath_1.alu_1.ALUInA [31])
);

INVX8 _12138_ (
    .A(ALUSrcB_1_bF$buf4),
    .Y(_3181_)
);

NAND3X1 _12139_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3182_)
);

INVX8 _12140_ (
    .A(ALUSrcB_0_bF$buf3),
    .Y(_3183_)
);

NAND3X1 _12141_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [0]),
    .C(_3183__bF$buf4),
    .Y(_3184_)
);

NOR2X1 _12142_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(ALUSrcB_1_bF$buf2),
    .Y(_3185_)
);

AND2X2 _12143_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(ALUSrcB_0_bF$buf1),
    .Y(_3186_)
);

AOI22X1 _12144_ (
    .A(_3185__bF$buf4),
    .B(_2_[0]),
    .C(gnd),
    .D(_3186__bF$buf4),
    .Y(_3187_)
);

NAND3X1 _12145_ (
    .A(_3184_),
    .B(_3182_),
    .C(_3187_),
    .Y(\datapath_1.alu_1.ALUInB [0])
);

NAND3X1 _12146_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3188_)
);

NAND3X1 _12147_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\aluControl_1.inst [1]),
    .C(_3183__bF$buf3),
    .Y(_3189_)
);

AOI22X1 _12148_ (
    .A(_3185__bF$buf3),
    .B(_2_[1]),
    .C(gnd),
    .D(_3186__bF$buf3),
    .Y(_3190_)
);

NAND3X1 _12149_ (
    .A(_3189_),
    .B(_3188_),
    .C(_3190_),
    .Y(\datapath_1.alu_1.ALUInB [1])
);

NAND3X1 _12150_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(vdd),
    .C(_3181__bF$buf2),
    .Y(_3191_)
);

NAND3X1 _12151_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\aluControl_1.inst [2]),
    .C(_3183__bF$buf2),
    .Y(_3192_)
);

AOI22X1 _12152_ (
    .A(_3185__bF$buf2),
    .B(_2_[2]),
    .C(\aluControl_1.inst [0]),
    .D(_3186__bF$buf2),
    .Y(_3193_)
);

NAND3X1 _12153_ (
    .A(_3192_),
    .B(_3191_),
    .C(_3193_),
    .Y(\datapath_1.alu_1.ALUInB [2])
);

NAND3X1 _12154_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3181__bF$buf1),
    .Y(_3194_)
);

NAND3X1 _12155_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [3]),
    .C(_3183__bF$buf1),
    .Y(_3195_)
);

AOI22X1 _12156_ (
    .A(_3185__bF$buf1),
    .B(_2_[3]),
    .C(\aluControl_1.inst [1]),
    .D(_3186__bF$buf1),
    .Y(_3196_)
);

NAND3X1 _12157_ (
    .A(_3195_),
    .B(_3194_),
    .C(_3196_),
    .Y(\datapath_1.alu_1.ALUInB [3])
);

NAND3X1 _12158_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3181__bF$buf0),
    .Y(_3197_)
);

NAND3X1 _12159_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\aluControl_1.inst [4]),
    .C(_3183__bF$buf0),
    .Y(_3198_)
);

AOI22X1 _12160_ (
    .A(_3185__bF$buf0),
    .B(_2_[4]),
    .C(\aluControl_1.inst [2]),
    .D(_3186__bF$buf0),
    .Y(_3199_)
);

NAND3X1 _12161_ (
    .A(_3198_),
    .B(_3197_),
    .C(_3199_),
    .Y(\datapath_1.alu_1.ALUInB [4])
);

NAND3X1 _12162_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3200_)
);

NAND3X1 _12163_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\aluControl_1.inst [5]),
    .C(_3183__bF$buf4),
    .Y(_3201_)
);

AOI22X1 _12164_ (
    .A(_3185__bF$buf4),
    .B(_2_[5]),
    .C(\aluControl_1.inst [3]),
    .D(_3186__bF$buf4),
    .Y(_3202_)
);

NAND3X1 _12165_ (
    .A(_3201_),
    .B(_3200_),
    .C(_3202_),
    .Y(\datapath_1.alu_1.ALUInB [5])
);

NAND3X1 _12166_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3203_)
);

NAND3X1 _12167_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [8]),
    .C(_3183__bF$buf3),
    .Y(_3204_)
);

AOI22X1 _12168_ (
    .A(_3185__bF$buf3),
    .B(_2_[6]),
    .C(\aluControl_1.inst [4]),
    .D(_3186__bF$buf3),
    .Y(_3205_)
);

NAND3X1 _12169_ (
    .A(_3204_),
    .B(_3203_),
    .C(_3205_),
    .Y(\datapath_1.alu_1.ALUInB [6])
);

NAND3X1 _12170_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3181__bF$buf2),
    .Y(_3206_)
);

NAND3X1 _12171_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [9]),
    .C(_3183__bF$buf2),
    .Y(_3207_)
);

AOI22X1 _12172_ (
    .A(_3185__bF$buf2),
    .B(_2_[7]),
    .C(\aluControl_1.inst [5]),
    .D(_3186__bF$buf2),
    .Y(_3208_)
);

NAND3X1 _12173_ (
    .A(_3207_),
    .B(_3206_),
    .C(_3208_),
    .Y(\datapath_1.alu_1.ALUInB [7])
);

NAND3X1 _12174_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3181__bF$buf1),
    .Y(_3209_)
);

NAND3X1 _12175_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump [10]),
    .C(_3183__bF$buf1),
    .Y(_3210_)
);

AOI22X1 _12176_ (
    .A(_3185__bF$buf1),
    .B(_2_[8]),
    .C(\datapath_1.PCJump [8]),
    .D(_3186__bF$buf1),
    .Y(_3211_)
);

NAND3X1 _12177_ (
    .A(_3210_),
    .B(_3209_),
    .C(_3211_),
    .Y(\datapath_1.alu_1.ALUInB [8])
);

NAND3X1 _12178_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3181__bF$buf0),
    .Y(_3212_)
);

NAND3X1 _12179_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump [11]),
    .C(_3183__bF$buf0),
    .Y(_3213_)
);

AOI22X1 _12180_ (
    .A(_3185__bF$buf0),
    .B(_2_[9]),
    .C(\datapath_1.PCJump [9]),
    .D(_3186__bF$buf0),
    .Y(_3214_)
);

NAND3X1 _12181_ (
    .A(_3213_),
    .B(_3212_),
    .C(_3214_),
    .Y(\datapath_1.alu_1.ALUInB [9])
);

NAND3X1 _12182_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3215_)
);

NAND3X1 _12183_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump [12]),
    .C(_3183__bF$buf4),
    .Y(_3216_)
);

AOI22X1 _12184_ (
    .A(_3185__bF$buf4),
    .B(_2_[10]),
    .C(\datapath_1.PCJump [10]),
    .D(_3186__bF$buf4),
    .Y(_3217_)
);

NAND3X1 _12185_ (
    .A(_3216_),
    .B(_3215_),
    .C(_3217_),
    .Y(\datapath_1.alu_1.ALUInB [10])
);

NAND3X1 _12186_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3218_)
);

NAND3X1 _12187_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [13]),
    .C(_3183__bF$buf3),
    .Y(_3219_)
);

AOI22X1 _12188_ (
    .A(_3185__bF$buf3),
    .B(_2_[11]),
    .C(\datapath_1.PCJump [11]),
    .D(_3186__bF$buf3),
    .Y(_3220_)
);

NAND3X1 _12189_ (
    .A(_3219_),
    .B(_3218_),
    .C(_3220_),
    .Y(\datapath_1.alu_1.ALUInB [11])
);

NAND3X1 _12190_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3181__bF$buf2),
    .Y(_3221_)
);

NAND3X1 _12191_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [14]),
    .C(_3183__bF$buf2),
    .Y(_3222_)
);

AOI22X1 _12192_ (
    .A(_3185__bF$buf2),
    .B(_2_[12]),
    .C(\datapath_1.PCJump [12]),
    .D(_3186__bF$buf2),
    .Y(_3223_)
);

NAND3X1 _12193_ (
    .A(_3222_),
    .B(_3221_),
    .C(_3223_),
    .Y(\datapath_1.alu_1.ALUInB [12])
);

NAND3X1 _12194_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3181__bF$buf1),
    .Y(_3224_)
);

NAND3X1 _12195_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump [15]),
    .C(_3183__bF$buf1),
    .Y(_3225_)
);

AOI22X1 _12196_ (
    .A(_3185__bF$buf1),
    .B(_2_[13]),
    .C(\datapath_1.PCJump [13]),
    .D(_3186__bF$buf1),
    .Y(_3226_)
);

NAND3X1 _12197_ (
    .A(_3225_),
    .B(_3224_),
    .C(_3226_),
    .Y(\datapath_1.alu_1.ALUInB [13])
);

NAND3X1 _12198_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3181__bF$buf0),
    .Y(_3227_)
);

NAND3X1 _12199_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump [16]),
    .C(_3183__bF$buf0),
    .Y(_3228_)
);

AOI22X1 _12200_ (
    .A(_3185__bF$buf0),
    .B(_2_[14]),
    .C(\datapath_1.PCJump [14]),
    .D(_3186__bF$buf0),
    .Y(_3229_)
);

NAND3X1 _12201_ (
    .A(_3228_),
    .B(_3227_),
    .C(_3229_),
    .Y(\datapath_1.alu_1.ALUInB [14])
);

NAND3X1 _12202_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3230_)
);

NAND3X1 _12203_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3183__bF$buf4),
    .Y(_3231_)
);

AOI22X1 _12204_ (
    .A(_3185__bF$buf4),
    .B(_2_[15]),
    .C(\datapath_1.PCJump [15]),
    .D(_3186__bF$buf4),
    .Y(_3232_)
);

NAND3X1 _12205_ (
    .A(_3231_),
    .B(_3230_),
    .C(_3232_),
    .Y(\datapath_1.alu_1.ALUInB [15])
);

NAND3X1 _12206_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3233_)
);

NAND3X1 _12207_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3183__bF$buf3),
    .Y(_3234_)
);

AOI22X1 _12208_ (
    .A(_3185__bF$buf3),
    .B(_2_[16]),
    .C(\datapath_1.PCJump [16]),
    .D(_3186__bF$buf3),
    .Y(_3235_)
);

NAND3X1 _12209_ (
    .A(_3234_),
    .B(_3233_),
    .C(_3235_),
    .Y(\datapath_1.alu_1.ALUInB [16])
);

NAND3X1 _12210_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3181__bF$buf2),
    .Y(_3236_)
);

NAND3X1 _12211_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3183__bF$buf2),
    .Y(_3237_)
);

AOI22X1 _12212_ (
    .A(_3185__bF$buf2),
    .B(_2_[17]),
    .C(\datapath_1.PCJump_17_bF$buf4 ),
    .D(_3186__bF$buf2),
    .Y(_3238_)
);

NAND3X1 _12213_ (
    .A(_3237_),
    .B(_3236_),
    .C(_3238_),
    .Y(\datapath_1.alu_1.ALUInB [17])
);

NAND3X1 _12214_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3181__bF$buf1),
    .Y(_3239_)
);

NAND3X1 _12215_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3183__bF$buf1),
    .Y(_3240_)
);

AOI22X1 _12216_ (
    .A(_3185__bF$buf1),
    .B(_2_[18]),
    .C(\datapath_1.PCJump_17_bF$buf2 ),
    .D(_3186__bF$buf1),
    .Y(_3241_)
);

NAND3X1 _12217_ (
    .A(_3240_),
    .B(_3239_),
    .C(_3241_),
    .Y(\datapath_1.alu_1.ALUInB [18])
);

NAND3X1 _12218_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3181__bF$buf0),
    .Y(_3242_)
);

NAND3X1 _12219_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3183__bF$buf0),
    .Y(_3243_)
);

AOI22X1 _12220_ (
    .A(_3185__bF$buf0),
    .B(_2_[19]),
    .C(\datapath_1.PCJump_17_bF$buf0 ),
    .D(_3186__bF$buf0),
    .Y(_3244_)
);

NAND3X1 _12221_ (
    .A(_3243_),
    .B(_3242_),
    .C(_3244_),
    .Y(\datapath_1.alu_1.ALUInB [19])
);

NAND3X1 _12222_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3245_)
);

NAND3X1 _12223_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3183__bF$buf4),
    .Y(_3246_)
);

AOI22X1 _12224_ (
    .A(_3185__bF$buf4),
    .B(_2_[20]),
    .C(\datapath_1.PCJump_17_bF$buf3 ),
    .D(_3186__bF$buf4),
    .Y(_3247_)
);

NAND3X1 _12225_ (
    .A(_3246_),
    .B(_3245_),
    .C(_3247_),
    .Y(\datapath_1.alu_1.ALUInB [20])
);

NAND3X1 _12226_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3248_)
);

NAND3X1 _12227_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3183__bF$buf3),
    .Y(_3249_)
);

AOI22X1 _12228_ (
    .A(_3185__bF$buf3),
    .B(_2_[21]),
    .C(\datapath_1.PCJump_17_bF$buf1 ),
    .D(_3186__bF$buf3),
    .Y(_3250_)
);

NAND3X1 _12229_ (
    .A(_3249_),
    .B(_3248_),
    .C(_3250_),
    .Y(\datapath_1.alu_1.ALUInB [21])
);

NAND3X1 _12230_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3181__bF$buf2),
    .Y(_3251_)
);

NAND3X1 _12231_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3183__bF$buf2),
    .Y(_3252_)
);

AOI22X1 _12232_ (
    .A(_3185__bF$buf2),
    .B(_2_[22]),
    .C(\datapath_1.PCJump_17_bF$buf4 ),
    .D(_3186__bF$buf2),
    .Y(_3253_)
);

NAND3X1 _12233_ (
    .A(_3252_),
    .B(_3251_),
    .C(_3253_),
    .Y(\datapath_1.alu_1.ALUInB [22])
);

NAND3X1 _12234_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3181__bF$buf1),
    .Y(_3254_)
);

NAND3X1 _12235_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3183__bF$buf1),
    .Y(_3255_)
);

AOI22X1 _12236_ (
    .A(_3185__bF$buf1),
    .B(_2_[23]),
    .C(\datapath_1.PCJump_17_bF$buf2 ),
    .D(_3186__bF$buf1),
    .Y(_3256_)
);

NAND3X1 _12237_ (
    .A(_3255_),
    .B(_3254_),
    .C(_3256_),
    .Y(\datapath_1.alu_1.ALUInB [23])
);

NAND3X1 _12238_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3181__bF$buf0),
    .Y(_3257_)
);

NAND3X1 _12239_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3183__bF$buf0),
    .Y(_3258_)
);

AOI22X1 _12240_ (
    .A(_3185__bF$buf0),
    .B(_2_[24]),
    .C(\datapath_1.PCJump_17_bF$buf0 ),
    .D(_3186__bF$buf0),
    .Y(_3259_)
);

NAND3X1 _12241_ (
    .A(_3258_),
    .B(_3257_),
    .C(_3259_),
    .Y(\datapath_1.alu_1.ALUInB [24])
);

NAND3X1 _12242_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3260_)
);

NAND3X1 _12243_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3183__bF$buf4),
    .Y(_3261_)
);

AOI22X1 _12244_ (
    .A(_3185__bF$buf4),
    .B(_2_[25]),
    .C(\datapath_1.PCJump_17_bF$buf3 ),
    .D(_3186__bF$buf4),
    .Y(_3262_)
);

NAND3X1 _12245_ (
    .A(_3261_),
    .B(_3260_),
    .C(_3262_),
    .Y(\datapath_1.alu_1.ALUInB [25])
);

NAND3X1 _12246_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3263_)
);

NAND3X1 _12247_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3183__bF$buf3),
    .Y(_3264_)
);

AOI22X1 _12248_ (
    .A(_3185__bF$buf3),
    .B(_2_[26]),
    .C(\datapath_1.PCJump_17_bF$buf1 ),
    .D(_3186__bF$buf3),
    .Y(_3265_)
);

NAND3X1 _12249_ (
    .A(_3264_),
    .B(_3263_),
    .C(_3265_),
    .Y(\datapath_1.alu_1.ALUInB [26])
);

NAND3X1 _12250_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3181__bF$buf2),
    .Y(_3266_)
);

NAND3X1 _12251_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3183__bF$buf2),
    .Y(_3267_)
);

AOI22X1 _12252_ (
    .A(_3185__bF$buf2),
    .B(_2_[27]),
    .C(\datapath_1.PCJump_17_bF$buf4 ),
    .D(_3186__bF$buf2),
    .Y(_3268_)
);

NAND3X1 _12253_ (
    .A(_3267_),
    .B(_3266_),
    .C(_3268_),
    .Y(\datapath_1.alu_1.ALUInB [27])
);

NAND3X1 _12254_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3181__bF$buf1),
    .Y(_3269_)
);

NAND3X1 _12255_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3183__bF$buf1),
    .Y(_3270_)
);

AOI22X1 _12256_ (
    .A(_3185__bF$buf1),
    .B(_2_[28]),
    .C(\datapath_1.PCJump_17_bF$buf2 ),
    .D(_3186__bF$buf1),
    .Y(_3271_)
);

NAND3X1 _12257_ (
    .A(_3270_),
    .B(_3269_),
    .C(_3271_),
    .Y(\datapath_1.alu_1.ALUInB [28])
);

NAND3X1 _12258_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3181__bF$buf0),
    .Y(_3272_)
);

NAND3X1 _12259_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3183__bF$buf0),
    .Y(_3273_)
);

AOI22X1 _12260_ (
    .A(_3185__bF$buf0),
    .B(_2_[29]),
    .C(\datapath_1.PCJump_17_bF$buf0 ),
    .D(_3186__bF$buf0),
    .Y(_3274_)
);

NAND3X1 _12261_ (
    .A(_3273_),
    .B(_3272_),
    .C(_3274_),
    .Y(\datapath_1.alu_1.ALUInB [29])
);

NAND3X1 _12262_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3181__bF$buf4),
    .Y(_3275_)
);

NAND3X1 _12263_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3183__bF$buf4),
    .Y(_3276_)
);

AOI22X1 _12264_ (
    .A(_3185__bF$buf4),
    .B(_2_[30]),
    .C(\datapath_1.PCJump_17_bF$buf3 ),
    .D(_3186__bF$buf4),
    .Y(_3277_)
);

NAND3X1 _12265_ (
    .A(_3276_),
    .B(_3275_),
    .C(_3277_),
    .Y(\datapath_1.alu_1.ALUInB [30])
);

NAND3X1 _12266_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3181__bF$buf3),
    .Y(_3278_)
);

NAND3X1 _12267_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3183__bF$buf3),
    .Y(_3279_)
);

AOI22X1 _12268_ (
    .A(_3185__bF$buf3),
    .B(_2_[31]),
    .C(\datapath_1.PCJump_17_bF$buf1 ),
    .D(_3186__bF$buf3),
    .Y(_3280_)
);

NAND3X1 _12269_ (
    .A(_3279_),
    .B(_3278_),
    .C(_3280_),
    .Y(\datapath_1.alu_1.ALUInB [31])
);

INVX1 _12270_ (
    .A(ALUOut[0]),
    .Y(_3343_)
);

NAND2X1 _12271_ (
    .A(\datapath_1.Data [0]),
    .B(MemToReg_bF$buf7),
    .Y(_3344_)
);

OAI21X1 _12272_ (
    .A(MemToReg_bF$buf6),
    .B(_3343_),
    .C(_3344_),
    .Y(\datapath_1.mux_wd3.dout [0])
);

INVX1 _12273_ (
    .A(ALUOut[1]),
    .Y(_3281_)
);

NAND2X1 _12274_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [1]),
    .Y(_3282_)
);

OAI21X1 _12275_ (
    .A(MemToReg_bF$buf4),
    .B(_3281_),
    .C(_3282_),
    .Y(\datapath_1.mux_wd3.dout [1])
);

INVX1 _12276_ (
    .A(ALUOut[2]),
    .Y(_3283_)
);

NAND2X1 _12277_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [2]),
    .Y(_3284_)
);

OAI21X1 _12278_ (
    .A(MemToReg_bF$buf2),
    .B(_3283_),
    .C(_3284_),
    .Y(\datapath_1.mux_wd3.dout [2])
);

INVX1 _12279_ (
    .A(ALUOut[3]),
    .Y(_3285_)
);

NAND2X1 _12280_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [3]),
    .Y(_3286_)
);

OAI21X1 _12281_ (
    .A(MemToReg_bF$buf0),
    .B(_3285_),
    .C(_3286_),
    .Y(\datapath_1.mux_wd3.dout [3])
);

INVX1 _12282_ (
    .A(ALUOut[4]),
    .Y(_3287_)
);

NAND2X1 _12283_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [4]),
    .Y(_3288_)
);

OAI21X1 _12284_ (
    .A(MemToReg_bF$buf6),
    .B(_3287_),
    .C(_3288_),
    .Y(\datapath_1.mux_wd3.dout [4])
);

INVX1 _12285_ (
    .A(ALUOut[5]),
    .Y(_3289_)
);

NAND2X1 _12286_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [5]),
    .Y(_3290_)
);

OAI21X1 _12287_ (
    .A(MemToReg_bF$buf4),
    .B(_3289_),
    .C(_3290_),
    .Y(\datapath_1.mux_wd3.dout [5])
);

INVX1 _12288_ (
    .A(ALUOut[6]),
    .Y(_3291_)
);

NAND2X1 _12289_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [6]),
    .Y(_3292_)
);

OAI21X1 _12290_ (
    .A(MemToReg_bF$buf2),
    .B(_3291_),
    .C(_3292_),
    .Y(\datapath_1.mux_wd3.dout [6])
);

INVX1 _12291_ (
    .A(ALUOut[7]),
    .Y(_3293_)
);

NAND2X1 _12292_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [7]),
    .Y(_3294_)
);

OAI21X1 _12293_ (
    .A(MemToReg_bF$buf0),
    .B(_3293_),
    .C(_3294_),
    .Y(\datapath_1.mux_wd3.dout [7])
);

INVX1 _12294_ (
    .A(ALUOut[8]),
    .Y(_3295_)
);

NAND2X1 _12295_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [8]),
    .Y(_3296_)
);

OAI21X1 _12296_ (
    .A(MemToReg_bF$buf6),
    .B(_3295_),
    .C(_3296_),
    .Y(\datapath_1.mux_wd3.dout [8])
);

INVX1 _12297_ (
    .A(ALUOut[9]),
    .Y(_3297_)
);

NAND2X1 _12298_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [9]),
    .Y(_3298_)
);

OAI21X1 _12299_ (
    .A(MemToReg_bF$buf4),
    .B(_3297_),
    .C(_3298_),
    .Y(\datapath_1.mux_wd3.dout [9])
);

INVX1 _12300_ (
    .A(ALUOut[10]),
    .Y(_3299_)
);

NAND2X1 _12301_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [10]),
    .Y(_3300_)
);

OAI21X1 _12302_ (
    .A(MemToReg_bF$buf2),
    .B(_3299_),
    .C(_3300_),
    .Y(\datapath_1.mux_wd3.dout [10])
);

INVX1 _12303_ (
    .A(ALUOut[11]),
    .Y(_3301_)
);

NAND2X1 _12304_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [11]),
    .Y(_3302_)
);

OAI21X1 _12305_ (
    .A(MemToReg_bF$buf0),
    .B(_3301_),
    .C(_3302_),
    .Y(\datapath_1.mux_wd3.dout [11])
);

INVX1 _12306_ (
    .A(ALUOut[12]),
    .Y(_3303_)
);

NAND2X1 _12307_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [12]),
    .Y(_3304_)
);

OAI21X1 _12308_ (
    .A(MemToReg_bF$buf6),
    .B(_3303_),
    .C(_3304_),
    .Y(\datapath_1.mux_wd3.dout [12])
);

INVX1 _12309_ (
    .A(ALUOut[13]),
    .Y(_3305_)
);

NAND2X1 _12310_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [13]),
    .Y(_3306_)
);

OAI21X1 _12311_ (
    .A(MemToReg_bF$buf4),
    .B(_3305_),
    .C(_3306_),
    .Y(\datapath_1.mux_wd3.dout [13])
);

INVX1 _12312_ (
    .A(ALUOut[14]),
    .Y(_3307_)
);

NAND2X1 _12313_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [14]),
    .Y(_3308_)
);

OAI21X1 _12314_ (
    .A(MemToReg_bF$buf2),
    .B(_3307_),
    .C(_3308_),
    .Y(\datapath_1.mux_wd3.dout [14])
);

INVX1 _12315_ (
    .A(ALUOut[15]),
    .Y(_3309_)
);

NAND2X1 _12316_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [15]),
    .Y(_3310_)
);

OAI21X1 _12317_ (
    .A(MemToReg_bF$buf0),
    .B(_3309_),
    .C(_3310_),
    .Y(\datapath_1.mux_wd3.dout [15])
);

INVX1 _12318_ (
    .A(ALUOut[16]),
    .Y(_3311_)
);

NAND2X1 _12319_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [16]),
    .Y(_3312_)
);

OAI21X1 _12320_ (
    .A(MemToReg_bF$buf6),
    .B(_3311_),
    .C(_3312_),
    .Y(\datapath_1.mux_wd3.dout [16])
);

INVX1 _12321_ (
    .A(ALUOut[17]),
    .Y(_3313_)
);

NAND2X1 _12322_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [17]),
    .Y(_3314_)
);

OAI21X1 _12323_ (
    .A(MemToReg_bF$buf4),
    .B(_3313_),
    .C(_3314_),
    .Y(\datapath_1.mux_wd3.dout [17])
);

INVX1 _12324_ (
    .A(ALUOut[18]),
    .Y(_3315_)
);

NAND2X1 _12325_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [18]),
    .Y(_3316_)
);

OAI21X1 _12326_ (
    .A(MemToReg_bF$buf2),
    .B(_3315_),
    .C(_3316_),
    .Y(\datapath_1.mux_wd3.dout [18])
);

INVX1 _12327_ (
    .A(ALUOut[19]),
    .Y(_3317_)
);

NAND2X1 _12328_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [19]),
    .Y(_3318_)
);

OAI21X1 _12329_ (
    .A(MemToReg_bF$buf0),
    .B(_3317_),
    .C(_3318_),
    .Y(\datapath_1.mux_wd3.dout [19])
);

INVX1 _12330_ (
    .A(ALUOut[20]),
    .Y(_3319_)
);

NAND2X1 _12331_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [20]),
    .Y(_3320_)
);

OAI21X1 _12332_ (
    .A(MemToReg_bF$buf6),
    .B(_3319_),
    .C(_3320_),
    .Y(\datapath_1.mux_wd3.dout [20])
);

INVX1 _12333_ (
    .A(ALUOut[21]),
    .Y(_3321_)
);

NAND2X1 _12334_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [21]),
    .Y(_3322_)
);

OAI21X1 _12335_ (
    .A(MemToReg_bF$buf4),
    .B(_3321_),
    .C(_3322_),
    .Y(\datapath_1.mux_wd3.dout [21])
);

INVX1 _12336_ (
    .A(ALUOut[22]),
    .Y(_3323_)
);

NAND2X1 _12337_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [22]),
    .Y(_3324_)
);

OAI21X1 _12338_ (
    .A(MemToReg_bF$buf2),
    .B(_3323_),
    .C(_3324_),
    .Y(\datapath_1.mux_wd3.dout [22])
);

INVX1 _12339_ (
    .A(ALUOut[23]),
    .Y(_3325_)
);

NAND2X1 _12340_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [23]),
    .Y(_3326_)
);

OAI21X1 _12341_ (
    .A(MemToReg_bF$buf0),
    .B(_3325_),
    .C(_3326_),
    .Y(\datapath_1.mux_wd3.dout [23])
);

INVX1 _12342_ (
    .A(ALUOut[24]),
    .Y(_3327_)
);

NAND2X1 _12343_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [24]),
    .Y(_3328_)
);

OAI21X1 _12344_ (
    .A(MemToReg_bF$buf6),
    .B(_3327_),
    .C(_3328_),
    .Y(\datapath_1.mux_wd3.dout [24])
);

INVX1 _12345_ (
    .A(ALUOut[25]),
    .Y(_3329_)
);

NAND2X1 _12346_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [25]),
    .Y(_3330_)
);

OAI21X1 _12347_ (
    .A(MemToReg_bF$buf4),
    .B(_3329_),
    .C(_3330_),
    .Y(\datapath_1.mux_wd3.dout [25])
);

INVX1 _12348_ (
    .A(ALUOut[26]),
    .Y(_3331_)
);

NAND2X1 _12349_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [26]),
    .Y(_3332_)
);

OAI21X1 _12350_ (
    .A(MemToReg_bF$buf2),
    .B(_3331_),
    .C(_3332_),
    .Y(\datapath_1.mux_wd3.dout [26])
);

INVX1 _12351_ (
    .A(ALUOut[27]),
    .Y(_3333_)
);

NAND2X1 _12352_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [27]),
    .Y(_3334_)
);

OAI21X1 _12353_ (
    .A(MemToReg_bF$buf0),
    .B(_3333_),
    .C(_3334_),
    .Y(\datapath_1.mux_wd3.dout [27])
);

INVX1 _12354_ (
    .A(ALUOut[28]),
    .Y(_3335_)
);

NAND2X1 _12355_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [28]),
    .Y(_3336_)
);

OAI21X1 _12356_ (
    .A(MemToReg_bF$buf6),
    .B(_3335_),
    .C(_3336_),
    .Y(\datapath_1.mux_wd3.dout [28])
);

INVX1 _12357_ (
    .A(ALUOut[29]),
    .Y(_3337_)
);

NAND2X1 _12358_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [29]),
    .Y(_3338_)
);

OAI21X1 _12359_ (
    .A(MemToReg_bF$buf4),
    .B(_3337_),
    .C(_3338_),
    .Y(\datapath_1.mux_wd3.dout [29])
);

INVX1 _12360_ (
    .A(ALUOut[30]),
    .Y(_3339_)
);

NAND2X1 _12361_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [30]),
    .Y(_3340_)
);

OAI21X1 _12362_ (
    .A(MemToReg_bF$buf2),
    .B(_3339_),
    .C(_3340_),
    .Y(\datapath_1.mux_wd3.dout [30])
);

INVX1 _12363_ (
    .A(ALUOut[31]),
    .Y(_3341_)
);

NAND2X1 _12364_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [31]),
    .Y(_3342_)
);

OAI21X1 _12365_ (
    .A(MemToReg_bF$buf0),
    .B(_3341_),
    .C(_3342_),
    .Y(\datapath_1.mux_wd3.dout [31])
);

INVX1 _12366_ (
    .A(ALUOut[0]),
    .Y(_3408_)
);

NAND2X1 _12367_ (
    .A(\datapath_1.ALUResult [0]),
    .B(vdd),
    .Y(_3409_)
);

OAI21X1 _12368_ (
    .A(vdd),
    .B(_3408_),
    .C(_3409_),
    .Y(_3345_[0])
);

INVX1 _12369_ (
    .A(ALUOut[1]),
    .Y(_3346_)
);

NAND2X1 _12370_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [1]),
    .Y(_3347_)
);

OAI21X1 _12371_ (
    .A(vdd),
    .B(_3346_),
    .C(_3347_),
    .Y(_3345_[1])
);

INVX1 _12372_ (
    .A(ALUOut[2]),
    .Y(_3348_)
);

NAND2X1 _12373_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [2]),
    .Y(_3349_)
);

OAI21X1 _12374_ (
    .A(vdd),
    .B(_3348_),
    .C(_3349_),
    .Y(_3345_[2])
);

INVX1 _12375_ (
    .A(ALUOut[3]),
    .Y(_3350_)
);

NAND2X1 _12376_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [3]),
    .Y(_3351_)
);

OAI21X1 _12377_ (
    .A(vdd),
    .B(_3350_),
    .C(_3351_),
    .Y(_3345_[3])
);

INVX1 _12378_ (
    .A(ALUOut[4]),
    .Y(_3352_)
);

NAND2X1 _12379_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [4]),
    .Y(_3353_)
);

OAI21X1 _12380_ (
    .A(vdd),
    .B(_3352_),
    .C(_3353_),
    .Y(_3345_[4])
);

INVX1 _12381_ (
    .A(ALUOut[5]),
    .Y(_3354_)
);

NAND2X1 _12382_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [5]),
    .Y(_3355_)
);

OAI21X1 _12383_ (
    .A(vdd),
    .B(_3354_),
    .C(_3355_),
    .Y(_3345_[5])
);

INVX1 _12384_ (
    .A(ALUOut[6]),
    .Y(_3356_)
);

NAND2X1 _12385_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [6]),
    .Y(_3357_)
);

OAI21X1 _12386_ (
    .A(vdd),
    .B(_3356_),
    .C(_3357_),
    .Y(_3345_[6])
);

INVX1 _12387_ (
    .A(ALUOut[7]),
    .Y(_3358_)
);

NAND2X1 _12388_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [7]),
    .Y(_3359_)
);

OAI21X1 _12389_ (
    .A(vdd),
    .B(_3358_),
    .C(_3359_),
    .Y(_3345_[7])
);

INVX1 _12390_ (
    .A(ALUOut[8]),
    .Y(_3360_)
);

NAND2X1 _12391_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [8]),
    .Y(_3361_)
);

OAI21X1 _12392_ (
    .A(vdd),
    .B(_3360_),
    .C(_3361_),
    .Y(_3345_[8])
);

INVX1 _12393_ (
    .A(ALUOut[9]),
    .Y(_3362_)
);

NAND2X1 _12394_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [9]),
    .Y(_3363_)
);

OAI21X1 _12395_ (
    .A(vdd),
    .B(_3362_),
    .C(_3363_),
    .Y(_3345_[9])
);

INVX1 _12396_ (
    .A(ALUOut[10]),
    .Y(_3364_)
);

NAND2X1 _12397_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [10]),
    .Y(_3365_)
);

OAI21X1 _12398_ (
    .A(vdd),
    .B(_3364_),
    .C(_3365_),
    .Y(_3345_[10])
);

INVX1 _12399_ (
    .A(ALUOut[11]),
    .Y(_3366_)
);

NAND2X1 _12400_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [11]),
    .Y(_3367_)
);

OAI21X1 _12401_ (
    .A(vdd),
    .B(_3366_),
    .C(_3367_),
    .Y(_3345_[11])
);

INVX1 _12402_ (
    .A(ALUOut[12]),
    .Y(_3368_)
);

NAND2X1 _12403_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [12]),
    .Y(_3369_)
);

OAI21X1 _12404_ (
    .A(vdd),
    .B(_3368_),
    .C(_3369_),
    .Y(_3345_[12])
);

INVX1 _12405_ (
    .A(ALUOut[13]),
    .Y(_3370_)
);

NAND2X1 _12406_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [13]),
    .Y(_3371_)
);

OAI21X1 _12407_ (
    .A(vdd),
    .B(_3370_),
    .C(_3371_),
    .Y(_3345_[13])
);

INVX1 _12408_ (
    .A(ALUOut[14]),
    .Y(_3372_)
);

NAND2X1 _12409_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [14]),
    .Y(_3373_)
);

OAI21X1 _12410_ (
    .A(vdd),
    .B(_3372_),
    .C(_3373_),
    .Y(_3345_[14])
);

INVX1 _12411_ (
    .A(ALUOut[15]),
    .Y(_3374_)
);

NAND2X1 _12412_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [15]),
    .Y(_3375_)
);

OAI21X1 _12413_ (
    .A(vdd),
    .B(_3374_),
    .C(_3375_),
    .Y(_3345_[15])
);

INVX1 _12414_ (
    .A(ALUOut[16]),
    .Y(_3376_)
);

NAND2X1 _12415_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [16]),
    .Y(_3377_)
);

OAI21X1 _12416_ (
    .A(vdd),
    .B(_3376_),
    .C(_3377_),
    .Y(_3345_[16])
);

INVX1 _12417_ (
    .A(ALUOut[17]),
    .Y(_3378_)
);

NAND2X1 _12418_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [17]),
    .Y(_3379_)
);

OAI21X1 _12419_ (
    .A(vdd),
    .B(_3378_),
    .C(_3379_),
    .Y(_3345_[17])
);

INVX1 _12420_ (
    .A(ALUOut[18]),
    .Y(_3380_)
);

NAND2X1 _12421_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [18]),
    .Y(_3381_)
);

OAI21X1 _12422_ (
    .A(vdd),
    .B(_3380_),
    .C(_3381_),
    .Y(_3345_[18])
);

INVX1 _12423_ (
    .A(ALUOut[19]),
    .Y(_3382_)
);

NAND2X1 _12424_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [19]),
    .Y(_3383_)
);

OAI21X1 _12425_ (
    .A(vdd),
    .B(_3382_),
    .C(_3383_),
    .Y(_3345_[19])
);

INVX1 _12426_ (
    .A(ALUOut[20]),
    .Y(_3384_)
);

NAND2X1 _12427_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [20]),
    .Y(_3385_)
);

OAI21X1 _12428_ (
    .A(vdd),
    .B(_3384_),
    .C(_3385_),
    .Y(_3345_[20])
);

INVX1 _12429_ (
    .A(ALUOut[21]),
    .Y(_3386_)
);

NAND2X1 _12430_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [21]),
    .Y(_3387_)
);

OAI21X1 _12431_ (
    .A(vdd),
    .B(_3386_),
    .C(_3387_),
    .Y(_3345_[21])
);

INVX1 _12432_ (
    .A(ALUOut[22]),
    .Y(_3388_)
);

NAND2X1 _12433_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [22]),
    .Y(_3389_)
);

OAI21X1 _12434_ (
    .A(vdd),
    .B(_3388_),
    .C(_3389_),
    .Y(_3345_[22])
);

INVX1 _12435_ (
    .A(ALUOut[23]),
    .Y(_3390_)
);

NAND2X1 _12436_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [23]),
    .Y(_3391_)
);

OAI21X1 _12437_ (
    .A(vdd),
    .B(_3390_),
    .C(_3391_),
    .Y(_3345_[23])
);

INVX1 _12438_ (
    .A(ALUOut[24]),
    .Y(_3392_)
);

NAND2X1 _12439_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [24]),
    .Y(_3393_)
);

OAI21X1 _12440_ (
    .A(vdd),
    .B(_3392_),
    .C(_3393_),
    .Y(_3345_[24])
);

INVX1 _12441_ (
    .A(ALUOut[25]),
    .Y(_3394_)
);

NAND2X1 _12442_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [25]),
    .Y(_3395_)
);

OAI21X1 _12443_ (
    .A(vdd),
    .B(_3394_),
    .C(_3395_),
    .Y(_3345_[25])
);

INVX1 _12444_ (
    .A(ALUOut[26]),
    .Y(_3396_)
);

NAND2X1 _12445_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [26]),
    .Y(_3397_)
);

OAI21X1 _12446_ (
    .A(vdd),
    .B(_3396_),
    .C(_3397_),
    .Y(_3345_[26])
);

INVX1 _12447_ (
    .A(ALUOut[27]),
    .Y(_3398_)
);

NAND2X1 _12448_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [27]),
    .Y(_3399_)
);

OAI21X1 _12449_ (
    .A(vdd),
    .B(_3398_),
    .C(_3399_),
    .Y(_3345_[27])
);

INVX1 _12450_ (
    .A(ALUOut[28]),
    .Y(_3400_)
);

NAND2X1 _12451_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [28]),
    .Y(_3401_)
);

OAI21X1 _12452_ (
    .A(vdd),
    .B(_3400_),
    .C(_3401_),
    .Y(_3345_[28])
);

INVX1 _12453_ (
    .A(ALUOut[29]),
    .Y(_3402_)
);

NAND2X1 _12454_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [29]),
    .Y(_3403_)
);

OAI21X1 _12455_ (
    .A(vdd),
    .B(_3402_),
    .C(_3403_),
    .Y(_3345_[29])
);

INVX1 _12456_ (
    .A(ALUOut[30]),
    .Y(_3404_)
);

NAND2X1 _12457_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [30]),
    .Y(_3405_)
);

OAI21X1 _12458_ (
    .A(vdd),
    .B(_3404_),
    .C(_3405_),
    .Y(_3345_[30])
);

INVX1 _12459_ (
    .A(ALUOut[31]),
    .Y(_3406_)
);

NAND2X1 _12460_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [31]),
    .Y(_3407_)
);

OAI21X1 _12461_ (
    .A(vdd),
    .B(_3406_),
    .C(_3407_),
    .Y(_3345_[31])
);

DFFSR _12462_ (
    .CLK(clk_bF$buf113),
    .D(_3345_[0]),
    .Q(ALUOut[0]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _12463_ (
    .CLK(clk_bF$buf112),
    .D(_3345_[1]),
    .Q(ALUOut[1]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _12464_ (
    .CLK(clk_bF$buf111),
    .D(_3345_[2]),
    .Q(ALUOut[2]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _12465_ (
    .CLK(clk_bF$buf110),
    .D(_3345_[3]),
    .Q(ALUOut[3]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _12466_ (
    .CLK(clk_bF$buf109),
    .D(_3345_[4]),
    .Q(ALUOut[4]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _12467_ (
    .CLK(clk_bF$buf108),
    .D(_3345_[5]),
    .Q(ALUOut[5]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _12468_ (
    .CLK(clk_bF$buf107),
    .D(_3345_[6]),
    .Q(ALUOut[6]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _12469_ (
    .CLK(clk_bF$buf106),
    .D(_3345_[7]),
    .Q(ALUOut[7]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _12470_ (
    .CLK(clk_bF$buf105),
    .D(_3345_[8]),
    .Q(ALUOut[8]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _12471_ (
    .CLK(clk_bF$buf104),
    .D(_3345_[9]),
    .Q(ALUOut[9]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _12472_ (
    .CLK(clk_bF$buf103),
    .D(_3345_[10]),
    .Q(ALUOut[10]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _12473_ (
    .CLK(clk_bF$buf102),
    .D(_3345_[11]),
    .Q(ALUOut[11]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _12474_ (
    .CLK(clk_bF$buf101),
    .D(_3345_[12]),
    .Q(ALUOut[12]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _12475_ (
    .CLK(clk_bF$buf100),
    .D(_3345_[13]),
    .Q(ALUOut[13]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _12476_ (
    .CLK(clk_bF$buf99),
    .D(_3345_[14]),
    .Q(ALUOut[14]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _12477_ (
    .CLK(clk_bF$buf98),
    .D(_3345_[15]),
    .Q(ALUOut[15]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _12478_ (
    .CLK(clk_bF$buf97),
    .D(_3345_[16]),
    .Q(ALUOut[16]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _12479_ (
    .CLK(clk_bF$buf96),
    .D(_3345_[17]),
    .Q(ALUOut[17]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _12480_ (
    .CLK(clk_bF$buf95),
    .D(_3345_[18]),
    .Q(ALUOut[18]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _12481_ (
    .CLK(clk_bF$buf94),
    .D(_3345_[19]),
    .Q(ALUOut[19]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _12482_ (
    .CLK(clk_bF$buf93),
    .D(_3345_[20]),
    .Q(ALUOut[20]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _12483_ (
    .CLK(clk_bF$buf92),
    .D(_3345_[21]),
    .Q(ALUOut[21]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _12484_ (
    .CLK(clk_bF$buf91),
    .D(_3345_[22]),
    .Q(ALUOut[22]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _12485_ (
    .CLK(clk_bF$buf90),
    .D(_3345_[23]),
    .Q(ALUOut[23]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _12486_ (
    .CLK(clk_bF$buf89),
    .D(_3345_[24]),
    .Q(ALUOut[24]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _12487_ (
    .CLK(clk_bF$buf88),
    .D(_3345_[25]),
    .Q(ALUOut[25]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _12488_ (
    .CLK(clk_bF$buf87),
    .D(_3345_[26]),
    .Q(ALUOut[26]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _12489_ (
    .CLK(clk_bF$buf86),
    .D(_3345_[27]),
    .Q(ALUOut[27]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _12490_ (
    .CLK(clk_bF$buf85),
    .D(_3345_[28]),
    .Q(ALUOut[28]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _12491_ (
    .CLK(clk_bF$buf84),
    .D(_3345_[29]),
    .Q(ALUOut[29]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _12492_ (
    .CLK(clk_bF$buf83),
    .D(_3345_[30]),
    .Q(ALUOut[30]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _12493_ (
    .CLK(clk_bF$buf82),
    .D(_3345_[31]),
    .Q(ALUOut[31]),
    .R(rst_bF$buf82),
    .S(vdd)
);

INVX1 _12494_ (
    .A(\datapath_1.Data [0]),
    .Y(_3473_)
);

NAND2X1 _12495_ (
    .A(memoryOutData[0]),
    .B(vdd),
    .Y(_3474_)
);

OAI21X1 _12496_ (
    .A(vdd),
    .B(_3473_),
    .C(_3474_),
    .Y(_3410_[0])
);

INVX1 _12497_ (
    .A(\datapath_1.Data [1]),
    .Y(_3411_)
);

NAND2X1 _12498_ (
    .A(vdd),
    .B(memoryOutData[1]),
    .Y(_3412_)
);

OAI21X1 _12499_ (
    .A(vdd),
    .B(_3411_),
    .C(_3412_),
    .Y(_3410_[1])
);

INVX1 _12500_ (
    .A(\datapath_1.Data [2]),
    .Y(_3413_)
);

NAND2X1 _12501_ (
    .A(vdd),
    .B(memoryOutData[2]),
    .Y(_3414_)
);

OAI21X1 _12502_ (
    .A(vdd),
    .B(_3413_),
    .C(_3414_),
    .Y(_3410_[2])
);

INVX1 _12503_ (
    .A(\datapath_1.Data [3]),
    .Y(_3415_)
);

NAND2X1 _12504_ (
    .A(vdd),
    .B(memoryOutData[3]),
    .Y(_3416_)
);

OAI21X1 _12505_ (
    .A(vdd),
    .B(_3415_),
    .C(_3416_),
    .Y(_3410_[3])
);

INVX1 _12506_ (
    .A(\datapath_1.Data [4]),
    .Y(_3417_)
);

NAND2X1 _12507_ (
    .A(vdd),
    .B(memoryOutData[4]),
    .Y(_3418_)
);

OAI21X1 _12508_ (
    .A(vdd),
    .B(_3417_),
    .C(_3418_),
    .Y(_3410_[4])
);

INVX1 _12509_ (
    .A(\datapath_1.Data [5]),
    .Y(_3419_)
);

NAND2X1 _12510_ (
    .A(vdd),
    .B(memoryOutData[5]),
    .Y(_3420_)
);

OAI21X1 _12511_ (
    .A(vdd),
    .B(_3419_),
    .C(_3420_),
    .Y(_3410_[5])
);

INVX1 _12512_ (
    .A(\datapath_1.Data [6]),
    .Y(_3421_)
);

NAND2X1 _12513_ (
    .A(vdd),
    .B(memoryOutData[6]),
    .Y(_3422_)
);

OAI21X1 _12514_ (
    .A(vdd),
    .B(_3421_),
    .C(_3422_),
    .Y(_3410_[6])
);

INVX1 _12515_ (
    .A(\datapath_1.Data [7]),
    .Y(_3423_)
);

NAND2X1 _12516_ (
    .A(vdd),
    .B(memoryOutData[7]),
    .Y(_3424_)
);

OAI21X1 _12517_ (
    .A(vdd),
    .B(_3423_),
    .C(_3424_),
    .Y(_3410_[7])
);

INVX1 _12518_ (
    .A(\datapath_1.Data [8]),
    .Y(_3425_)
);

NAND2X1 _12519_ (
    .A(vdd),
    .B(memoryOutData[8]),
    .Y(_3426_)
);

OAI21X1 _12520_ (
    .A(vdd),
    .B(_3425_),
    .C(_3426_),
    .Y(_3410_[8])
);

INVX1 _12521_ (
    .A(\datapath_1.Data [9]),
    .Y(_3427_)
);

NAND2X1 _12522_ (
    .A(vdd),
    .B(memoryOutData[9]),
    .Y(_3428_)
);

OAI21X1 _12523_ (
    .A(vdd),
    .B(_3427_),
    .C(_3428_),
    .Y(_3410_[9])
);

INVX1 _12524_ (
    .A(\datapath_1.Data [10]),
    .Y(_3429_)
);

NAND2X1 _12525_ (
    .A(vdd),
    .B(memoryOutData[10]),
    .Y(_3430_)
);

OAI21X1 _12526_ (
    .A(vdd),
    .B(_3429_),
    .C(_3430_),
    .Y(_3410_[10])
);

INVX1 _12527_ (
    .A(\datapath_1.Data [11]),
    .Y(_3431_)
);

NAND2X1 _12528_ (
    .A(vdd),
    .B(memoryOutData[11]),
    .Y(_3432_)
);

OAI21X1 _12529_ (
    .A(vdd),
    .B(_3431_),
    .C(_3432_),
    .Y(_3410_[11])
);

INVX1 _12530_ (
    .A(\datapath_1.Data [12]),
    .Y(_3433_)
);

NAND2X1 _12531_ (
    .A(vdd),
    .B(memoryOutData[12]),
    .Y(_3434_)
);

OAI21X1 _12532_ (
    .A(vdd),
    .B(_3433_),
    .C(_3434_),
    .Y(_3410_[12])
);

INVX1 _12533_ (
    .A(\datapath_1.Data [13]),
    .Y(_3435_)
);

NAND2X1 _12534_ (
    .A(vdd),
    .B(memoryOutData[13]),
    .Y(_3436_)
);

OAI21X1 _12535_ (
    .A(vdd),
    .B(_3435_),
    .C(_3436_),
    .Y(_3410_[13])
);

INVX1 _12536_ (
    .A(\datapath_1.Data [14]),
    .Y(_3437_)
);

NAND2X1 _12537_ (
    .A(vdd),
    .B(memoryOutData[14]),
    .Y(_3438_)
);

OAI21X1 _12538_ (
    .A(vdd),
    .B(_3437_),
    .C(_3438_),
    .Y(_3410_[14])
);

INVX1 _12539_ (
    .A(\datapath_1.Data [15]),
    .Y(_3439_)
);

NAND2X1 _12540_ (
    .A(vdd),
    .B(memoryOutData[15]),
    .Y(_3440_)
);

OAI21X1 _12541_ (
    .A(vdd),
    .B(_3439_),
    .C(_3440_),
    .Y(_3410_[15])
);

INVX1 _12542_ (
    .A(\datapath_1.Data [16]),
    .Y(_3441_)
);

NAND2X1 _12543_ (
    .A(vdd),
    .B(memoryOutData[16]),
    .Y(_3442_)
);

OAI21X1 _12544_ (
    .A(vdd),
    .B(_3441_),
    .C(_3442_),
    .Y(_3410_[16])
);

INVX1 _12545_ (
    .A(\datapath_1.Data [17]),
    .Y(_3443_)
);

NAND2X1 _12546_ (
    .A(vdd),
    .B(memoryOutData[17]),
    .Y(_3444_)
);

OAI21X1 _12547_ (
    .A(vdd),
    .B(_3443_),
    .C(_3444_),
    .Y(_3410_[17])
);

INVX1 _12548_ (
    .A(\datapath_1.Data [18]),
    .Y(_3445_)
);

NAND2X1 _12549_ (
    .A(vdd),
    .B(memoryOutData[18]),
    .Y(_3446_)
);

OAI21X1 _12550_ (
    .A(vdd),
    .B(_3445_),
    .C(_3446_),
    .Y(_3410_[18])
);

INVX1 _12551_ (
    .A(\datapath_1.Data [19]),
    .Y(_3447_)
);

NAND2X1 _12552_ (
    .A(vdd),
    .B(memoryOutData[19]),
    .Y(_3448_)
);

OAI21X1 _12553_ (
    .A(vdd),
    .B(_3447_),
    .C(_3448_),
    .Y(_3410_[19])
);

INVX1 _12554_ (
    .A(\datapath_1.Data [20]),
    .Y(_3449_)
);

NAND2X1 _12555_ (
    .A(vdd),
    .B(memoryOutData[20]),
    .Y(_3450_)
);

OAI21X1 _12556_ (
    .A(vdd),
    .B(_3449_),
    .C(_3450_),
    .Y(_3410_[20])
);

INVX1 _12557_ (
    .A(\datapath_1.Data [21]),
    .Y(_3451_)
);

NAND2X1 _12558_ (
    .A(vdd),
    .B(memoryOutData[21]),
    .Y(_3452_)
);

OAI21X1 _12559_ (
    .A(vdd),
    .B(_3451_),
    .C(_3452_),
    .Y(_3410_[21])
);

INVX1 _12560_ (
    .A(\datapath_1.Data [22]),
    .Y(_3453_)
);

NAND2X1 _12561_ (
    .A(vdd),
    .B(memoryOutData[22]),
    .Y(_3454_)
);

OAI21X1 _12562_ (
    .A(vdd),
    .B(_3453_),
    .C(_3454_),
    .Y(_3410_[22])
);

INVX1 _12563_ (
    .A(\datapath_1.Data [23]),
    .Y(_3455_)
);

NAND2X1 _12564_ (
    .A(vdd),
    .B(memoryOutData[23]),
    .Y(_3456_)
);

OAI21X1 _12565_ (
    .A(vdd),
    .B(_3455_),
    .C(_3456_),
    .Y(_3410_[23])
);

INVX1 _12566_ (
    .A(\datapath_1.Data [24]),
    .Y(_3457_)
);

NAND2X1 _12567_ (
    .A(vdd),
    .B(memoryOutData[24]),
    .Y(_3458_)
);

OAI21X1 _12568_ (
    .A(vdd),
    .B(_3457_),
    .C(_3458_),
    .Y(_3410_[24])
);

INVX1 _12569_ (
    .A(\datapath_1.Data [25]),
    .Y(_3459_)
);

NAND2X1 _12570_ (
    .A(vdd),
    .B(memoryOutData[25]),
    .Y(_3460_)
);

OAI21X1 _12571_ (
    .A(vdd),
    .B(_3459_),
    .C(_3460_),
    .Y(_3410_[25])
);

INVX1 _12572_ (
    .A(\datapath_1.Data [26]),
    .Y(_3461_)
);

NAND2X1 _12573_ (
    .A(vdd),
    .B(memoryOutData[26]),
    .Y(_3462_)
);

OAI21X1 _12574_ (
    .A(vdd),
    .B(_3461_),
    .C(_3462_),
    .Y(_3410_[26])
);

INVX1 _12575_ (
    .A(\datapath_1.Data [27]),
    .Y(_3463_)
);

NAND2X1 _12576_ (
    .A(vdd),
    .B(memoryOutData[27]),
    .Y(_3464_)
);

OAI21X1 _12577_ (
    .A(vdd),
    .B(_3463_),
    .C(_3464_),
    .Y(_3410_[27])
);

INVX1 _12578_ (
    .A(\datapath_1.Data [28]),
    .Y(_3465_)
);

NAND2X1 _12579_ (
    .A(vdd),
    .B(memoryOutData[28]),
    .Y(_3466_)
);

OAI21X1 _12580_ (
    .A(vdd),
    .B(_3465_),
    .C(_3466_),
    .Y(_3410_[28])
);

INVX1 _12581_ (
    .A(\datapath_1.Data [29]),
    .Y(_3467_)
);

NAND2X1 _12582_ (
    .A(vdd),
    .B(memoryOutData[29]),
    .Y(_3468_)
);

OAI21X1 _12583_ (
    .A(vdd),
    .B(_3467_),
    .C(_3468_),
    .Y(_3410_[29])
);

INVX1 _12584_ (
    .A(\datapath_1.Data [30]),
    .Y(_3469_)
);

NAND2X1 _12585_ (
    .A(vdd),
    .B(memoryOutData[30]),
    .Y(_3470_)
);

OAI21X1 _12586_ (
    .A(vdd),
    .B(_3469_),
    .C(_3470_),
    .Y(_3410_[30])
);

INVX1 _12587_ (
    .A(\datapath_1.Data [31]),
    .Y(_3471_)
);

NAND2X1 _12588_ (
    .A(vdd),
    .B(memoryOutData[31]),
    .Y(_3472_)
);

OAI21X1 _12589_ (
    .A(vdd),
    .B(_3471_),
    .C(_3472_),
    .Y(_3410_[31])
);

DFFSR _12590_ (
    .CLK(clk_bF$buf81),
    .D(_3410_[0]),
    .Q(\datapath_1.Data [0]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _12591_ (
    .CLK(clk_bF$buf80),
    .D(_3410_[1]),
    .Q(\datapath_1.Data [1]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _12592_ (
    .CLK(clk_bF$buf79),
    .D(_3410_[2]),
    .Q(\datapath_1.Data [2]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _12593_ (
    .CLK(clk_bF$buf78),
    .D(_3410_[3]),
    .Q(\datapath_1.Data [3]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _12594_ (
    .CLK(clk_bF$buf77),
    .D(_3410_[4]),
    .Q(\datapath_1.Data [4]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _12595_ (
    .CLK(clk_bF$buf76),
    .D(_3410_[5]),
    .Q(\datapath_1.Data [5]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _12596_ (
    .CLK(clk_bF$buf75),
    .D(_3410_[6]),
    .Q(\datapath_1.Data [6]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _12597_ (
    .CLK(clk_bF$buf74),
    .D(_3410_[7]),
    .Q(\datapath_1.Data [7]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _12598_ (
    .CLK(clk_bF$buf73),
    .D(_3410_[8]),
    .Q(\datapath_1.Data [8]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _12599_ (
    .CLK(clk_bF$buf72),
    .D(_3410_[9]),
    .Q(\datapath_1.Data [9]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _12600_ (
    .CLK(clk_bF$buf71),
    .D(_3410_[10]),
    .Q(\datapath_1.Data [10]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _12601_ (
    .CLK(clk_bF$buf70),
    .D(_3410_[11]),
    .Q(\datapath_1.Data [11]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _12602_ (
    .CLK(clk_bF$buf69),
    .D(_3410_[12]),
    .Q(\datapath_1.Data [12]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _12603_ (
    .CLK(clk_bF$buf68),
    .D(_3410_[13]),
    .Q(\datapath_1.Data [13]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _12604_ (
    .CLK(clk_bF$buf67),
    .D(_3410_[14]),
    .Q(\datapath_1.Data [14]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _12605_ (
    .CLK(clk_bF$buf66),
    .D(_3410_[15]),
    .Q(\datapath_1.Data [15]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _12606_ (
    .CLK(clk_bF$buf65),
    .D(_3410_[16]),
    .Q(\datapath_1.Data [16]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _12607_ (
    .CLK(clk_bF$buf64),
    .D(_3410_[17]),
    .Q(\datapath_1.Data [17]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _12608_ (
    .CLK(clk_bF$buf63),
    .D(_3410_[18]),
    .Q(\datapath_1.Data [18]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _12609_ (
    .CLK(clk_bF$buf62),
    .D(_3410_[19]),
    .Q(\datapath_1.Data [19]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _12610_ (
    .CLK(clk_bF$buf61),
    .D(_3410_[20]),
    .Q(\datapath_1.Data [20]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _12611_ (
    .CLK(clk_bF$buf60),
    .D(_3410_[21]),
    .Q(\datapath_1.Data [21]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _12612_ (
    .CLK(clk_bF$buf59),
    .D(_3410_[22]),
    .Q(\datapath_1.Data [22]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _12613_ (
    .CLK(clk_bF$buf58),
    .D(_3410_[23]),
    .Q(\datapath_1.Data [23]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _12614_ (
    .CLK(clk_bF$buf57),
    .D(_3410_[24]),
    .Q(\datapath_1.Data [24]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _12615_ (
    .CLK(clk_bF$buf56),
    .D(_3410_[25]),
    .Q(\datapath_1.Data [25]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _12616_ (
    .CLK(clk_bF$buf55),
    .D(_3410_[26]),
    .Q(\datapath_1.Data [26]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _12617_ (
    .CLK(clk_bF$buf54),
    .D(_3410_[27]),
    .Q(\datapath_1.Data [27]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _12618_ (
    .CLK(clk_bF$buf53),
    .D(_3410_[28]),
    .Q(\datapath_1.Data [28]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _12619_ (
    .CLK(clk_bF$buf52),
    .D(_3410_[29]),
    .Q(\datapath_1.Data [29]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _12620_ (
    .CLK(clk_bF$buf51),
    .D(_3410_[30]),
    .Q(\datapath_1.Data [30]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _12621_ (
    .CLK(clk_bF$buf50),
    .D(_3410_[31]),
    .Q(\datapath_1.Data [31]),
    .R(rst_bF$buf50),
    .S(vdd)
);

INVX1 _12622_ (
    .A(\aluControl_1.inst [0]),
    .Y(_3538_)
);

NAND2X1 _12623_ (
    .A(memoryOutData[0]),
    .B(IRWrite_bF$buf6),
    .Y(_3539_)
);

OAI21X1 _12624_ (
    .A(IRWrite_bF$buf5),
    .B(_3538_),
    .C(_3539_),
    .Y(_3475_[0])
);

INVX1 _12625_ (
    .A(\aluControl_1.inst [1]),
    .Y(_3476_)
);

NAND2X1 _12626_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[1]),
    .Y(_3477_)
);

OAI21X1 _12627_ (
    .A(IRWrite_bF$buf3),
    .B(_3476_),
    .C(_3477_),
    .Y(_3475_[1])
);

INVX1 _12628_ (
    .A(\aluControl_1.inst [2]),
    .Y(_3478_)
);

NAND2X1 _12629_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[2]),
    .Y(_3479_)
);

OAI21X1 _12630_ (
    .A(IRWrite_bF$buf1),
    .B(_3478_),
    .C(_3479_),
    .Y(_3475_[2])
);

INVX1 _12631_ (
    .A(\aluControl_1.inst [3]),
    .Y(_3480_)
);

NAND2X1 _12632_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[3]),
    .Y(_3481_)
);

OAI21X1 _12633_ (
    .A(IRWrite_bF$buf7),
    .B(_3480_),
    .C(_3481_),
    .Y(_3475_[3])
);

INVX1 _12634_ (
    .A(\aluControl_1.inst [4]),
    .Y(_3482_)
);

NAND2X1 _12635_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[4]),
    .Y(_3483_)
);

OAI21X1 _12636_ (
    .A(IRWrite_bF$buf5),
    .B(_3482_),
    .C(_3483_),
    .Y(_3475_[4])
);

INVX1 _12637_ (
    .A(\aluControl_1.inst [5]),
    .Y(_3484_)
);

NAND2X1 _12638_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[5]),
    .Y(_3485_)
);

OAI21X1 _12639_ (
    .A(IRWrite_bF$buf3),
    .B(_3484_),
    .C(_3485_),
    .Y(_3475_[5])
);

INVX1 _12640_ (
    .A(\datapath_1.PCJump [8]),
    .Y(_3486_)
);

NAND2X1 _12641_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[6]),
    .Y(_3487_)
);

OAI21X1 _12642_ (
    .A(IRWrite_bF$buf1),
    .B(_3486_),
    .C(_3487_),
    .Y(_3475_[6])
);

INVX1 _12643_ (
    .A(\datapath_1.PCJump [9]),
    .Y(_3488_)
);

NAND2X1 _12644_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[7]),
    .Y(_3489_)
);

OAI21X1 _12645_ (
    .A(IRWrite_bF$buf7),
    .B(_3488_),
    .C(_3489_),
    .Y(_3475_[7])
);

INVX1 _12646_ (
    .A(\datapath_1.PCJump [10]),
    .Y(_3490_)
);

NAND2X1 _12647_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[8]),
    .Y(_3491_)
);

OAI21X1 _12648_ (
    .A(IRWrite_bF$buf5),
    .B(_3490_),
    .C(_3491_),
    .Y(_3475_[8])
);

INVX1 _12649_ (
    .A(\datapath_1.PCJump [11]),
    .Y(_3492_)
);

NAND2X1 _12650_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[9]),
    .Y(_3493_)
);

OAI21X1 _12651_ (
    .A(IRWrite_bF$buf3),
    .B(_3492_),
    .C(_3493_),
    .Y(_3475_[9])
);

INVX1 _12652_ (
    .A(\datapath_1.PCJump [12]),
    .Y(_3494_)
);

NAND2X1 _12653_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[10]),
    .Y(_3495_)
);

OAI21X1 _12654_ (
    .A(IRWrite_bF$buf1),
    .B(_3494_),
    .C(_3495_),
    .Y(_3475_[10])
);

INVX1 _12655_ (
    .A(\datapath_1.PCJump [13]),
    .Y(_3496_)
);

NAND2X1 _12656_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[11]),
    .Y(_3497_)
);

OAI21X1 _12657_ (
    .A(IRWrite_bF$buf7),
    .B(_3496_),
    .C(_3497_),
    .Y(_3475_[11])
);

INVX1 _12658_ (
    .A(\datapath_1.PCJump [14]),
    .Y(_3498_)
);

NAND2X1 _12659_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[12]),
    .Y(_3499_)
);

OAI21X1 _12660_ (
    .A(IRWrite_bF$buf5),
    .B(_3498_),
    .C(_3499_),
    .Y(_3475_[12])
);

INVX1 _12661_ (
    .A(\datapath_1.PCJump [15]),
    .Y(_3500_)
);

NAND2X1 _12662_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[13]),
    .Y(_3501_)
);

OAI21X1 _12663_ (
    .A(IRWrite_bF$buf3),
    .B(_3500_),
    .C(_3501_),
    .Y(_3475_[13])
);

INVX1 _12664_ (
    .A(\datapath_1.PCJump [16]),
    .Y(_3502_)
);

NAND2X1 _12665_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[14]),
    .Y(_3503_)
);

OAI21X1 _12666_ (
    .A(IRWrite_bF$buf1),
    .B(_3502_),
    .C(_3503_),
    .Y(_3475_[14])
);

INVX1 _12667_ (
    .A(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3504_)
);

NAND2X1 _12668_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[15]),
    .Y(_3505_)
);

OAI21X1 _12669_ (
    .A(IRWrite_bF$buf7),
    .B(_3504_),
    .C(_3505_),
    .Y(_3475_[15])
);

INVX1 _12670_ (
    .A(\datapath_1.PCJump [18]),
    .Y(_3506_)
);

NAND2X1 _12671_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[16]),
    .Y(_3507_)
);

OAI21X1 _12672_ (
    .A(IRWrite_bF$buf5),
    .B(_3506_),
    .C(_3507_),
    .Y(_3475_[16])
);

INVX1 _12673_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_3508_)
);

NAND2X1 _12674_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[17]),
    .Y(_3509_)
);

OAI21X1 _12675_ (
    .A(IRWrite_bF$buf3),
    .B(_3508_),
    .C(_3509_),
    .Y(_3475_[17])
);

INVX1 _12676_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_3510_)
);

NAND2X1 _12677_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[18]),
    .Y(_3511_)
);

OAI21X1 _12678_ (
    .A(IRWrite_bF$buf1),
    .B(_3510_),
    .C(_3511_),
    .Y(_3475_[18])
);

INVX1 _12679_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_3512_)
);

NAND2X1 _12680_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[19]),
    .Y(_3513_)
);

OAI21X1 _12681_ (
    .A(IRWrite_bF$buf7),
    .B(_3512_),
    .C(_3513_),
    .Y(_3475_[19])
);

INVX1 _12682_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_3514_)
);

NAND2X1 _12683_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[20]),
    .Y(_3515_)
);

OAI21X1 _12684_ (
    .A(IRWrite_bF$buf5),
    .B(_3514_),
    .C(_3515_),
    .Y(_3475_[20])
);

INVX1 _12685_ (
    .A(\datapath_1.PCJump [23]),
    .Y(_3516_)
);

NAND2X1 _12686_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[21]),
    .Y(_3517_)
);

OAI21X1 _12687_ (
    .A(IRWrite_bF$buf3),
    .B(_3516_),
    .C(_3517_),
    .Y(_3475_[21])
);

INVX1 _12688_ (
    .A(\datapath_1.PCJump [24]),
    .Y(_3518_)
);

NAND2X1 _12689_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[22]),
    .Y(_3519_)
);

OAI21X1 _12690_ (
    .A(IRWrite_bF$buf1),
    .B(_3518_),
    .C(_3519_),
    .Y(_3475_[22])
);

INVX1 _12691_ (
    .A(\datapath_1.PCJump [25]),
    .Y(_3520_)
);

NAND2X1 _12692_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[23]),
    .Y(_3521_)
);

OAI21X1 _12693_ (
    .A(IRWrite_bF$buf7),
    .B(_3520_),
    .C(_3521_),
    .Y(_3475_[23])
);

INVX1 _12694_ (
    .A(\datapath_1.PCJump [26]),
    .Y(_3522_)
);

NAND2X1 _12695_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[24]),
    .Y(_3523_)
);

OAI21X1 _12696_ (
    .A(IRWrite_bF$buf5),
    .B(_3522_),
    .C(_3523_),
    .Y(_3475_[24])
);

INVX1 _12697_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_3524_)
);

NAND2X1 _12698_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[25]),
    .Y(_3525_)
);

OAI21X1 _12699_ (
    .A(IRWrite_bF$buf3),
    .B(_3524_),
    .C(_3525_),
    .Y(_3475_[25])
);

INVX1 _12700_ (
    .A(\control_1.op [0]),
    .Y(_3526_)
);

NAND2X1 _12701_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[26]),
    .Y(_3527_)
);

OAI21X1 _12702_ (
    .A(IRWrite_bF$buf1),
    .B(_3526_),
    .C(_3527_),
    .Y(_3475_[26])
);

INVX1 _12703_ (
    .A(\control_1.op [1]),
    .Y(_3528_)
);

NAND2X1 _12704_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[27]),
    .Y(_3529_)
);

OAI21X1 _12705_ (
    .A(IRWrite_bF$buf7),
    .B(_3528_),
    .C(_3529_),
    .Y(_3475_[27])
);

INVX1 _12706_ (
    .A(\control_1.op [2]),
    .Y(_3530_)
);

NAND2X1 _12707_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[28]),
    .Y(_3531_)
);

OAI21X1 _12708_ (
    .A(IRWrite_bF$buf5),
    .B(_3530_),
    .C(_3531_),
    .Y(_3475_[28])
);

INVX1 _12709_ (
    .A(\control_1.op [3]),
    .Y(_3532_)
);

NAND2X1 _12710_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[29]),
    .Y(_3533_)
);

OAI21X1 _12711_ (
    .A(IRWrite_bF$buf3),
    .B(_3532_),
    .C(_3533_),
    .Y(_3475_[29])
);

INVX1 _12712_ (
    .A(\control_1.op [4]),
    .Y(_3534_)
);

NAND2X1 _12713_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[30]),
    .Y(_3535_)
);

OAI21X1 _12714_ (
    .A(IRWrite_bF$buf1),
    .B(_3534_),
    .C(_3535_),
    .Y(_3475_[30])
);

INVX1 _12715_ (
    .A(\control_1.op [5]),
    .Y(_3536_)
);

NAND2X1 _12716_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[31]),
    .Y(_3537_)
);

OAI21X1 _12717_ (
    .A(IRWrite_bF$buf7),
    .B(_3536_),
    .C(_3537_),
    .Y(_3475_[31])
);

DFFSR _12718_ (
    .CLK(clk_bF$buf49),
    .D(_3475_[0]),
    .Q(\aluControl_1.inst [0]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _12719_ (
    .CLK(clk_bF$buf48),
    .D(_3475_[1]),
    .Q(\aluControl_1.inst [1]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _12720_ (
    .CLK(clk_bF$buf47),
    .D(_3475_[2]),
    .Q(\aluControl_1.inst [2]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _12721_ (
    .CLK(clk_bF$buf46),
    .D(_3475_[3]),
    .Q(\aluControl_1.inst [3]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _12722_ (
    .CLK(clk_bF$buf45),
    .D(_3475_[4]),
    .Q(\aluControl_1.inst [4]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _12723_ (
    .CLK(clk_bF$buf44),
    .D(_3475_[5]),
    .Q(\aluControl_1.inst [5]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _12724_ (
    .CLK(clk_bF$buf43),
    .D(_3475_[6]),
    .Q(\datapath_1.PCJump [8]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _12725_ (
    .CLK(clk_bF$buf42),
    .D(_3475_[7]),
    .Q(\datapath_1.PCJump [9]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _12726_ (
    .CLK(clk_bF$buf41),
    .D(_3475_[8]),
    .Q(\datapath_1.PCJump [10]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _12727_ (
    .CLK(clk_bF$buf40),
    .D(_3475_[9]),
    .Q(\datapath_1.PCJump [11]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _12728_ (
    .CLK(clk_bF$buf39),
    .D(_3475_[10]),
    .Q(\datapath_1.PCJump [12]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _12729_ (
    .CLK(clk_bF$buf38),
    .D(_3475_[11]),
    .Q(\datapath_1.PCJump [13]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _12730_ (
    .CLK(clk_bF$buf37),
    .D(_3475_[12]),
    .Q(\datapath_1.PCJump [14]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _12731_ (
    .CLK(clk_bF$buf36),
    .D(_3475_[13]),
    .Q(\datapath_1.PCJump [15]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _12732_ (
    .CLK(clk_bF$buf35),
    .D(_3475_[14]),
    .Q(\datapath_1.PCJump [16]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _12733_ (
    .CLK(clk_bF$buf34),
    .D(_3475_[15]),
    .Q(\datapath_1.PCJump [17]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _12734_ (
    .CLK(clk_bF$buf33),
    .D(_3475_[16]),
    .Q(\datapath_1.PCJump [18]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _12735_ (
    .CLK(clk_bF$buf32),
    .D(_3475_[17]),
    .Q(\datapath_1.PCJump [19]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _12736_ (
    .CLK(clk_bF$buf31),
    .D(_3475_[18]),
    .Q(\datapath_1.PCJump [20]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _12737_ (
    .CLK(clk_bF$buf30),
    .D(_3475_[19]),
    .Q(\datapath_1.PCJump [21]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _12738_ (
    .CLK(clk_bF$buf29),
    .D(_3475_[20]),
    .Q(\datapath_1.PCJump [22]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _12739_ (
    .CLK(clk_bF$buf28),
    .D(_3475_[21]),
    .Q(\datapath_1.PCJump [23]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _12740_ (
    .CLK(clk_bF$buf27),
    .D(_3475_[22]),
    .Q(\datapath_1.PCJump [24]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _12741_ (
    .CLK(clk_bF$buf26),
    .D(_3475_[23]),
    .Q(\datapath_1.PCJump [25]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _12742_ (
    .CLK(clk_bF$buf25),
    .D(_3475_[24]),
    .Q(\datapath_1.PCJump [26]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _12743_ (
    .CLK(clk_bF$buf24),
    .D(_3475_[25]),
    .Q(\datapath_1.PCJump [27]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _12744_ (
    .CLK(clk_bF$buf23),
    .D(_3475_[26]),
    .Q(\control_1.op [0]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _12745_ (
    .CLK(clk_bF$buf22),
    .D(_3475_[27]),
    .Q(\control_1.op [1]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _12746_ (
    .CLK(clk_bF$buf21),
    .D(_3475_[28]),
    .Q(\control_1.op [2]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _12747_ (
    .CLK(clk_bF$buf20),
    .D(_3475_[29]),
    .Q(\control_1.op [3]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _12748_ (
    .CLK(clk_bF$buf19),
    .D(_3475_[30]),
    .Q(\control_1.op [4]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _12749_ (
    .CLK(clk_bF$buf18),
    .D(_3475_[31]),
    .Q(\control_1.op [5]),
    .R(rst_bF$buf18),
    .S(vdd)
);

INVX1 _12750_ (
    .A(\datapath_1.a [0]),
    .Y(_3603_)
);

NAND2X1 _12751_ (
    .A(\datapath_1.rd1 [0]),
    .B(vdd),
    .Y(_3604_)
);

OAI21X1 _12752_ (
    .A(vdd),
    .B(_3603_),
    .C(_3604_),
    .Y(_3540_[0])
);

INVX1 _12753_ (
    .A(\datapath_1.a [1]),
    .Y(_3541_)
);

NAND2X1 _12754_ (
    .A(vdd),
    .B(\datapath_1.rd1 [1]),
    .Y(_3542_)
);

OAI21X1 _12755_ (
    .A(vdd),
    .B(_3541_),
    .C(_3542_),
    .Y(_3540_[1])
);

INVX1 _12756_ (
    .A(\datapath_1.a [2]),
    .Y(_3543_)
);

NAND2X1 _12757_ (
    .A(vdd),
    .B(\datapath_1.rd1 [2]),
    .Y(_3544_)
);

OAI21X1 _12758_ (
    .A(vdd),
    .B(_3543_),
    .C(_3544_),
    .Y(_3540_[2])
);

INVX1 _12759_ (
    .A(\datapath_1.a [3]),
    .Y(_3545_)
);

NAND2X1 _12760_ (
    .A(vdd),
    .B(\datapath_1.rd1 [3]),
    .Y(_3546_)
);

OAI21X1 _12761_ (
    .A(vdd),
    .B(_3545_),
    .C(_3546_),
    .Y(_3540_[3])
);

INVX1 _12762_ (
    .A(\datapath_1.a [4]),
    .Y(_3547_)
);

NAND2X1 _12763_ (
    .A(vdd),
    .B(\datapath_1.rd1 [4]),
    .Y(_3548_)
);

OAI21X1 _12764_ (
    .A(vdd),
    .B(_3547_),
    .C(_3548_),
    .Y(_3540_[4])
);

INVX1 _12765_ (
    .A(\datapath_1.a [5]),
    .Y(_3549_)
);

NAND2X1 _12766_ (
    .A(vdd),
    .B(\datapath_1.rd1 [5]),
    .Y(_3550_)
);

OAI21X1 _12767_ (
    .A(vdd),
    .B(_3549_),
    .C(_3550_),
    .Y(_3540_[5])
);

INVX1 _12768_ (
    .A(\datapath_1.a [6]),
    .Y(_3551_)
);

NAND2X1 _12769_ (
    .A(vdd),
    .B(\datapath_1.rd1 [6]),
    .Y(_3552_)
);

OAI21X1 _12770_ (
    .A(vdd),
    .B(_3551_),
    .C(_3552_),
    .Y(_3540_[6])
);

INVX1 _12771_ (
    .A(\datapath_1.a [7]),
    .Y(_3553_)
);

NAND2X1 _12772_ (
    .A(vdd),
    .B(\datapath_1.rd1 [7]),
    .Y(_3554_)
);

OAI21X1 _12773_ (
    .A(vdd),
    .B(_3553_),
    .C(_3554_),
    .Y(_3540_[7])
);

INVX1 _12774_ (
    .A(\datapath_1.a [8]),
    .Y(_3555_)
);

NAND2X1 _12775_ (
    .A(vdd),
    .B(\datapath_1.rd1 [8]),
    .Y(_3556_)
);

OAI21X1 _12776_ (
    .A(vdd),
    .B(_3555_),
    .C(_3556_),
    .Y(_3540_[8])
);

INVX1 _12777_ (
    .A(\datapath_1.a [9]),
    .Y(_3557_)
);

NAND2X1 _12778_ (
    .A(vdd),
    .B(\datapath_1.rd1 [9]),
    .Y(_3558_)
);

OAI21X1 _12779_ (
    .A(vdd),
    .B(_3557_),
    .C(_3558_),
    .Y(_3540_[9])
);

INVX1 _12780_ (
    .A(\datapath_1.a [10]),
    .Y(_3559_)
);

NAND2X1 _12781_ (
    .A(vdd),
    .B(\datapath_1.rd1 [10]),
    .Y(_3560_)
);

OAI21X1 _12782_ (
    .A(vdd),
    .B(_3559_),
    .C(_3560_),
    .Y(_3540_[10])
);

INVX1 _12783_ (
    .A(\datapath_1.a [11]),
    .Y(_3561_)
);

NAND2X1 _12784_ (
    .A(vdd),
    .B(\datapath_1.rd1 [11]),
    .Y(_3562_)
);

OAI21X1 _12785_ (
    .A(vdd),
    .B(_3561_),
    .C(_3562_),
    .Y(_3540_[11])
);

INVX1 _12786_ (
    .A(\datapath_1.a [12]),
    .Y(_3563_)
);

NAND2X1 _12787_ (
    .A(vdd),
    .B(\datapath_1.rd1 [12]),
    .Y(_3564_)
);

OAI21X1 _12788_ (
    .A(vdd),
    .B(_3563_),
    .C(_3564_),
    .Y(_3540_[12])
);

INVX1 _12789_ (
    .A(\datapath_1.a [13]),
    .Y(_3565_)
);

NAND2X1 _12790_ (
    .A(vdd),
    .B(\datapath_1.rd1 [13]),
    .Y(_3566_)
);

OAI21X1 _12791_ (
    .A(vdd),
    .B(_3565_),
    .C(_3566_),
    .Y(_3540_[13])
);

INVX1 _12792_ (
    .A(\datapath_1.a [14]),
    .Y(_3567_)
);

NAND2X1 _12793_ (
    .A(vdd),
    .B(\datapath_1.rd1 [14]),
    .Y(_3568_)
);

OAI21X1 _12794_ (
    .A(vdd),
    .B(_3567_),
    .C(_3568_),
    .Y(_3540_[14])
);

INVX1 _12795_ (
    .A(\datapath_1.a [15]),
    .Y(_3569_)
);

NAND2X1 _12796_ (
    .A(vdd),
    .B(\datapath_1.rd1 [15]),
    .Y(_3570_)
);

OAI21X1 _12797_ (
    .A(vdd),
    .B(_3569_),
    .C(_3570_),
    .Y(_3540_[15])
);

INVX1 _12798_ (
    .A(\datapath_1.a [16]),
    .Y(_3571_)
);

NAND2X1 _12799_ (
    .A(vdd),
    .B(\datapath_1.rd1 [16]),
    .Y(_3572_)
);

OAI21X1 _12800_ (
    .A(vdd),
    .B(_3571_),
    .C(_3572_),
    .Y(_3540_[16])
);

INVX1 _12801_ (
    .A(\datapath_1.a [17]),
    .Y(_3573_)
);

NAND2X1 _12802_ (
    .A(vdd),
    .B(\datapath_1.rd1 [17]),
    .Y(_3574_)
);

OAI21X1 _12803_ (
    .A(vdd),
    .B(_3573_),
    .C(_3574_),
    .Y(_3540_[17])
);

INVX1 _12804_ (
    .A(\datapath_1.a [18]),
    .Y(_3575_)
);

NAND2X1 _12805_ (
    .A(vdd),
    .B(\datapath_1.rd1 [18]),
    .Y(_3576_)
);

OAI21X1 _12806_ (
    .A(vdd),
    .B(_3575_),
    .C(_3576_),
    .Y(_3540_[18])
);

INVX1 _12807_ (
    .A(\datapath_1.a [19]),
    .Y(_3577_)
);

NAND2X1 _12808_ (
    .A(vdd),
    .B(\datapath_1.rd1 [19]),
    .Y(_3578_)
);

OAI21X1 _12809_ (
    .A(vdd),
    .B(_3577_),
    .C(_3578_),
    .Y(_3540_[19])
);

INVX1 _12810_ (
    .A(\datapath_1.a [20]),
    .Y(_3579_)
);

NAND2X1 _12811_ (
    .A(vdd),
    .B(\datapath_1.rd1 [20]),
    .Y(_3580_)
);

OAI21X1 _12812_ (
    .A(vdd),
    .B(_3579_),
    .C(_3580_),
    .Y(_3540_[20])
);

INVX1 _12813_ (
    .A(\datapath_1.a [21]),
    .Y(_3581_)
);

NAND2X1 _12814_ (
    .A(vdd),
    .B(\datapath_1.rd1 [21]),
    .Y(_3582_)
);

OAI21X1 _12815_ (
    .A(vdd),
    .B(_3581_),
    .C(_3582_),
    .Y(_3540_[21])
);

INVX1 _12816_ (
    .A(\datapath_1.a [22]),
    .Y(_3583_)
);

NAND2X1 _12817_ (
    .A(vdd),
    .B(\datapath_1.rd1 [22]),
    .Y(_3584_)
);

OAI21X1 _12818_ (
    .A(vdd),
    .B(_3583_),
    .C(_3584_),
    .Y(_3540_[22])
);

INVX1 _12819_ (
    .A(\datapath_1.a [23]),
    .Y(_3585_)
);

NAND2X1 _12820_ (
    .A(vdd),
    .B(\datapath_1.rd1 [23]),
    .Y(_3586_)
);

OAI21X1 _12821_ (
    .A(vdd),
    .B(_3585_),
    .C(_3586_),
    .Y(_3540_[23])
);

INVX1 _12822_ (
    .A(\datapath_1.a [24]),
    .Y(_3587_)
);

NAND2X1 _12823_ (
    .A(vdd),
    .B(\datapath_1.rd1 [24]),
    .Y(_3588_)
);

OAI21X1 _12824_ (
    .A(vdd),
    .B(_3587_),
    .C(_3588_),
    .Y(_3540_[24])
);

INVX1 _12825_ (
    .A(\datapath_1.a [25]),
    .Y(_3589_)
);

NAND2X1 _12826_ (
    .A(vdd),
    .B(\datapath_1.rd1 [25]),
    .Y(_3590_)
);

OAI21X1 _12827_ (
    .A(vdd),
    .B(_3589_),
    .C(_3590_),
    .Y(_3540_[25])
);

INVX1 _12828_ (
    .A(\datapath_1.a [26]),
    .Y(_3591_)
);

NAND2X1 _12829_ (
    .A(vdd),
    .B(\datapath_1.rd1 [26]),
    .Y(_3592_)
);

OAI21X1 _12830_ (
    .A(vdd),
    .B(_3591_),
    .C(_3592_),
    .Y(_3540_[26])
);

INVX1 _12831_ (
    .A(\datapath_1.a [27]),
    .Y(_3593_)
);

NAND2X1 _12832_ (
    .A(vdd),
    .B(\datapath_1.rd1 [27]),
    .Y(_3594_)
);

OAI21X1 _12833_ (
    .A(vdd),
    .B(_3593_),
    .C(_3594_),
    .Y(_3540_[27])
);

INVX1 _12834_ (
    .A(\datapath_1.a [28]),
    .Y(_3595_)
);

NAND2X1 _12835_ (
    .A(vdd),
    .B(\datapath_1.rd1 [28]),
    .Y(_3596_)
);

OAI21X1 _12836_ (
    .A(vdd),
    .B(_3595_),
    .C(_3596_),
    .Y(_3540_[28])
);

INVX1 _12837_ (
    .A(\datapath_1.a [29]),
    .Y(_3597_)
);

NAND2X1 _12838_ (
    .A(vdd),
    .B(\datapath_1.rd1 [29]),
    .Y(_3598_)
);

OAI21X1 _12839_ (
    .A(vdd),
    .B(_3597_),
    .C(_3598_),
    .Y(_3540_[29])
);

INVX1 _12840_ (
    .A(\datapath_1.a [30]),
    .Y(_3599_)
);

NAND2X1 _12841_ (
    .A(vdd),
    .B(\datapath_1.rd1 [30]),
    .Y(_3600_)
);

OAI21X1 _12842_ (
    .A(vdd),
    .B(_3599_),
    .C(_3600_),
    .Y(_3540_[30])
);

INVX1 _12843_ (
    .A(\datapath_1.a [31]),
    .Y(_3601_)
);

NAND2X1 _12844_ (
    .A(vdd),
    .B(\datapath_1.rd1 [31]),
    .Y(_3602_)
);

OAI21X1 _12845_ (
    .A(vdd),
    .B(_3601_),
    .C(_3602_),
    .Y(_3540_[31])
);

DFFSR _12846_ (
    .CLK(clk_bF$buf17),
    .D(_3540_[0]),
    .Q(\datapath_1.a [0]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _12847_ (
    .CLK(clk_bF$buf16),
    .D(_3540_[1]),
    .Q(\datapath_1.a [1]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _12848_ (
    .CLK(clk_bF$buf15),
    .D(_3540_[2]),
    .Q(\datapath_1.a [2]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _12849_ (
    .CLK(clk_bF$buf14),
    .D(_3540_[3]),
    .Q(\datapath_1.a [3]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _12850_ (
    .CLK(clk_bF$buf13),
    .D(_3540_[4]),
    .Q(\datapath_1.a [4]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _12851_ (
    .CLK(clk_bF$buf12),
    .D(_3540_[5]),
    .Q(\datapath_1.a [5]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _12852_ (
    .CLK(clk_bF$buf11),
    .D(_3540_[6]),
    .Q(\datapath_1.a [6]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _12853_ (
    .CLK(clk_bF$buf10),
    .D(_3540_[7]),
    .Q(\datapath_1.a [7]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _12854_ (
    .CLK(clk_bF$buf9),
    .D(_3540_[8]),
    .Q(\datapath_1.a [8]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _12855_ (
    .CLK(clk_bF$buf8),
    .D(_3540_[9]),
    .Q(\datapath_1.a [9]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _12856_ (
    .CLK(clk_bF$buf7),
    .D(_3540_[10]),
    .Q(\datapath_1.a [10]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _12857_ (
    .CLK(clk_bF$buf6),
    .D(_3540_[11]),
    .Q(\datapath_1.a [11]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _12858_ (
    .CLK(clk_bF$buf5),
    .D(_3540_[12]),
    .Q(\datapath_1.a [12]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _12859_ (
    .CLK(clk_bF$buf4),
    .D(_3540_[13]),
    .Q(\datapath_1.a [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _12860_ (
    .CLK(clk_bF$buf3),
    .D(_3540_[14]),
    .Q(\datapath_1.a [14]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _12861_ (
    .CLK(clk_bF$buf2),
    .D(_3540_[15]),
    .Q(\datapath_1.a [15]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _12862_ (
    .CLK(clk_bF$buf1),
    .D(_3540_[16]),
    .Q(\datapath_1.a [16]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _12863_ (
    .CLK(clk_bF$buf0),
    .D(_3540_[17]),
    .Q(\datapath_1.a [17]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _12864_ (
    .CLK(clk_bF$buf113),
    .D(_3540_[18]),
    .Q(\datapath_1.a [18]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _12865_ (
    .CLK(clk_bF$buf112),
    .D(_3540_[19]),
    .Q(\datapath_1.a [19]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _12866_ (
    .CLK(clk_bF$buf111),
    .D(_3540_[20]),
    .Q(\datapath_1.a [20]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _12867_ (
    .CLK(clk_bF$buf110),
    .D(_3540_[21]),
    .Q(\datapath_1.a [21]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _12868_ (
    .CLK(clk_bF$buf109),
    .D(_3540_[22]),
    .Q(\datapath_1.a [22]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _12869_ (
    .CLK(clk_bF$buf108),
    .D(_3540_[23]),
    .Q(\datapath_1.a [23]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _12870_ (
    .CLK(clk_bF$buf107),
    .D(_3540_[24]),
    .Q(\datapath_1.a [24]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _12871_ (
    .CLK(clk_bF$buf106),
    .D(_3540_[25]),
    .Q(\datapath_1.a [25]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _12872_ (
    .CLK(clk_bF$buf105),
    .D(_3540_[26]),
    .Q(\datapath_1.a [26]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _12873_ (
    .CLK(clk_bF$buf104),
    .D(_3540_[27]),
    .Q(\datapath_1.a [27]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _12874_ (
    .CLK(clk_bF$buf103),
    .D(_3540_[28]),
    .Q(\datapath_1.a [28]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _12875_ (
    .CLK(clk_bF$buf102),
    .D(_3540_[29]),
    .Q(\datapath_1.a [29]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _12876_ (
    .CLK(clk_bF$buf101),
    .D(_3540_[30]),
    .Q(\datapath_1.a [30]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _12877_ (
    .CLK(clk_bF$buf100),
    .D(_3540_[31]),
    .Q(\datapath_1.a [31]),
    .R(rst_bF$buf100),
    .S(vdd)
);

INVX1 _12878_ (
    .A(_2_[0]),
    .Y(_3668_)
);

NAND2X1 _12879_ (
    .A(\datapath_1.rd2 [0]),
    .B(vdd),
    .Y(_3669_)
);

OAI21X1 _12880_ (
    .A(vdd),
    .B(_3668_),
    .C(_3669_),
    .Y(_3605_[0])
);

INVX1 _12881_ (
    .A(_2_[1]),
    .Y(_3606_)
);

NAND2X1 _12882_ (
    .A(vdd),
    .B(\datapath_1.rd2 [1]),
    .Y(_3607_)
);

OAI21X1 _12883_ (
    .A(vdd),
    .B(_3606_),
    .C(_3607_),
    .Y(_3605_[1])
);

INVX1 _12884_ (
    .A(_2_[2]),
    .Y(_3608_)
);

NAND2X1 _12885_ (
    .A(vdd),
    .B(\datapath_1.rd2 [2]),
    .Y(_3609_)
);

OAI21X1 _12886_ (
    .A(vdd),
    .B(_3608_),
    .C(_3609_),
    .Y(_3605_[2])
);

INVX1 _12887_ (
    .A(_2_[3]),
    .Y(_3610_)
);

NAND2X1 _12888_ (
    .A(vdd),
    .B(\datapath_1.rd2 [3]),
    .Y(_3611_)
);

OAI21X1 _12889_ (
    .A(vdd),
    .B(_3610_),
    .C(_3611_),
    .Y(_3605_[3])
);

INVX1 _12890_ (
    .A(_2_[4]),
    .Y(_3612_)
);

NAND2X1 _12891_ (
    .A(vdd),
    .B(\datapath_1.rd2 [4]),
    .Y(_3613_)
);

OAI21X1 _12892_ (
    .A(vdd),
    .B(_3612_),
    .C(_3613_),
    .Y(_3605_[4])
);

INVX1 _12893_ (
    .A(_2_[5]),
    .Y(_3614_)
);

NAND2X1 _12894_ (
    .A(vdd),
    .B(\datapath_1.rd2 [5]),
    .Y(_3615_)
);

OAI21X1 _12895_ (
    .A(vdd),
    .B(_3614_),
    .C(_3615_),
    .Y(_3605_[5])
);

INVX1 _12896_ (
    .A(_2_[6]),
    .Y(_3616_)
);

NAND2X1 _12897_ (
    .A(vdd),
    .B(\datapath_1.rd2 [6]),
    .Y(_3617_)
);

OAI21X1 _12898_ (
    .A(vdd),
    .B(_3616_),
    .C(_3617_),
    .Y(_3605_[6])
);

INVX1 _12899_ (
    .A(_2_[7]),
    .Y(_3618_)
);

NAND2X1 _12900_ (
    .A(vdd),
    .B(\datapath_1.rd2 [7]),
    .Y(_3619_)
);

OAI21X1 _12901_ (
    .A(vdd),
    .B(_3618_),
    .C(_3619_),
    .Y(_3605_[7])
);

INVX1 _12902_ (
    .A(_2_[8]),
    .Y(_3620_)
);

NAND2X1 _12903_ (
    .A(vdd),
    .B(\datapath_1.rd2 [8]),
    .Y(_3621_)
);

OAI21X1 _12904_ (
    .A(vdd),
    .B(_3620_),
    .C(_3621_),
    .Y(_3605_[8])
);

INVX1 _12905_ (
    .A(_2_[9]),
    .Y(_3622_)
);

NAND2X1 _12906_ (
    .A(vdd),
    .B(\datapath_1.rd2 [9]),
    .Y(_3623_)
);

OAI21X1 _12907_ (
    .A(vdd),
    .B(_3622_),
    .C(_3623_),
    .Y(_3605_[9])
);

INVX1 _12908_ (
    .A(_2_[10]),
    .Y(_3624_)
);

NAND2X1 _12909_ (
    .A(vdd),
    .B(\datapath_1.rd2 [10]),
    .Y(_3625_)
);

OAI21X1 _12910_ (
    .A(vdd),
    .B(_3624_),
    .C(_3625_),
    .Y(_3605_[10])
);

INVX1 _12911_ (
    .A(_2_[11]),
    .Y(_3626_)
);

NAND2X1 _12912_ (
    .A(vdd),
    .B(\datapath_1.rd2 [11]),
    .Y(_3627_)
);

OAI21X1 _12913_ (
    .A(vdd),
    .B(_3626_),
    .C(_3627_),
    .Y(_3605_[11])
);

INVX1 _12914_ (
    .A(_2_[12]),
    .Y(_3628_)
);

NAND2X1 _12915_ (
    .A(vdd),
    .B(\datapath_1.rd2 [12]),
    .Y(_3629_)
);

OAI21X1 _12916_ (
    .A(vdd),
    .B(_3628_),
    .C(_3629_),
    .Y(_3605_[12])
);

INVX1 _12917_ (
    .A(_2_[13]),
    .Y(_3630_)
);

NAND2X1 _12918_ (
    .A(vdd),
    .B(\datapath_1.rd2 [13]),
    .Y(_3631_)
);

OAI21X1 _12919_ (
    .A(vdd),
    .B(_3630_),
    .C(_3631_),
    .Y(_3605_[13])
);

INVX1 _12920_ (
    .A(_2_[14]),
    .Y(_3632_)
);

NAND2X1 _12921_ (
    .A(vdd),
    .B(\datapath_1.rd2 [14]),
    .Y(_3633_)
);

OAI21X1 _12922_ (
    .A(vdd),
    .B(_3632_),
    .C(_3633_),
    .Y(_3605_[14])
);

INVX1 _12923_ (
    .A(_2_[15]),
    .Y(_3634_)
);

NAND2X1 _12924_ (
    .A(vdd),
    .B(\datapath_1.rd2 [15]),
    .Y(_3635_)
);

OAI21X1 _12925_ (
    .A(vdd),
    .B(_3634_),
    .C(_3635_),
    .Y(_3605_[15])
);

INVX1 _12926_ (
    .A(_2_[16]),
    .Y(_3636_)
);

NAND2X1 _12927_ (
    .A(vdd),
    .B(\datapath_1.rd2 [16]),
    .Y(_3637_)
);

OAI21X1 _12928_ (
    .A(vdd),
    .B(_3636_),
    .C(_3637_),
    .Y(_3605_[16])
);

INVX1 _12929_ (
    .A(_2_[17]),
    .Y(_3638_)
);

NAND2X1 _12930_ (
    .A(vdd),
    .B(\datapath_1.rd2 [17]),
    .Y(_3639_)
);

OAI21X1 _12931_ (
    .A(vdd),
    .B(_3638_),
    .C(_3639_),
    .Y(_3605_[17])
);

INVX1 _12932_ (
    .A(_2_[18]),
    .Y(_3640_)
);

NAND2X1 _12933_ (
    .A(vdd),
    .B(\datapath_1.rd2 [18]),
    .Y(_3641_)
);

OAI21X1 _12934_ (
    .A(vdd),
    .B(_3640_),
    .C(_3641_),
    .Y(_3605_[18])
);

INVX1 _12935_ (
    .A(_2_[19]),
    .Y(_3642_)
);

NAND2X1 _12936_ (
    .A(vdd),
    .B(\datapath_1.rd2 [19]),
    .Y(_3643_)
);

OAI21X1 _12937_ (
    .A(vdd),
    .B(_3642_),
    .C(_3643_),
    .Y(_3605_[19])
);

INVX1 _12938_ (
    .A(_2_[20]),
    .Y(_3644_)
);

NAND2X1 _12939_ (
    .A(vdd),
    .B(\datapath_1.rd2 [20]),
    .Y(_3645_)
);

OAI21X1 _12940_ (
    .A(vdd),
    .B(_3644_),
    .C(_3645_),
    .Y(_3605_[20])
);

INVX1 _12941_ (
    .A(_2_[21]),
    .Y(_3646_)
);

NAND2X1 _12942_ (
    .A(vdd),
    .B(\datapath_1.rd2 [21]),
    .Y(_3647_)
);

OAI21X1 _12943_ (
    .A(vdd),
    .B(_3646_),
    .C(_3647_),
    .Y(_3605_[21])
);

INVX1 _12944_ (
    .A(_2_[22]),
    .Y(_3648_)
);

NAND2X1 _12945_ (
    .A(vdd),
    .B(\datapath_1.rd2 [22]),
    .Y(_3649_)
);

OAI21X1 _12946_ (
    .A(vdd),
    .B(_3648_),
    .C(_3649_),
    .Y(_3605_[22])
);

INVX1 _12947_ (
    .A(_2_[23]),
    .Y(_3650_)
);

NAND2X1 _12948_ (
    .A(vdd),
    .B(\datapath_1.rd2 [23]),
    .Y(_3651_)
);

OAI21X1 _12949_ (
    .A(vdd),
    .B(_3650_),
    .C(_3651_),
    .Y(_3605_[23])
);

INVX1 _12950_ (
    .A(_2_[24]),
    .Y(_3652_)
);

NAND2X1 _12951_ (
    .A(vdd),
    .B(\datapath_1.rd2 [24]),
    .Y(_3653_)
);

OAI21X1 _12952_ (
    .A(vdd),
    .B(_3652_),
    .C(_3653_),
    .Y(_3605_[24])
);

INVX1 _12953_ (
    .A(_2_[25]),
    .Y(_3654_)
);

NAND2X1 _12954_ (
    .A(vdd),
    .B(\datapath_1.rd2 [25]),
    .Y(_3655_)
);

OAI21X1 _12955_ (
    .A(vdd),
    .B(_3654_),
    .C(_3655_),
    .Y(_3605_[25])
);

INVX1 _12956_ (
    .A(_2_[26]),
    .Y(_3656_)
);

NAND2X1 _12957_ (
    .A(vdd),
    .B(\datapath_1.rd2 [26]),
    .Y(_3657_)
);

OAI21X1 _12958_ (
    .A(vdd),
    .B(_3656_),
    .C(_3657_),
    .Y(_3605_[26])
);

INVX1 _12959_ (
    .A(_2_[27]),
    .Y(_3658_)
);

NAND2X1 _12960_ (
    .A(vdd),
    .B(\datapath_1.rd2 [27]),
    .Y(_3659_)
);

OAI21X1 _12961_ (
    .A(vdd),
    .B(_3658_),
    .C(_3659_),
    .Y(_3605_[27])
);

INVX1 _12962_ (
    .A(_2_[28]),
    .Y(_3660_)
);

NAND2X1 _12963_ (
    .A(vdd),
    .B(\datapath_1.rd2 [28]),
    .Y(_3661_)
);

OAI21X1 _12964_ (
    .A(vdd),
    .B(_3660_),
    .C(_3661_),
    .Y(_3605_[28])
);

INVX1 _12965_ (
    .A(_2_[29]),
    .Y(_3662_)
);

NAND2X1 _12966_ (
    .A(vdd),
    .B(\datapath_1.rd2 [29]),
    .Y(_3663_)
);

OAI21X1 _12967_ (
    .A(vdd),
    .B(_3662_),
    .C(_3663_),
    .Y(_3605_[29])
);

INVX1 _12968_ (
    .A(_2_[30]),
    .Y(_3664_)
);

NAND2X1 _12969_ (
    .A(vdd),
    .B(\datapath_1.rd2 [30]),
    .Y(_3665_)
);

OAI21X1 _12970_ (
    .A(vdd),
    .B(_3664_),
    .C(_3665_),
    .Y(_3605_[30])
);

INVX1 _12971_ (
    .A(_2_[31]),
    .Y(_3666_)
);

NAND2X1 _12972_ (
    .A(vdd),
    .B(\datapath_1.rd2 [31]),
    .Y(_3667_)
);

OAI21X1 _12973_ (
    .A(vdd),
    .B(_3666_),
    .C(_3667_),
    .Y(_3605_[31])
);

DFFSR _12974_ (
    .CLK(clk_bF$buf99),
    .D(_3605_[0]),
    .Q(_2_[0]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _12975_ (
    .CLK(clk_bF$buf98),
    .D(_3605_[1]),
    .Q(_2_[1]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _12976_ (
    .CLK(clk_bF$buf97),
    .D(_3605_[2]),
    .Q(_2_[2]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _12977_ (
    .CLK(clk_bF$buf96),
    .D(_3605_[3]),
    .Q(_2_[3]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _12978_ (
    .CLK(clk_bF$buf95),
    .D(_3605_[4]),
    .Q(_2_[4]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _12979_ (
    .CLK(clk_bF$buf94),
    .D(_3605_[5]),
    .Q(_2_[5]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _12980_ (
    .CLK(clk_bF$buf93),
    .D(_3605_[6]),
    .Q(_2_[6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _12981_ (
    .CLK(clk_bF$buf92),
    .D(_3605_[7]),
    .Q(_2_[7]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _12982_ (
    .CLK(clk_bF$buf91),
    .D(_3605_[8]),
    .Q(_2_[8]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _12983_ (
    .CLK(clk_bF$buf90),
    .D(_3605_[9]),
    .Q(_2_[9]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _12984_ (
    .CLK(clk_bF$buf89),
    .D(_3605_[10]),
    .Q(_2_[10]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _12985_ (
    .CLK(clk_bF$buf88),
    .D(_3605_[11]),
    .Q(_2_[11]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _12986_ (
    .CLK(clk_bF$buf87),
    .D(_3605_[12]),
    .Q(_2_[12]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _12987_ (
    .CLK(clk_bF$buf86),
    .D(_3605_[13]),
    .Q(_2_[13]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _12988_ (
    .CLK(clk_bF$buf85),
    .D(_3605_[14]),
    .Q(_2_[14]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _12989_ (
    .CLK(clk_bF$buf84),
    .D(_3605_[15]),
    .Q(_2_[15]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _12990_ (
    .CLK(clk_bF$buf83),
    .D(_3605_[16]),
    .Q(_2_[16]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _12991_ (
    .CLK(clk_bF$buf82),
    .D(_3605_[17]),
    .Q(_2_[17]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _12992_ (
    .CLK(clk_bF$buf81),
    .D(_3605_[18]),
    .Q(_2_[18]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _12993_ (
    .CLK(clk_bF$buf80),
    .D(_3605_[19]),
    .Q(_2_[19]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _12994_ (
    .CLK(clk_bF$buf79),
    .D(_3605_[20]),
    .Q(_2_[20]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _12995_ (
    .CLK(clk_bF$buf78),
    .D(_3605_[21]),
    .Q(_2_[21]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _12996_ (
    .CLK(clk_bF$buf77),
    .D(_3605_[22]),
    .Q(_2_[22]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _12997_ (
    .CLK(clk_bF$buf76),
    .D(_3605_[23]),
    .Q(_2_[23]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _12998_ (
    .CLK(clk_bF$buf75),
    .D(_3605_[24]),
    .Q(_2_[24]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _12999_ (
    .CLK(clk_bF$buf74),
    .D(_3605_[25]),
    .Q(_2_[25]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _13000_ (
    .CLK(clk_bF$buf73),
    .D(_3605_[26]),
    .Q(_2_[26]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _13001_ (
    .CLK(clk_bF$buf72),
    .D(_3605_[27]),
    .Q(_2_[27]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _13002_ (
    .CLK(clk_bF$buf71),
    .D(_3605_[28]),
    .Q(_2_[28]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _13003_ (
    .CLK(clk_bF$buf70),
    .D(_3605_[29]),
    .Q(_2_[29]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _13004_ (
    .CLK(clk_bF$buf69),
    .D(_3605_[30]),
    .Q(_2_[30]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _13005_ (
    .CLK(clk_bF$buf68),
    .D(_3605_[31]),
    .Q(_2_[31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

INVX1 _13006_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3733_)
);

NAND2X1 _13007_ (
    .A(\datapath_1.mux_pcsrc.dout [0]),
    .B(PCEn_bF$buf7),
    .Y(_3734_)
);

OAI21X1 _13008_ (
    .A(PCEn_bF$buf6),
    .B(_3733_),
    .C(_3734_),
    .Y(_3670_[0])
);

INVX1 _13009_ (
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_3671_)
);

NAND2X1 _13010_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [1]),
    .Y(_3672_)
);

OAI21X1 _13011_ (
    .A(PCEn_bF$buf4),
    .B(_3671_),
    .C(_3672_),
    .Y(_3670_[1])
);

INVX1 _13012_ (
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_3673_)
);

NAND2X1 _13013_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [2]),
    .Y(_3674_)
);

OAI21X1 _13014_ (
    .A(PCEn_bF$buf2),
    .B(_3673_),
    .C(_3674_),
    .Y(_3670_[2])
);

INVX1 _13015_ (
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_3675_)
);

NAND2X1 _13016_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [3]),
    .Y(_3676_)
);

OAI21X1 _13017_ (
    .A(PCEn_bF$buf0),
    .B(_3675_),
    .C(_3676_),
    .Y(_3670_[3])
);

INVX1 _13018_ (
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_3677_)
);

NAND2X1 _13019_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [4]),
    .Y(_3678_)
);

OAI21X1 _13020_ (
    .A(PCEn_bF$buf6),
    .B(_3677_),
    .C(_3678_),
    .Y(_3670_[4])
);

INVX1 _13021_ (
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_3679_)
);

NAND2X1 _13022_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [5]),
    .Y(_3680_)
);

OAI21X1 _13023_ (
    .A(PCEn_bF$buf4),
    .B(_3679_),
    .C(_3680_),
    .Y(_3670_[5])
);

INVX1 _13024_ (
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_3681_)
);

NAND2X1 _13025_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [6]),
    .Y(_3682_)
);

OAI21X1 _13026_ (
    .A(PCEn_bF$buf2),
    .B(_3681_),
    .C(_3682_),
    .Y(_3670_[6])
);

INVX1 _13027_ (
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_3683_)
);

NAND2X1 _13028_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [7]),
    .Y(_3684_)
);

OAI21X1 _13029_ (
    .A(PCEn_bF$buf0),
    .B(_3683_),
    .C(_3684_),
    .Y(_3670_[7])
);

INVX1 _13030_ (
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_3685_)
);

NAND2X1 _13031_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [8]),
    .Y(_3686_)
);

OAI21X1 _13032_ (
    .A(PCEn_bF$buf6),
    .B(_3685_),
    .C(_3686_),
    .Y(_3670_[8])
);

INVX1 _13033_ (
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_3687_)
);

NAND2X1 _13034_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [9]),
    .Y(_3688_)
);

OAI21X1 _13035_ (
    .A(PCEn_bF$buf4),
    .B(_3687_),
    .C(_3688_),
    .Y(_3670_[9])
);

INVX1 _13036_ (
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_3689_)
);

NAND2X1 _13037_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [10]),
    .Y(_3690_)
);

OAI21X1 _13038_ (
    .A(PCEn_bF$buf2),
    .B(_3689_),
    .C(_3690_),
    .Y(_3670_[10])
);

INVX1 _13039_ (
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_3691_)
);

NAND2X1 _13040_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [11]),
    .Y(_3692_)
);

OAI21X1 _13041_ (
    .A(PCEn_bF$buf0),
    .B(_3691_),
    .C(_3692_),
    .Y(_3670_[11])
);

INVX1 _13042_ (
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_3693_)
);

NAND2X1 _13043_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [12]),
    .Y(_3694_)
);

OAI21X1 _13044_ (
    .A(PCEn_bF$buf6),
    .B(_3693_),
    .C(_3694_),
    .Y(_3670_[12])
);

INVX1 _13045_ (
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_3695_)
);

NAND2X1 _13046_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [13]),
    .Y(_3696_)
);

OAI21X1 _13047_ (
    .A(PCEn_bF$buf4),
    .B(_3695_),
    .C(_3696_),
    .Y(_3670_[13])
);

INVX1 _13048_ (
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_3697_)
);

NAND2X1 _13049_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [14]),
    .Y(_3698_)
);

OAI21X1 _13050_ (
    .A(PCEn_bF$buf2),
    .B(_3697_),
    .C(_3698_),
    .Y(_3670_[14])
);

INVX1 _13051_ (
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_3699_)
);

NAND2X1 _13052_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [15]),
    .Y(_3700_)
);

OAI21X1 _13053_ (
    .A(PCEn_bF$buf0),
    .B(_3699_),
    .C(_3700_),
    .Y(_3670_[15])
);

INVX1 _13054_ (
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_3701_)
);

NAND2X1 _13055_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [16]),
    .Y(_3702_)
);

OAI21X1 _13056_ (
    .A(PCEn_bF$buf6),
    .B(_3701_),
    .C(_3702_),
    .Y(_3670_[16])
);

INVX1 _13057_ (
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3703_)
);

NAND2X1 _13058_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [17]),
    .Y(_3704_)
);

OAI21X1 _13059_ (
    .A(PCEn_bF$buf4),
    .B(_3703_),
    .C(_3704_),
    .Y(_3670_[17])
);

INVX1 _13060_ (
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3705_)
);

NAND2X1 _13061_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [18]),
    .Y(_3706_)
);

OAI21X1 _13062_ (
    .A(PCEn_bF$buf2),
    .B(_3705_),
    .C(_3706_),
    .Y(_3670_[18])
);

INVX1 _13063_ (
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3707_)
);

NAND2X1 _13064_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [19]),
    .Y(_3708_)
);

OAI21X1 _13065_ (
    .A(PCEn_bF$buf0),
    .B(_3707_),
    .C(_3708_),
    .Y(_3670_[19])
);

INVX1 _13066_ (
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3709_)
);

NAND2X1 _13067_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [20]),
    .Y(_3710_)
);

OAI21X1 _13068_ (
    .A(PCEn_bF$buf6),
    .B(_3709_),
    .C(_3710_),
    .Y(_3670_[20])
);

INVX1 _13069_ (
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3711_)
);

NAND2X1 _13070_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [21]),
    .Y(_3712_)
);

OAI21X1 _13071_ (
    .A(PCEn_bF$buf4),
    .B(_3711_),
    .C(_3712_),
    .Y(_3670_[21])
);

INVX1 _13072_ (
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3713_)
);

NAND2X1 _13073_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [22]),
    .Y(_3714_)
);

OAI21X1 _13074_ (
    .A(PCEn_bF$buf2),
    .B(_3713_),
    .C(_3714_),
    .Y(_3670_[22])
);

INVX1 _13075_ (
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3715_)
);

NAND2X1 _13076_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [23]),
    .Y(_3716_)
);

OAI21X1 _13077_ (
    .A(PCEn_bF$buf0),
    .B(_3715_),
    .C(_3716_),
    .Y(_3670_[23])
);

INVX1 _13078_ (
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3717_)
);

NAND2X1 _13079_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [24]),
    .Y(_3718_)
);

OAI21X1 _13080_ (
    .A(PCEn_bF$buf6),
    .B(_3717_),
    .C(_3718_),
    .Y(_3670_[24])
);

INVX1 _13081_ (
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3719_)
);

NAND2X1 _13082_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [25]),
    .Y(_3720_)
);

OAI21X1 _13083_ (
    .A(PCEn_bF$buf4),
    .B(_3719_),
    .C(_3720_),
    .Y(_3670_[25])
);

INVX1 _13084_ (
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3721_)
);

NAND2X1 _13085_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [26]),
    .Y(_3722_)
);

OAI21X1 _13086_ (
    .A(PCEn_bF$buf2),
    .B(_3721_),
    .C(_3722_),
    .Y(_3670_[26])
);

INVX1 _13087_ (
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3723_)
);

NAND2X1 _13088_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [27]),
    .Y(_3724_)
);

OAI21X1 _13089_ (
    .A(PCEn_bF$buf0),
    .B(_3723_),
    .C(_3724_),
    .Y(_3670_[27])
);

INVX1 _13090_ (
    .A(\datapath_1.PCJump [28]),
    .Y(_3725_)
);

NAND2X1 _13091_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [28]),
    .Y(_3726_)
);

OAI21X1 _13092_ (
    .A(PCEn_bF$buf6),
    .B(_3725_),
    .C(_3726_),
    .Y(_3670_[28])
);

INVX1 _13093_ (
    .A(\datapath_1.PCJump [29]),
    .Y(_3727_)
);

NAND2X1 _13094_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [29]),
    .Y(_3728_)
);

OAI21X1 _13095_ (
    .A(PCEn_bF$buf4),
    .B(_3727_),
    .C(_3728_),
    .Y(_3670_[29])
);

INVX1 _13096_ (
    .A(\datapath_1.PCJump [30]),
    .Y(_3729_)
);

NAND2X1 _13097_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [30]),
    .Y(_3730_)
);

OAI21X1 _13098_ (
    .A(PCEn_bF$buf2),
    .B(_3729_),
    .C(_3730_),
    .Y(_3670_[30])
);

INVX1 _13099_ (
    .A(\datapath_1.PCJump [31]),
    .Y(_3731_)
);

NAND2X1 _13100_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [31]),
    .Y(_3732_)
);

OAI21X1 _13101_ (
    .A(PCEn_bF$buf0),
    .B(_3731_),
    .C(_3732_),
    .Y(_3670_[31])
);

DFFSR _13102_ (
    .CLK(clk_bF$buf67),
    .D(_3670_[0]),
    .Q(\datapath_1.mux_iord.din0 [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _13103_ (
    .CLK(clk_bF$buf66),
    .D(_3670_[1]),
    .Q(\datapath_1.mux_iord.din0 [1]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _13104_ (
    .CLK(clk_bF$buf65),
    .D(_3670_[2]),
    .Q(\datapath_1.mux_iord.din0 [2]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _13105_ (
    .CLK(clk_bF$buf64),
    .D(_3670_[3]),
    .Q(\datapath_1.mux_iord.din0 [3]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _13106_ (
    .CLK(clk_bF$buf63),
    .D(_3670_[4]),
    .Q(\datapath_1.mux_iord.din0 [4]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _13107_ (
    .CLK(clk_bF$buf62),
    .D(_3670_[5]),
    .Q(\datapath_1.mux_iord.din0 [5]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _13108_ (
    .CLK(clk_bF$buf61),
    .D(_3670_[6]),
    .Q(\datapath_1.mux_iord.din0 [6]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _13109_ (
    .CLK(clk_bF$buf60),
    .D(_3670_[7]),
    .Q(\datapath_1.mux_iord.din0 [7]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _13110_ (
    .CLK(clk_bF$buf59),
    .D(_3670_[8]),
    .Q(\datapath_1.mux_iord.din0 [8]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _13111_ (
    .CLK(clk_bF$buf58),
    .D(_3670_[9]),
    .Q(\datapath_1.mux_iord.din0 [9]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _13112_ (
    .CLK(clk_bF$buf57),
    .D(_3670_[10]),
    .Q(\datapath_1.mux_iord.din0 [10]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _13113_ (
    .CLK(clk_bF$buf56),
    .D(_3670_[11]),
    .Q(\datapath_1.mux_iord.din0 [11]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _13114_ (
    .CLK(clk_bF$buf55),
    .D(_3670_[12]),
    .Q(\datapath_1.mux_iord.din0 [12]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _13115_ (
    .CLK(clk_bF$buf54),
    .D(_3670_[13]),
    .Q(\datapath_1.mux_iord.din0 [13]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _13116_ (
    .CLK(clk_bF$buf53),
    .D(_3670_[14]),
    .Q(\datapath_1.mux_iord.din0 [14]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _13117_ (
    .CLK(clk_bF$buf52),
    .D(_3670_[15]),
    .Q(\datapath_1.mux_iord.din0 [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _13118_ (
    .CLK(clk_bF$buf51),
    .D(_3670_[16]),
    .Q(\datapath_1.mux_iord.din0 [16]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _13119_ (
    .CLK(clk_bF$buf50),
    .D(_3670_[17]),
    .Q(\datapath_1.mux_iord.din0 [17]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _13120_ (
    .CLK(clk_bF$buf49),
    .D(_3670_[18]),
    .Q(\datapath_1.mux_iord.din0 [18]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _13121_ (
    .CLK(clk_bF$buf48),
    .D(_3670_[19]),
    .Q(\datapath_1.mux_iord.din0 [19]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _13122_ (
    .CLK(clk_bF$buf47),
    .D(_3670_[20]),
    .Q(\datapath_1.mux_iord.din0 [20]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _13123_ (
    .CLK(clk_bF$buf46),
    .D(_3670_[21]),
    .Q(\datapath_1.mux_iord.din0 [21]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _13124_ (
    .CLK(clk_bF$buf45),
    .D(_3670_[22]),
    .Q(\datapath_1.mux_iord.din0 [22]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _13125_ (
    .CLK(clk_bF$buf44),
    .D(_3670_[23]),
    .Q(\datapath_1.mux_iord.din0 [23]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _13126_ (
    .CLK(clk_bF$buf43),
    .D(_3670_[24]),
    .Q(\datapath_1.mux_iord.din0 [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _13127_ (
    .CLK(clk_bF$buf42),
    .D(_3670_[25]),
    .Q(\datapath_1.mux_iord.din0 [25]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _13128_ (
    .CLK(clk_bF$buf41),
    .D(_3670_[26]),
    .Q(\datapath_1.mux_iord.din0 [26]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _13129_ (
    .CLK(clk_bF$buf40),
    .D(_3670_[27]),
    .Q(\datapath_1.mux_iord.din0 [27]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _13130_ (
    .CLK(clk_bF$buf39),
    .D(_3670_[28]),
    .Q(\datapath_1.PCJump [28]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _13131_ (
    .CLK(clk_bF$buf38),
    .D(_3670_[29]),
    .Q(\datapath_1.PCJump [29]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _13132_ (
    .CLK(clk_bF$buf37),
    .D(_3670_[30]),
    .Q(\datapath_1.PCJump [30]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _13133_ (
    .CLK(clk_bF$buf36),
    .D(_3670_[31]),
    .Q(\datapath_1.PCJump [31]),
    .R(rst_bF$buf36),
    .S(vdd)
);

INVX4 _13134_ (
    .A(\datapath_1.a3 [4]),
    .Y(_3735_)
);

INVX1 _13135_ (
    .A(\datapath_1.a3 [0]),
    .Y(_3736_)
);

NOR2X1 _13136_ (
    .A(\datapath_1.a3 [1]),
    .B(_3736_),
    .Y(_3737_)
);

NAND2X1 _13137_ (
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_3738_)
);

INVX1 _13138_ (
    .A(_3738_),
    .Y(_3739_)
);

NAND2X1 _13139_ (
    .A(_3739_),
    .B(_3737_),
    .Y(_3740_)
);

INVX1 _13140_ (
    .A(\datapath_1.a3 [3]),
    .Y(_3741_)
);

NOR2X1 _13141_ (
    .A(\datapath_1.a3 [2]),
    .B(_3741_),
    .Y(_3742_)
);

NAND2X1 _13142_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_3743_)
);

INVX1 _13143_ (
    .A(_3743_),
    .Y(_3744_)
);

NAND2X1 _13144_ (
    .A(_3744_),
    .B(_3742_),
    .Y(_3745_)
);

AOI21X1 _13145_ (
    .A(_3740_),
    .B(_3745_),
    .C(_3735_),
    .Y(_3746_)
);

INVX2 _13146_ (
    .A(\datapath_1.a3 [1]),
    .Y(_3747_)
);

NOR2X1 _13147_ (
    .A(\datapath_1.a3 [0]),
    .B(_3747_),
    .Y(_3748_)
);

NOR2X1 _13148_ (
    .A(_3748_),
    .B(_3737_),
    .Y(_3749_)
);

NAND2X1 _13149_ (
    .A(\datapath_1.a3 [4]),
    .B(_3742_),
    .Y(_3750_)
);

NAND2X1 _13150_ (
    .A(\datapath_1.a3 [4]),
    .B(_3739_),
    .Y(_3751_)
);

OAI22X1 _13151_ (
    .A(_3737_),
    .B(_3751_),
    .C(_3750_),
    .D(_3749_),
    .Y(_3752_)
);

NOR2X1 _13152_ (
    .A(_3746_),
    .B(_3752_),
    .Y(_3753_)
);

NOR2X1 _13153_ (
    .A(\datapath_1.a3 [0]),
    .B(\datapath_1.a3 [1]),
    .Y(_3754_)
);

INVX1 _13154_ (
    .A(\datapath_1.a3 [2]),
    .Y(_3755_)
);

NOR2X1 _13155_ (
    .A(\datapath_1.a3 [3]),
    .B(_3755_),
    .Y(_3756_)
);

INVX2 _13156_ (
    .A(_3756_),
    .Y(_3757_)
);

NAND2X1 _13157_ (
    .A(_3754_),
    .B(_3742_),
    .Y(_3758_)
);

OAI21X1 _13158_ (
    .A(_3754_),
    .B(_3757_),
    .C(_3758_),
    .Y(_3759_)
);

INVX1 _13159_ (
    .A(_3754_),
    .Y(_3760_)
);

NAND2X1 _13160_ (
    .A(_3741_),
    .B(_3755_),
    .Y(_3761_)
);

INVX1 _13161_ (
    .A(_3761_),
    .Y(_3762_)
);

OAI21X1 _13162_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .C(_3762_),
    .Y(_3763_)
);

OAI21X1 _13163_ (
    .A(_3760_),
    .B(_3757_),
    .C(_3763_),
    .Y(_3764_)
);

OAI21X1 _13164_ (
    .A(_3759_),
    .B(_3764_),
    .C(\datapath_1.a3 [4]),
    .Y(_3765_)
);

NAND2X1 _13165_ (
    .A(_3753_),
    .B(_3765_),
    .Y(_3766_)
);

NOR2X1 _13166_ (
    .A(_3738_),
    .B(_3743_),
    .Y(_3767_)
);

NOR2X1 _13167_ (
    .A(_3761_),
    .B(_3760_),
    .Y(_3768_)
);

MUX2X1 _13168_ (
    .A(_3768_),
    .B(_3767_),
    .S(\datapath_1.a3 [4]),
    .Y(_3769_)
);

NAND2X1 _13169_ (
    .A(_3735_),
    .B(_3739_),
    .Y(_3770_)
);

OR2X2 _13170_ (
    .A(_3749_),
    .B(_3770_),
    .Y(_3771_)
);

AND2X2 _13171_ (
    .A(_3771_),
    .B(_3769_),
    .Y(_3772_)
);

INVX1 _13172_ (
    .A(_3749_),
    .Y(_3773_)
);

INVX1 _13173_ (
    .A(_3742_),
    .Y(_3774_)
);

NOR2X1 _13174_ (
    .A(\datapath_1.a3 [4]),
    .B(_3774_),
    .Y(_3775_)
);

NAND2X1 _13175_ (
    .A(_3754_),
    .B(_3739_),
    .Y(_3776_)
);

AOI21X1 _13176_ (
    .A(_3745_),
    .B(_3776_),
    .C(\datapath_1.a3 [4]),
    .Y(_3777_)
);

AOI21X1 _13177_ (
    .A(_3773_),
    .B(_3775_),
    .C(_3777_),
    .Y(_3778_)
);

NAND2X1 _13178_ (
    .A(_3778_),
    .B(_3772_),
    .Y(_3779_)
);

INVX2 _13179_ (
    .A(RegWrite_bF$buf7),
    .Y(_3780_)
);

NAND2X1 _13180_ (
    .A(\datapath_1.a3 [4]),
    .B(RegWrite_bF$buf6),
    .Y(_3781_)
);

NAND2X1 _13181_ (
    .A(_3754_),
    .B(_3756_),
    .Y(_3782_)
);

OAI21X1 _13182_ (
    .A(_3743_),
    .B(_3761_),
    .C(_3782_),
    .Y(_3783_)
);

OAI21X1 _13183_ (
    .A(_3780_),
    .B(_3783_),
    .C(_3781_),
    .Y(_3784_)
);

NAND2X1 _13184_ (
    .A(_3735_),
    .B(_3759_),
    .Y(_3785_)
);

INVX1 _13185_ (
    .A(_3748_),
    .Y(_3786_)
);

NOR2X1 _13186_ (
    .A(_3761_),
    .B(_3786_),
    .Y(_3787_)
);

OAI21X1 _13187_ (
    .A(_3768_),
    .B(_3787_),
    .C(_3735_),
    .Y(_3788_)
);

NAND3X1 _13188_ (
    .A(_3785_),
    .B(_3788_),
    .C(_3784_),
    .Y(_3789_)
);

OR2X2 _13189_ (
    .A(_3779_),
    .B(_3789_),
    .Y(_3790_)
);

NOR2X1 _13190_ (
    .A(_3766_),
    .B(_3790_),
    .Y(\datapath_1.regfile_1.regEn [1])
);

NOR2X1 _13191_ (
    .A(\datapath_1.a3 [4]),
    .B(_3761_),
    .Y(_3791_)
);

AOI22X1 _13192_ (
    .A(_3747_),
    .B(_3791_),
    .C(_3735_),
    .D(_3759_),
    .Y(_3792_)
);

NAND2X1 _13193_ (
    .A(_3784_),
    .B(_3792_),
    .Y(_3793_)
);

OR2X2 _13194_ (
    .A(_3779_),
    .B(_3793_),
    .Y(_3794_)
);

NOR2X1 _13195_ (
    .A(_3766_),
    .B(_3794_),
    .Y(\datapath_1.regfile_1.regEn [2])
);

INVX1 _13196_ (
    .A(_3782_),
    .Y(_3795_)
);

OAI21X1 _13197_ (
    .A(_3795_),
    .B(_3787_),
    .C(_3735_),
    .Y(_3796_)
);

NAND3X1 _13198_ (
    .A(RegWrite_bF$buf5),
    .B(_3796_),
    .C(_3792_),
    .Y(_3797_)
);

OR2X2 _13199_ (
    .A(_3779_),
    .B(_3797_),
    .Y(_3798_)
);

NOR2X1 _13200_ (
    .A(_3766_),
    .B(_3798_),
    .Y(\datapath_1.regfile_1.regEn [3])
);

NOR2X1 _13201_ (
    .A(_3780_),
    .B(_3791_),
    .Y(_3799_)
);

NAND2X1 _13202_ (
    .A(_3799_),
    .B(_3785_),
    .Y(_3800_)
);

OR2X2 _13203_ (
    .A(_3779_),
    .B(_3800_),
    .Y(_3801_)
);

NOR2X1 _13204_ (
    .A(_3766_),
    .B(_3801_),
    .Y(\datapath_1.regfile_1.regEn [4])
);

OAI21X1 _13205_ (
    .A(_3743_),
    .B(_3757_),
    .C(_3758_),
    .Y(_3802_)
);

NOR2X1 _13206_ (
    .A(_3757_),
    .B(_3786_),
    .Y(_3803_)
);

OAI21X1 _13207_ (
    .A(_3795_),
    .B(_3803_),
    .C(_3735_),
    .Y(_3804_)
);

NAND2X1 _13208_ (
    .A(_3799_),
    .B(_3804_),
    .Y(_3805_)
);

AOI21X1 _13209_ (
    .A(_3735_),
    .B(_3802_),
    .C(_3805_),
    .Y(_3806_)
);

NOR2X1 _13210_ (
    .A(_3766_),
    .B(_3779_),
    .Y(_3807_)
);

AND2X2 _13211_ (
    .A(_3807_),
    .B(_3806_),
    .Y(\datapath_1.regfile_1.regEn [5])
);

INVX1 _13212_ (
    .A(_3802_),
    .Y(_3808_)
);

NAND3X1 _13213_ (
    .A(_3735_),
    .B(_3747_),
    .C(_3756_),
    .Y(_3809_)
);

AND2X2 _13214_ (
    .A(_3799_),
    .B(_3809_),
    .Y(_3810_)
);

OAI21X1 _13215_ (
    .A(\datapath_1.a3 [4]),
    .B(_3808_),
    .C(_3810_),
    .Y(_3811_)
);

OR2X2 _13216_ (
    .A(_3779_),
    .B(_3811_),
    .Y(_3812_)
);

NOR2X1 _13217_ (
    .A(_3766_),
    .B(_3812_),
    .Y(\datapath_1.regfile_1.regEn [6])
);

INVX1 _13218_ (
    .A(_3758_),
    .Y(_3813_)
);

OAI21X1 _13219_ (
    .A(_3813_),
    .B(_3803_),
    .C(_3735_),
    .Y(_3814_)
);

AND2X2 _13220_ (
    .A(_3810_),
    .B(_3814_),
    .Y(_3815_)
);

AND2X2 _13221_ (
    .A(_3807_),
    .B(_3815_),
    .Y(\datapath_1.regfile_1.regEn [7])
);

OAI21X1 _13222_ (
    .A(_3741_),
    .B(_3780_),
    .C(_3781_),
    .Y(_3816_)
);

INVX1 _13223_ (
    .A(_3816_),
    .Y(_3817_)
);

OR2X2 _13224_ (
    .A(_3766_),
    .B(_3817_),
    .Y(_3818_)
);

NOR2X1 _13225_ (
    .A(_3779_),
    .B(_3818_),
    .Y(\datapath_1.regfile_1.regEn [8])
);

OAI21X1 _13226_ (
    .A(_3749_),
    .B(_3770_),
    .C(_3769_),
    .Y(_3819_)
);

NOR2X1 _13227_ (
    .A(_3777_),
    .B(_3819_),
    .Y(_3820_)
);

NOR2X1 _13228_ (
    .A(_3774_),
    .B(_3786_),
    .Y(_3821_)
);

OAI21X1 _13229_ (
    .A(_3813_),
    .B(_3821_),
    .C(_3735_),
    .Y(_3822_)
);

NAND2X1 _13230_ (
    .A(_3822_),
    .B(_3820_),
    .Y(_3823_)
);

NOR2X1 _13231_ (
    .A(_3823_),
    .B(_3818_),
    .Y(\datapath_1.regfile_1.regEn [9])
);

AOI21X1 _13232_ (
    .A(_3775_),
    .B(_3747_),
    .C(_3817_),
    .Y(_3824_)
);

NAND2X1 _13233_ (
    .A(_3824_),
    .B(_3820_),
    .Y(_3825_)
);

NOR2X1 _13234_ (
    .A(_3766_),
    .B(_3825_),
    .Y(\datapath_1.regfile_1.regEn [10])
);

INVX1 _13235_ (
    .A(_3776_),
    .Y(_3826_)
);

OAI21X1 _13236_ (
    .A(_3826_),
    .B(_3821_),
    .C(_3735_),
    .Y(_3827_)
);

NAND3X1 _13237_ (
    .A(_3824_),
    .B(_3827_),
    .C(_3772_),
    .Y(_3828_)
);

NOR2X1 _13238_ (
    .A(_3766_),
    .B(_3828_),
    .Y(\datapath_1.regfile_1.regEn [11])
);

NAND2X1 _13239_ (
    .A(_3816_),
    .B(_3769_),
    .Y(_3829_)
);

NOR2X1 _13240_ (
    .A(_3775_),
    .B(_3829_),
    .Y(_3830_)
);

OAI21X1 _13241_ (
    .A(_3749_),
    .B(_3770_),
    .C(_3830_),
    .Y(_3831_)
);

NOR2X1 _13242_ (
    .A(_3766_),
    .B(_3831_),
    .Y(\datapath_1.regfile_1.regEn [12])
);

OAI21X1 _13243_ (
    .A(\datapath_1.a3 [0]),
    .B(_3770_),
    .C(_3830_),
    .Y(_3832_)
);

NOR2X1 _13244_ (
    .A(_3766_),
    .B(_3832_),
    .Y(\datapath_1.regfile_1.regEn [13])
);

NOR2X1 _13245_ (
    .A(\datapath_1.a3 [1]),
    .B(_3738_),
    .Y(_3833_)
);

INVX1 _13246_ (
    .A(_3833_),
    .Y(_3834_)
);

OAI21X1 _13247_ (
    .A(\datapath_1.a3 [4]),
    .B(_3834_),
    .C(_3830_),
    .Y(_3835_)
);

NOR2X1 _13248_ (
    .A(_3766_),
    .B(_3835_),
    .Y(\datapath_1.regfile_1.regEn [14])
);

NAND2X1 _13249_ (
    .A(_3735_),
    .B(_3767_),
    .Y(_3836_)
);

NOR2X1 _13250_ (
    .A(_3780_),
    .B(_3836_),
    .Y(\datapath_1.regfile_1.regEn [15])
);

INVX2 _13251_ (
    .A(_3781_),
    .Y(_3837_)
);

NAND2X1 _13252_ (
    .A(_3837_),
    .B(_3768_),
    .Y(_3838_)
);

INVX8 _13253_ (
    .A(_3838_),
    .Y(\datapath_1.regfile_1.regEn [16])
);

NAND2X1 _13254_ (
    .A(_3737_),
    .B(_3762_),
    .Y(_3839_)
);

NOR2X1 _13255_ (
    .A(_3781_),
    .B(_3839_),
    .Y(\datapath_1.regfile_1.regEn [17])
);

AND2X2 _13256_ (
    .A(_3787_),
    .B(_3837_),
    .Y(\datapath_1.regfile_1.regEn [18])
);

NAND2X1 _13257_ (
    .A(_3744_),
    .B(_3762_),
    .Y(_3840_)
);

NOR2X1 _13258_ (
    .A(_3781_),
    .B(_3840_),
    .Y(\datapath_1.regfile_1.regEn [19])
);

NOR2X1 _13259_ (
    .A(_3781_),
    .B(_3782_),
    .Y(\datapath_1.regfile_1.regEn [20])
);

INVX1 _13260_ (
    .A(_3753_),
    .Y(_3841_)
);

AOI21X1 _13261_ (
    .A(_3736_),
    .B(_3756_),
    .C(_3802_),
    .Y(_3842_)
);

NAND3X1 _13262_ (
    .A(_3837_),
    .B(_3761_),
    .C(_3842_),
    .Y(_3843_)
);

NOR2X1 _13263_ (
    .A(_3843_),
    .B(_3841_),
    .Y(\datapath_1.regfile_1.regEn [21])
);

NAND2X1 _13264_ (
    .A(\datapath_1.a3 [4]),
    .B(_3803_),
    .Y(_3844_)
);

NOR2X1 _13265_ (
    .A(_3780_),
    .B(_3844_),
    .Y(\datapath_1.regfile_1.regEn [22])
);

OAI21X1 _13266_ (
    .A(_3760_),
    .B(_3774_),
    .C(_3837_),
    .Y(_3845_)
);

INVX1 _13267_ (
    .A(_3845_),
    .Y(_3846_)
);

AOI22X1 _13268_ (
    .A(\datapath_1.a3 [4]),
    .B(_3762_),
    .C(_3747_),
    .D(_3756_),
    .Y(_3847_)
);

NAND3X1 _13269_ (
    .A(_3847_),
    .B(_3846_),
    .C(_3844_),
    .Y(_3848_)
);

NOR2X1 _13270_ (
    .A(_3848_),
    .B(_3841_),
    .Y(\datapath_1.regfile_1.regEn [23])
);

NOR2X1 _13271_ (
    .A(_3781_),
    .B(_3758_),
    .Y(\datapath_1.regfile_1.regEn [24])
);

INVX1 _13272_ (
    .A(_3821_),
    .Y(_3849_)
);

AOI21X1 _13273_ (
    .A(_3849_),
    .B(\datapath_1.a3 [3]),
    .C(_3735_),
    .Y(_3850_)
);

OR2X2 _13274_ (
    .A(_3850_),
    .B(_3746_),
    .Y(_3851_)
);

OAI21X1 _13275_ (
    .A(_3737_),
    .B(_3751_),
    .C(_3846_),
    .Y(_3852_)
);

NOR2X1 _13276_ (
    .A(_3852_),
    .B(_3851_),
    .Y(\datapath_1.regfile_1.regEn [25])
);

NOR2X1 _13277_ (
    .A(_3781_),
    .B(_3849_),
    .Y(\datapath_1.regfile_1.regEn [26])
);

NAND3X1 _13278_ (
    .A(_3837_),
    .B(\datapath_1.a3 [3]),
    .C(_3751_),
    .Y(_3853_)
);

OR2X2 _13279_ (
    .A(_3821_),
    .B(_3853_),
    .Y(_3854_)
);

OAI21X1 _13280_ (
    .A(\datapath_1.a3 [1]),
    .B(_3750_),
    .C(_3740_),
    .Y(_3855_)
);

NOR2X1 _13281_ (
    .A(_3855_),
    .B(_3854_),
    .Y(\datapath_1.regfile_1.regEn [27])
);

NAND2X1 _13282_ (
    .A(\datapath_1.a3 [4]),
    .B(_3767_),
    .Y(_3856_)
);

NAND2X1 _13283_ (
    .A(RegWrite_bF$buf4),
    .B(_3856_),
    .Y(_3857_)
);

INVX1 _13284_ (
    .A(_3751_),
    .Y(_3858_)
);

OAI21X1 _13285_ (
    .A(_3738_),
    .B(_3749_),
    .C(_3858_),
    .Y(_3859_)
);

NOR2X1 _13286_ (
    .A(_3857_),
    .B(_3859_),
    .Y(\datapath_1.regfile_1.regEn [28])
);

NOR2X1 _13287_ (
    .A(_3781_),
    .B(_3740_),
    .Y(\datapath_1.regfile_1.regEn [29])
);

NAND2X1 _13288_ (
    .A(\datapath_1.a3 [1]),
    .B(_3858_),
    .Y(_3860_)
);

NOR2X1 _13289_ (
    .A(_3857_),
    .B(_3860_),
    .Y(\datapath_1.regfile_1.regEn [30])
);

NOR2X1 _13290_ (
    .A(_3780_),
    .B(_3856_),
    .Y(\datapath_1.regfile_1.regEn [31])
);

INVX1 _13291_ (
    .A(\datapath_1.PCJump [18]),
    .Y(_3861_)
);

NOR2X1 _13292_ (
    .A(\datapath_1.PCJump [19]),
    .B(_3861_),
    .Y(_3862_)
);

NAND2X1 _13293_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3863_)
);

INVX2 _13294_ (
    .A(_3863_),
    .Y(_3864_)
);

NAND3X1 _13295_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3864_),
    .C(_3862_),
    .Y(_3865_)
);

INVX8 _13296_ (
    .A(_3865_),
    .Y(_3866_)
);

INVX1 _13297_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_3867_)
);

NOR2X1 _13298_ (
    .A(\datapath_1.PCJump [18]),
    .B(_3867_),
    .Y(_3868_)
);

NAND3X1 _13299_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3864_),
    .C(_3868_),
    .Y(_3869_)
);

INVX8 _13300_ (
    .A(_3869_),
    .Y(_3870_)
);

AOI22X1 _13301_ (
    .A(_3870__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [0]),
    .C(_3866__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_3871_)
);

INVX1 _13302_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_3872_)
);

NOR2X1 _13303_ (
    .A(\datapath_1.PCJump [21]),
    .B(_3872_),
    .Y(_3873_)
);

NOR3X1 _13304_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(\datapath_1.PCJump [18]),
    .C(\datapath_1.PCJump [19]),
    .Y(_3874_)
);

NAND2X1 _13305_ (
    .A(_3874_),
    .B(_3873_),
    .Y(_3875_)
);

INVX8 _13306_ (
    .A(_3875__bF$buf3),
    .Y(_3876_)
);

NOR2X1 _13307_ (
    .A(\datapath_1.PCJump [18]),
    .B(\datapath_1.PCJump [19]),
    .Y(_3877_)
);

AND2X2 _13308_ (
    .A(_3877_),
    .B(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_3878_)
);

AND2X2 _13309_ (
    .A(_3878_),
    .B(_3864_),
    .Y(_3879_)
);

AOI22X1 _13310_ (
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .B(_3876_),
    .C(\datapath_1.regfile_1.regOut[28] [0]),
    .D(_3879__bF$buf3),
    .Y(_3880_)
);

INVX1 _13311_ (
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_3881_)
);

INVX1 _13312_ (
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_3882_)
);

INVX4 _13313_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .Y(_3883_)
);

NAND2X1 _13314_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3884_)
);

NOR2X1 _13315_ (
    .A(_3884_),
    .B(_3863_),
    .Y(_3885_)
);

NAND2X1 _13316_ (
    .A(_3883_),
    .B(_3885_),
    .Y(_3886_)
);

AND2X2 _13317_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3887_)
);

NOR2X1 _13318_ (
    .A(\datapath_1.PCJump [20]),
    .B(\datapath_1.PCJump [21]),
    .Y(_3888_)
);

NAND3X1 _13319_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3888_),
    .C(_3887_),
    .Y(_3889_)
);

OAI22X1 _13320_ (
    .A(_3889__bF$buf4),
    .B(_3881_),
    .C(_3882_),
    .D(_3886__bF$buf3),
    .Y(_3890_)
);

INVX1 _13321_ (
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_3891_)
);

INVX1 _13322_ (
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_3892_)
);

NAND3X1 _13323_ (
    .A(_3883_),
    .B(_3873_),
    .C(_3868_),
    .Y(_3893_)
);

NAND2X1 _13324_ (
    .A(_3864_),
    .B(_3874_),
    .Y(_3894_)
);

OAI22X1 _13325_ (
    .A(_3894__bF$buf4),
    .B(_3891_),
    .C(_3892_),
    .D(_3893_),
    .Y(_3895_)
);

NOR2X1 _13326_ (
    .A(_3895_),
    .B(_3890_),
    .Y(_3896_)
);

NAND3X1 _13327_ (
    .A(_3880_),
    .B(_3871_),
    .C(_3896_),
    .Y(_3897_)
);

NAND3X1 _13328_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3887_),
    .C(_3873_),
    .Y(_3898_)
);

INVX8 _13329_ (
    .A(_3898_),
    .Y(_3899_)
);

INVX1 _13330_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_3900_)
);

NOR2X1 _13331_ (
    .A(\datapath_1.PCJump [20]),
    .B(_3900_),
    .Y(_3901_)
);

AND2X2 _13332_ (
    .A(_3878_),
    .B(_3901_),
    .Y(_3902_)
);

AOI22X1 _13333_ (
    .A(_3899__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [0]),
    .C(\datapath_1.regfile_1.regOut[24] [0]),
    .D(_3902__bF$buf4),
    .Y(_3903_)
);

AND2X2 _13334_ (
    .A(_3878_),
    .B(_3873_),
    .Y(_3904_)
);

NAND2X1 _13335_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3885_),
    .Y(_3905_)
);

INVX8 _13336_ (
    .A(_3905_),
    .Y(_3906_)
);

AOI22X1 _13337_ (
    .A(_3904__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [0]),
    .C(\datapath_1.regfile_1.regOut[31] [0]),
    .D(_3906__bF$buf3),
    .Y(_3907_)
);

INVX1 _13338_ (
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_3908_)
);

INVX1 _13339_ (
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_3909_)
);

NAND2X1 _13340_ (
    .A(_3888_),
    .B(_3874_),
    .Y(_3910_)
);

NAND2X1 _13341_ (
    .A(_3874_),
    .B(_3901_),
    .Y(_3911_)
);

OAI22X1 _13342_ (
    .A(_3908_),
    .B(_3910__bF$buf3),
    .C(_3909_),
    .D(_3911_),
    .Y(_3912_)
);

INVX1 _13343_ (
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_3913_)
);

INVX1 _13344_ (
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_3914_)
);

NAND3X1 _13345_ (
    .A(_3883_),
    .B(_3901_),
    .C(_3868_),
    .Y(_3915_)
);

NAND3X1 _13346_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3888_),
    .C(_3877_),
    .Y(_3916_)
);

OAI22X1 _13347_ (
    .A(_3916__bF$buf4),
    .B(_3913_),
    .C(_3914_),
    .D(_3915__bF$buf3),
    .Y(_3917_)
);

NOR2X1 _13348_ (
    .A(_3912_),
    .B(_3917_),
    .Y(_3918_)
);

NAND3X1 _13349_ (
    .A(_3907_),
    .B(_3903_),
    .C(_3918_),
    .Y(_3919_)
);

NOR2X1 _13350_ (
    .A(_3919_),
    .B(_3897_),
    .Y(_3920_)
);

INVX1 _13351_ (
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_3921_)
);

INVX1 _13352_ (
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .Y(_3922_)
);

NAND3X1 _13353_ (
    .A(_3883_),
    .B(_3888_),
    .C(_3887_),
    .Y(_3923_)
);

NAND3X1 _13354_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3901_),
    .C(_3868_),
    .Y(_3924_)
);

OAI22X1 _13355_ (
    .A(_3923__bF$buf4),
    .B(_3922_),
    .C(_3921_),
    .D(_3924__bF$buf3),
    .Y(_3925_)
);

INVX1 _13356_ (
    .A(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_3926_)
);

INVX1 _13357_ (
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .Y(_3927_)
);

NAND3X1 _13358_ (
    .A(_3883_),
    .B(_3887_),
    .C(_3873_),
    .Y(_3928_)
);

NAND3X1 _13359_ (
    .A(_3887_),
    .B(_3883_),
    .C(_3901_),
    .Y(_3929_)
);

OAI22X1 _13360_ (
    .A(_3927_),
    .B(_3928_),
    .C(_3929__bF$buf4),
    .D(_3926_),
    .Y(_3930_)
);

NOR2X1 _13361_ (
    .A(_3930_),
    .B(_3925_),
    .Y(_3931_)
);

INVX1 _13362_ (
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_3932_)
);

INVX1 _13363_ (
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_3933_)
);

NAND3X1 _13364_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3873_),
    .C(_3862_),
    .Y(_3934_)
);

NAND3X1 _13365_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3873_),
    .C(_3868_),
    .Y(_3935_)
);

OAI22X1 _13366_ (
    .A(_3933_),
    .B(_3934__bF$buf3),
    .C(_3935__bF$buf3),
    .D(_3932_),
    .Y(_3936_)
);

INVX1 _13367_ (
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_3937_)
);

INVX1 _13368_ (
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_3938_)
);

NAND3X1 _13369_ (
    .A(_3883_),
    .B(_3888_),
    .C(_3862_),
    .Y(_3939_)
);

NAND3X1 _13370_ (
    .A(_3883_),
    .B(_3888_),
    .C(_3868_),
    .Y(_3940_)
);

OAI22X1 _13371_ (
    .A(_3938_),
    .B(_3940__bF$buf3),
    .C(_3939__bF$buf4),
    .D(_3937_),
    .Y(_3941_)
);

NOR2X1 _13372_ (
    .A(_3941_),
    .B(_3936_),
    .Y(_3942_)
);

NAND2X1 _13373_ (
    .A(_3931_),
    .B(_3942_),
    .Y(_3943_)
);

NAND3X1 _13374_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3901_),
    .C(_3862_),
    .Y(_3944_)
);

INVX8 _13375_ (
    .A(_3944__bF$buf3),
    .Y(_3945_)
);

NAND3X1 _13376_ (
    .A(_3887_),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .C(_3901_),
    .Y(_3946_)
);

INVX8 _13377_ (
    .A(_3946_),
    .Y(_3947_)
);

AOI22X1 _13378_ (
    .A(_3947__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [0]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_3948_)
);

NAND3X1 _13379_ (
    .A(_3883_),
    .B(_3901_),
    .C(_3862_),
    .Y(_3949_)
);

INVX8 _13380_ (
    .A(_3949_),
    .Y(_3950_)
);

NAND3X1 _13381_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3888_),
    .C(_3868_),
    .Y(_3951_)
);

INVX8 _13382_ (
    .A(_3951_),
    .Y(_3952_)
);

AOI22X1 _13383_ (
    .A(_3952__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [0]),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_3953_)
);

INVX1 _13384_ (
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_3954_)
);

INVX1 _13385_ (
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_3955_)
);

NAND3X1 _13386_ (
    .A(_3883_),
    .B(_3873_),
    .C(_3862_),
    .Y(_3956_)
);

NAND3X1 _13387_ (
    .A(_3883_),
    .B(_3864_),
    .C(_3862_),
    .Y(_3957_)
);

OAI22X1 _13388_ (
    .A(_3957__bF$buf4),
    .B(_3954_),
    .C(_3955_),
    .D(_3956__bF$buf4),
    .Y(_3958_)
);

INVX1 _13389_ (
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_3959_)
);

INVX1 _13390_ (
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_3960_)
);

NAND3X1 _13391_ (
    .A(_3883_),
    .B(_3864_),
    .C(_3868_),
    .Y(_3961_)
);

NAND3X1 _13392_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3888_),
    .C(_3862_),
    .Y(_3962_)
);

OAI22X1 _13393_ (
    .A(_3960_),
    .B(_3961__bF$buf4),
    .C(_3962__bF$buf3),
    .D(_3959_),
    .Y(_3963_)
);

NOR2X1 _13394_ (
    .A(_3963_),
    .B(_3958_),
    .Y(_3964_)
);

NAND3X1 _13395_ (
    .A(_3953_),
    .B(_3948_),
    .C(_3964_),
    .Y(_3965_)
);

NOR2X1 _13396_ (
    .A(_3943_),
    .B(_3965_),
    .Y(_3966_)
);

AOI21X1 _13397_ (
    .A(_3920_),
    .B(_3966_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [0])
);

INVX1 _13398_ (
    .A(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_3967_)
);

INVX1 _13399_ (
    .A(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_3968_)
);

OAI22X1 _13400_ (
    .A(_3968_),
    .B(_3929__bF$buf3),
    .C(_3962__bF$buf2),
    .D(_3967_),
    .Y(_3969_)
);

INVX1 _13401_ (
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_3970_)
);

INVX1 _13402_ (
    .A(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_3971_)
);

OAI22X1 _13403_ (
    .A(_3916__bF$buf3),
    .B(_3970_),
    .C(_3971_),
    .D(_3915__bF$buf2),
    .Y(_3972_)
);

NOR2X1 _13404_ (
    .A(_3969_),
    .B(_3972_),
    .Y(_3973_)
);

AOI22X1 _13405_ (
    .A(_3866__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [1]),
    .C(\datapath_1.regfile_1.regOut[31] [1]),
    .D(_3906__bF$buf2),
    .Y(_3974_)
);

INVX4 _13406_ (
    .A(_3940__bF$buf2),
    .Y(_3975_)
);

INVX1 _13407_ (
    .A(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_3976_)
);

NOR2X1 _13408_ (
    .A(_3976_),
    .B(_3939__bF$buf3),
    .Y(_3977_)
);

AOI21X1 _13409_ (
    .A(_3975_),
    .B(\datapath_1.regfile_1.regOut[2] [1]),
    .C(_3977_),
    .Y(_3978_)
);

NAND3X1 _13410_ (
    .A(_3974_),
    .B(_3978_),
    .C(_3973_),
    .Y(_3979_)
);

INVX1 _13411_ (
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_3980_)
);

INVX1 _13412_ (
    .A(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_3981_)
);

OAI22X1 _13413_ (
    .A(_3981_),
    .B(_3956__bF$buf3),
    .C(_3893_),
    .D(_3980_),
    .Y(_3982_)
);

INVX1 _13414_ (
    .A(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_3983_)
);

INVX1 _13415_ (
    .A(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_3984_)
);

OAI22X1 _13416_ (
    .A(_3984_),
    .B(_3923__bF$buf3),
    .C(_3983_),
    .D(_3894__bF$buf3),
    .Y(_3985_)
);

NOR2X1 _13417_ (
    .A(_3985_),
    .B(_3982_),
    .Y(_3986_)
);

INVX8 _13418_ (
    .A(_3910__bF$buf2),
    .Y(_3987_)
);

AOI22X1 _13419_ (
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[27] [1]),
    .D(_3947__bF$buf2),
    .Y(_3988_)
);

AND2X2 _13420_ (
    .A(_3885_),
    .B(_3883_),
    .Y(_3989_)
);

INVX4 _13421_ (
    .A(_3934__bF$buf2),
    .Y(_3990_)
);

AOI22X1 _13422_ (
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[21] [1]),
    .D(_3990_),
    .Y(_3991_)
);

NAND3X1 _13423_ (
    .A(_3988_),
    .B(_3991_),
    .C(_3986_),
    .Y(_3992_)
);

NOR2X1 _13424_ (
    .A(_3992_),
    .B(_3979_),
    .Y(_3993_)
);

AOI22X1 _13425_ (
    .A(_3904__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [1]),
    .C(\datapath_1.regfile_1.regOut[9] [1]),
    .D(_3950__bF$buf2),
    .Y(_3994_)
);

AOI22X1 _13426_ (
    .A(_3952__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [1]),
    .C(\datapath_1.regfile_1.regOut[24] [1]),
    .D(_3902__bF$buf3),
    .Y(_3995_)
);

INVX1 _13427_ (
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_3996_)
);

INVX1 _13428_ (
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_3997_)
);

OAI22X1 _13429_ (
    .A(_3997_),
    .B(_3875__bF$buf2),
    .C(_3911_),
    .D(_3996_),
    .Y(_3998_)
);

INVX1 _13430_ (
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_3999_)
);

INVX1 _13431_ (
    .A(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_4000_)
);

OAI22X1 _13432_ (
    .A(_3889__bF$buf3),
    .B(_4000_),
    .C(_3999_),
    .D(_3935__bF$buf2),
    .Y(_4001_)
);

NOR2X1 _13433_ (
    .A(_3998_),
    .B(_4001_),
    .Y(_4002_)
);

NAND3X1 _13434_ (
    .A(_3995_),
    .B(_3994_),
    .C(_4002_),
    .Y(_4003_)
);

INVX1 _13435_ (
    .A(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_4004_)
);

INVX1 _13436_ (
    .A(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_4005_)
);

OAI22X1 _13437_ (
    .A(_4005_),
    .B(_3957__bF$buf3),
    .C(_3961__bF$buf3),
    .D(_4004_),
    .Y(_4006_)
);

INVX1 _13438_ (
    .A(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_4007_)
);

INVX1 _13439_ (
    .A(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_4008_)
);

OAI22X1 _13440_ (
    .A(_4008_),
    .B(_3928_),
    .C(_4007_),
    .D(_3924__bF$buf2),
    .Y(_4009_)
);

NOR2X1 _13441_ (
    .A(_4006_),
    .B(_4009_),
    .Y(_4010_)
);

AOI22X1 _13442_ (
    .A(_3899__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [1]),
    .C(\datapath_1.regfile_1.regOut[28] [1]),
    .D(_3879__bF$buf2),
    .Y(_4011_)
);

AOI22X1 _13443_ (
    .A(_3870__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [1]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_4012_)
);

NAND3X1 _13444_ (
    .A(_4011_),
    .B(_4012_),
    .C(_4010_),
    .Y(_4013_)
);

NOR2X1 _13445_ (
    .A(_4003_),
    .B(_4013_),
    .Y(_4014_)
);

AOI21X1 _13446_ (
    .A(_3993_),
    .B(_4014_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [1])
);

INVX1 _13447_ (
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_4015_)
);

INVX1 _13448_ (
    .A(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_4016_)
);

OAI22X1 _13449_ (
    .A(_3894__bF$buf2),
    .B(_4015_),
    .C(_4016_),
    .D(_3915__bF$buf1),
    .Y(_4017_)
);

INVX1 _13450_ (
    .A(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_4018_)
);

INVX1 _13451_ (
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_4019_)
);

OAI22X1 _13452_ (
    .A(_3946_),
    .B(_4018_),
    .C(_4019_),
    .D(_3886__bF$buf2),
    .Y(_4020_)
);

NOR2X1 _13453_ (
    .A(_4017_),
    .B(_4020_),
    .Y(_4021_)
);

INVX1 _13454_ (
    .A(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_4022_)
);

INVX1 _13455_ (
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_4023_)
);

OAI22X1 _13456_ (
    .A(_3875__bF$buf1),
    .B(_4023_),
    .C(_4022_),
    .D(_3957__bF$buf2),
    .Y(_4024_)
);

INVX1 _13457_ (
    .A(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_4025_)
);

INVX1 _13458_ (
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_4026_)
);

OAI22X1 _13459_ (
    .A(_3923__bF$buf2),
    .B(_4026_),
    .C(_4025_),
    .D(_3929__bF$buf2),
    .Y(_4027_)
);

NOR2X1 _13460_ (
    .A(_4027_),
    .B(_4024_),
    .Y(_4028_)
);

NAND2X1 _13461_ (
    .A(_4028_),
    .B(_4021_),
    .Y(_4029_)
);

INVX1 _13462_ (
    .A(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_4030_)
);

INVX1 _13463_ (
    .A(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_4031_)
);

OAI22X1 _13464_ (
    .A(_3961__bF$buf2),
    .B(_4030_),
    .C(_4031_),
    .D(_3949_),
    .Y(_4032_)
);

INVX1 _13465_ (
    .A(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_4033_)
);

INVX1 _13466_ (
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_4034_)
);

OAI22X1 _13467_ (
    .A(_3910__bF$buf1),
    .B(_4033_),
    .C(_4034_),
    .D(_3934__bF$buf1),
    .Y(_4035_)
);

NOR2X1 _13468_ (
    .A(_4035_),
    .B(_4032_),
    .Y(_4036_)
);

AOI22X1 _13469_ (
    .A(_3866__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [2]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_4037_)
);

INVX8 _13470_ (
    .A(_3935__bF$buf1),
    .Y(_4038_)
);

AOI22X1 _13471_ (
    .A(_3904__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [2]),
    .C(\datapath_1.regfile_1.regOut[22] [2]),
    .D(_4038_),
    .Y(_4039_)
);

NAND3X1 _13472_ (
    .A(_4037_),
    .B(_4039_),
    .C(_4036_),
    .Y(_4040_)
);

NOR2X1 _13473_ (
    .A(_4029_),
    .B(_4040_),
    .Y(_4041_)
);

INVX1 _13474_ (
    .A(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_4042_)
);

INVX1 _13475_ (
    .A(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_4043_)
);

NAND3X1 _13476_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3877_),
    .C(_3864_),
    .Y(_4044_)
);

OAI22X1 _13477_ (
    .A(_4044_),
    .B(_4042_),
    .C(_4043_),
    .D(_3951_),
    .Y(_4045_)
);

INVX1 _13478_ (
    .A(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_4046_)
);

INVX1 _13479_ (
    .A(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_4047_)
);

OAI22X1 _13480_ (
    .A(_3889__bF$buf2),
    .B(_4046_),
    .C(_4047_),
    .D(_3893_),
    .Y(_4048_)
);

NOR2X1 _13481_ (
    .A(_4045_),
    .B(_4048_),
    .Y(_4049_)
);

AOI22X1 _13482_ (
    .A(_3870__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .C(_3906__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_4050_)
);

AOI22X1 _13483_ (
    .A(_3899__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [2]),
    .C(\datapath_1.regfile_1.regOut[24] [2]),
    .D(_3902__bF$buf2),
    .Y(_4051_)
);

NAND3X1 _13484_ (
    .A(_4050_),
    .B(_4051_),
    .C(_4049_),
    .Y(_4052_)
);

INVX1 _13485_ (
    .A(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_4053_)
);

INVX1 _13486_ (
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_4054_)
);

OAI22X1 _13487_ (
    .A(_3916__bF$buf2),
    .B(_4054_),
    .C(_4053_),
    .D(_3924__bF$buf1),
    .Y(_4055_)
);

INVX1 _13488_ (
    .A(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_4056_)
);

INVX1 _13489_ (
    .A(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_4057_)
);

OAI22X1 _13490_ (
    .A(_3962__bF$buf1),
    .B(_4056_),
    .C(_4057_),
    .D(_3956__bF$buf2),
    .Y(_4058_)
);

NOR2X1 _13491_ (
    .A(_4058_),
    .B(_4055_),
    .Y(_4059_)
);

INVX8 _13492_ (
    .A(_3928_),
    .Y(_4060_)
);

AOI22X1 _13493_ (
    .A(_4060__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [2]),
    .C(_3975_),
    .D(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_4061_)
);

INVX8 _13494_ (
    .A(_3911_),
    .Y(_4062_)
);

INVX1 _13495_ (
    .A(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_4063_)
);

NOR2X1 _13496_ (
    .A(_4063_),
    .B(_3939__bF$buf2),
    .Y(_4064_)
);

AOI21X1 _13497_ (
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .B(_4062__bF$buf3),
    .C(_4064_),
    .Y(_4065_)
);

NAND3X1 _13498_ (
    .A(_4061_),
    .B(_4065_),
    .C(_4059_),
    .Y(_4066_)
);

NOR2X1 _13499_ (
    .A(_4052_),
    .B(_4066_),
    .Y(_4067_)
);

AOI21X1 _13500_ (
    .A(_4067_),
    .B(_4041_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [2])
);

INVX8 _13501_ (
    .A(_3893_),
    .Y(_4068_)
);

AOI22X1 _13502_ (
    .A(_4060__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [3]),
    .C(\datapath_1.regfile_1.regOut[6] [3]),
    .D(_4068__bF$buf3),
    .Y(_4069_)
);

INVX8 _13503_ (
    .A(_3924__bF$buf0),
    .Y(_4070_)
);

AOI22X1 _13504_ (
    .A(_4070_),
    .B(\datapath_1.regfile_1.regOut[26] [3]),
    .C(_4038_),
    .D(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_4071_)
);

INVX1 _13505_ (
    .A(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_4072_)
);

INVX1 _13506_ (
    .A(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_4073_)
);

OAI22X1 _13507_ (
    .A(_4073_),
    .B(_3940__bF$buf1),
    .C(_3929__bF$buf1),
    .D(_4072_),
    .Y(_4074_)
);

INVX1 _13508_ (
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_4075_)
);

INVX1 _13509_ (
    .A(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_4076_)
);

OAI22X1 _13510_ (
    .A(_3910__bF$buf0),
    .B(_4075_),
    .C(_4076_),
    .D(_3939__bF$buf1),
    .Y(_4077_)
);

NOR2X1 _13511_ (
    .A(_4077_),
    .B(_4074_),
    .Y(_4078_)
);

NAND3X1 _13512_ (
    .A(_4069_),
    .B(_4071_),
    .C(_4078_),
    .Y(_4079_)
);

INVX1 _13513_ (
    .A(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_4080_)
);

INVX1 _13514_ (
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_4081_)
);

OAI22X1 _13515_ (
    .A(_3916__bF$buf1),
    .B(_4081_),
    .C(_4080_),
    .D(_3944__bF$buf2),
    .Y(_4082_)
);

INVX1 _13516_ (
    .A(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_4083_)
);

INVX1 _13517_ (
    .A(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_4084_)
);

OAI22X1 _13518_ (
    .A(_3889__bF$buf1),
    .B(_4083_),
    .C(_4084_),
    .D(_3956__bF$buf1),
    .Y(_4085_)
);

NOR2X1 _13519_ (
    .A(_4085_),
    .B(_4082_),
    .Y(_4086_)
);

INVX4 _13520_ (
    .A(_3915__bF$buf0),
    .Y(_4087_)
);

AOI22X1 _13521_ (
    .A(_3879__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [3]),
    .C(_4087_),
    .D(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_4088_)
);

AOI22X1 _13522_ (
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[21] [3]),
    .D(_3990_),
    .Y(_4089_)
);

NAND3X1 _13523_ (
    .A(_4088_),
    .B(_4089_),
    .C(_4086_),
    .Y(_4090_)
);

NOR2X1 _13524_ (
    .A(_4079_),
    .B(_4090_),
    .Y(_4091_)
);

INVX1 _13525_ (
    .A(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_4092_)
);

INVX1 _13526_ (
    .A(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_4093_)
);

OAI22X1 _13527_ (
    .A(_3894__bF$buf1),
    .B(_4093_),
    .C(_4092_),
    .D(_3961__bF$buf1),
    .Y(_4094_)
);

INVX1 _13528_ (
    .A(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_4095_)
);

INVX1 _13529_ (
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_4096_)
);

OAI22X1 _13530_ (
    .A(_4096_),
    .B(_3875__bF$buf0),
    .C(_3911_),
    .D(_4095_),
    .Y(_4097_)
);

NOR2X1 _13531_ (
    .A(_4097_),
    .B(_4094_),
    .Y(_4098_)
);

INVX4 _13532_ (
    .A(_3957__bF$buf1),
    .Y(_4099_)
);

INVX1 _13533_ (
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_4100_)
);

NOR2X1 _13534_ (
    .A(_4100_),
    .B(_3923__bF$buf1),
    .Y(_4101_)
);

AOI21X1 _13535_ (
    .A(_4099_),
    .B(\datapath_1.regfile_1.regOut[13] [3]),
    .C(_4101_),
    .Y(_4102_)
);

AOI22X1 _13536_ (
    .A(_3947__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [3]),
    .C(_3902__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_4103_)
);

NAND3X1 _13537_ (
    .A(_4102_),
    .B(_4103_),
    .C(_4098_),
    .Y(_4104_)
);

INVX1 _13538_ (
    .A(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_4105_)
);

INVX1 _13539_ (
    .A(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_4106_)
);

OAI22X1 _13540_ (
    .A(_4106_),
    .B(_3962__bF$buf0),
    .C(_3898_),
    .D(_4105_),
    .Y(_4107_)
);

INVX1 _13541_ (
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_4108_)
);

INVX1 _13542_ (
    .A(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_4109_)
);

OAI22X1 _13543_ (
    .A(_4109_),
    .B(_3951_),
    .C(_4108_),
    .D(_3869_),
    .Y(_4110_)
);

NOR2X1 _13544_ (
    .A(_4107_),
    .B(_4110_),
    .Y(_4111_)
);

AOI22X1 _13545_ (
    .A(_3866__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [3]),
    .C(\datapath_1.regfile_1.regOut[31] [3]),
    .D(_3906__bF$buf0),
    .Y(_4112_)
);

AOI22X1 _13546_ (
    .A(_3904__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [3]),
    .C(\datapath_1.regfile_1.regOut[9] [3]),
    .D(_3950__bF$buf1),
    .Y(_4113_)
);

NAND3X1 _13547_ (
    .A(_4112_),
    .B(_4113_),
    .C(_4111_),
    .Y(_4114_)
);

NOR2X1 _13548_ (
    .A(_4104_),
    .B(_4114_),
    .Y(_4115_)
);

AOI21X1 _13549_ (
    .A(_4091_),
    .B(_4115_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [3])
);

AOI22X1 _13550_ (
    .A(_4038_),
    .B(\datapath_1.regfile_1.regOut[22] [4]),
    .C(_3990_),
    .D(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_4116_)
);

INVX1 _13551_ (
    .A(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_4117_)
);

INVX1 _13552_ (
    .A(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_4118_)
);

OAI22X1 _13553_ (
    .A(_4118_),
    .B(_3949_),
    .C(_3915__bF$buf3),
    .D(_4117_),
    .Y(_4119_)
);

INVX1 _13554_ (
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_4120_)
);

INVX1 _13555_ (
    .A(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_4121_)
);

OAI22X1 _13556_ (
    .A(_3916__bF$buf0),
    .B(_4120_),
    .C(_4121_),
    .D(_3886__bF$buf1),
    .Y(_4122_)
);

NOR2X1 _13557_ (
    .A(_4122_),
    .B(_4119_),
    .Y(_4123_)
);

INVX1 _13558_ (
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_4124_)
);

NOR2X1 _13559_ (
    .A(_4124_),
    .B(_3889__bF$buf0),
    .Y(_4125_)
);

AOI21X1 _13560_ (
    .A(_3904__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [4]),
    .C(_4125_),
    .Y(_4126_)
);

NAND3X1 _13561_ (
    .A(_4116_),
    .B(_4126_),
    .C(_4123_),
    .Y(_4127_)
);

INVX1 _13562_ (
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_4128_)
);

INVX1 _13563_ (
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_4129_)
);

OAI22X1 _13564_ (
    .A(_4128_),
    .B(_3894__bF$buf0),
    .C(_4129_),
    .D(_3929__bF$buf0),
    .Y(_4130_)
);

INVX1 _13565_ (
    .A(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_4131_)
);

INVX1 _13566_ (
    .A(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_4132_)
);

OAI22X1 _13567_ (
    .A(_4132_),
    .B(_3957__bF$buf0),
    .C(_3961__bF$buf0),
    .D(_4131_),
    .Y(_4133_)
);

NOR2X1 _13568_ (
    .A(_4130_),
    .B(_4133_),
    .Y(_4134_)
);

INVX4 _13569_ (
    .A(_3962__bF$buf3),
    .Y(_4135_)
);

AOI22X1 _13570_ (
    .A(_3952__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [4]),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_4136_)
);

AOI22X1 _13571_ (
    .A(_3899__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [4]),
    .C(\datapath_1.regfile_1.regOut[24] [4]),
    .D(_3902__bF$buf0),
    .Y(_4137_)
);

NAND3X1 _13572_ (
    .A(_4136_),
    .B(_4137_),
    .C(_4134_),
    .Y(_4138_)
);

NOR2X1 _13573_ (
    .A(_4138_),
    .B(_4127_),
    .Y(_4139_)
);

AOI22X1 _13574_ (
    .A(_4060__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [4]),
    .C(\datapath_1.regfile_1.regOut[6] [4]),
    .D(_4068__bF$buf2),
    .Y(_4140_)
);

AOI22X1 _13575_ (
    .A(_3870__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [4]),
    .C(_3906__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_4141_)
);

INVX1 _13576_ (
    .A(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_4142_)
);

INVX1 _13577_ (
    .A(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_4143_)
);

OAI22X1 _13578_ (
    .A(_3923__bF$buf0),
    .B(_4143_),
    .C(_4142_),
    .D(_3940__bF$buf0),
    .Y(_4144_)
);

INVX1 _13579_ (
    .A(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_4145_)
);

INVX1 _13580_ (
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_4146_)
);

OAI22X1 _13581_ (
    .A(_3939__bF$buf0),
    .B(_4146_),
    .C(_4145_),
    .D(_3924__bF$buf3),
    .Y(_4147_)
);

NOR2X1 _13582_ (
    .A(_4144_),
    .B(_4147_),
    .Y(_4148_)
);

NAND3X1 _13583_ (
    .A(_4141_),
    .B(_4140_),
    .C(_4148_),
    .Y(_4149_)
);

INVX1 _13584_ (
    .A(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_4150_)
);

INVX1 _13585_ (
    .A(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_4151_)
);

OAI22X1 _13586_ (
    .A(_3911_),
    .B(_4150_),
    .C(_4151_),
    .D(_3956__bF$buf0),
    .Y(_4152_)
);

INVX1 _13587_ (
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_4153_)
);

INVX1 _13588_ (
    .A(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_4154_)
);

OAI22X1 _13589_ (
    .A(_4044_),
    .B(_4153_),
    .C(_4154_),
    .D(_3946_),
    .Y(_4155_)
);

NOR2X1 _13590_ (
    .A(_4155_),
    .B(_4152_),
    .Y(_4156_)
);

AOI22X1 _13591_ (
    .A(_3866__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [4]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_4157_)
);

AOI22X1 _13592_ (
    .A(_3987_),
    .B(\datapath_1.regfile_1.regOut[0] [4]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_4158_)
);

NAND3X1 _13593_ (
    .A(_4157_),
    .B(_4158_),
    .C(_4156_),
    .Y(_4159_)
);

NOR2X1 _13594_ (
    .A(_4149_),
    .B(_4159_),
    .Y(_4160_)
);

AOI21X1 _13595_ (
    .A(_4139_),
    .B(_4160_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [4])
);

AOI22X1 _13596_ (
    .A(_4060__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [5]),
    .C(\datapath_1.regfile_1.regOut[31] [5]),
    .D(_3906__bF$buf2),
    .Y(_4161_)
);

AOI22X1 _13597_ (
    .A(_4087_),
    .B(\datapath_1.regfile_1.regOut[10] [5]),
    .C(_4068__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_4162_)
);

INVX1 _13598_ (
    .A(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_4163_)
);

INVX1 _13599_ (
    .A(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_4164_)
);

OAI22X1 _13600_ (
    .A(_4164_),
    .B(_3939__bF$buf4),
    .C(_3898_),
    .D(_4163_),
    .Y(_4165_)
);

INVX1 _13601_ (
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_4166_)
);

INVX1 _13602_ (
    .A(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_4167_)
);

OAI22X1 _13603_ (
    .A(_4044_),
    .B(_4166_),
    .C(_4167_),
    .D(_3944__bF$buf1),
    .Y(_4168_)
);

NOR2X1 _13604_ (
    .A(_4165_),
    .B(_4168_),
    .Y(_4169_)
);

NAND3X1 _13605_ (
    .A(_4161_),
    .B(_4162_),
    .C(_4169_),
    .Y(_4170_)
);

AOI22X1 _13606_ (
    .A(_3947__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [5]),
    .C(\datapath_1.regfile_1.regOut[26] [5]),
    .D(_4070_),
    .Y(_4171_)
);

AOI22X1 _13607_ (
    .A(_3870__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [5]),
    .C(_4038_),
    .D(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_4172_)
);

INVX1 _13608_ (
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_4173_)
);

INVX1 _13609_ (
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_4174_)
);

OAI22X1 _13610_ (
    .A(_4173_),
    .B(_3934__bF$buf0),
    .C(_3886__bF$buf0),
    .D(_4174_),
    .Y(_4175_)
);

INVX1 _13611_ (
    .A(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_4176_)
);

INVX1 _13612_ (
    .A(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_4177_)
);

OAI22X1 _13613_ (
    .A(_4177_),
    .B(_3940__bF$buf3),
    .C(_3962__bF$buf2),
    .D(_4176_),
    .Y(_4178_)
);

NOR2X1 _13614_ (
    .A(_4178_),
    .B(_4175_),
    .Y(_4179_)
);

NAND3X1 _13615_ (
    .A(_4171_),
    .B(_4172_),
    .C(_4179_),
    .Y(_4180_)
);

NOR2X1 _13616_ (
    .A(_4180_),
    .B(_4170_),
    .Y(_4181_)
);

AOI22X1 _13617_ (
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .B(_4062__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[9] [5]),
    .D(_3950__bF$buf0),
    .Y(_4182_)
);

INVX1 _13618_ (
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_4183_)
);

NOR2X1 _13619_ (
    .A(_4183_),
    .B(_3923__bF$buf4),
    .Y(_4184_)
);

AOI21X1 _13620_ (
    .A(_3904__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [5]),
    .C(_4184_),
    .Y(_4185_)
);

INVX1 _13621_ (
    .A(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_4186_)
);

INVX1 _13622_ (
    .A(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_4187_)
);

OAI22X1 _13623_ (
    .A(_3894__bF$buf4),
    .B(_4186_),
    .C(_4187_),
    .D(_3957__bF$buf4),
    .Y(_4188_)
);

INVX1 _13624_ (
    .A(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_4189_)
);

INVX1 _13625_ (
    .A(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_4190_)
);

OAI22X1 _13626_ (
    .A(_4190_),
    .B(_3929__bF$buf4),
    .C(_4189_),
    .D(_3865_),
    .Y(_4191_)
);

NOR2X1 _13627_ (
    .A(_4188_),
    .B(_4191_),
    .Y(_4192_)
);

NAND3X1 _13628_ (
    .A(_4185_),
    .B(_4182_),
    .C(_4192_),
    .Y(_4193_)
);

INVX1 _13629_ (
    .A(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_4194_)
);

INVX1 _13630_ (
    .A(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_4195_)
);

OAI22X1 _13631_ (
    .A(_3889__bF$buf4),
    .B(_4194_),
    .C(_4195_),
    .D(_3956__bF$buf4),
    .Y(_4196_)
);

INVX1 _13632_ (
    .A(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_4197_)
);

INVX1 _13633_ (
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_4198_)
);

OAI22X1 _13634_ (
    .A(_3916__bF$buf4),
    .B(_4198_),
    .C(_4197_),
    .D(_3951_),
    .Y(_4199_)
);

NOR2X1 _13635_ (
    .A(_4199_),
    .B(_4196_),
    .Y(_4200_)
);

INVX1 _13636_ (
    .A(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_4201_)
);

NOR2X1 _13637_ (
    .A(_4201_),
    .B(_3961__bF$buf4),
    .Y(_4202_)
);

AOI21X1 _13638_ (
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .B(_3876_),
    .C(_4202_),
    .Y(_4203_)
);

AOI22X1 _13639_ (
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[24] [5]),
    .D(_3902__bF$buf4),
    .Y(_4204_)
);

NAND3X1 _13640_ (
    .A(_4203_),
    .B(_4204_),
    .C(_4200_),
    .Y(_4205_)
);

NOR2X1 _13641_ (
    .A(_4205_),
    .B(_4193_),
    .Y(_4206_)
);

AOI21X1 _13642_ (
    .A(_4181_),
    .B(_4206_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [5])
);

INVX1 _13643_ (
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_4207_)
);

INVX1 _13644_ (
    .A(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_4208_)
);

OAI22X1 _13645_ (
    .A(_3889__bF$buf3),
    .B(_4207_),
    .C(_4208_),
    .D(_3894__bF$buf3),
    .Y(_4209_)
);

INVX1 _13646_ (
    .A(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_4210_)
);

INVX1 _13647_ (
    .A(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_4211_)
);

OAI22X1 _13648_ (
    .A(_4211_),
    .B(_3961__bF$buf3),
    .C(_4210_),
    .D(_3905_),
    .Y(_4212_)
);

NOR2X1 _13649_ (
    .A(_4209_),
    .B(_4212_),
    .Y(_4213_)
);

AOI22X1 _13650_ (
    .A(_3975_),
    .B(\datapath_1.regfile_1.regOut[2] [6]),
    .C(\datapath_1.regfile_1.regOut[26] [6]),
    .D(_4070_),
    .Y(_4214_)
);

AOI22X1 _13651_ (
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[25] [6]),
    .D(_3945_),
    .Y(_4215_)
);

NAND3X1 _13652_ (
    .A(_4215_),
    .B(_4214_),
    .C(_4213_),
    .Y(_4216_)
);

AOI22X1 _13653_ (
    .A(_3899__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [6]),
    .C(\datapath_1.regfile_1.regOut[24] [6]),
    .D(_3902__bF$buf3),
    .Y(_4217_)
);

AOI22X1 _13654_ (
    .A(_3952__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [6]),
    .C(\datapath_1.regfile_1.regOut[28] [6]),
    .D(_3879__bF$buf0),
    .Y(_4218_)
);

INVX1 _13655_ (
    .A(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_4219_)
);

INVX1 _13656_ (
    .A(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_4220_)
);

OAI22X1 _13657_ (
    .A(_4220_),
    .B(_3929__bF$buf3),
    .C(_3962__bF$buf1),
    .D(_4219_),
    .Y(_4221_)
);

INVX1 _13658_ (
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_4222_)
);

INVX1 _13659_ (
    .A(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_4223_)
);

OAI22X1 _13660_ (
    .A(_3869_),
    .B(_4222_),
    .C(_4223_),
    .D(_3956__bF$buf3),
    .Y(_4224_)
);

NOR2X1 _13661_ (
    .A(_4221_),
    .B(_4224_),
    .Y(_4225_)
);

NAND3X1 _13662_ (
    .A(_4218_),
    .B(_4217_),
    .C(_4225_),
    .Y(_4226_)
);

NOR2X1 _13663_ (
    .A(_4216_),
    .B(_4226_),
    .Y(_4227_)
);

INVX1 _13664_ (
    .A(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_4228_)
);

INVX1 _13665_ (
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_4229_)
);

OAI22X1 _13666_ (
    .A(_3911_),
    .B(_4228_),
    .C(_4229_),
    .D(_3939__bF$buf3),
    .Y(_4230_)
);

INVX1 _13667_ (
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_4231_)
);

INVX1 _13668_ (
    .A(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_4232_)
);

OAI22X1 _13669_ (
    .A(_4232_),
    .B(_3923__bF$buf3),
    .C(_4231_),
    .D(_3910__bF$buf3),
    .Y(_4233_)
);

NOR2X1 _13670_ (
    .A(_4233_),
    .B(_4230_),
    .Y(_4234_)
);

AOI22X1 _13671_ (
    .A(_4060__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [6]),
    .C(\datapath_1.regfile_1.regOut[6] [6]),
    .D(_4068__bF$buf0),
    .Y(_4235_)
);

AOI22X1 _13672_ (
    .A(_4099_),
    .B(\datapath_1.regfile_1.regOut[13] [6]),
    .C(\datapath_1.regfile_1.regOut[29] [6]),
    .D(_3866__bF$buf2),
    .Y(_4236_)
);

NAND3X1 _13673_ (
    .A(_4236_),
    .B(_4235_),
    .C(_4234_),
    .Y(_4237_)
);

INVX1 _13674_ (
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_4238_)
);

NOR2X1 _13675_ (
    .A(_4238_),
    .B(_3916__bF$buf3),
    .Y(_4239_)
);

AOI21X1 _13676_ (
    .A(_3950__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[9] [6]),
    .C(_4239_),
    .Y(_4240_)
);

AOI22X1 _13677_ (
    .A(_3904__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [6]),
    .C(\datapath_1.regfile_1.regOut[10] [6]),
    .D(_4087_),
    .Y(_4241_)
);

INVX1 _13678_ (
    .A(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_4242_)
);

INVX1 _13679_ (
    .A(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_4243_)
);

OAI22X1 _13680_ (
    .A(_4243_),
    .B(_3934__bF$buf3),
    .C(_3935__bF$buf0),
    .D(_4242_),
    .Y(_4244_)
);

INVX1 _13681_ (
    .A(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_4245_)
);

INVX1 _13682_ (
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_4246_)
);

OAI22X1 _13683_ (
    .A(_3875__bF$buf3),
    .B(_4246_),
    .C(_4245_),
    .D(_3946_),
    .Y(_4247_)
);

NOR2X1 _13684_ (
    .A(_4247_),
    .B(_4244_),
    .Y(_4248_)
);

NAND3X1 _13685_ (
    .A(_4241_),
    .B(_4240_),
    .C(_4248_),
    .Y(_4249_)
);

NOR2X1 _13686_ (
    .A(_4237_),
    .B(_4249_),
    .Y(_4250_)
);

AOI21X1 _13687_ (
    .A(_4227_),
    .B(_4250_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [6])
);

AOI22X1 _13688_ (
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[27] [7]),
    .D(_3947__bF$buf3),
    .Y(_4251_)
);

AOI22X1 _13689_ (
    .A(_3952__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [7]),
    .C(\datapath_1.regfile_1.regOut[24] [7]),
    .D(_3902__bF$buf2),
    .Y(_4252_)
);

INVX1 _13690_ (
    .A(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_4253_)
);

INVX1 _13691_ (
    .A(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_4254_)
);

OAI22X1 _13692_ (
    .A(_4253_),
    .B(_3894__bF$buf2),
    .C(_4254_),
    .D(_3929__bF$buf2),
    .Y(_4255_)
);

INVX1 _13693_ (
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_4256_)
);

INVX1 _13694_ (
    .A(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_4257_)
);

OAI22X1 _13695_ (
    .A(_3889__bF$buf2),
    .B(_4256_),
    .C(_4257_),
    .D(_3886__bF$buf3),
    .Y(_4258_)
);

NOR2X1 _13696_ (
    .A(_4255_),
    .B(_4258_),
    .Y(_4259_)
);

NAND3X1 _13697_ (
    .A(_4252_),
    .B(_4251_),
    .C(_4259_),
    .Y(_4260_)
);

AOI22X1 _13698_ (
    .A(_3879__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [7]),
    .C(_3904__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_4261_)
);

AOI22X1 _13699_ (
    .A(_3899__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [7]),
    .C(\datapath_1.regfile_1.regOut[29] [7]),
    .D(_3866__bF$buf1),
    .Y(_4262_)
);

INVX1 _13700_ (
    .A(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_4263_)
);

INVX1 _13701_ (
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_4264_)
);

OAI22X1 _13702_ (
    .A(_3939__bF$buf2),
    .B(_4264_),
    .C(_4263_),
    .D(_3924__bF$buf2),
    .Y(_4265_)
);

INVX1 _13703_ (
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_4266_)
);

INVX1 _13704_ (
    .A(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_4267_)
);

OAI22X1 _13705_ (
    .A(_3916__bF$buf2),
    .B(_4266_),
    .C(_4267_),
    .D(_3915__bF$buf2),
    .Y(_4268_)
);

NOR2X1 _13706_ (
    .A(_4265_),
    .B(_4268_),
    .Y(_4269_)
);

NAND3X1 _13707_ (
    .A(_4262_),
    .B(_4261_),
    .C(_4269_),
    .Y(_4270_)
);

NOR2X1 _13708_ (
    .A(_4260_),
    .B(_4270_),
    .Y(_4271_)
);

AOI22X1 _13709_ (
    .A(_4060__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [7]),
    .C(\datapath_1.regfile_1.regOut[6] [7]),
    .D(_4068__bF$buf3),
    .Y(_4272_)
);

AOI22X1 _13710_ (
    .A(_4062__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [7]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_4273_)
);

INVX1 _13711_ (
    .A(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_4274_)
);

INVX1 _13712_ (
    .A(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_4275_)
);

OAI22X1 _13713_ (
    .A(_3923__bF$buf2),
    .B(_4275_),
    .C(_4274_),
    .D(_3940__bF$buf2),
    .Y(_4276_)
);

INVX1 _13714_ (
    .A(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_4277_)
);

INVX1 _13715_ (
    .A(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_4278_)
);

OAI22X1 _13716_ (
    .A(_4278_),
    .B(_3934__bF$buf2),
    .C(_3935__bF$buf3),
    .D(_4277_),
    .Y(_4279_)
);

NOR2X1 _13717_ (
    .A(_4276_),
    .B(_4279_),
    .Y(_4280_)
);

NAND3X1 _13718_ (
    .A(_4273_),
    .B(_4272_),
    .C(_4280_),
    .Y(_4281_)
);

AOI22X1 _13719_ (
    .A(_3870__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [7]),
    .C(_3906__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_4282_)
);

AOI22X1 _13720_ (
    .A(_3945_),
    .B(\datapath_1.regfile_1.regOut[25] [7]),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_4283_)
);

INVX1 _13721_ (
    .A(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_4284_)
);

INVX1 _13722_ (
    .A(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_4285_)
);

OAI22X1 _13723_ (
    .A(_3957__bF$buf3),
    .B(_4284_),
    .C(_4285_),
    .D(_3956__bF$buf2),
    .Y(_4286_)
);

INVX1 _13724_ (
    .A(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_4287_)
);

INVX1 _13725_ (
    .A(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_4288_)
);

OAI22X1 _13726_ (
    .A(_4288_),
    .B(_3961__bF$buf2),
    .C(_3962__bF$buf0),
    .D(_4287_),
    .Y(_4289_)
);

NOR2X1 _13727_ (
    .A(_4289_),
    .B(_4286_),
    .Y(_4290_)
);

NAND3X1 _13728_ (
    .A(_4283_),
    .B(_4282_),
    .C(_4290_),
    .Y(_4291_)
);

NOR2X1 _13729_ (
    .A(_4281_),
    .B(_4291_),
    .Y(_4292_)
);

AOI21X1 _13730_ (
    .A(_4292_),
    .B(_4271_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [7])
);

INVX1 _13731_ (
    .A(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_4293_)
);

NOR2X1 _13732_ (
    .A(_4293_),
    .B(_3923__bF$buf1),
    .Y(_4294_)
);

AOI21X1 _13733_ (
    .A(_3876_),
    .B(\datapath_1.regfile_1.regOut[4] [8]),
    .C(_4294_),
    .Y(_4295_)
);

AOI22X1 _13734_ (
    .A(_4070_),
    .B(\datapath_1.regfile_1.regOut[26] [8]),
    .C(_4038_),
    .D(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_4296_)
);

INVX1 _13735_ (
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_4297_)
);

INVX1 _13736_ (
    .A(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_4298_)
);

OAI22X1 _13737_ (
    .A(_3894__bF$buf1),
    .B(_4297_),
    .C(_4298_),
    .D(_3893_),
    .Y(_4299_)
);

INVX1 _13738_ (
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_4300_)
);

INVX1 _13739_ (
    .A(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_4301_)
);

OAI22X1 _13740_ (
    .A(_4044_),
    .B(_4300_),
    .C(_4301_),
    .D(_3956__bF$buf1),
    .Y(_4302_)
);

NOR2X1 _13741_ (
    .A(_4299_),
    .B(_4302_),
    .Y(_4303_)
);

NAND3X1 _13742_ (
    .A(_4296_),
    .B(_4295_),
    .C(_4303_),
    .Y(_4304_)
);

INVX1 _13743_ (
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_4305_)
);

INVX1 _13744_ (
    .A(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_4306_)
);

OAI22X1 _13745_ (
    .A(_4306_),
    .B(_3939__bF$buf1),
    .C(_4305_),
    .D(_3886__bF$buf2),
    .Y(_4307_)
);

INVX1 _13746_ (
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_4308_)
);

INVX1 _13747_ (
    .A(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_4309_)
);

OAI22X1 _13748_ (
    .A(_3889__bF$buf1),
    .B(_4308_),
    .C(_4309_),
    .D(_3940__bF$buf1),
    .Y(_4310_)
);

NOR2X1 _13749_ (
    .A(_4310_),
    .B(_4307_),
    .Y(_4311_)
);

AOI22X1 _13750_ (
    .A(_3945_),
    .B(\datapath_1.regfile_1.regOut[25] [8]),
    .C(_4087_),
    .D(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_4312_)
);

INVX1 _13751_ (
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_4313_)
);

NOR2X1 _13752_ (
    .A(_4313_),
    .B(_3916__bF$buf1),
    .Y(_4314_)
);

AOI21X1 _13753_ (
    .A(_3990_),
    .B(\datapath_1.regfile_1.regOut[21] [8]),
    .C(_4314_),
    .Y(_4315_)
);

NAND3X1 _13754_ (
    .A(_4315_),
    .B(_4312_),
    .C(_4311_),
    .Y(_4316_)
);

NOR2X1 _13755_ (
    .A(_4316_),
    .B(_4304_),
    .Y(_4317_)
);

INVX1 _13756_ (
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_4318_)
);

NOR2X1 _13757_ (
    .A(_4318_),
    .B(_3961__bF$buf1),
    .Y(_4319_)
);

AOI21X1 _13758_ (
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .B(_4099_),
    .C(_4319_),
    .Y(_4320_)
);

AOI22X1 _13759_ (
    .A(_4062__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [8]),
    .C(\datapath_1.regfile_1.regOut[7] [8]),
    .D(_4060__bF$buf1),
    .Y(_4321_)
);

INVX1 _13760_ (
    .A(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_4322_)
);

INVX1 _13761_ (
    .A(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_4323_)
);

OAI22X1 _13762_ (
    .A(_4323_),
    .B(_3929__bF$buf1),
    .C(_3962__bF$buf3),
    .D(_4322_),
    .Y(_4324_)
);

INVX1 _13763_ (
    .A(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_4325_)
);

INVX1 _13764_ (
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_4326_)
);

OAI22X1 _13765_ (
    .A(_4326_),
    .B(_3946_),
    .C(_4325_),
    .D(_3869_),
    .Y(_4327_)
);

NOR2X1 _13766_ (
    .A(_4324_),
    .B(_4327_),
    .Y(_4328_)
);

NAND3X1 _13767_ (
    .A(_4321_),
    .B(_4320_),
    .C(_4328_),
    .Y(_4329_)
);

INVX1 _13768_ (
    .A(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_4330_)
);

INVX1 _13769_ (
    .A(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_4331_)
);

NAND2X1 _13770_ (
    .A(_3901_),
    .B(_3878_),
    .Y(_4332_)
);

OAI22X1 _13771_ (
    .A(_4331_),
    .B(_3951_),
    .C(_4330_),
    .D(_4332_),
    .Y(_4333_)
);

INVX1 _13772_ (
    .A(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_4334_)
);

INVX1 _13773_ (
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_4335_)
);

OAI22X1 _13774_ (
    .A(_4335_),
    .B(_3898_),
    .C(_4334_),
    .D(_3865_),
    .Y(_4336_)
);

NOR2X1 _13775_ (
    .A(_4336_),
    .B(_4333_),
    .Y(_4337_)
);

INVX1 _13776_ (
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_4338_)
);

INVX1 _13777_ (
    .A(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_4339_)
);

NAND2X1 _13778_ (
    .A(_3873_),
    .B(_3878_),
    .Y(_4340_)
);

OAI22X1 _13779_ (
    .A(_4339_),
    .B(_3949_),
    .C(_4338_),
    .D(_4340_),
    .Y(_4341_)
);

INVX1 _13780_ (
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_4342_)
);

INVX1 _13781_ (
    .A(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_4343_)
);

OAI22X1 _13782_ (
    .A(_3910__bF$buf2),
    .B(_4342_),
    .C(_4343_),
    .D(_3905_),
    .Y(_4344_)
);

NOR2X1 _13783_ (
    .A(_4344_),
    .B(_4341_),
    .Y(_4345_)
);

NAND2X1 _13784_ (
    .A(_4337_),
    .B(_4345_),
    .Y(_4346_)
);

NOR2X1 _13785_ (
    .A(_4329_),
    .B(_4346_),
    .Y(_4347_)
);

AOI21X1 _13786_ (
    .A(_4347_),
    .B(_4317_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [8])
);

AOI22X1 _13787_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [9]),
    .C(\datapath_1.regfile_1.regOut[24] [9]),
    .D(_3902__bF$buf1),
    .Y(_4348_)
);

AOI22X1 _13788_ (
    .A(_3879__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[28] [9]),
    .C(_4070_),
    .D(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_4349_)
);

INVX1 _13789_ (
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_4350_)
);

INVX1 _13790_ (
    .A(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_4351_)
);

OAI22X1 _13791_ (
    .A(_3889__bF$buf0),
    .B(_4350_),
    .C(_4351_),
    .D(_3886__bF$buf1),
    .Y(_4352_)
);

INVX1 _13792_ (
    .A(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_4353_)
);

INVX1 _13793_ (
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_4354_)
);

OAI22X1 _13794_ (
    .A(_3923__bF$buf0),
    .B(_4354_),
    .C(_4353_),
    .D(_3929__bF$buf0),
    .Y(_4355_)
);

NOR2X1 _13795_ (
    .A(_4355_),
    .B(_4352_),
    .Y(_4356_)
);

NAND3X1 _13796_ (
    .A(_4349_),
    .B(_4348_),
    .C(_4356_),
    .Y(_4357_)
);

AOI22X1 _13797_ (
    .A(_3870__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [9]),
    .C(_3904__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_4358_)
);

AOI22X1 _13798_ (
    .A(_3899__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [9]),
    .C(_3952__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_4359_)
);

INVX1 _13799_ (
    .A(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_4360_)
);

INVX1 _13800_ (
    .A(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_4361_)
);

OAI22X1 _13801_ (
    .A(_3911_),
    .B(_4361_),
    .C(_4360_),
    .D(_3944__bF$buf0),
    .Y(_4362_)
);

INVX1 _13802_ (
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_4363_)
);

INVX1 _13803_ (
    .A(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_4364_)
);

OAI22X1 _13804_ (
    .A(_3916__bF$buf0),
    .B(_4363_),
    .C(_4364_),
    .D(_3915__bF$buf1),
    .Y(_4365_)
);

NOR2X1 _13805_ (
    .A(_4362_),
    .B(_4365_),
    .Y(_4366_)
);

NAND3X1 _13806_ (
    .A(_4359_),
    .B(_4358_),
    .C(_4366_),
    .Y(_4367_)
);

NOR2X1 _13807_ (
    .A(_4357_),
    .B(_4367_),
    .Y(_4368_)
);

AOI22X1 _13808_ (
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[6] [9]),
    .D(_4068__bF$buf2),
    .Y(_4369_)
);

AOI22X1 _13809_ (
    .A(_3876_),
    .B(\datapath_1.regfile_1.regOut[4] [9]),
    .C(\datapath_1.regfile_1.regOut[2] [9]),
    .D(_3975_),
    .Y(_4370_)
);

INVX1 _13810_ (
    .A(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_4371_)
);

INVX1 _13811_ (
    .A(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_4372_)
);

OAI22X1 _13812_ (
    .A(_4372_),
    .B(_3934__bF$buf1),
    .C(_3935__bF$buf2),
    .D(_4371_),
    .Y(_4373_)
);

INVX1 _13813_ (
    .A(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_4374_)
);

INVX1 _13814_ (
    .A(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_4375_)
);

OAI22X1 _13815_ (
    .A(_3928_),
    .B(_4374_),
    .C(_4375_),
    .D(_3956__bF$buf0),
    .Y(_4376_)
);

NOR2X1 _13816_ (
    .A(_4376_),
    .B(_4373_),
    .Y(_4377_)
);

NAND3X1 _13817_ (
    .A(_4370_),
    .B(_4369_),
    .C(_4377_),
    .Y(_4378_)
);

AOI22X1 _13818_ (
    .A(_3947__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [9]),
    .C(\datapath_1.regfile_1.regOut[29] [9]),
    .D(_3866__bF$buf0),
    .Y(_4379_)
);

AOI22X1 _13819_ (
    .A(_3950__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[9] [9]),
    .C(\datapath_1.regfile_1.regOut[31] [9]),
    .D(_3906__bF$buf0),
    .Y(_4380_)
);

INVX1 _13820_ (
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_4381_)
);

INVX1 _13821_ (
    .A(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_4382_)
);

OAI22X1 _13822_ (
    .A(_4382_),
    .B(_3957__bF$buf2),
    .C(_3961__bF$buf0),
    .D(_4381_),
    .Y(_4383_)
);

INVX1 _13823_ (
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_4384_)
);

INVX1 _13824_ (
    .A(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_4385_)
);

OAI22X1 _13825_ (
    .A(_4384_),
    .B(_3894__bF$buf0),
    .C(_4385_),
    .D(_3939__bF$buf0),
    .Y(_4386_)
);

NOR2X1 _13826_ (
    .A(_4386_),
    .B(_4383_),
    .Y(_4387_)
);

NAND3X1 _13827_ (
    .A(_4380_),
    .B(_4379_),
    .C(_4387_),
    .Y(_4388_)
);

NOR2X1 _13828_ (
    .A(_4388_),
    .B(_4378_),
    .Y(_4389_)
);

AOI21X1 _13829_ (
    .A(_4368_),
    .B(_4389_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [9])
);

INVX1 _13830_ (
    .A(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_4390_)
);

INVX1 _13831_ (
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_4391_)
);

OAI22X1 _13832_ (
    .A(_3923__bF$buf4),
    .B(_4391_),
    .C(_4390_),
    .D(_3929__bF$buf4),
    .Y(_4392_)
);

INVX1 _13833_ (
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_4393_)
);

INVX1 _13834_ (
    .A(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_4394_)
);

OAI22X1 _13835_ (
    .A(_3910__bF$buf1),
    .B(_4393_),
    .C(_4394_),
    .D(_3924__bF$buf1),
    .Y(_4395_)
);

NOR2X1 _13836_ (
    .A(_4392_),
    .B(_4395_),
    .Y(_4396_)
);

AOI22X1 _13837_ (
    .A(_4060__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [10]),
    .C(\datapath_1.regfile_1.regOut[21] [10]),
    .D(_3990_),
    .Y(_4397_)
);

INVX1 _13838_ (
    .A(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_4398_)
);

NOR2X1 _13839_ (
    .A(_4398_),
    .B(_3956__bF$buf4),
    .Y(_4399_)
);

AOI21X1 _13840_ (
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .B(_4062__bF$buf3),
    .C(_4399_),
    .Y(_4400_)
);

NAND3X1 _13841_ (
    .A(_4400_),
    .B(_4397_),
    .C(_4396_),
    .Y(_4401_)
);

INVX1 _13842_ (
    .A(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_4402_)
);

INVX1 _13843_ (
    .A(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_4403_)
);

OAI22X1 _13844_ (
    .A(_3865_),
    .B(_4402_),
    .C(_4403_),
    .D(_3893_),
    .Y(_4404_)
);

INVX1 _13845_ (
    .A(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_4405_)
);

INVX1 _13846_ (
    .A(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_4406_)
);

OAI22X1 _13847_ (
    .A(_4406_),
    .B(_3951_),
    .C(_4405_),
    .D(_4332_),
    .Y(_4407_)
);

NOR2X1 _13848_ (
    .A(_4404_),
    .B(_4407_),
    .Y(_4408_)
);

INVX1 _13849_ (
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_4409_)
);

INVX1 _13850_ (
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_4410_)
);

OAI22X1 _13851_ (
    .A(_3889__bF$buf4),
    .B(_4410_),
    .C(_4409_),
    .D(_3946_),
    .Y(_4411_)
);

INVX1 _13852_ (
    .A(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_4412_)
);

INVX1 _13853_ (
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_4413_)
);

OAI22X1 _13854_ (
    .A(_3944__bF$buf3),
    .B(_4412_),
    .C(_4413_),
    .D(_4340_),
    .Y(_4414_)
);

NOR2X1 _13855_ (
    .A(_4411_),
    .B(_4414_),
    .Y(_4415_)
);

NAND2X1 _13856_ (
    .A(_4408_),
    .B(_4415_),
    .Y(_4416_)
);

NOR2X1 _13857_ (
    .A(_4401_),
    .B(_4416_),
    .Y(_4417_)
);

INVX1 _13858_ (
    .A(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_4418_)
);

INVX1 _13859_ (
    .A(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_4419_)
);

OAI22X1 _13860_ (
    .A(_4419_),
    .B(_3949_),
    .C(_3886__bF$buf0),
    .D(_4418_),
    .Y(_4420_)
);

INVX1 _13861_ (
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_4421_)
);

INVX1 _13862_ (
    .A(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_4422_)
);

OAI22X1 _13863_ (
    .A(_3916__bF$buf4),
    .B(_4421_),
    .C(_4422_),
    .D(_3915__bF$buf0),
    .Y(_4423_)
);

NOR2X1 _13864_ (
    .A(_4423_),
    .B(_4420_),
    .Y(_4424_)
);

INVX1 _13865_ (
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_4425_)
);

INVX1 _13866_ (
    .A(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_4426_)
);

OAI22X1 _13867_ (
    .A(_3875__bF$buf2),
    .B(_4425_),
    .C(_4426_),
    .D(_3940__bF$buf0),
    .Y(_4427_)
);

INVX1 _13868_ (
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_4428_)
);

INVX1 _13869_ (
    .A(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_4429_)
);

OAI22X1 _13870_ (
    .A(_4428_),
    .B(_3894__bF$buf4),
    .C(_4429_),
    .D(_3939__bF$buf4),
    .Y(_4430_)
);

NOR2X1 _13871_ (
    .A(_4430_),
    .B(_4427_),
    .Y(_4431_)
);

NAND2X1 _13872_ (
    .A(_4431_),
    .B(_4424_),
    .Y(_4432_)
);

AOI22X1 _13873_ (
    .A(_3899__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [10]),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_4433_)
);

AOI22X1 _13874_ (
    .A(_3870__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [10]),
    .C(_4038_),
    .D(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_4434_)
);

INVX1 _13875_ (
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_4435_)
);

INVX1 _13876_ (
    .A(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_4436_)
);

OAI22X1 _13877_ (
    .A(_4436_),
    .B(_3957__bF$buf1),
    .C(_3961__bF$buf4),
    .D(_4435_),
    .Y(_4437_)
);

INVX1 _13878_ (
    .A(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_4438_)
);

INVX1 _13879_ (
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_4439_)
);

OAI22X1 _13880_ (
    .A(_4044_),
    .B(_4439_),
    .C(_4438_),
    .D(_3905_),
    .Y(_4440_)
);

NOR2X1 _13881_ (
    .A(_4437_),
    .B(_4440_),
    .Y(_4441_)
);

NAND3X1 _13882_ (
    .A(_4434_),
    .B(_4433_),
    .C(_4441_),
    .Y(_4442_)
);

NOR2X1 _13883_ (
    .A(_4432_),
    .B(_4442_),
    .Y(_4443_)
);

AOI21X1 _13884_ (
    .A(_4417_),
    .B(_4443_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [10])
);

INVX1 _13885_ (
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_4444_)
);

INVX1 _13886_ (
    .A(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_4445_)
);

OAI22X1 _13887_ (
    .A(_3875__bF$buf1),
    .B(_4444_),
    .C(_4445_),
    .D(_3940__bF$buf3),
    .Y(_4446_)
);

INVX1 _13888_ (
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_4447_)
);

INVX1 _13889_ (
    .A(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_4448_)
);

OAI22X1 _13890_ (
    .A(_4448_),
    .B(_3915__bF$buf3),
    .C(_3886__bF$buf3),
    .D(_4447_),
    .Y(_4449_)
);

NOR2X1 _13891_ (
    .A(_4446_),
    .B(_4449_),
    .Y(_4450_)
);

INVX1 _13892_ (
    .A(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_4451_)
);

NOR2X1 _13893_ (
    .A(_4451_),
    .B(_3956__bF$buf3),
    .Y(_4452_)
);

AOI21X1 _13894_ (
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .B(_3987_),
    .C(_4452_),
    .Y(_4453_)
);

AOI22X1 _13895_ (
    .A(_3899__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [11]),
    .C(\datapath_1.regfile_1.regOut[29] [11]),
    .D(_3866__bF$buf3),
    .Y(_4454_)
);

NAND3X1 _13896_ (
    .A(_4453_),
    .B(_4454_),
    .C(_4450_),
    .Y(_4455_)
);

INVX1 _13897_ (
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_4456_)
);

INVX1 _13898_ (
    .A(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_4457_)
);

OAI22X1 _13899_ (
    .A(_3894__bF$buf3),
    .B(_4456_),
    .C(_4457_),
    .D(_3893_),
    .Y(_4458_)
);

INVX1 _13900_ (
    .A(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_4459_)
);

INVX1 _13901_ (
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_4460_)
);

OAI22X1 _13902_ (
    .A(_4460_),
    .B(_3923__bF$buf3),
    .C(_4459_),
    .D(_3939__bF$buf3),
    .Y(_4461_)
);

NOR2X1 _13903_ (
    .A(_4461_),
    .B(_4458_),
    .Y(_4462_)
);

INVX1 _13904_ (
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_4463_)
);

NOR2X1 _13905_ (
    .A(_4463_),
    .B(_3916__bF$buf3),
    .Y(_4464_)
);

AOI21X1 _13906_ (
    .A(_4038_),
    .B(\datapath_1.regfile_1.regOut[22] [11]),
    .C(_4464_),
    .Y(_4465_)
);

AOI22X1 _13907_ (
    .A(_3879__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [11]),
    .C(_4070_),
    .D(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_4466_)
);

NAND3X1 _13908_ (
    .A(_4465_),
    .B(_4466_),
    .C(_4462_),
    .Y(_4467_)
);

NOR2X1 _13909_ (
    .A(_4467_),
    .B(_4455_),
    .Y(_4468_)
);

AOI22X1 _13910_ (
    .A(_3904__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [11]),
    .C(\datapath_1.regfile_1.regOut[9] [11]),
    .D(_3950__bF$buf0),
    .Y(_4469_)
);

AOI22X1 _13911_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [11]),
    .C(\datapath_1.regfile_1.regOut[24] [11]),
    .D(_3902__bF$buf0),
    .Y(_4470_)
);

INVX1 _13912_ (
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_4471_)
);

INVX1 _13913_ (
    .A(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_4472_)
);

OAI22X1 _13914_ (
    .A(_3911_),
    .B(_4471_),
    .C(_4472_),
    .D(_3928_),
    .Y(_4473_)
);

INVX1 _13915_ (
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_4474_)
);

INVX1 _13916_ (
    .A(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_4475_)
);

OAI22X1 _13917_ (
    .A(_3889__bF$buf3),
    .B(_4475_),
    .C(_4474_),
    .D(_3934__bF$buf0),
    .Y(_4476_)
);

NOR2X1 _13918_ (
    .A(_4473_),
    .B(_4476_),
    .Y(_4477_)
);

NAND3X1 _13919_ (
    .A(_4470_),
    .B(_4469_),
    .C(_4477_),
    .Y(_4478_)
);

INVX1 _13920_ (
    .A(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_4479_)
);

INVX1 _13921_ (
    .A(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_4480_)
);

OAI22X1 _13922_ (
    .A(_4480_),
    .B(_3929__bF$buf3),
    .C(_3957__bF$buf0),
    .D(_4479_),
    .Y(_4481_)
);

INVX1 _13923_ (
    .A(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_4482_)
);

INVX1 _13924_ (
    .A(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_4483_)
);

OAI22X1 _13925_ (
    .A(_4483_),
    .B(_3961__bF$buf3),
    .C(_4482_),
    .D(_3944__bF$buf2),
    .Y(_4484_)
);

NOR2X1 _13926_ (
    .A(_4481_),
    .B(_4484_),
    .Y(_4485_)
);

AOI22X1 _13927_ (
    .A(_3947__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [11]),
    .C(\datapath_1.regfile_1.regOut[30] [11]),
    .D(_3870__bF$buf3),
    .Y(_4486_)
);

AOI22X1 _13928_ (
    .A(_3952__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [11]),
    .C(\datapath_1.regfile_1.regOut[31] [11]),
    .D(_3906__bF$buf3),
    .Y(_4487_)
);

NAND3X1 _13929_ (
    .A(_4486_),
    .B(_4487_),
    .C(_4485_),
    .Y(_4488_)
);

NOR2X1 _13930_ (
    .A(_4478_),
    .B(_4488_),
    .Y(_4489_)
);

AOI21X1 _13931_ (
    .A(_4489_),
    .B(_4468_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [11])
);

INVX1 _13932_ (
    .A(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_4490_)
);

INVX1 _13933_ (
    .A(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_4491_)
);

OAI22X1 _13934_ (
    .A(_4491_),
    .B(_3956__bF$buf2),
    .C(_3905_),
    .D(_4490_),
    .Y(_4492_)
);

INVX1 _13935_ (
    .A(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_4493_)
);

INVX1 _13936_ (
    .A(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_4494_)
);

OAI22X1 _13937_ (
    .A(_4494_),
    .B(_3961__bF$buf2),
    .C(_4493_),
    .D(_3944__bF$buf1),
    .Y(_4495_)
);

NOR2X1 _13938_ (
    .A(_4495_),
    .B(_4492_),
    .Y(_4496_)
);

AOI22X1 _13939_ (
    .A(_4062__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [12]),
    .C(\datapath_1.regfile_1.regOut[7] [12]),
    .D(_4060__bF$buf3),
    .Y(_4497_)
);

AOI22X1 _13940_ (
    .A(_3902__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [12]),
    .C(\datapath_1.regfile_1.regOut[26] [12]),
    .D(_4070_),
    .Y(_4498_)
);

NAND3X1 _13941_ (
    .A(_4497_),
    .B(_4498_),
    .C(_4496_),
    .Y(_4499_)
);

INVX1 _13942_ (
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_4500_)
);

INVX1 _13943_ (
    .A(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_4501_)
);

OAI22X1 _13944_ (
    .A(_4500_),
    .B(_3894__bF$buf2),
    .C(_4501_),
    .D(_3939__bF$buf2),
    .Y(_4502_)
);

INVX1 _13945_ (
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_4503_)
);

INVX1 _13946_ (
    .A(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_4504_)
);

OAI22X1 _13947_ (
    .A(_4504_),
    .B(_3957__bF$buf4),
    .C(_3869_),
    .D(_4503_),
    .Y(_4505_)
);

NOR2X1 _13948_ (
    .A(_4502_),
    .B(_4505_),
    .Y(_4506_)
);

AOI22X1 _13949_ (
    .A(_3876_),
    .B(\datapath_1.regfile_1.regOut[4] [12]),
    .C(\datapath_1.regfile_1.regOut[2] [12]),
    .D(_3975_),
    .Y(_4507_)
);

INVX1 _13950_ (
    .A(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_4508_)
);

NOR2X1 _13951_ (
    .A(_4508_),
    .B(_3923__bF$buf2),
    .Y(_4509_)
);

AOI21X1 _13952_ (
    .A(_3987_),
    .B(\datapath_1.regfile_1.regOut[0] [12]),
    .C(_4509_),
    .Y(_4510_)
);

NAND3X1 _13953_ (
    .A(_4507_),
    .B(_4510_),
    .C(_4506_),
    .Y(_4511_)
);

NOR2X1 _13954_ (
    .A(_4511_),
    .B(_4499_),
    .Y(_4512_)
);

AOI22X1 _13955_ (
    .A(_3904__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [12]),
    .C(\datapath_1.regfile_1.regOut[21] [12]),
    .D(_3990_),
    .Y(_4513_)
);

AOI22X1 _13956_ (
    .A(_3899__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [12]),
    .C(_4087_),
    .D(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_4514_)
);

INVX1 _13957_ (
    .A(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_4515_)
);

INVX1 _13958_ (
    .A(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_4516_)
);

OAI22X1 _13959_ (
    .A(_3889__bF$buf2),
    .B(_4516_),
    .C(_4515_),
    .D(_3951_),
    .Y(_4517_)
);

INVX1 _13960_ (
    .A(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_4518_)
);

INVX1 _13961_ (
    .A(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_4519_)
);

OAI22X1 _13962_ (
    .A(_4519_),
    .B(_3962__bF$buf2),
    .C(_4518_),
    .D(_3935__bF$buf1),
    .Y(_4520_)
);

NOR2X1 _13963_ (
    .A(_4517_),
    .B(_4520_),
    .Y(_4521_)
);

NAND3X1 _13964_ (
    .A(_4513_),
    .B(_4514_),
    .C(_4521_),
    .Y(_4522_)
);

AOI22X1 _13965_ (
    .A(_3947__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .C(_4068__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_4523_)
);

INVX1 _13966_ (
    .A(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_4524_)
);

NOR2X1 _13967_ (
    .A(_4524_),
    .B(_3929__bF$buf2),
    .Y(_4525_)
);

AOI21X1 _13968_ (
    .A(_3866__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [12]),
    .C(_4525_),
    .Y(_4526_)
);

INVX1 _13969_ (
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_4527_)
);

INVX1 _13970_ (
    .A(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_4528_)
);

OAI22X1 _13971_ (
    .A(_3916__bF$buf2),
    .B(_4527_),
    .C(_4528_),
    .D(_3886__bF$buf2),
    .Y(_4529_)
);

INVX1 _13972_ (
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_4530_)
);

INVX1 _13973_ (
    .A(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_4531_)
);

OAI22X1 _13974_ (
    .A(_4044_),
    .B(_4530_),
    .C(_4531_),
    .D(_3949_),
    .Y(_4532_)
);

NOR2X1 _13975_ (
    .A(_4532_),
    .B(_4529_),
    .Y(_4533_)
);

NAND3X1 _13976_ (
    .A(_4526_),
    .B(_4523_),
    .C(_4533_),
    .Y(_4534_)
);

NOR2X1 _13977_ (
    .A(_4522_),
    .B(_4534_),
    .Y(_4535_)
);

AOI21X1 _13978_ (
    .A(_4512_),
    .B(_4535_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [12])
);

INVX1 _13979_ (
    .A(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_4536_)
);

INVX1 _13980_ (
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_4537_)
);

OAI22X1 _13981_ (
    .A(_3894__bF$buf1),
    .B(_4537_),
    .C(_4536_),
    .D(_3961__bF$buf1),
    .Y(_4538_)
);

INVX1 _13982_ (
    .A(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_4539_)
);

INVX1 _13983_ (
    .A(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_4540_)
);

OAI22X1 _13984_ (
    .A(_4540_),
    .B(_3940__bF$buf2),
    .C(_3946_),
    .D(_4539_),
    .Y(_4541_)
);

NOR2X1 _13985_ (
    .A(_4538_),
    .B(_4541_),
    .Y(_4542_)
);

INVX1 _13986_ (
    .A(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_4543_)
);

NOR2X1 _13987_ (
    .A(_4543_),
    .B(_3956__bF$buf1),
    .Y(_4544_)
);

AOI21X1 _13988_ (
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .B(_3879__bF$buf0),
    .C(_4544_),
    .Y(_4545_)
);

AOI22X1 _13989_ (
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .B(_3876_),
    .C(\datapath_1.regfile_1.regOut[26] [13]),
    .D(_4070_),
    .Y(_4546_)
);

NAND3X1 _13990_ (
    .A(_4545_),
    .B(_4546_),
    .C(_4542_),
    .Y(_4547_)
);

INVX1 _13991_ (
    .A(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_4548_)
);

INVX1 _13992_ (
    .A(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_4549_)
);

OAI22X1 _13993_ (
    .A(_4549_),
    .B(_3923__bF$buf1),
    .C(_4548_),
    .D(_3898_),
    .Y(_4550_)
);

INVX1 _13994_ (
    .A(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_4551_)
);

INVX1 _13995_ (
    .A(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_4552_)
);

OAI22X1 _13996_ (
    .A(_4552_),
    .B(_3929__bF$buf1),
    .C(_4551_),
    .D(_3865_),
    .Y(_4553_)
);

NOR2X1 _13997_ (
    .A(_4550_),
    .B(_4553_),
    .Y(_4554_)
);

INVX1 _13998_ (
    .A(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_4555_)
);

NOR2X1 _13999_ (
    .A(_4555_),
    .B(_3939__bF$buf1),
    .Y(_4556_)
);

AOI21X1 _14000_ (
    .A(_3952__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [13]),
    .C(_4556_),
    .Y(_4557_)
);

AOI22X1 _14001_ (
    .A(_3870__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [13]),
    .C(_3902__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_4558_)
);

NAND3X1 _14002_ (
    .A(_4557_),
    .B(_4558_),
    .C(_4554_),
    .Y(_4559_)
);

NOR2X1 _14003_ (
    .A(_4547_),
    .B(_4559_),
    .Y(_4560_)
);

AOI22X1 _14004_ (
    .A(_4060__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [13]),
    .C(\datapath_1.regfile_1.regOut[6] [13]),
    .D(_4068__bF$buf0),
    .Y(_4561_)
);

AOI22X1 _14005_ (
    .A(_4099_),
    .B(\datapath_1.regfile_1.regOut[13] [13]),
    .C(\datapath_1.regfile_1.regOut[25] [13]),
    .D(_3945_),
    .Y(_4562_)
);

INVX1 _14006_ (
    .A(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_4563_)
);

INVX1 _14007_ (
    .A(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_4564_)
);

OAI22X1 _14008_ (
    .A(_4563_),
    .B(_3910__bF$buf0),
    .C(_4564_),
    .D(_3911_),
    .Y(_4565_)
);

INVX1 _14009_ (
    .A(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_4566_)
);

INVX1 _14010_ (
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_4567_)
);

OAI22X1 _14011_ (
    .A(_4567_),
    .B(_3916__bF$buf1),
    .C(_3889__bF$buf1),
    .D(_4566_),
    .Y(_4568_)
);

NOR2X1 _14012_ (
    .A(_4568_),
    .B(_4565_),
    .Y(_4569_)
);

NAND3X1 _14013_ (
    .A(_4562_),
    .B(_4561_),
    .C(_4569_),
    .Y(_4570_)
);

AOI22X1 _14014_ (
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[9] [13]),
    .D(_3950__bF$buf3),
    .Y(_4571_)
);

AOI22X1 _14015_ (
    .A(_3904__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [13]),
    .C(\datapath_1.regfile_1.regOut[10] [13]),
    .D(_4087_),
    .Y(_4572_)
);

NAND2X1 _14016_ (
    .A(_4571_),
    .B(_4572_),
    .Y(_4573_)
);

AOI22X1 _14017_ (
    .A(_4038_),
    .B(\datapath_1.regfile_1.regOut[22] [13]),
    .C(_3990_),
    .D(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_4574_)
);

AOI22X1 _14018_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [13]),
    .C(\datapath_1.regfile_1.regOut[31] [13]),
    .D(_3906__bF$buf2),
    .Y(_4575_)
);

NAND2X1 _14019_ (
    .A(_4575_),
    .B(_4574_),
    .Y(_4576_)
);

NOR3X1 _14020_ (
    .A(_4573_),
    .B(_4576_),
    .C(_4570_),
    .Y(_4577_)
);

AOI21X1 _14021_ (
    .A(_4577_),
    .B(_4560_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [13])
);

AOI22X1 _14022_ (
    .A(_4070_),
    .B(\datapath_1.regfile_1.regOut[26] [14]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_4578_)
);

AOI22X1 _14023_ (
    .A(_3952__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [14]),
    .C(\datapath_1.regfile_1.regOut[24] [14]),
    .D(_3902__bF$buf2),
    .Y(_4579_)
);

INVX1 _14024_ (
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_4580_)
);

INVX1 _14025_ (
    .A(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_4581_)
);

OAI22X1 _14026_ (
    .A(_4580_),
    .B(_3894__bF$buf0),
    .C(_4581_),
    .D(_3929__bF$buf0),
    .Y(_4582_)
);

INVX1 _14027_ (
    .A(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_4583_)
);

INVX1 _14028_ (
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_4584_)
);

OAI22X1 _14029_ (
    .A(_4584_),
    .B(_3916__bF$buf0),
    .C(_3889__bF$buf0),
    .D(_4583_),
    .Y(_4585_)
);

NOR2X1 _14030_ (
    .A(_4585_),
    .B(_4582_),
    .Y(_4586_)
);

NAND3X1 _14031_ (
    .A(_4579_),
    .B(_4578_),
    .C(_4586_),
    .Y(_4587_)
);

AOI22X1 _14032_ (
    .A(_3866__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [14]),
    .C(_3904__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_4588_)
);

AOI22X1 _14033_ (
    .A(_3947__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [14]),
    .C(_3899__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_4589_)
);

INVX1 _14034_ (
    .A(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_4590_)
);

INVX1 _14035_ (
    .A(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_4591_)
);

OAI22X1 _14036_ (
    .A(_3911_),
    .B(_4590_),
    .C(_4591_),
    .D(_3939__bF$buf0),
    .Y(_4592_)
);

INVX1 _14037_ (
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_4593_)
);

INVX1 _14038_ (
    .A(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_4594_)
);

OAI22X1 _14039_ (
    .A(_4594_),
    .B(_3915__bF$buf2),
    .C(_3886__bF$buf1),
    .D(_4593_),
    .Y(_4595_)
);

NOR2X1 _14040_ (
    .A(_4592_),
    .B(_4595_),
    .Y(_4596_)
);

NAND3X1 _14041_ (
    .A(_4589_),
    .B(_4588_),
    .C(_4596_),
    .Y(_4597_)
);

NOR2X1 _14042_ (
    .A(_4587_),
    .B(_4597_),
    .Y(_4598_)
);

INVX1 _14043_ (
    .A(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_4599_)
);

INVX1 _14044_ (
    .A(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_4600_)
);

OAI22X1 _14045_ (
    .A(_4600_),
    .B(_3928_),
    .C(_4599_),
    .D(_3893_),
    .Y(_4601_)
);

INVX1 _14046_ (
    .A(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_4602_)
);

INVX1 _14047_ (
    .A(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_4603_)
);

OAI22X1 _14048_ (
    .A(_4603_),
    .B(_3923__bF$buf0),
    .C(_4602_),
    .D(_4044_),
    .Y(_4604_)
);

NOR2X1 _14049_ (
    .A(_4604_),
    .B(_4601_),
    .Y(_4605_)
);

AOI22X1 _14050_ (
    .A(_4038_),
    .B(\datapath_1.regfile_1.regOut[22] [14]),
    .C(_3990_),
    .D(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_4606_)
);

AOI22X1 _14051_ (
    .A(_3876_),
    .B(\datapath_1.regfile_1.regOut[4] [14]),
    .C(\datapath_1.regfile_1.regOut[2] [14]),
    .D(_3975_),
    .Y(_4607_)
);

NAND3X1 _14052_ (
    .A(_4606_),
    .B(_4607_),
    .C(_4605_),
    .Y(_4608_)
);

AOI22X1 _14053_ (
    .A(_3870__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[30] [14]),
    .C(_3906__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_4609_)
);

AOI22X1 _14054_ (
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[9] [14]),
    .D(_3950__bF$buf2),
    .Y(_4610_)
);

INVX1 _14055_ (
    .A(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_4611_)
);

INVX1 _14056_ (
    .A(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_4612_)
);

OAI22X1 _14057_ (
    .A(_3957__bF$buf3),
    .B(_4611_),
    .C(_4612_),
    .D(_3956__bF$buf0),
    .Y(_4613_)
);

INVX1 _14058_ (
    .A(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_4614_)
);

INVX1 _14059_ (
    .A(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_4615_)
);

OAI22X1 _14060_ (
    .A(_4615_),
    .B(_3961__bF$buf0),
    .C(_3962__bF$buf1),
    .D(_4614_),
    .Y(_4616_)
);

NOR2X1 _14061_ (
    .A(_4616_),
    .B(_4613_),
    .Y(_4617_)
);

NAND3X1 _14062_ (
    .A(_4610_),
    .B(_4609_),
    .C(_4617_),
    .Y(_4618_)
);

NOR2X1 _14063_ (
    .A(_4608_),
    .B(_4618_),
    .Y(_4619_)
);

AOI21X1 _14064_ (
    .A(_4619_),
    .B(_4598_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [14])
);

INVX1 _14065_ (
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_4620_)
);

INVX1 _14066_ (
    .A(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_4621_)
);

OAI22X1 _14067_ (
    .A(_4620_),
    .B(_3910__bF$buf3),
    .C(_4621_),
    .D(_4044_),
    .Y(_4622_)
);

INVX1 _14068_ (
    .A(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_4623_)
);

INVX1 _14069_ (
    .A(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_4624_)
);

OAI22X1 _14070_ (
    .A(_4624_),
    .B(_3929__bF$buf4),
    .C(_3962__bF$buf0),
    .D(_4623_),
    .Y(_4625_)
);

NOR2X1 _14071_ (
    .A(_4622_),
    .B(_4625_),
    .Y(_4626_)
);

AOI22X1 _14072_ (
    .A(_3866__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [15]),
    .C(\datapath_1.regfile_1.regOut[31] [15]),
    .D(_3906__bF$buf0),
    .Y(_4627_)
);

INVX1 _14073_ (
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_4628_)
);

NOR2X1 _14074_ (
    .A(_4628_),
    .B(_3889__bF$buf4),
    .Y(_4629_)
);

AOI21X1 _14075_ (
    .A(_3989_),
    .B(\datapath_1.regfile_1.regOut[15] [15]),
    .C(_4629_),
    .Y(_4630_)
);

NAND3X1 _14076_ (
    .A(_4627_),
    .B(_4630_),
    .C(_4626_),
    .Y(_4631_)
);

INVX1 _14077_ (
    .A(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_4632_)
);

NOR2X1 _14078_ (
    .A(_4632_),
    .B(_3956__bF$buf4),
    .Y(_4633_)
);

AOI21X1 _14079_ (
    .A(\datapath_1.regfile_1.regOut[6] [15]),
    .B(_4068__bF$buf3),
    .C(_4633_),
    .Y(_4634_)
);

INVX1 _14080_ (
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_4635_)
);

NOR2X1 _14081_ (
    .A(_4635_),
    .B(_3894__bF$buf4),
    .Y(_4636_)
);

AOI21X1 _14082_ (
    .A(_3904__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [15]),
    .C(_4636_),
    .Y(_4637_)
);

INVX1 _14083_ (
    .A(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_4638_)
);

INVX1 _14084_ (
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_4639_)
);

OAI22X1 _14085_ (
    .A(_3939__bF$buf4),
    .B(_4639_),
    .C(_4638_),
    .D(_3924__bF$buf0),
    .Y(_4640_)
);

INVX1 _14086_ (
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_4641_)
);

INVX1 _14087_ (
    .A(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_4642_)
);

OAI22X1 _14088_ (
    .A(_3916__bF$buf4),
    .B(_4641_),
    .C(_4642_),
    .D(_3915__bF$buf1),
    .Y(_4643_)
);

NOR2X1 _14089_ (
    .A(_4640_),
    .B(_4643_),
    .Y(_4644_)
);

NAND3X1 _14090_ (
    .A(_4637_),
    .B(_4634_),
    .C(_4644_),
    .Y(_4645_)
);

NOR2X1 _14091_ (
    .A(_4631_),
    .B(_4645_),
    .Y(_4646_)
);

AOI22X1 _14092_ (
    .A(_4062__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [15]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_4647_)
);

AOI22X1 _14093_ (
    .A(_3952__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [15]),
    .C(\datapath_1.regfile_1.regOut[24] [15]),
    .D(_3902__bF$buf1),
    .Y(_4648_)
);

INVX1 _14094_ (
    .A(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_4649_)
);

INVX1 _14095_ (
    .A(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_4650_)
);

OAI22X1 _14096_ (
    .A(_3923__bF$buf4),
    .B(_4650_),
    .C(_4649_),
    .D(_3940__bF$buf1),
    .Y(_4651_)
);

INVX1 _14097_ (
    .A(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_4652_)
);

INVX1 _14098_ (
    .A(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_4653_)
);

OAI22X1 _14099_ (
    .A(_4653_),
    .B(_3934__bF$buf3),
    .C(_3935__bF$buf0),
    .D(_4652_),
    .Y(_4654_)
);

NOR2X1 _14100_ (
    .A(_4651_),
    .B(_4654_),
    .Y(_4655_)
);

NAND3X1 _14101_ (
    .A(_4648_),
    .B(_4647_),
    .C(_4655_),
    .Y(_4656_)
);

INVX1 _14102_ (
    .A(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_4657_)
);

INVX1 _14103_ (
    .A(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_4658_)
);

OAI22X1 _14104_ (
    .A(_4658_),
    .B(_3957__bF$buf2),
    .C(_3961__bF$buf4),
    .D(_4657_),
    .Y(_4659_)
);

INVX1 _14105_ (
    .A(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_4660_)
);

INVX1 _14106_ (
    .A(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_4661_)
);

OAI22X1 _14107_ (
    .A(_3928_),
    .B(_4661_),
    .C(_4660_),
    .D(_3949_),
    .Y(_4662_)
);

NOR2X1 _14108_ (
    .A(_4659_),
    .B(_4662_),
    .Y(_4663_)
);

AOI22X1 _14109_ (
    .A(_3947__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [15]),
    .C(_3899__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_4664_)
);

AOI22X1 _14110_ (
    .A(_3870__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [15]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_4665_)
);

NAND3X1 _14111_ (
    .A(_4664_),
    .B(_4665_),
    .C(_4663_),
    .Y(_4666_)
);

NOR2X1 _14112_ (
    .A(_4656_),
    .B(_4666_),
    .Y(_4667_)
);

AOI21X1 _14113_ (
    .A(_4667_),
    .B(_4646_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [15])
);

INVX1 _14114_ (
    .A(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_4668_)
);

INVX1 _14115_ (
    .A(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_4669_)
);

OAI22X1 _14116_ (
    .A(_3894__bF$buf3),
    .B(_4668_),
    .C(_4669_),
    .D(_3915__bF$buf0),
    .Y(_4670_)
);

INVX1 _14117_ (
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_4671_)
);

INVX1 _14118_ (
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_4672_)
);

OAI22X1 _14119_ (
    .A(_3916__bF$buf3),
    .B(_4672_),
    .C(_4671_),
    .D(_3946_),
    .Y(_4673_)
);

NOR2X1 _14120_ (
    .A(_4673_),
    .B(_4670_),
    .Y(_4674_)
);

INVX1 _14121_ (
    .A(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_4675_)
);

INVX1 _14122_ (
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_4676_)
);

OAI22X1 _14123_ (
    .A(_3875__bF$buf0),
    .B(_4676_),
    .C(_4675_),
    .D(_3957__bF$buf1),
    .Y(_4677_)
);

INVX1 _14124_ (
    .A(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_4678_)
);

INVX1 _14125_ (
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_4679_)
);

OAI22X1 _14126_ (
    .A(_3923__bF$buf3),
    .B(_4679_),
    .C(_4678_),
    .D(_3929__bF$buf3),
    .Y(_4680_)
);

NOR2X1 _14127_ (
    .A(_4680_),
    .B(_4677_),
    .Y(_4681_)
);

NAND2X1 _14128_ (
    .A(_4674_),
    .B(_4681_),
    .Y(_4682_)
);

INVX1 _14129_ (
    .A(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_4683_)
);

INVX1 _14130_ (
    .A(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_4684_)
);

OAI22X1 _14131_ (
    .A(_3961__bF$buf3),
    .B(_4683_),
    .C(_4684_),
    .D(_3949_),
    .Y(_4685_)
);

INVX1 _14132_ (
    .A(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_4686_)
);

INVX1 _14133_ (
    .A(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_4687_)
);

OAI22X1 _14134_ (
    .A(_3939__bF$buf3),
    .B(_4687_),
    .C(_4686_),
    .D(_3934__bF$buf2),
    .Y(_4688_)
);

NOR2X1 _14135_ (
    .A(_4688_),
    .B(_4685_),
    .Y(_4689_)
);

AOI22X1 _14136_ (
    .A(_3952__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [16]),
    .C(\datapath_1.regfile_1.regOut[24] [16]),
    .D(_3902__bF$buf0),
    .Y(_4690_)
);

AOI22X1 _14137_ (
    .A(_3904__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [16]),
    .C(\datapath_1.regfile_1.regOut[22] [16]),
    .D(_4038_),
    .Y(_4691_)
);

NAND3X1 _14138_ (
    .A(_4690_),
    .B(_4691_),
    .C(_4689_),
    .Y(_4692_)
);

NOR2X1 _14139_ (
    .A(_4682_),
    .B(_4692_),
    .Y(_4693_)
);

INVX1 _14140_ (
    .A(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_4694_)
);

INVX1 _14141_ (
    .A(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_4695_)
);

OAI22X1 _14142_ (
    .A(_3869_),
    .B(_4694_),
    .C(_4695_),
    .D(_3944__bF$buf0),
    .Y(_4696_)
);

INVX1 _14143_ (
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_4697_)
);

INVX1 _14144_ (
    .A(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_4698_)
);

OAI22X1 _14145_ (
    .A(_3889__bF$buf3),
    .B(_4697_),
    .C(_4698_),
    .D(_3893_),
    .Y(_4699_)
);

NOR2X1 _14146_ (
    .A(_4699_),
    .B(_4696_),
    .Y(_4700_)
);

AOI22X1 _14147_ (
    .A(_3899__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [16]),
    .C(\datapath_1.regfile_1.regOut[29] [16]),
    .D(_3866__bF$buf3),
    .Y(_4701_)
);

AOI22X1 _14148_ (
    .A(_3879__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [16]),
    .C(\datapath_1.regfile_1.regOut[31] [16]),
    .D(_3906__bF$buf3),
    .Y(_4702_)
);

NAND3X1 _14149_ (
    .A(_4701_),
    .B(_4702_),
    .C(_4700_),
    .Y(_4703_)
);

INVX1 _14150_ (
    .A(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_4704_)
);

INVX1 _14151_ (
    .A(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_4705_)
);

OAI22X1 _14152_ (
    .A(_4704_),
    .B(_3924__bF$buf3),
    .C(_3886__bF$buf0),
    .D(_4705_),
    .Y(_4706_)
);

INVX1 _14153_ (
    .A(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_4707_)
);

INVX1 _14154_ (
    .A(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_4708_)
);

OAI22X1 _14155_ (
    .A(_3962__bF$buf3),
    .B(_4707_),
    .C(_4708_),
    .D(_3956__bF$buf3),
    .Y(_4709_)
);

NOR2X1 _14156_ (
    .A(_4709_),
    .B(_4706_),
    .Y(_4710_)
);

AOI22X1 _14157_ (
    .A(_4060__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [16]),
    .C(_3975_),
    .D(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_4711_)
);

AOI22X1 _14158_ (
    .A(_3987_),
    .B(\datapath_1.regfile_1.regOut[0] [16]),
    .C(_4062__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_4712_)
);

NAND3X1 _14159_ (
    .A(_4711_),
    .B(_4712_),
    .C(_4710_),
    .Y(_4713_)
);

NOR2X1 _14160_ (
    .A(_4713_),
    .B(_4703_),
    .Y(_4714_)
);

AOI21X1 _14161_ (
    .A(_4714_),
    .B(_4693_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [16])
);

INVX1 _14162_ (
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_4715_)
);

INVX1 _14163_ (
    .A(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_4716_)
);

OAI22X1 _14164_ (
    .A(_3894__bF$buf2),
    .B(_4715_),
    .C(_4716_),
    .D(_3915__bF$buf3),
    .Y(_4717_)
);

INVX1 _14165_ (
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_4718_)
);

INVX1 _14166_ (
    .A(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_4719_)
);

OAI22X1 _14167_ (
    .A(_4718_),
    .B(_3944__bF$buf3),
    .C(_3886__bF$buf3),
    .D(_4719_),
    .Y(_4720_)
);

NOR2X1 _14168_ (
    .A(_4717_),
    .B(_4720_),
    .Y(_4721_)
);

INVX1 _14169_ (
    .A(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_4722_)
);

INVX1 _14170_ (
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_4723_)
);

OAI22X1 _14171_ (
    .A(_3875__bF$buf3),
    .B(_4723_),
    .C(_4722_),
    .D(_3957__bF$buf0),
    .Y(_4724_)
);

INVX1 _14172_ (
    .A(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_4725_)
);

INVX1 _14173_ (
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_4726_)
);

OAI22X1 _14174_ (
    .A(_3923__bF$buf2),
    .B(_4726_),
    .C(_4725_),
    .D(_3929__bF$buf2),
    .Y(_4727_)
);

NOR2X1 _14175_ (
    .A(_4727_),
    .B(_4724_),
    .Y(_4728_)
);

NAND2X1 _14176_ (
    .A(_4728_),
    .B(_4721_),
    .Y(_4729_)
);

INVX1 _14177_ (
    .A(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_4730_)
);

INVX1 _14178_ (
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_4731_)
);

OAI22X1 _14179_ (
    .A(_3961__bF$buf2),
    .B(_4730_),
    .C(_4731_),
    .D(_3949_),
    .Y(_4732_)
);

INVX1 _14180_ (
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_4733_)
);

INVX1 _14181_ (
    .A(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_4734_)
);

OAI22X1 _14182_ (
    .A(_3939__bF$buf2),
    .B(_4734_),
    .C(_4733_),
    .D(_3934__bF$buf1),
    .Y(_4735_)
);

NOR2X1 _14183_ (
    .A(_4735_),
    .B(_4732_),
    .Y(_4736_)
);

AOI22X1 _14184_ (
    .A(_3952__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [17]),
    .C(\datapath_1.regfile_1.regOut[24] [17]),
    .D(_3902__bF$buf4),
    .Y(_4737_)
);

AOI22X1 _14185_ (
    .A(_3904__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [17]),
    .C(\datapath_1.regfile_1.regOut[22] [17]),
    .D(_4038_),
    .Y(_4738_)
);

NAND3X1 _14186_ (
    .A(_4737_),
    .B(_4738_),
    .C(_4736_),
    .Y(_4739_)
);

NOR2X1 _14187_ (
    .A(_4729_),
    .B(_4739_),
    .Y(_4740_)
);

INVX1 _14188_ (
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_4741_)
);

INVX1 _14189_ (
    .A(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_4742_)
);

OAI22X1 _14190_ (
    .A(_3910__bF$buf2),
    .B(_4741_),
    .C(_4742_),
    .D(_3905_),
    .Y(_4743_)
);

INVX1 _14191_ (
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_4744_)
);

INVX1 _14192_ (
    .A(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_4745_)
);

OAI22X1 _14193_ (
    .A(_3889__bF$buf2),
    .B(_4744_),
    .C(_4745_),
    .D(_3893_),
    .Y(_4746_)
);

NOR2X1 _14194_ (
    .A(_4746_),
    .B(_4743_),
    .Y(_4747_)
);

AOI22X1 _14195_ (
    .A(_3899__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [17]),
    .C(\datapath_1.regfile_1.regOut[28] [17]),
    .D(_3879__bF$buf2),
    .Y(_4748_)
);

AOI22X1 _14196_ (
    .A(_3870__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[30] [17]),
    .C(_3866__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_4749_)
);

NAND3X1 _14197_ (
    .A(_4748_),
    .B(_4749_),
    .C(_4747_),
    .Y(_4750_)
);

INVX1 _14198_ (
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_4751_)
);

INVX1 _14199_ (
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_4752_)
);

OAI22X1 _14200_ (
    .A(_3916__bF$buf2),
    .B(_4752_),
    .C(_4751_),
    .D(_3946_),
    .Y(_4753_)
);

INVX1 _14201_ (
    .A(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_4754_)
);

INVX1 _14202_ (
    .A(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_4755_)
);

OAI22X1 _14203_ (
    .A(_3962__bF$buf2),
    .B(_4754_),
    .C(_4755_),
    .D(_3956__bF$buf2),
    .Y(_4756_)
);

NOR2X1 _14204_ (
    .A(_4753_),
    .B(_4756_),
    .Y(_4757_)
);

AOI22X1 _14205_ (
    .A(_4060__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [17]),
    .C(_3975_),
    .D(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_4758_)
);

AOI22X1 _14206_ (
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .B(_4062__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[26] [17]),
    .D(_4070_),
    .Y(_4759_)
);

NAND3X1 _14207_ (
    .A(_4759_),
    .B(_4758_),
    .C(_4757_),
    .Y(_4760_)
);

NOR2X1 _14208_ (
    .A(_4760_),
    .B(_4750_),
    .Y(_4761_)
);

AOI21X1 _14209_ (
    .A(_4761_),
    .B(_4740_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [17])
);

INVX1 _14210_ (
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_4762_)
);

NOR2X1 _14211_ (
    .A(_4762_),
    .B(_3961__bF$buf1),
    .Y(_4763_)
);

AOI21X1 _14212_ (
    .A(\datapath_1.regfile_1.regOut[13] [18]),
    .B(_4099_),
    .C(_4763_),
    .Y(_4764_)
);

AOI22X1 _14213_ (
    .A(_3945_),
    .B(\datapath_1.regfile_1.regOut[25] [18]),
    .C(_4068__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_4765_)
);

INVX1 _14214_ (
    .A(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_4766_)
);

INVX1 _14215_ (
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_4767_)
);

OAI22X1 _14216_ (
    .A(_4767_),
    .B(_3916__bF$buf1),
    .C(_3889__bF$buf1),
    .D(_4766_),
    .Y(_4768_)
);

INVX1 _14217_ (
    .A(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_4769_)
);

INVX1 _14218_ (
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_4770_)
);

OAI22X1 _14219_ (
    .A(_4770_),
    .B(_3928_),
    .C(_4769_),
    .D(_3915__bF$buf2),
    .Y(_4771_)
);

NOR2X1 _14220_ (
    .A(_4768_),
    .B(_4771_),
    .Y(_4772_)
);

NAND3X1 _14221_ (
    .A(_4764_),
    .B(_4765_),
    .C(_4772_),
    .Y(_4773_)
);

INVX1 _14222_ (
    .A(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_4774_)
);

INVX1 _14223_ (
    .A(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_4775_)
);

OAI22X1 _14224_ (
    .A(_4775_),
    .B(_3929__bF$buf1),
    .C(_4774_),
    .D(_3865_),
    .Y(_4776_)
);

INVX1 _14225_ (
    .A(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_4777_)
);

INVX1 _14226_ (
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_4778_)
);

OAI22X1 _14227_ (
    .A(_3894__bF$buf1),
    .B(_4778_),
    .C(_4777_),
    .D(_3905_),
    .Y(_4779_)
);

NOR2X1 _14228_ (
    .A(_4776_),
    .B(_4779_),
    .Y(_4780_)
);

INVX1 _14229_ (
    .A(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_4781_)
);

NOR2X1 _14230_ (
    .A(_4781_),
    .B(_3956__bF$buf1),
    .Y(_4782_)
);

AOI21X1 _14231_ (
    .A(\datapath_1.regfile_1.regOut[23] [18]),
    .B(_3899__bF$buf0),
    .C(_4782_),
    .Y(_4783_)
);

AOI22X1 _14232_ (
    .A(_3870__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [18]),
    .C(_3902__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_4784_)
);

NAND3X1 _14233_ (
    .A(_4783_),
    .B(_4784_),
    .C(_4780_),
    .Y(_4785_)
);

NOR2X1 _14234_ (
    .A(_4773_),
    .B(_4785_),
    .Y(_4786_)
);

AOI22X1 _14235_ (
    .A(_3904__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [18]),
    .C(\datapath_1.regfile_1.regOut[22] [18]),
    .D(_4038_),
    .Y(_4787_)
);

AOI22X1 _14236_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [18]),
    .C(_3950__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_4788_)
);

INVX1 _14237_ (
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_4789_)
);

INVX1 _14238_ (
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_4790_)
);

OAI22X1 _14239_ (
    .A(_4789_),
    .B(_3934__bF$buf0),
    .C(_3886__bF$buf2),
    .D(_4790_),
    .Y(_4791_)
);

INVX1 _14240_ (
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_4792_)
);

INVX1 _14241_ (
    .A(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_4793_)
);

OAI22X1 _14242_ (
    .A(_3910__bF$buf1),
    .B(_4792_),
    .C(_4793_),
    .D(_3940__bF$buf0),
    .Y(_4794_)
);

NOR2X1 _14243_ (
    .A(_4794_),
    .B(_4791_),
    .Y(_4795_)
);

NAND3X1 _14244_ (
    .A(_4788_),
    .B(_4787_),
    .C(_4795_),
    .Y(_4796_)
);

INVX1 _14245_ (
    .A(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_4797_)
);

INVX1 _14246_ (
    .A(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_4798_)
);

OAI22X1 _14247_ (
    .A(_3939__bF$buf1),
    .B(_4798_),
    .C(_4797_),
    .D(_3924__bF$buf2),
    .Y(_4799_)
);

INVX1 _14248_ (
    .A(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_4800_)
);

INVX1 _14249_ (
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_4801_)
);

OAI22X1 _14250_ (
    .A(_3923__bF$buf1),
    .B(_4801_),
    .C(_4800_),
    .D(_3946_),
    .Y(_4802_)
);

NOR2X1 _14251_ (
    .A(_4802_),
    .B(_4799_),
    .Y(_4803_)
);

AOI22X1 _14252_ (
    .A(_4062__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [18]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_4804_)
);

AOI22X1 _14253_ (
    .A(_3952__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [18]),
    .C(\datapath_1.regfile_1.regOut[28] [18]),
    .D(_3879__bF$buf1),
    .Y(_4805_)
);

NAND3X1 _14254_ (
    .A(_4804_),
    .B(_4805_),
    .C(_4803_),
    .Y(_4806_)
);

NOR2X1 _14255_ (
    .A(_4806_),
    .B(_4796_),
    .Y(_4807_)
);

AOI21X1 _14256_ (
    .A(_4807_),
    .B(_4786_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [18])
);

AOI22X1 _14257_ (
    .A(_3866__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [19]),
    .C(\datapath_1.regfile_1.regOut[31] [19]),
    .D(_3906__bF$buf2),
    .Y(_4808_)
);

AOI22X1 _14258_ (
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[27] [19]),
    .D(_3947__bF$buf1),
    .Y(_4809_)
);

INVX1 _14259_ (
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_4810_)
);

INVX1 _14260_ (
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_4811_)
);

OAI22X1 _14261_ (
    .A(_3875__bF$buf2),
    .B(_4811_),
    .C(_4810_),
    .D(_3935__bF$buf3),
    .Y(_4812_)
);

INVX1 _14262_ (
    .A(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_4813_)
);

INVX1 _14263_ (
    .A(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_4814_)
);

OAI22X1 _14264_ (
    .A(_3911_),
    .B(_4813_),
    .C(_4814_),
    .D(_3940__bF$buf3),
    .Y(_4815_)
);

NOR2X1 _14265_ (
    .A(_4815_),
    .B(_4812_),
    .Y(_4816_)
);

NAND3X1 _14266_ (
    .A(_4809_),
    .B(_4808_),
    .C(_4816_),
    .Y(_4817_)
);

INVX1 _14267_ (
    .A(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_4818_)
);

INVX1 _14268_ (
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_4819_)
);

OAI22X1 _14269_ (
    .A(_3923__bF$buf0),
    .B(_4819_),
    .C(_4818_),
    .D(_3957__bF$buf4),
    .Y(_4820_)
);

INVX1 _14270_ (
    .A(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_4821_)
);

INVX1 _14271_ (
    .A(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_4822_)
);

OAI22X1 _14272_ (
    .A(_3929__bF$buf0),
    .B(_4821_),
    .C(_4822_),
    .D(_3956__bF$buf0),
    .Y(_4823_)
);

NOR2X1 _14273_ (
    .A(_4820_),
    .B(_4823_),
    .Y(_4824_)
);

INVX1 _14274_ (
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_4825_)
);

INVX1 _14275_ (
    .A(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_4826_)
);

OAI22X1 _14276_ (
    .A(_3889__bF$buf0),
    .B(_4825_),
    .C(_4826_),
    .D(_3939__bF$buf0),
    .Y(_4827_)
);

INVX1 _14277_ (
    .A(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_4828_)
);

INVX1 _14278_ (
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_4829_)
);

OAI22X1 _14279_ (
    .A(_3924__bF$buf1),
    .B(_4828_),
    .C(_4829_),
    .D(_4340_),
    .Y(_4830_)
);

NOR2X1 _14280_ (
    .A(_4827_),
    .B(_4830_),
    .Y(_4831_)
);

NAND2X1 _14281_ (
    .A(_4824_),
    .B(_4831_),
    .Y(_4832_)
);

NOR2X1 _14282_ (
    .A(_4817_),
    .B(_4832_),
    .Y(_4833_)
);

INVX1 _14283_ (
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_4834_)
);

INVX1 _14284_ (
    .A(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_4835_)
);

OAI22X1 _14285_ (
    .A(_4835_),
    .B(_3949_),
    .C(_3886__bF$buf1),
    .D(_4834_),
    .Y(_4836_)
);

INVX1 _14286_ (
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_4837_)
);

INVX1 _14287_ (
    .A(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_4838_)
);

OAI22X1 _14288_ (
    .A(_3916__bF$buf0),
    .B(_4837_),
    .C(_4838_),
    .D(_3915__bF$buf1),
    .Y(_4839_)
);

NOR2X1 _14289_ (
    .A(_4839_),
    .B(_4836_),
    .Y(_4840_)
);

AOI22X1 _14290_ (
    .A(_3952__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [19]),
    .C(\datapath_1.regfile_1.regOut[24] [19]),
    .D(_3902__bF$buf2),
    .Y(_4841_)
);

AOI22X1 _14291_ (
    .A(_3899__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .C(\datapath_1.regfile_1.regOut[28] [19]),
    .D(_3879__bF$buf0),
    .Y(_4842_)
);

NAND3X1 _14292_ (
    .A(_4841_),
    .B(_4842_),
    .C(_4840_),
    .Y(_4843_)
);

AOI22X1 _14293_ (
    .A(_4060__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[7] [19]),
    .C(\datapath_1.regfile_1.regOut[6] [19]),
    .D(_4068__bF$buf1),
    .Y(_4844_)
);

AOI22X1 _14294_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [19]),
    .C(\datapath_1.regfile_1.regOut[21] [19]),
    .D(_3990_),
    .Y(_4845_)
);

INVX1 _14295_ (
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_4846_)
);

INVX1 _14296_ (
    .A(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_4847_)
);

OAI22X1 _14297_ (
    .A(_3869_),
    .B(_4846_),
    .C(_4847_),
    .D(_3944__bF$buf2),
    .Y(_4848_)
);

INVX1 _14298_ (
    .A(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_4849_)
);

INVX1 _14299_ (
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_4850_)
);

OAI22X1 _14300_ (
    .A(_3894__bF$buf0),
    .B(_4850_),
    .C(_4849_),
    .D(_3961__bF$buf0),
    .Y(_4851_)
);

NOR2X1 _14301_ (
    .A(_4851_),
    .B(_4848_),
    .Y(_4852_)
);

NAND3X1 _14302_ (
    .A(_4845_),
    .B(_4844_),
    .C(_4852_),
    .Y(_4853_)
);

NOR2X1 _14303_ (
    .A(_4853_),
    .B(_4843_),
    .Y(_4854_)
);

AOI21X1 _14304_ (
    .A(_4833_),
    .B(_4854_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [19])
);

INVX1 _14305_ (
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_4855_)
);

NOR2X1 _14306_ (
    .A(_4855_),
    .B(_3961__bF$buf4),
    .Y(_4856_)
);

AOI21X1 _14307_ (
    .A(\datapath_1.regfile_1.regOut[13] [20]),
    .B(_4099_),
    .C(_4856_),
    .Y(_4857_)
);

AOI22X1 _14308_ (
    .A(_4068__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [20]),
    .C(\datapath_1.regfile_1.regOut[31] [20]),
    .D(_3906__bF$buf1),
    .Y(_4858_)
);

INVX1 _14309_ (
    .A(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_4859_)
);

INVX1 _14310_ (
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_4860_)
);

OAI22X1 _14311_ (
    .A(_4860_),
    .B(_3916__bF$buf4),
    .C(_3889__bF$buf4),
    .D(_4859_),
    .Y(_4861_)
);

INVX1 _14312_ (
    .A(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_4862_)
);

INVX1 _14313_ (
    .A(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_4863_)
);

OAI22X1 _14314_ (
    .A(_4863_),
    .B(_3928_),
    .C(_4862_),
    .D(_3915__bF$buf0),
    .Y(_4864_)
);

NOR2X1 _14315_ (
    .A(_4861_),
    .B(_4864_),
    .Y(_4865_)
);

NAND3X1 _14316_ (
    .A(_4858_),
    .B(_4857_),
    .C(_4865_),
    .Y(_4866_)
);

INVX1 _14317_ (
    .A(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_4867_)
);

INVX1 _14318_ (
    .A(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_4868_)
);

OAI22X1 _14319_ (
    .A(_4868_),
    .B(_3929__bF$buf4),
    .C(_3946_),
    .D(_4867_),
    .Y(_4869_)
);

INVX1 _14320_ (
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_4870_)
);

INVX1 _14321_ (
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_4871_)
);

OAI22X1 _14322_ (
    .A(_4871_),
    .B(_3894__bF$buf4),
    .C(_4870_),
    .D(_3869_),
    .Y(_4872_)
);

NOR2X1 _14323_ (
    .A(_4872_),
    .B(_4869_),
    .Y(_4873_)
);

INVX1 _14324_ (
    .A(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_4874_)
);

NOR2X1 _14325_ (
    .A(_4874_),
    .B(_3956__bF$buf4),
    .Y(_4875_)
);

AOI21X1 _14326_ (
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .B(_3899__bF$buf3),
    .C(_4875_),
    .Y(_4876_)
);

AOI22X1 _14327_ (
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[24] [20]),
    .D(_3902__bF$buf1),
    .Y(_4877_)
);

NAND3X1 _14328_ (
    .A(_4876_),
    .B(_4877_),
    .C(_4873_),
    .Y(_4878_)
);

NOR2X1 _14329_ (
    .A(_4866_),
    .B(_4878_),
    .Y(_4879_)
);

AOI22X1 _14330_ (
    .A(_3904__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[20] [20]),
    .C(\datapath_1.regfile_1.regOut[22] [20]),
    .D(_4038_),
    .Y(_4880_)
);

AOI22X1 _14331_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [20]),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_4881_)
);

INVX1 _14332_ (
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_4882_)
);

INVX1 _14333_ (
    .A(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_4883_)
);

OAI22X1 _14334_ (
    .A(_4882_),
    .B(_3934__bF$buf3),
    .C(_3886__bF$buf0),
    .D(_4883_),
    .Y(_4884_)
);

INVX1 _14335_ (
    .A(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_4885_)
);

INVX1 _14336_ (
    .A(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_4886_)
);

OAI22X1 _14337_ (
    .A(_4886_),
    .B(_3940__bF$buf2),
    .C(_4885_),
    .D(_3924__bF$buf0),
    .Y(_4887_)
);

NOR2X1 _14338_ (
    .A(_4887_),
    .B(_4884_),
    .Y(_4888_)
);

NAND3X1 _14339_ (
    .A(_4881_),
    .B(_4880_),
    .C(_4888_),
    .Y(_4889_)
);

INVX1 _14340_ (
    .A(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_4890_)
);

INVX1 _14341_ (
    .A(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_4891_)
);

OAI22X1 _14342_ (
    .A(_4044_),
    .B(_4890_),
    .C(_4891_),
    .D(_3939__bF$buf4),
    .Y(_4892_)
);

INVX1 _14343_ (
    .A(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_4893_)
);

INVX1 _14344_ (
    .A(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_4894_)
);

OAI22X1 _14345_ (
    .A(_3923__bF$buf4),
    .B(_4894_),
    .C(_4893_),
    .D(_3944__bF$buf1),
    .Y(_4895_)
);

NOR2X1 _14346_ (
    .A(_4892_),
    .B(_4895_),
    .Y(_4896_)
);

AOI22X1 _14347_ (
    .A(_4062__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [20]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_4897_)
);

AOI22X1 _14348_ (
    .A(_3952__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [20]),
    .C(\datapath_1.regfile_1.regOut[29] [20]),
    .D(_3866__bF$buf0),
    .Y(_4898_)
);

NAND3X1 _14349_ (
    .A(_4897_),
    .B(_4898_),
    .C(_4896_),
    .Y(_4899_)
);

NOR2X1 _14350_ (
    .A(_4899_),
    .B(_4889_),
    .Y(_4900_)
);

AOI21X1 _14351_ (
    .A(_4900_),
    .B(_4879_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [20])
);

INVX1 _14352_ (
    .A(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_4901_)
);

INVX1 _14353_ (
    .A(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_4902_)
);

OAI22X1 _14354_ (
    .A(_4902_),
    .B(_3957__bF$buf3),
    .C(_3961__bF$buf3),
    .D(_4901_),
    .Y(_4903_)
);

INVX1 _14355_ (
    .A(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_4904_)
);

INVX1 _14356_ (
    .A(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_4905_)
);

OAI22X1 _14357_ (
    .A(_3865_),
    .B(_4904_),
    .C(_4905_),
    .D(_3893_),
    .Y(_4906_)
);

NOR2X1 _14358_ (
    .A(_4903_),
    .B(_4906_),
    .Y(_4907_)
);

INVX1 _14359_ (
    .A(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_4908_)
);

NOR2X1 _14360_ (
    .A(_4908_),
    .B(_3923__bF$buf3),
    .Y(_4909_)
);

AOI21X1 _14361_ (
    .A(_3987_),
    .B(\datapath_1.regfile_1.regOut[0] [21]),
    .C(_4909_),
    .Y(_4910_)
);

AOI22X1 _14362_ (
    .A(_4060__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[7] [21]),
    .C(\datapath_1.regfile_1.regOut[30] [21]),
    .D(_3870__bF$buf1),
    .Y(_4911_)
);

NAND3X1 _14363_ (
    .A(_4910_),
    .B(_4911_),
    .C(_4907_),
    .Y(_4912_)
);

INVX1 _14364_ (
    .A(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_4913_)
);

INVX1 _14365_ (
    .A(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_4914_)
);

OAI22X1 _14366_ (
    .A(_3929__bF$buf3),
    .B(_4914_),
    .C(_4913_),
    .D(_3944__bF$buf0),
    .Y(_4915_)
);

INVX1 _14367_ (
    .A(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_4916_)
);

INVX1 _14368_ (
    .A(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_4917_)
);

OAI22X1 _14369_ (
    .A(_3894__bF$buf3),
    .B(_4917_),
    .C(_4916_),
    .D(_3924__bF$buf3),
    .Y(_4918_)
);

NOR2X1 _14370_ (
    .A(_4918_),
    .B(_4915_),
    .Y(_4919_)
);

INVX1 _14371_ (
    .A(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_4920_)
);

NOR2X1 _14372_ (
    .A(_4920_),
    .B(_3956__bF$buf3),
    .Y(_4921_)
);

AOI21X1 _14373_ (
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .B(_3899__bF$buf2),
    .C(_4921_),
    .Y(_4922_)
);

AOI22X1 _14374_ (
    .A(_3879__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [21]),
    .C(_3902__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_4923_)
);

NAND3X1 _14375_ (
    .A(_4922_),
    .B(_4923_),
    .C(_4919_),
    .Y(_4924_)
);

NOR2X1 _14376_ (
    .A(_4912_),
    .B(_4924_),
    .Y(_4925_)
);

AOI22X1 _14377_ (
    .A(_3876_),
    .B(\datapath_1.regfile_1.regOut[4] [21]),
    .C(\datapath_1.regfile_1.regOut[2] [21]),
    .D(_3975_),
    .Y(_4926_)
);

AOI22X1 _14378_ (
    .A(_4062__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [21]),
    .C(\datapath_1.regfile_1.regOut[17] [21]),
    .D(_4135_),
    .Y(_4927_)
);

INVX1 _14379_ (
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_4928_)
);

INVX1 _14380_ (
    .A(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_4929_)
);

OAI22X1 _14381_ (
    .A(_4929_),
    .B(_3939__bF$buf3),
    .C(_4928_),
    .D(_3905_),
    .Y(_4930_)
);

INVX1 _14382_ (
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_4931_)
);

INVX1 _14383_ (
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_4932_)
);

OAI22X1 _14384_ (
    .A(_4932_),
    .B(_3916__bF$buf3),
    .C(_3889__bF$buf3),
    .D(_4931_),
    .Y(_4933_)
);

NOR2X1 _14385_ (
    .A(_4933_),
    .B(_4930_),
    .Y(_4934_)
);

NAND3X1 _14386_ (
    .A(_4927_),
    .B(_4926_),
    .C(_4934_),
    .Y(_4935_)
);

AOI22X1 _14387_ (
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[9] [21]),
    .D(_3950__bF$buf3),
    .Y(_4936_)
);

AOI22X1 _14388_ (
    .A(_3904__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[20] [21]),
    .C(\datapath_1.regfile_1.regOut[10] [21]),
    .D(_4087_),
    .Y(_4937_)
);

INVX1 _14389_ (
    .A(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_4938_)
);

INVX1 _14390_ (
    .A(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_4939_)
);

OAI22X1 _14391_ (
    .A(_4939_),
    .B(_3934__bF$buf2),
    .C(_3935__bF$buf2),
    .D(_4938_),
    .Y(_4940_)
);

INVX1 _14392_ (
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_4941_)
);

INVX1 _14393_ (
    .A(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_4942_)
);

OAI22X1 _14394_ (
    .A(_4942_),
    .B(_3951_),
    .C(_3946_),
    .D(_4941_),
    .Y(_4943_)
);

NOR2X1 _14395_ (
    .A(_4943_),
    .B(_4940_),
    .Y(_4944_)
);

NAND3X1 _14396_ (
    .A(_4937_),
    .B(_4936_),
    .C(_4944_),
    .Y(_4945_)
);

NOR2X1 _14397_ (
    .A(_4935_),
    .B(_4945_),
    .Y(_4946_)
);

AOI21X1 _14398_ (
    .A(_4925_),
    .B(_4946_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [21])
);

INVX1 _14399_ (
    .A(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_4947_)
);

INVX1 _14400_ (
    .A(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_4948_)
);

OAI22X1 _14401_ (
    .A(_4948_),
    .B(_3928_),
    .C(_4947_),
    .D(_3893_),
    .Y(_4949_)
);

INVX1 _14402_ (
    .A(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_4950_)
);

INVX1 _14403_ (
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_4951_)
);

OAI22X1 _14404_ (
    .A(_3869_),
    .B(_4950_),
    .C(_4951_),
    .D(_3935__bF$buf1),
    .Y(_4952_)
);

NOR2X1 _14405_ (
    .A(_4949_),
    .B(_4952_),
    .Y(_4953_)
);

AOI22X1 _14406_ (
    .A(_3902__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[24] [22]),
    .C(\datapath_1.regfile_1.regOut[26] [22]),
    .D(_4070_),
    .Y(_4954_)
);

AOI22X1 _14407_ (
    .A(_3952__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [22]),
    .C(\datapath_1.regfile_1.regOut[29] [22]),
    .D(_3866__bF$buf3),
    .Y(_4955_)
);

NAND3X1 _14408_ (
    .A(_4954_),
    .B(_4955_),
    .C(_4953_),
    .Y(_4956_)
);

INVX1 _14409_ (
    .A(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_4957_)
);

INVX1 _14410_ (
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_4958_)
);

OAI22X1 _14411_ (
    .A(_4958_),
    .B(_3916__bF$buf2),
    .C(_4957_),
    .D(_3910__bF$buf0),
    .Y(_4959_)
);

INVX1 _14412_ (
    .A(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_4960_)
);

INVX1 _14413_ (
    .A(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_4961_)
);

OAI22X1 _14414_ (
    .A(_3889__bF$buf2),
    .B(_4960_),
    .C(_4961_),
    .D(_3956__bF$buf2),
    .Y(_4962_)
);

NOR2X1 _14415_ (
    .A(_4959_),
    .B(_4962_),
    .Y(_4963_)
);

AOI22X1 _14416_ (
    .A(_4087_),
    .B(\datapath_1.regfile_1.regOut[10] [22]),
    .C(\datapath_1.regfile_1.regOut[31] [22]),
    .D(_3906__bF$buf0),
    .Y(_4964_)
);

AOI22X1 _14417_ (
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[21] [22]),
    .D(_3990_),
    .Y(_4965_)
);

NAND3X1 _14418_ (
    .A(_4964_),
    .B(_4965_),
    .C(_4963_),
    .Y(_4966_)
);

NOR2X1 _14419_ (
    .A(_4966_),
    .B(_4956_),
    .Y(_4967_)
);

AOI22X1 _14420_ (
    .A(_3947__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [22]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_4968_)
);

AOI22X1 _14421_ (
    .A(_4062__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [22]),
    .C(\datapath_1.regfile_1.regOut[28] [22]),
    .D(_3879__bF$buf2),
    .Y(_4969_)
);

INVX1 _14422_ (
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_4970_)
);

INVX1 _14423_ (
    .A(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_4971_)
);

OAI22X1 _14424_ (
    .A(_4971_),
    .B(_3962__bF$buf1),
    .C(_3898_),
    .D(_4970_),
    .Y(_4972_)
);

INVX1 _14425_ (
    .A(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_4973_)
);

INVX1 _14426_ (
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_4974_)
);

OAI22X1 _14427_ (
    .A(_3923__bF$buf2),
    .B(_4974_),
    .C(_4973_),
    .D(_3929__bF$buf2),
    .Y(_4975_)
);

NOR2X1 _14428_ (
    .A(_4975_),
    .B(_4972_),
    .Y(_4976_)
);

NAND3X1 _14429_ (
    .A(_4969_),
    .B(_4968_),
    .C(_4976_),
    .Y(_4977_)
);

INVX1 _14430_ (
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_4978_)
);

INVX1 _14431_ (
    .A(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_4979_)
);

OAI22X1 _14432_ (
    .A(_3875__bF$buf1),
    .B(_4978_),
    .C(_4979_),
    .D(_3940__bF$buf1),
    .Y(_4980_)
);

INVX1 _14433_ (
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_4981_)
);

INVX1 _14434_ (
    .A(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_4982_)
);

OAI22X1 _14435_ (
    .A(_4981_),
    .B(_3894__bF$buf2),
    .C(_4982_),
    .D(_3939__bF$buf2),
    .Y(_4983_)
);

NOR2X1 _14436_ (
    .A(_4983_),
    .B(_4980_),
    .Y(_4984_)
);

INVX1 _14437_ (
    .A(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_4985_)
);

INVX1 _14438_ (
    .A(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_4986_)
);

OAI22X1 _14439_ (
    .A(_4986_),
    .B(_3957__bF$buf2),
    .C(_3961__bF$buf2),
    .D(_4985_),
    .Y(_4987_)
);

INVX1 _14440_ (
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_4988_)
);

INVX1 _14441_ (
    .A(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_4989_)
);

OAI22X1 _14442_ (
    .A(_4989_),
    .B(_3949_),
    .C(_4988_),
    .D(_4340_),
    .Y(_4990_)
);

NOR2X1 _14443_ (
    .A(_4987_),
    .B(_4990_),
    .Y(_4991_)
);

NAND2X1 _14444_ (
    .A(_4984_),
    .B(_4991_),
    .Y(_4992_)
);

NOR2X1 _14445_ (
    .A(_4977_),
    .B(_4992_),
    .Y(_4993_)
);

AOI21X1 _14446_ (
    .A(_4993_),
    .B(_4967_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [22])
);

AOI22X1 _14447_ (
    .A(_3952__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [23]),
    .C(\datapath_1.regfile_1.regOut[24] [23]),
    .D(_3902__bF$buf3),
    .Y(_4994_)
);

INVX1 _14448_ (
    .A(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_4995_)
);

NOR2X1 _14449_ (
    .A(_4995_),
    .B(_3939__bF$buf1),
    .Y(_4996_)
);

AOI21X1 _14450_ (
    .A(_3870__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [23]),
    .C(_4996_),
    .Y(_4997_)
);

INVX1 _14451_ (
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_4998_)
);

INVX1 _14452_ (
    .A(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_4999_)
);

OAI22X1 _14453_ (
    .A(_4998_),
    .B(_3894__bF$buf1),
    .C(_4999_),
    .D(_3929__bF$buf1),
    .Y(_5000_)
);

INVX1 _14454_ (
    .A(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_5001_)
);

INVX1 _14455_ (
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_5002_)
);

OAI22X1 _14456_ (
    .A(_5002_),
    .B(_3916__bF$buf1),
    .C(_3889__bF$buf1),
    .D(_5001_),
    .Y(_5003_)
);

NOR2X1 _14457_ (
    .A(_5003_),
    .B(_5000_),
    .Y(_5004_)
);

NAND3X1 _14458_ (
    .A(_4994_),
    .B(_4997_),
    .C(_5004_),
    .Y(_5005_)
);

AOI22X1 _14459_ (
    .A(_3947__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [23]),
    .C(_3904__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_5006_)
);

AOI22X1 _14460_ (
    .A(_3899__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [23]),
    .C(\datapath_1.regfile_1.regOut[25] [23]),
    .D(_3945_),
    .Y(_5007_)
);

INVX1 _14461_ (
    .A(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_5008_)
);

INVX1 _14462_ (
    .A(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_5009_)
);

OAI22X1 _14463_ (
    .A(_5008_),
    .B(_3910__bF$buf3),
    .C(_5009_),
    .D(_3911_),
    .Y(_5010_)
);

INVX1 _14464_ (
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_5011_)
);

INVX1 _14465_ (
    .A(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_5012_)
);

OAI22X1 _14466_ (
    .A(_5012_),
    .B(_3915__bF$buf3),
    .C(_3886__bF$buf3),
    .D(_5011_),
    .Y(_5013_)
);

NOR2X1 _14467_ (
    .A(_5010_),
    .B(_5013_),
    .Y(_5014_)
);

NAND3X1 _14468_ (
    .A(_5007_),
    .B(_5006_),
    .C(_5014_),
    .Y(_5015_)
);

NOR2X1 _14469_ (
    .A(_5005_),
    .B(_5015_),
    .Y(_5016_)
);

AOI22X1 _14470_ (
    .A(_4060__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[7] [23]),
    .C(\datapath_1.regfile_1.regOut[6] [23]),
    .D(_4068__bF$buf3),
    .Y(_5017_)
);

INVX1 _14471_ (
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_5018_)
);

NOR2X1 _14472_ (
    .A(_5018_),
    .B(_3923__bF$buf1),
    .Y(_5019_)
);

AOI21X1 _14473_ (
    .A(_3906__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[31] [23]),
    .C(_5019_),
    .Y(_5020_)
);

INVX1 _14474_ (
    .A(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_5021_)
);

INVX1 _14475_ (
    .A(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_5022_)
);

OAI22X1 _14476_ (
    .A(_5022_),
    .B(_3934__bF$buf1),
    .C(_3935__bF$buf0),
    .D(_5021_),
    .Y(_5023_)
);

INVX1 _14477_ (
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_5024_)
);

INVX1 _14478_ (
    .A(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_5025_)
);

OAI22X1 _14479_ (
    .A(_3875__bF$buf0),
    .B(_5024_),
    .C(_5025_),
    .D(_3940__bF$buf0),
    .Y(_5026_)
);

NOR2X1 _14480_ (
    .A(_5026_),
    .B(_5023_),
    .Y(_5027_)
);

NAND3X1 _14481_ (
    .A(_5020_),
    .B(_5017_),
    .C(_5027_),
    .Y(_5028_)
);

AOI22X1 _14482_ (
    .A(_3879__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[28] [23]),
    .C(_4070_),
    .D(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_5029_)
);

AOI22X1 _14483_ (
    .A(_3866__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [23]),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_5030_)
);

INVX1 _14484_ (
    .A(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_5031_)
);

INVX1 _14485_ (
    .A(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_5032_)
);

OAI22X1 _14486_ (
    .A(_3957__bF$buf1),
    .B(_5031_),
    .C(_5032_),
    .D(_3956__bF$buf1),
    .Y(_5033_)
);

INVX1 _14487_ (
    .A(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_5034_)
);

INVX1 _14488_ (
    .A(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_5035_)
);

OAI22X1 _14489_ (
    .A(_5035_),
    .B(_3961__bF$buf1),
    .C(_3962__bF$buf0),
    .D(_5034_),
    .Y(_5036_)
);

NOR2X1 _14490_ (
    .A(_5036_),
    .B(_5033_),
    .Y(_5037_)
);

NAND3X1 _14491_ (
    .A(_5030_),
    .B(_5029_),
    .C(_5037_),
    .Y(_5038_)
);

NOR2X1 _14492_ (
    .A(_5028_),
    .B(_5038_),
    .Y(_5039_)
);

AOI21X1 _14493_ (
    .A(_5039_),
    .B(_5016_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [23])
);

INVX1 _14494_ (
    .A(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_5040_)
);

INVX1 _14495_ (
    .A(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_5041_)
);

OAI22X1 _14496_ (
    .A(_5041_),
    .B(_3865_),
    .C(_3869_),
    .D(_5040_),
    .Y(_5042_)
);

INVX1 _14497_ (
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_5043_)
);

INVX1 _14498_ (
    .A(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_5044_)
);

OAI22X1 _14499_ (
    .A(_3916__bF$buf0),
    .B(_5043_),
    .C(_5044_),
    .D(_3915__bF$buf2),
    .Y(_5045_)
);

NOR2X1 _14500_ (
    .A(_5042_),
    .B(_5045_),
    .Y(_5046_)
);

INVX1 _14501_ (
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_5047_)
);

INVX1 _14502_ (
    .A(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_5048_)
);

OAI22X1 _14503_ (
    .A(_5047_),
    .B(_3894__bF$buf0),
    .C(_5048_),
    .D(_3929__bF$buf0),
    .Y(_5049_)
);

INVX1 _14504_ (
    .A(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_5050_)
);

INVX1 _14505_ (
    .A(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_5051_)
);

OAI22X1 _14506_ (
    .A(_5051_),
    .B(_3940__bF$buf3),
    .C(_3939__bF$buf0),
    .D(_5050_),
    .Y(_5052_)
);

NOR2X1 _14507_ (
    .A(_5049_),
    .B(_5052_),
    .Y(_5053_)
);

NAND2X1 _14508_ (
    .A(_5053_),
    .B(_5046_),
    .Y(_5054_)
);

AOI22X1 _14509_ (
    .A(_3899__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [24]),
    .C(\datapath_1.regfile_1.regOut[24] [24]),
    .D(_3902__bF$buf2),
    .Y(_5055_)
);

INVX1 _14510_ (
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_5056_)
);

NOR2X1 _14511_ (
    .A(_5056_),
    .B(_3923__bF$buf0),
    .Y(_5057_)
);

AOI21X1 _14512_ (
    .A(_3906__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [24]),
    .C(_5057_),
    .Y(_5058_)
);

INVX1 _14513_ (
    .A(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_5059_)
);

INVX1 _14514_ (
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_5060_)
);

OAI22X1 _14515_ (
    .A(_5059_),
    .B(_3910__bF$buf2),
    .C(_5060_),
    .D(_4044_),
    .Y(_5061_)
);

INVX1 _14516_ (
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_5062_)
);

INVX1 _14517_ (
    .A(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_5063_)
);

OAI22X1 _14518_ (
    .A(_5062_),
    .B(_3934__bF$buf0),
    .C(_3886__bF$buf2),
    .D(_5063_),
    .Y(_5064_)
);

NOR2X1 _14519_ (
    .A(_5061_),
    .B(_5064_),
    .Y(_5065_)
);

NAND3X1 _14520_ (
    .A(_5058_),
    .B(_5055_),
    .C(_5065_),
    .Y(_5066_)
);

NOR2X1 _14521_ (
    .A(_5054_),
    .B(_5066_),
    .Y(_5067_)
);

AOI22X1 _14522_ (
    .A(_4060__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[7] [24]),
    .C(\datapath_1.regfile_1.regOut[6] [24]),
    .D(_4068__bF$buf2),
    .Y(_5068_)
);

AOI22X1 _14523_ (
    .A(_3904__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [24]),
    .C(\datapath_1.regfile_1.regOut[9] [24]),
    .D(_3950__bF$buf1),
    .Y(_5069_)
);

INVX1 _14524_ (
    .A(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_5070_)
);

INVX1 _14525_ (
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_5071_)
);

OAI22X1 _14526_ (
    .A(_5071_),
    .B(_3875__bF$buf3),
    .C(_3911_),
    .D(_5070_),
    .Y(_5072_)
);

INVX1 _14527_ (
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_5073_)
);

INVX1 _14528_ (
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_5074_)
);

OAI22X1 _14529_ (
    .A(_3889__bF$buf0),
    .B(_5074_),
    .C(_5073_),
    .D(_3935__bF$buf3),
    .Y(_5075_)
);

NOR2X1 _14530_ (
    .A(_5072_),
    .B(_5075_),
    .Y(_5076_)
);

NAND3X1 _14531_ (
    .A(_5069_),
    .B(_5068_),
    .C(_5076_),
    .Y(_5077_)
);

AOI22X1 _14532_ (
    .A(_3947__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [24]),
    .C(_3945_),
    .D(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_5078_)
);

AOI22X1 _14533_ (
    .A(_3952__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[18] [24]),
    .C(\datapath_1.regfile_1.regOut[26] [24]),
    .D(_4070_),
    .Y(_5079_)
);

INVX1 _14534_ (
    .A(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_5080_)
);

INVX1 _14535_ (
    .A(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_5081_)
);

OAI22X1 _14536_ (
    .A(_3957__bF$buf0),
    .B(_5080_),
    .C(_5081_),
    .D(_3956__bF$buf0),
    .Y(_5082_)
);

INVX1 _14537_ (
    .A(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_5083_)
);

INVX1 _14538_ (
    .A(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_5084_)
);

OAI22X1 _14539_ (
    .A(_5084_),
    .B(_3961__bF$buf0),
    .C(_3962__bF$buf3),
    .D(_5083_),
    .Y(_5085_)
);

NOR2X1 _14540_ (
    .A(_5085_),
    .B(_5082_),
    .Y(_5086_)
);

NAND3X1 _14541_ (
    .A(_5079_),
    .B(_5078_),
    .C(_5086_),
    .Y(_5087_)
);

NOR2X1 _14542_ (
    .A(_5077_),
    .B(_5087_),
    .Y(_5088_)
);

AOI21X1 _14543_ (
    .A(_5088_),
    .B(_5067_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [24])
);

INVX1 _14544_ (
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_5089_)
);

INVX1 _14545_ (
    .A(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_5090_)
);

OAI22X1 _14546_ (
    .A(_3875__bF$buf2),
    .B(_5089_),
    .C(_5090_),
    .D(_3940__bF$buf2),
    .Y(_5091_)
);

INVX1 _14547_ (
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_5092_)
);

INVX1 _14548_ (
    .A(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_5093_)
);

OAI22X1 _14549_ (
    .A(_4044_),
    .B(_5092_),
    .C(_5093_),
    .D(_3924__bF$buf2),
    .Y(_5094_)
);

NOR2X1 _14550_ (
    .A(_5091_),
    .B(_5094_),
    .Y(_5095_)
);

INVX1 _14551_ (
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_5096_)
);

INVX1 _14552_ (
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_5097_)
);

OAI22X1 _14553_ (
    .A(_5097_),
    .B(_3916__bF$buf4),
    .C(_3889__bF$buf4),
    .D(_5096_),
    .Y(_5098_)
);

INVX1 _14554_ (
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_5099_)
);

INVX1 _14555_ (
    .A(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_5100_)
);

OAI22X1 _14556_ (
    .A(_3946_),
    .B(_5099_),
    .C(_5100_),
    .D(_4332_),
    .Y(_5101_)
);

NOR2X1 _14557_ (
    .A(_5098_),
    .B(_5101_),
    .Y(_5102_)
);

NAND2X1 _14558_ (
    .A(_5095_),
    .B(_5102_),
    .Y(_5103_)
);

INVX1 _14559_ (
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_5104_)
);

INVX1 _14560_ (
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_5105_)
);

OAI22X1 _14561_ (
    .A(_3894__bF$buf4),
    .B(_5105_),
    .C(_5104_),
    .D(_4340_),
    .Y(_5106_)
);

INVX1 _14562_ (
    .A(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_5107_)
);

INVX1 _14563_ (
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_5108_)
);

OAI22X1 _14564_ (
    .A(_5108_),
    .B(_3923__bF$buf4),
    .C(_5107_),
    .D(_3939__bF$buf4),
    .Y(_5109_)
);

NOR2X1 _14565_ (
    .A(_5109_),
    .B(_5106_),
    .Y(_5110_)
);

INVX1 _14566_ (
    .A(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_5111_)
);

INVX1 _14567_ (
    .A(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_5112_)
);

OAI22X1 _14568_ (
    .A(_3911_),
    .B(_5112_),
    .C(_5111_),
    .D(_3944__bF$buf3),
    .Y(_5113_)
);

INVX1 _14569_ (
    .A(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_5114_)
);

INVX1 _14570_ (
    .A(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_5115_)
);

OAI22X1 _14571_ (
    .A(_5115_),
    .B(_3915__bF$buf1),
    .C(_3886__bF$buf1),
    .D(_5114_),
    .Y(_5116_)
);

NOR2X1 _14572_ (
    .A(_5113_),
    .B(_5116_),
    .Y(_5117_)
);

NAND2X1 _14573_ (
    .A(_5117_),
    .B(_5110_),
    .Y(_5118_)
);

NOR2X1 _14574_ (
    .A(_5118_),
    .B(_5103_),
    .Y(_5119_)
);

AOI22X1 _14575_ (
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[6] [25]),
    .D(_4068__bF$buf1),
    .Y(_5120_)
);

AOI22X1 _14576_ (
    .A(_3899__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [25]),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_5121_)
);

INVX1 _14577_ (
    .A(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_5122_)
);

INVX1 _14578_ (
    .A(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_5123_)
);

OAI22X1 _14579_ (
    .A(_5123_),
    .B(_3934__bF$buf3),
    .C(_3935__bF$buf2),
    .D(_5122_),
    .Y(_5124_)
);

INVX1 _14580_ (
    .A(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_5125_)
);

INVX1 _14581_ (
    .A(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_5126_)
);

OAI22X1 _14582_ (
    .A(_3928_),
    .B(_5125_),
    .C(_5126_),
    .D(_3956__bF$buf4),
    .Y(_5127_)
);

NOR2X1 _14583_ (
    .A(_5127_),
    .B(_5124_),
    .Y(_5128_)
);

NAND3X1 _14584_ (
    .A(_5121_),
    .B(_5120_),
    .C(_5128_),
    .Y(_5129_)
);

INVX1 _14585_ (
    .A(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_5130_)
);

INVX1 _14586_ (
    .A(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_5131_)
);

OAI22X1 _14587_ (
    .A(_5131_),
    .B(_3929__bF$buf4),
    .C(_3957__bF$buf4),
    .D(_5130_),
    .Y(_5132_)
);

INVX1 _14588_ (
    .A(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_5133_)
);

INVX1 _14589_ (
    .A(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_5134_)
);

OAI22X1 _14590_ (
    .A(_3961__bF$buf4),
    .B(_5133_),
    .C(_5134_),
    .D(_3949_),
    .Y(_5135_)
);

NOR2X1 _14591_ (
    .A(_5132_),
    .B(_5135_),
    .Y(_5136_)
);

AOI22X1 _14592_ (
    .A(_3866__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [25]),
    .C(\datapath_1.regfile_1.regOut[31] [25]),
    .D(_3906__bF$buf1),
    .Y(_5137_)
);

AOI22X1 _14593_ (
    .A(_3952__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [25]),
    .C(\datapath_1.regfile_1.regOut[30] [25]),
    .D(_3870__bF$buf3),
    .Y(_5138_)
);

NAND3X1 _14594_ (
    .A(_5137_),
    .B(_5138_),
    .C(_5136_),
    .Y(_5139_)
);

NOR2X1 _14595_ (
    .A(_5139_),
    .B(_5129_),
    .Y(_5140_)
);

AOI21X1 _14596_ (
    .A(_5119_),
    .B(_5140_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [25])
);

INVX1 _14597_ (
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_5141_)
);

NOR2X1 _14598_ (
    .A(_5141_),
    .B(_3961__bF$buf3),
    .Y(_5142_)
);

AOI21X1 _14599_ (
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .B(_4099_),
    .C(_5142_),
    .Y(_5143_)
);

AOI22X1 _14600_ (
    .A(_4068__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .C(\datapath_1.regfile_1.regOut[31] [26]),
    .D(_3906__bF$buf0),
    .Y(_5144_)
);

INVX1 _14601_ (
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_5145_)
);

INVX1 _14602_ (
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_5146_)
);

OAI22X1 _14603_ (
    .A(_5146_),
    .B(_3916__bF$buf3),
    .C(_3889__bF$buf3),
    .D(_5145_),
    .Y(_5147_)
);

INVX1 _14604_ (
    .A(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_5148_)
);

INVX1 _14605_ (
    .A(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_5149_)
);

OAI22X1 _14606_ (
    .A(_5149_),
    .B(_3928_),
    .C(_5148_),
    .D(_3915__bF$buf0),
    .Y(_5150_)
);

NOR2X1 _14607_ (
    .A(_5147_),
    .B(_5150_),
    .Y(_5151_)
);

NAND3X1 _14608_ (
    .A(_5144_),
    .B(_5143_),
    .C(_5151_),
    .Y(_5152_)
);

INVX1 _14609_ (
    .A(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_5153_)
);

INVX1 _14610_ (
    .A(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_5154_)
);

OAI22X1 _14611_ (
    .A(_5154_),
    .B(_3929__bF$buf3),
    .C(_3946_),
    .D(_5153_),
    .Y(_5155_)
);

INVX1 _14612_ (
    .A(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_5156_)
);

INVX1 _14613_ (
    .A(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_5157_)
);

OAI22X1 _14614_ (
    .A(_5157_),
    .B(_3894__bF$buf3),
    .C(_5156_),
    .D(_3869_),
    .Y(_5158_)
);

NOR2X1 _14615_ (
    .A(_5158_),
    .B(_5155_),
    .Y(_5159_)
);

INVX1 _14616_ (
    .A(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_5160_)
);

NOR2X1 _14617_ (
    .A(_5160_),
    .B(_3956__bF$buf3),
    .Y(_5161_)
);

AOI21X1 _14618_ (
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .B(_3899__bF$buf3),
    .C(_5161_),
    .Y(_5162_)
);

AOI22X1 _14619_ (
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[24] [26]),
    .D(_3902__bF$buf1),
    .Y(_5163_)
);

NAND3X1 _14620_ (
    .A(_5162_),
    .B(_5163_),
    .C(_5159_),
    .Y(_5164_)
);

NOR2X1 _14621_ (
    .A(_5152_),
    .B(_5164_),
    .Y(_5165_)
);

AOI22X1 _14622_ (
    .A(_3904__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[20] [26]),
    .C(\datapath_1.regfile_1.regOut[21] [26]),
    .D(_3990_),
    .Y(_5166_)
);

AOI22X1 _14623_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [26]),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_5167_)
);

INVX1 _14624_ (
    .A(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_5168_)
);

INVX1 _14625_ (
    .A(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_5169_)
);

OAI22X1 _14626_ (
    .A(_5168_),
    .B(_3935__bF$buf1),
    .C(_3886__bF$buf0),
    .D(_5169_),
    .Y(_5170_)
);

INVX1 _14627_ (
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_5171_)
);

INVX1 _14628_ (
    .A(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_5172_)
);

OAI22X1 _14629_ (
    .A(_5172_),
    .B(_3940__bF$buf1),
    .C(_3939__bF$buf3),
    .D(_5171_),
    .Y(_5173_)
);

NOR2X1 _14630_ (
    .A(_5173_),
    .B(_5170_),
    .Y(_5174_)
);

NAND3X1 _14631_ (
    .A(_5167_),
    .B(_5166_),
    .C(_5174_),
    .Y(_5175_)
);

INVX1 _14632_ (
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_5176_)
);

INVX1 _14633_ (
    .A(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_5177_)
);

OAI22X1 _14634_ (
    .A(_4044_),
    .B(_5176_),
    .C(_5177_),
    .D(_3924__bF$buf1),
    .Y(_5178_)
);

INVX1 _14635_ (
    .A(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_5179_)
);

INVX1 _14636_ (
    .A(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_5180_)
);

OAI22X1 _14637_ (
    .A(_3923__bF$buf3),
    .B(_5180_),
    .C(_5179_),
    .D(_3944__bF$buf2),
    .Y(_5181_)
);

NOR2X1 _14638_ (
    .A(_5181_),
    .B(_5178_),
    .Y(_5182_)
);

AOI22X1 _14639_ (
    .A(_4062__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[8] [26]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_5183_)
);

AOI22X1 _14640_ (
    .A(_3952__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[18] [26]),
    .C(\datapath_1.regfile_1.regOut[29] [26]),
    .D(_3866__bF$buf0),
    .Y(_5184_)
);

NAND3X1 _14641_ (
    .A(_5183_),
    .B(_5184_),
    .C(_5182_),
    .Y(_5185_)
);

NOR2X1 _14642_ (
    .A(_5175_),
    .B(_5185_),
    .Y(_5186_)
);

AOI21X1 _14643_ (
    .A(_5186_),
    .B(_5165_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [26])
);

INVX1 _14644_ (
    .A(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_5187_)
);

INVX1 _14645_ (
    .A(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_5188_)
);

OAI22X1 _14646_ (
    .A(_3929__bF$buf2),
    .B(_5187_),
    .C(_5188_),
    .D(_3956__bF$buf2),
    .Y(_5189_)
);

INVX1 _14647_ (
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_5190_)
);

INVX1 _14648_ (
    .A(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_5191_)
);

OAI22X1 _14649_ (
    .A(_4044_),
    .B(_5190_),
    .C(_5191_),
    .D(_3957__bF$buf3),
    .Y(_5192_)
);

NOR2X1 _14650_ (
    .A(_5192_),
    .B(_5189_),
    .Y(_5193_)
);

INVX1 _14651_ (
    .A(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_5194_)
);

INVX1 _14652_ (
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_5195_)
);

OAI22X1 _14653_ (
    .A(_5195_),
    .B(_3916__bF$buf2),
    .C(_3889__bF$buf2),
    .D(_5194_),
    .Y(_5196_)
);

INVX1 _14654_ (
    .A(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_5197_)
);

INVX1 _14655_ (
    .A(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_5198_)
);

OAI22X1 _14656_ (
    .A(_3946_),
    .B(_5197_),
    .C(_5198_),
    .D(_3915__bF$buf3),
    .Y(_5199_)
);

NOR2X1 _14657_ (
    .A(_5196_),
    .B(_5199_),
    .Y(_5200_)
);

NAND2X1 _14658_ (
    .A(_5200_),
    .B(_5193_),
    .Y(_5201_)
);

AOI22X1 _14659_ (
    .A(_3899__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_5202_)
);

AOI22X1 _14660_ (
    .A(_3952__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[18] [27]),
    .C(\datapath_1.regfile_1.regOut[24] [27]),
    .D(_3902__bF$buf0),
    .Y(_5203_)
);

INVX1 _14661_ (
    .A(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_5204_)
);

INVX1 _14662_ (
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_5205_)
);

OAI22X1 _14663_ (
    .A(_3923__bF$buf2),
    .B(_5205_),
    .C(_5204_),
    .D(_3961__bF$buf2),
    .Y(_5206_)
);

INVX1 _14664_ (
    .A(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_5207_)
);

INVX1 _14665_ (
    .A(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_5208_)
);

OAI22X1 _14666_ (
    .A(_5208_),
    .B(_3939__bF$buf2),
    .C(_5207_),
    .D(_3865_),
    .Y(_5209_)
);

NOR2X1 _14667_ (
    .A(_5206_),
    .B(_5209_),
    .Y(_5210_)
);

NAND3X1 _14668_ (
    .A(_5203_),
    .B(_5202_),
    .C(_5210_),
    .Y(_5211_)
);

NOR2X1 _14669_ (
    .A(_5201_),
    .B(_5211_),
    .Y(_5212_)
);

AOI22X1 _14670_ (
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[22] [27]),
    .D(_4038_),
    .Y(_5213_)
);

AOI22X1 _14671_ (
    .A(_3870__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[30] [27]),
    .C(_3904__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_5214_)
);

INVX1 _14672_ (
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_5215_)
);

INVX1 _14673_ (
    .A(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_5216_)
);

OAI22X1 _14674_ (
    .A(_3875__bF$buf1),
    .B(_5215_),
    .C(_5216_),
    .D(_3940__bF$buf0),
    .Y(_5217_)
);

INVX1 _14675_ (
    .A(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_5218_)
);

INVX1 _14676_ (
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_5219_)
);

OAI22X1 _14677_ (
    .A(_3894__bF$buf2),
    .B(_5219_),
    .C(_5218_),
    .D(_3905_),
    .Y(_5220_)
);

NOR2X1 _14678_ (
    .A(_5217_),
    .B(_5220_),
    .Y(_5221_)
);

NAND3X1 _14679_ (
    .A(_5214_),
    .B(_5213_),
    .C(_5221_),
    .Y(_5222_)
);

INVX1 _14680_ (
    .A(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_5223_)
);

INVX1 _14681_ (
    .A(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_5224_)
);

OAI22X1 _14682_ (
    .A(_3910__bF$buf1),
    .B(_5223_),
    .C(_5224_),
    .D(_3944__bF$buf1),
    .Y(_5225_)
);

INVX1 _14683_ (
    .A(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_5226_)
);

INVX1 _14684_ (
    .A(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_5227_)
);

OAI22X1 _14685_ (
    .A(_5227_),
    .B(_3893_),
    .C(_3924__bF$buf0),
    .D(_5226_),
    .Y(_5228_)
);

NOR2X1 _14686_ (
    .A(_5225_),
    .B(_5228_),
    .Y(_5229_)
);

AOI22X1 _14687_ (
    .A(_4062__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[8] [27]),
    .C(\datapath_1.regfile_1.regOut[7] [27]),
    .D(_4060__bF$buf3),
    .Y(_5230_)
);

AOI22X1 _14688_ (
    .A(_3990_),
    .B(\datapath_1.regfile_1.regOut[21] [27]),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_5231_)
);

NAND3X1 _14689_ (
    .A(_5230_),
    .B(_5231_),
    .C(_5229_),
    .Y(_5232_)
);

NOR2X1 _14690_ (
    .A(_5222_),
    .B(_5232_),
    .Y(_5233_)
);

AOI21X1 _14691_ (
    .A(_5233_),
    .B(_5212_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [27])
);

INVX1 _14692_ (
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_5234_)
);

INVX1 _14693_ (
    .A(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_5235_)
);

OAI22X1 _14694_ (
    .A(_5234_),
    .B(_3894__bF$buf1),
    .C(_5235_),
    .D(_3940__bF$buf3),
    .Y(_5236_)
);

INVX1 _14695_ (
    .A(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_5237_)
);

INVX1 _14696_ (
    .A(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_5238_)
);

OAI22X1 _14697_ (
    .A(_5238_),
    .B(_3961__bF$buf1),
    .C(_5237_),
    .D(_3905_),
    .Y(_5239_)
);

NOR2X1 _14698_ (
    .A(_5236_),
    .B(_5239_),
    .Y(_5240_)
);

INVX1 _14699_ (
    .A(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_5241_)
);

INVX1 _14700_ (
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_5242_)
);

OAI22X1 _14701_ (
    .A(_5242_),
    .B(_3916__bF$buf1),
    .C(_3889__bF$buf1),
    .D(_5241_),
    .Y(_5243_)
);

INVX1 _14702_ (
    .A(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_5244_)
);

INVX1 _14703_ (
    .A(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_5245_)
);

OAI22X1 _14704_ (
    .A(_5245_),
    .B(_3915__bF$buf2),
    .C(_3924__bF$buf3),
    .D(_5244_),
    .Y(_5246_)
);

NOR2X1 _14705_ (
    .A(_5243_),
    .B(_5246_),
    .Y(_5247_)
);

NAND2X1 _14706_ (
    .A(_5240_),
    .B(_5247_),
    .Y(_5248_)
);

AOI22X1 _14707_ (
    .A(_3899__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [28]),
    .C(\datapath_1.regfile_1.regOut[24] [28]),
    .D(_3902__bF$buf4),
    .Y(_5249_)
);

AOI22X1 _14708_ (
    .A(_3947__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .C(_3952__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_5250_)
);

INVX1 _14709_ (
    .A(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_5251_)
);

INVX1 _14710_ (
    .A(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_5252_)
);

OAI22X1 _14711_ (
    .A(_5252_),
    .B(_3929__bF$buf1),
    .C(_3962__bF$buf2),
    .D(_5251_),
    .Y(_5253_)
);

INVX1 _14712_ (
    .A(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_5254_)
);

INVX1 _14713_ (
    .A(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_5255_)
);

OAI22X1 _14714_ (
    .A(_3869_),
    .B(_5254_),
    .C(_5255_),
    .D(_3956__bF$buf1),
    .Y(_5256_)
);

NOR2X1 _14715_ (
    .A(_5253_),
    .B(_5256_),
    .Y(_5257_)
);

NAND3X1 _14716_ (
    .A(_5250_),
    .B(_5249_),
    .C(_5257_),
    .Y(_5258_)
);

NOR2X1 _14717_ (
    .A(_5248_),
    .B(_5258_),
    .Y(_5259_)
);

AOI22X1 _14718_ (
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .B(_3989_),
    .C(\datapath_1.regfile_1.regOut[21] [28]),
    .D(_3990_),
    .Y(_5260_)
);

AOI22X1 _14719_ (
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[20] [28]),
    .D(_3904__bF$buf1),
    .Y(_5261_)
);

INVX1 _14720_ (
    .A(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_5262_)
);

INVX1 _14721_ (
    .A(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_5263_)
);

OAI22X1 _14722_ (
    .A(_5263_),
    .B(_3928_),
    .C(_5262_),
    .D(_3893_),
    .Y(_5264_)
);

INVX1 _14723_ (
    .A(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_5265_)
);

INVX1 _14724_ (
    .A(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_5266_)
);

OAI22X1 _14725_ (
    .A(_5266_),
    .B(_3957__bF$buf2),
    .C(_3865_),
    .D(_5265_),
    .Y(_5267_)
);

NOR2X1 _14726_ (
    .A(_5267_),
    .B(_5264_),
    .Y(_5268_)
);

NAND3X1 _14727_ (
    .A(_5261_),
    .B(_5260_),
    .C(_5268_),
    .Y(_5269_)
);

INVX1 _14728_ (
    .A(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_5270_)
);

INVX1 _14729_ (
    .A(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_5271_)
);

OAI22X1 _14730_ (
    .A(_4044_),
    .B(_5270_),
    .C(_5271_),
    .D(_3939__bF$buf1),
    .Y(_5272_)
);

INVX1 _14731_ (
    .A(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_5273_)
);

INVX1 _14732_ (
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_5274_)
);

OAI22X1 _14733_ (
    .A(_3923__bF$buf1),
    .B(_5274_),
    .C(_5273_),
    .D(_3944__bF$buf0),
    .Y(_5275_)
);

NOR2X1 _14734_ (
    .A(_5272_),
    .B(_5275_),
    .Y(_5276_)
);

AOI22X1 _14735_ (
    .A(_4062__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[8] [28]),
    .C(_3876_),
    .D(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_5277_)
);

AOI22X1 _14736_ (
    .A(_4038_),
    .B(\datapath_1.regfile_1.regOut[22] [28]),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_5278_)
);

NAND3X1 _14737_ (
    .A(_5277_),
    .B(_5278_),
    .C(_5276_),
    .Y(_5279_)
);

NOR2X1 _14738_ (
    .A(_5279_),
    .B(_5269_),
    .Y(_5280_)
);

AOI21X1 _14739_ (
    .A(_5280_),
    .B(_5259_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [28])
);

INVX1 _14740_ (
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_5281_)
);

INVX1 _14741_ (
    .A(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_5282_)
);

OAI22X1 _14742_ (
    .A(_5282_),
    .B(_3923__bF$buf0),
    .C(_5281_),
    .D(_3875__bF$buf0),
    .Y(_5283_)
);

INVX1 _14743_ (
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_5284_)
);

INVX1 _14744_ (
    .A(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_5285_)
);

OAI22X1 _14745_ (
    .A(_5285_),
    .B(_3915__bF$buf1),
    .C(_3886__bF$buf3),
    .D(_5284_),
    .Y(_5286_)
);

NOR2X1 _14746_ (
    .A(_5283_),
    .B(_5286_),
    .Y(_5287_)
);

AOI22X1 _14747_ (
    .A(_4070_),
    .B(\datapath_1.regfile_1.regOut[26] [29]),
    .C(_3990_),
    .D(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_5288_)
);

INVX1 _14748_ (
    .A(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_5289_)
);

NOR2X1 _14749_ (
    .A(_5289_),
    .B(_3939__bF$buf0),
    .Y(_5290_)
);

AOI21X1 _14750_ (
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .B(_3879__bF$buf0),
    .C(_5290_),
    .Y(_5291_)
);

NAND3X1 _14751_ (
    .A(_5291_),
    .B(_5288_),
    .C(_5287_),
    .Y(_5292_)
);

AOI22X1 _14752_ (
    .A(_4062__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[8] [29]),
    .C(\datapath_1.regfile_1.regOut[2] [29]),
    .D(_3975_),
    .Y(_5293_)
);

AOI22X1 _14753_ (
    .A(_3904__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[20] [29]),
    .C(\datapath_1.regfile_1.regOut[9] [29]),
    .D(_3950__bF$buf1),
    .Y(_5294_)
);

INVX1 _14754_ (
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_5295_)
);

INVX1 _14755_ (
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_5296_)
);

OAI22X1 _14756_ (
    .A(_3916__bF$buf0),
    .B(_5296_),
    .C(_5295_),
    .D(_3935__bF$buf0),
    .Y(_5297_)
);

INVX1 _14757_ (
    .A(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_5298_)
);

INVX1 _14758_ (
    .A(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_5299_)
);

OAI22X1 _14759_ (
    .A(_3889__bF$buf0),
    .B(_5299_),
    .C(_5298_),
    .D(_3910__bF$buf0),
    .Y(_5300_)
);

NOR2X1 _14760_ (
    .A(_5300_),
    .B(_5297_),
    .Y(_5301_)
);

NAND3X1 _14761_ (
    .A(_5294_),
    .B(_5293_),
    .C(_5301_),
    .Y(_5302_)
);

NOR2X1 _14762_ (
    .A(_5302_),
    .B(_5292_),
    .Y(_5303_)
);

INVX1 _14763_ (
    .A(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_5304_)
);

INVX1 _14764_ (
    .A(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_5305_)
);

OAI22X1 _14765_ (
    .A(_5305_),
    .B(_3961__bF$buf0),
    .C(_3962__bF$buf1),
    .D(_5304_),
    .Y(_5306_)
);

INVX1 _14766_ (
    .A(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_5307_)
);

INVX1 _14767_ (
    .A(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_5308_)
);

OAI22X1 _14768_ (
    .A(_3894__bF$buf0),
    .B(_5307_),
    .C(_5308_),
    .D(_3956__bF$buf0),
    .Y(_5309_)
);

NOR2X1 _14769_ (
    .A(_5306_),
    .B(_5309_),
    .Y(_5310_)
);

AOI22X1 _14770_ (
    .A(_3899__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [29]),
    .C(\datapath_1.regfile_1.regOut[24] [29]),
    .D(_3902__bF$buf3),
    .Y(_5311_)
);

AOI22X1 _14771_ (
    .A(_3952__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[18] [29]),
    .C(\datapath_1.regfile_1.regOut[30] [29]),
    .D(_3870__bF$buf1),
    .Y(_5312_)
);

NAND3X1 _14772_ (
    .A(_5311_),
    .B(_5312_),
    .C(_5310_),
    .Y(_5313_)
);

INVX1 _14773_ (
    .A(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_5314_)
);

INVX1 _14774_ (
    .A(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_5315_)
);

OAI22X1 _14775_ (
    .A(_3928_),
    .B(_5315_),
    .C(_5314_),
    .D(_3944__bF$buf3),
    .Y(_5316_)
);

INVX1 _14776_ (
    .A(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_5317_)
);

INVX1 _14777_ (
    .A(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_5318_)
);

OAI22X1 _14778_ (
    .A(_5318_),
    .B(_3957__bF$buf1),
    .C(_3946_),
    .D(_5317_),
    .Y(_5319_)
);

NOR2X1 _14779_ (
    .A(_5319_),
    .B(_5316_),
    .Y(_5320_)
);

INVX1 _14780_ (
    .A(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_5321_)
);

NOR2X1 _14781_ (
    .A(_5321_),
    .B(_3929__bF$buf0),
    .Y(_5322_)
);

AOI21X1 _14782_ (
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .B(_3906__bF$buf3),
    .C(_5322_),
    .Y(_5323_)
);

AOI22X1 _14783_ (
    .A(_3866__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [29]),
    .C(_4068__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_5324_)
);

NAND3X1 _14784_ (
    .A(_5323_),
    .B(_5324_),
    .C(_5320_),
    .Y(_5325_)
);

NOR2X1 _14785_ (
    .A(_5325_),
    .B(_5313_),
    .Y(_5326_)
);

AOI21X1 _14786_ (
    .A(_5326_),
    .B(_5303_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [29])
);

AOI22X1 _14787_ (
    .A(_3870__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[30] [30]),
    .C(_3906__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_5327_)
);

AOI22X1 _14788_ (
    .A(_3947__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [30]),
    .C(_3902__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_5328_)
);

INVX1 _14789_ (
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_5329_)
);

INVX1 _14790_ (
    .A(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_5330_)
);

OAI22X1 _14791_ (
    .A(_3889__bF$buf4),
    .B(_5329_),
    .C(_5330_),
    .D(_3886__bF$buf2),
    .Y(_5331_)
);

INVX1 _14792_ (
    .A(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_5332_)
);

INVX1 _14793_ (
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_5333_)
);

OAI22X1 _14794_ (
    .A(_3923__bF$buf4),
    .B(_5333_),
    .C(_5332_),
    .D(_3929__bF$buf4),
    .Y(_5334_)
);

NOR2X1 _14795_ (
    .A(_5334_),
    .B(_5331_),
    .Y(_5335_)
);

NAND3X1 _14796_ (
    .A(_5328_),
    .B(_5327_),
    .C(_5335_),
    .Y(_5336_)
);

AOI22X1 _14797_ (
    .A(_3904__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[20] [30]),
    .C(\datapath_1.regfile_1.regOut[25] [30]),
    .D(_3945_),
    .Y(_5337_)
);

AOI22X1 _14798_ (
    .A(_3899__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[23] [30]),
    .C(_3952__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_5338_)
);

INVX1 _14799_ (
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_5339_)
);

INVX1 _14800_ (
    .A(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_5340_)
);

OAI22X1 _14801_ (
    .A(_5339_),
    .B(_3910__bF$buf3),
    .C(_5340_),
    .D(_3911_),
    .Y(_5341_)
);

INVX1 _14802_ (
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_5342_)
);

INVX1 _14803_ (
    .A(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_5343_)
);

OAI22X1 _14804_ (
    .A(_3916__bF$buf4),
    .B(_5342_),
    .C(_5343_),
    .D(_3915__bF$buf0),
    .Y(_5344_)
);

NOR2X1 _14805_ (
    .A(_5341_),
    .B(_5344_),
    .Y(_5345_)
);

NAND3X1 _14806_ (
    .A(_5337_),
    .B(_5338_),
    .C(_5345_),
    .Y(_5346_)
);

NOR2X1 _14807_ (
    .A(_5346_),
    .B(_5336_),
    .Y(_5347_)
);

AOI22X1 _14808_ (
    .A(_3866__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [30]),
    .C(_4068__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_5348_)
);

AOI22X1 _14809_ (
    .A(_3876_),
    .B(\datapath_1.regfile_1.regOut[4] [30]),
    .C(\datapath_1.regfile_1.regOut[2] [30]),
    .D(_3975_),
    .Y(_5349_)
);

INVX1 _14810_ (
    .A(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_5350_)
);

INVX1 _14811_ (
    .A(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_5351_)
);

OAI22X1 _14812_ (
    .A(_5351_),
    .B(_3934__bF$buf2),
    .C(_3935__bF$buf3),
    .D(_5350_),
    .Y(_5352_)
);

INVX1 _14813_ (
    .A(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_5353_)
);

INVX1 _14814_ (
    .A(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_5354_)
);

OAI22X1 _14815_ (
    .A(_3928_),
    .B(_5353_),
    .C(_5354_),
    .D(_3956__bF$buf4),
    .Y(_5355_)
);

NOR2X1 _14816_ (
    .A(_5355_),
    .B(_5352_),
    .Y(_5356_)
);

NAND3X1 _14817_ (
    .A(_5349_),
    .B(_5348_),
    .C(_5356_),
    .Y(_5357_)
);

AOI22X1 _14818_ (
    .A(_3879__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[28] [30]),
    .C(_4070_),
    .D(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_5358_)
);

AOI22X1 _14819_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[17] [30]),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_5359_)
);

INVX1 _14820_ (
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_5360_)
);

INVX1 _14821_ (
    .A(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_5361_)
);

OAI22X1 _14822_ (
    .A(_5361_),
    .B(_3957__bF$buf0),
    .C(_3961__bF$buf4),
    .D(_5360_),
    .Y(_5362_)
);

INVX1 _14823_ (
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_5363_)
);

INVX1 _14824_ (
    .A(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_5364_)
);

OAI22X1 _14825_ (
    .A(_5363_),
    .B(_3894__bF$buf4),
    .C(_5364_),
    .D(_3939__bF$buf4),
    .Y(_5365_)
);

NOR2X1 _14826_ (
    .A(_5365_),
    .B(_5362_),
    .Y(_5366_)
);

NAND3X1 _14827_ (
    .A(_5359_),
    .B(_5358_),
    .C(_5366_),
    .Y(_5367_)
);

NOR2X1 _14828_ (
    .A(_5367_),
    .B(_5357_),
    .Y(_5368_)
);

AOI21X1 _14829_ (
    .A(_5368_),
    .B(_5347_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [30])
);

INVX1 _14830_ (
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_5369_)
);

INVX1 _14831_ (
    .A(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_5370_)
);

OAI22X1 _14832_ (
    .A(_5370_),
    .B(_3957__bF$buf4),
    .C(_5369_),
    .D(_4340_),
    .Y(_5371_)
);

INVX1 _14833_ (
    .A(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_5372_)
);

INVX1 _14834_ (
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_5373_)
);

OAI22X1 _14835_ (
    .A(_5373_),
    .B(_3894__bF$buf3),
    .C(_5372_),
    .D(_3951_),
    .Y(_5374_)
);

NOR2X1 _14836_ (
    .A(_5374_),
    .B(_5371_),
    .Y(_5375_)
);

INVX1 _14837_ (
    .A(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_5376_)
);

INVX1 _14838_ (
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_5377_)
);

OAI22X1 _14839_ (
    .A(_3916__bF$buf3),
    .B(_5377_),
    .C(_5376_),
    .D(_3924__bF$buf2),
    .Y(_5378_)
);

INVX1 _14840_ (
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_5379_)
);

INVX1 _14841_ (
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_5380_)
);

OAI22X1 _14842_ (
    .A(_3875__bF$buf3),
    .B(_5380_),
    .C(_5379_),
    .D(_3934__bF$buf1),
    .Y(_5381_)
);

NOR2X1 _14843_ (
    .A(_5381_),
    .B(_5378_),
    .Y(_5382_)
);

NAND2X1 _14844_ (
    .A(_5382_),
    .B(_5375_),
    .Y(_5383_)
);

INVX1 _14845_ (
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_5384_)
);

INVX1 _14846_ (
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_5385_)
);

OAI22X1 _14847_ (
    .A(_4044_),
    .B(_5384_),
    .C(_5385_),
    .D(_3935__bF$buf2),
    .Y(_5386_)
);

INVX1 _14848_ (
    .A(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_5387_)
);

INVX1 _14849_ (
    .A(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_5388_)
);

OAI22X1 _14850_ (
    .A(_5388_),
    .B(_3940__bF$buf2),
    .C(_3939__bF$buf3),
    .D(_5387_),
    .Y(_5389_)
);

NOR2X1 _14851_ (
    .A(_5389_),
    .B(_5386_),
    .Y(_5390_)
);

AOI22X1 _14852_ (
    .A(_3899__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [31]),
    .C(\datapath_1.regfile_1.regOut[30] [31]),
    .D(_3870__bF$buf3),
    .Y(_5391_)
);

AOI22X1 _14853_ (
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .B(_3987_),
    .C(\datapath_1.regfile_1.regOut[9] [31]),
    .D(_3950__bF$buf3),
    .Y(_5392_)
);

NAND3X1 _14854_ (
    .A(_5391_),
    .B(_5392_),
    .C(_5390_),
    .Y(_5393_)
);

NOR2X1 _14855_ (
    .A(_5393_),
    .B(_5383_),
    .Y(_5394_)
);

INVX1 _14856_ (
    .A(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_5395_)
);

NOR2X1 _14857_ (
    .A(_5395_),
    .B(_3961__bF$buf3),
    .Y(_5396_)
);

AOI21X1 _14858_ (
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .B(_4135_),
    .C(_5396_),
    .Y(_5397_)
);

AOI22X1 _14859_ (
    .A(_3947__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[27] [31]),
    .C(\datapath_1.regfile_1.regOut[31] [31]),
    .D(_3906__bF$buf1),
    .Y(_5398_)
);

INVX1 _14860_ (
    .A(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_5399_)
);

INVX1 _14861_ (
    .A(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_5400_)
);

OAI22X1 _14862_ (
    .A(_5400_),
    .B(_3928_),
    .C(_5399_),
    .D(_3893_),
    .Y(_5401_)
);

INVX1 _14863_ (
    .A(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_5402_)
);

INVX1 _14864_ (
    .A(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_5403_)
);

OAI22X1 _14865_ (
    .A(_3889__bF$buf3),
    .B(_5402_),
    .C(_5403_),
    .D(_3956__bF$buf3),
    .Y(_5404_)
);

NOR2X1 _14866_ (
    .A(_5404_),
    .B(_5401_),
    .Y(_5405_)
);

NAND3X1 _14867_ (
    .A(_5398_),
    .B(_5397_),
    .C(_5405_),
    .Y(_5406_)
);

INVX1 _14868_ (
    .A(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_5407_)
);

NOR2X1 _14869_ (
    .A(_5407_),
    .B(_3929__bF$buf3),
    .Y(_5408_)
);

AOI21X1 _14870_ (
    .A(_3866__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [31]),
    .C(_5408_),
    .Y(_5409_)
);

AOI22X1 _14871_ (
    .A(_3902__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[24] [31]),
    .C(\datapath_1.regfile_1.regOut[10] [31]),
    .D(_4087_),
    .Y(_5410_)
);

INVX1 _14872_ (
    .A(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_5411_)
);

INVX1 _14873_ (
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_5412_)
);

OAI22X1 _14874_ (
    .A(_3911_),
    .B(_5412_),
    .C(_5411_),
    .D(_3944__bF$buf2),
    .Y(_5413_)
);

INVX1 _14875_ (
    .A(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_5414_)
);

INVX1 _14876_ (
    .A(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_5415_)
);

OAI22X1 _14877_ (
    .A(_5415_),
    .B(_3923__bF$buf3),
    .C(_5414_),
    .D(_3886__bF$buf1),
    .Y(_5416_)
);

NOR2X1 _14878_ (
    .A(_5413_),
    .B(_5416_),
    .Y(_5417_)
);

NAND3X1 _14879_ (
    .A(_5410_),
    .B(_5409_),
    .C(_5417_),
    .Y(_5418_)
);

NOR2X1 _14880_ (
    .A(_5406_),
    .B(_5418_),
    .Y(_5419_)
);

AOI21X1 _14881_ (
    .A(_5419_),
    .B(_5394_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [31])
);

INVX1 _14882_ (
    .A(\datapath_1.PCJump [26]),
    .Y(_5420_)
);

NAND2X1 _14883_ (
    .A(\datapath_1.PCJump [25]),
    .B(_5420_),
    .Y(_5421_)
);

NOR2X1 _14884_ (
    .A(\datapath_1.PCJump [23]),
    .B(\datapath_1.PCJump [24]),
    .Y(_5422_)
);

NAND2X1 _14885_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5422_),
    .Y(_5423_)
);

NOR2X1 _14886_ (
    .A(_5421__bF$buf3),
    .B(_5423__bF$buf3),
    .Y(_5424_)
);

NAND2X1 _14887_ (
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .B(_5424_),
    .Y(_5425_)
);

AND2X2 _14888_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5426_)
);

NOR2X1 _14889_ (
    .A(\datapath_1.PCJump [25]),
    .B(\datapath_1.PCJump [26]),
    .Y(_5427_)
);

NAND3X1 _14890_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5427_),
    .C(_5426_),
    .Y(_5428_)
);

INVX4 _14891_ (
    .A(_5428__bF$buf3),
    .Y(_5429_)
);

INVX1 _14892_ (
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_5430_)
);

INVX1 _14893_ (
    .A(\datapath_1.PCJump [23]),
    .Y(_5431_)
);

NOR2X1 _14894_ (
    .A(\datapath_1.PCJump [24]),
    .B(_5431_),
    .Y(_5432_)
);

NAND3X1 _14895_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5427_),
    .C(_5432_),
    .Y(_5433_)
);

INVX1 _14896_ (
    .A(\datapath_1.PCJump [24]),
    .Y(_5434_)
);

NOR2X1 _14897_ (
    .A(\datapath_1.PCJump [23]),
    .B(_5434_),
    .Y(_5435_)
);

NAND3X1 _14898_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5427_),
    .C(_5435_),
    .Y(_5436_)
);

OAI22X1 _14899_ (
    .A(_3959_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_5430_),
    .Y(_5437_)
);

AOI21X1 _14900_ (
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .B(_5429_),
    .C(_5437_),
    .Y(_5438_)
);

INVX1 _14901_ (
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_5439_)
);

INVX1 _14902_ (
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_5440_)
);

INVX1 _14903_ (
    .A(\datapath_1.PCJump [25]),
    .Y(_5441_)
);

NOR2X1 _14904_ (
    .A(\datapath_1.PCJump [26]),
    .B(_5441_),
    .Y(_5442_)
);

NAND3X1 _14905_ (
    .A(_5426_),
    .B(\datapath_1.PCJump_27_bF$buf3 ),
    .C(_5442_),
    .Y(_5443_)
);

NOR2X1 _14906_ (
    .A(\datapath_1.PCJump [25]),
    .B(_5420_),
    .Y(_5444_)
);

INVX4 _14907_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_5445_)
);

NOR3X1 _14908_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .C(_5445_),
    .Y(_5446_)
);

NAND2X1 _14909_ (
    .A(_5444_),
    .B(_5446_),
    .Y(_5447_)
);

OAI22X1 _14910_ (
    .A(_5443_),
    .B(_5440_),
    .C(_5439_),
    .D(_5447_),
    .Y(_5448_)
);

NAND3X1 _14911_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5442_),
    .C(_5432_),
    .Y(_5449_)
);

NAND3X1 _14912_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5435_),
    .C(_5442_),
    .Y(_5450_)
);

OAI22X1 _14913_ (
    .A(_3933_),
    .B(_5449_),
    .C(_5450_),
    .D(_3932_),
    .Y(_5451_)
);

NOR2X1 _14914_ (
    .A(_5451_),
    .B(_5448_),
    .Y(_5452_)
);

NAND3X1 _14915_ (
    .A(_5438_),
    .B(_5425_),
    .C(_5452_),
    .Y(_5453_)
);

NAND3X1 _14916_ (
    .A(_5445_),
    .B(_5427_),
    .C(_5432_),
    .Y(_5454_)
);

INVX8 _14917_ (
    .A(_5454_),
    .Y(_5455_)
);

NOR3X1 _14918_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(\datapath_1.PCJump [23]),
    .C(\datapath_1.PCJump [24]),
    .Y(_5456_)
);

AND2X2 _14919_ (
    .A(_5442_),
    .B(_5456_),
    .Y(_5457_)
);

AOI22X1 _14920_ (
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [0]),
    .D(_5455__bF$buf4),
    .Y(_5458_)
);

NAND2X1 _14921_ (
    .A(_5442_),
    .B(_5435_),
    .Y(_5459_)
);

NOR2X1 _14922_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(_5459_),
    .Y(_5460_)
);

NAND2X1 _14923_ (
    .A(_5432_),
    .B(_5442_),
    .Y(_5461_)
);

NOR2X1 _14924_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5461_),
    .Y(_5462_)
);

AOI22X1 _14925_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [0]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_5463_)
);

INVX1 _14926_ (
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_5464_)
);

NAND3X1 _14927_ (
    .A(_5445_),
    .B(_5444_),
    .C(_5432_),
    .Y(_5465_)
);

NAND3X1 _14928_ (
    .A(_5445_),
    .B(_5435_),
    .C(_5444_),
    .Y(_5466_)
);

OAI22X1 _14929_ (
    .A(_5464_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_3914_),
    .Y(_5467_)
);

NAND2X1 _14930_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5468_)
);

NAND2X1 _14931_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5469_)
);

NOR2X1 _14932_ (
    .A(_5469_),
    .B(_5468_),
    .Y(_5470_)
);

NAND2X1 _14933_ (
    .A(_5445_),
    .B(_5470_),
    .Y(_5471_)
);

NAND2X1 _14934_ (
    .A(_5427_),
    .B(_5446_),
    .Y(_5472_)
);

OAI22X1 _14935_ (
    .A(_3882_),
    .B(_5471__bF$buf4),
    .C(_3913_),
    .D(_5472__bF$buf4),
    .Y(_5473_)
);

NOR2X1 _14936_ (
    .A(_5467_),
    .B(_5473_),
    .Y(_5474_)
);

NAND3X1 _14937_ (
    .A(_5463_),
    .B(_5458_),
    .C(_5474_),
    .Y(_5475_)
);

NOR2X1 _14938_ (
    .A(_5453_),
    .B(_5475_),
    .Y(_5476_)
);

NAND3X1 _14939_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5426_),
    .C(_5444_),
    .Y(_5477_)
);

INVX4 _14940_ (
    .A(_5477_),
    .Y(_5478_)
);

NAND2X1 _14941_ (
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .B(_5478__bF$buf3),
    .Y(_5479_)
);

INVX2 _14942_ (
    .A(_5468_),
    .Y(_5480_)
);

NAND3X1 _14943_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5422_),
    .C(_5480_),
    .Y(_5481_)
);

INVX8 _14944_ (
    .A(_5481_),
    .Y(_5482_)
);

INVX1 _14945_ (
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_5483_)
);

NAND3X1 _14946_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5444_),
    .C(_5432_),
    .Y(_5484_)
);

NAND3X1 _14947_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(_5435_),
    .C(_5444_),
    .Y(_5485_)
);

OAI22X1 _14948_ (
    .A(_5483_),
    .B(_5484__bF$buf4),
    .C(_5485__bF$buf4),
    .D(_3921_),
    .Y(_5486_)
);

AOI21X1 _14949_ (
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .B(_5482__bF$buf3),
    .C(_5486_),
    .Y(_5487_)
);

NAND3X1 _14950_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5480_),
    .C(_5435_),
    .Y(_5488_)
);

INVX4 _14951_ (
    .A(_5488__bF$buf3),
    .Y(_5489_)
);

INVX1 _14952_ (
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_5490_)
);

INVX1 _14953_ (
    .A(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_5491_)
);

NAND3X1 _14954_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5480_),
    .C(_5432_),
    .Y(_5492_)
);

NAND2X1 _14955_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5470_),
    .Y(_5493_)
);

OAI22X1 _14956_ (
    .A(_5492__bF$buf4),
    .B(_5491_),
    .C(_5490_),
    .D(_5493__bF$buf3),
    .Y(_5494_)
);

AOI21X1 _14957_ (
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .B(_5489_),
    .C(_5494_),
    .Y(_5495_)
);

NAND3X1 _14958_ (
    .A(_5479_),
    .B(_5495_),
    .C(_5487_),
    .Y(_5496_)
);

NAND2X1 _14959_ (
    .A(\datapath_1.PCJump [24]),
    .B(_5431_),
    .Y(_5497_)
);

AOI21X1 _14960_ (
    .A(_5497_),
    .B(_5469_),
    .C(_5421__bF$buf2),
    .Y(_5498_)
);

NAND2X1 _14961_ (
    .A(\datapath_1.PCJump [23]),
    .B(_5434_),
    .Y(_5499_)
);

NAND2X1 _14962_ (
    .A(_5434_),
    .B(_5431_),
    .Y(_5500_)
);

AOI21X1 _14963_ (
    .A(_5500_),
    .B(_5499_),
    .C(_5421__bF$buf1),
    .Y(_5501_)
);

OAI21X1 _14964_ (
    .A(_5498_),
    .B(_5501_),
    .C(_5445_),
    .Y(_5502_)
);

INVX1 _14965_ (
    .A(_5427_),
    .Y(_5503_)
);

NOR2X1 _14966_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump_27_bF$buf4 ),
    .Y(_5504_)
);

OAI21X1 _14967_ (
    .A(_5497_),
    .B(_5503_),
    .C(_5504_),
    .Y(_5505_)
);

NAND3X1 _14968_ (
    .A(_5445_),
    .B(_5427_),
    .C(_5426_),
    .Y(_5506_)
);

NAND3X1 _14969_ (
    .A(\datapath_1.PCJump [23]),
    .B(_5434_),
    .C(_5427_),
    .Y(_5507_)
);

OAI21X1 _14970_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(_5507_),
    .C(_5506__bF$buf4),
    .Y(_5508_)
);

NOR2X1 _14971_ (
    .A(_5505_),
    .B(_5508_),
    .Y(_5509_)
);

NAND3X1 _14972_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [0]),
    .C(_5509_),
    .Y(_5510_)
);

NAND3X1 _14973_ (
    .A(_5445_),
    .B(_5427_),
    .C(_5435_),
    .Y(_5511_)
);

OAI22X1 _14974_ (
    .A(_3922_),
    .B(_5506__bF$buf3),
    .C(_3938_),
    .D(_5511__bF$buf4),
    .Y(_5512_)
);

NAND3X1 _14975_ (
    .A(_5426_),
    .B(_5445_),
    .C(_5442_),
    .Y(_5513_)
);

NAND2X1 _14976_ (
    .A(_5456_),
    .B(_5444_),
    .Y(_5514_)
);

OAI22X1 _14977_ (
    .A(_5514__bF$buf4),
    .B(_3909_),
    .C(_3927_),
    .D(_5513__bF$buf4),
    .Y(_5515_)
);

NOR2X1 _14978_ (
    .A(_5515_),
    .B(_5512_),
    .Y(_5516_)
);

NAND3X1 _14979_ (
    .A(_5445_),
    .B(_5426_),
    .C(_5444_),
    .Y(_5517_)
);

NAND2X1 _14980_ (
    .A(_5480_),
    .B(_5456_),
    .Y(_5518_)
);

OAI22X1 _14981_ (
    .A(_5518__bF$buf4),
    .B(_3891_),
    .C(_3926_),
    .D(_5517__bF$buf4),
    .Y(_5519_)
);

NAND3X1 _14982_ (
    .A(_5445_),
    .B(_5480_),
    .C(_5432_),
    .Y(_5520_)
);

NAND3X1 _14983_ (
    .A(_5445_),
    .B(_5480_),
    .C(_5435_),
    .Y(_5521_)
);

OAI22X1 _14984_ (
    .A(_3954_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_3960_),
    .Y(_5522_)
);

NOR2X1 _14985_ (
    .A(_5519_),
    .B(_5522_),
    .Y(_5523_)
);

NAND3X1 _14986_ (
    .A(_5516_),
    .B(_5523_),
    .C(_5510_),
    .Y(_5524_)
);

NOR2X1 _14987_ (
    .A(_5496_),
    .B(_5524_),
    .Y(_5525_)
);

AOI21X1 _14988_ (
    .A(_5525_),
    .B(_5476_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [0])
);

INVX1 _14989_ (
    .A(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_5526_)
);

OAI22X1 _14990_ (
    .A(_3967_),
    .B(_5433__bF$buf3),
    .C(_5436__bF$buf3),
    .D(_5526_),
    .Y(_5527_)
);

NOR2X1 _14991_ (
    .A(_4000_),
    .B(_5428__bF$buf2),
    .Y(_5528_)
);

INVX1 _14992_ (
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_5529_)
);

NOR3X1 _14993_ (
    .A(_5421__bF$buf0),
    .B(_5529_),
    .C(_5423__bF$buf2),
    .Y(_5530_)
);

NOR3X1 _14994_ (
    .A(_5528_),
    .B(_5530_),
    .C(_5527_),
    .Y(_5531_)
);

INVX1 _14995_ (
    .A(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_5532_)
);

OAI22X1 _14996_ (
    .A(_5532_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_4007_),
    .Y(_5533_)
);

AOI21X1 _14997_ (
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .B(_5482__bF$buf2),
    .C(_5533_),
    .Y(_5534_)
);

INVX1 _14998_ (
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_5535_)
);

INVX1 _14999_ (
    .A(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_5536_)
);

OAI22X1 _15000_ (
    .A(_5492__bF$buf3),
    .B(_5536_),
    .C(_5535_),
    .D(_5493__bF$buf2),
    .Y(_5537_)
);

INVX1 _15001_ (
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_5538_)
);

INVX1 _15002_ (
    .A(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_5539_)
);

OAI22X1 _15003_ (
    .A(_5539_),
    .B(_5477_),
    .C(_5488__bF$buf2),
    .D(_5538_),
    .Y(_5540_)
);

NOR2X1 _15004_ (
    .A(_5540_),
    .B(_5537_),
    .Y(_5541_)
);

NAND3X1 _15005_ (
    .A(_5534_),
    .B(_5541_),
    .C(_5531_),
    .Y(_5542_)
);

AOI22X1 _15006_ (
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [1]),
    .D(_5455__bF$buf3),
    .Y(_5543_)
);

AOI22X1 _15007_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [1]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_5544_)
);

INVX1 _15008_ (
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_5545_)
);

OAI22X1 _15009_ (
    .A(_5545_),
    .B(_5471__bF$buf3),
    .C(_3970_),
    .D(_5472__bF$buf3),
    .Y(_5546_)
);

INVX1 _15010_ (
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_5547_)
);

OAI22X1 _15011_ (
    .A(_5547_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_3971_),
    .Y(_5548_)
);

NOR2X1 _15012_ (
    .A(_5548_),
    .B(_5546_),
    .Y(_5549_)
);

NAND3X1 _15013_ (
    .A(_5544_),
    .B(_5543_),
    .C(_5549_),
    .Y(_5550_)
);

NOR2X1 _15014_ (
    .A(_5550_),
    .B(_5542_),
    .Y(_5551_)
);

INVX1 _15015_ (
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_5552_)
);

OAI21X1 _15016_ (
    .A(_5426_),
    .B(_5435_),
    .C(_5442_),
    .Y(_5553_)
);

OAI21X1 _15017_ (
    .A(_5422_),
    .B(_5432_),
    .C(_5442_),
    .Y(_5554_)
);

AOI21X1 _15018_ (
    .A(_5553_),
    .B(_5554_),
    .C(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_5555_)
);

INVX1 _15019_ (
    .A(_5504_),
    .Y(_5556_)
);

AOI21X1 _15020_ (
    .A(_5435_),
    .B(_5427_),
    .C(_5556_),
    .Y(_5557_)
);

NAND3X1 _15021_ (
    .A(_5454_),
    .B(_5506__bF$buf2),
    .C(_5557_),
    .Y(_5558_)
);

NOR3X1 _15022_ (
    .A(_5552_),
    .B(_5558__bF$buf3),
    .C(_5555__bF$buf3),
    .Y(_5559_)
);

NOR3X1 _15023_ (
    .A(_5469_),
    .B(_5445_),
    .C(_5421__bF$buf3),
    .Y(_5560_)
);

AND2X2 _15024_ (
    .A(_5446_),
    .B(_5444_),
    .Y(_5561_)
);

AOI22X1 _15025_ (
    .A(_5560__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [1]),
    .C(\datapath_1.regfile_1.regOut[24] [1]),
    .D(_5561__bF$buf3),
    .Y(_5562_)
);

INVX8 _15026_ (
    .A(_5450_),
    .Y(_5563_)
);

NAND2X1 _15027_ (
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .B(_5563__bF$buf3),
    .Y(_5564_)
);

INVX8 _15028_ (
    .A(_5449_),
    .Y(_5565_)
);

NAND2X1 _15029_ (
    .A(\datapath_1.regfile_1.regOut[21] [1]),
    .B(_5565__bF$buf3),
    .Y(_5566_)
);

NAND3X1 _15030_ (
    .A(_5564_),
    .B(_5562_),
    .C(_5566_),
    .Y(_5567_)
);

INVX1 _15031_ (
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_5568_)
);

OAI22X1 _15032_ (
    .A(_3984_),
    .B(_5506__bF$buf1),
    .C(_5568_),
    .D(_5511__bF$buf3),
    .Y(_5569_)
);

OAI22X1 _15033_ (
    .A(_5514__bF$buf3),
    .B(_3996_),
    .C(_4008_),
    .D(_5513__bF$buf3),
    .Y(_5570_)
);

NOR2X1 _15034_ (
    .A(_5570_),
    .B(_5569_),
    .Y(_5571_)
);

OAI22X1 _15035_ (
    .A(_5518__bF$buf3),
    .B(_3983_),
    .C(_3968_),
    .D(_5517__bF$buf3),
    .Y(_5572_)
);

OAI22X1 _15036_ (
    .A(_4005_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_4004_),
    .Y(_5573_)
);

NOR2X1 _15037_ (
    .A(_5572_),
    .B(_5573_),
    .Y(_5574_)
);

NAND2X1 _15038_ (
    .A(_5571_),
    .B(_5574_),
    .Y(_5575_)
);

NOR3X1 _15039_ (
    .A(_5567_),
    .B(_5559_),
    .C(_5575_),
    .Y(_5576_)
);

AOI21X1 _15040_ (
    .A(_5551_),
    .B(_5576_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [1])
);

NOR2X1 _15041_ (
    .A(_4046_),
    .B(_5428__bF$buf1),
    .Y(_5577_)
);

INVX1 _15042_ (
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_5578_)
);

NOR3X1 _15043_ (
    .A(_5421__bF$buf2),
    .B(_5578_),
    .C(_5423__bF$buf1),
    .Y(_5579_)
);

OAI22X1 _15044_ (
    .A(_4056_),
    .B(_5433__bF$buf2),
    .C(_5436__bF$buf2),
    .D(_4043_),
    .Y(_5580_)
);

NOR3X1 _15045_ (
    .A(_5579_),
    .B(_5577_),
    .C(_5580_),
    .Y(_5581_)
);

INVX1 _15046_ (
    .A(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_5582_)
);

INVX1 _15047_ (
    .A(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_5583_)
);

OAI22X1 _15048_ (
    .A(_5492__bF$buf2),
    .B(_5583_),
    .C(_5582_),
    .D(_5493__bF$buf1),
    .Y(_5584_)
);

AOI21X1 _15049_ (
    .A(\datapath_1.regfile_1.regOut[30] [2]),
    .B(_5489_),
    .C(_5584_),
    .Y(_5585_)
);

INVX1 _15050_ (
    .A(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_5586_)
);

OAI22X1 _15051_ (
    .A(_5586_),
    .B(_5484__bF$buf2),
    .C(_5485__bF$buf2),
    .D(_4053_),
    .Y(_5587_)
);

OAI22X1 _15052_ (
    .A(_5481_),
    .B(_4042_),
    .C(_4018_),
    .D(_5477_),
    .Y(_5588_)
);

NOR2X1 _15053_ (
    .A(_5588_),
    .B(_5587_),
    .Y(_5589_)
);

NAND3X1 _15054_ (
    .A(_5585_),
    .B(_5589_),
    .C(_5581_),
    .Y(_5590_)
);

AOI22X1 _15055_ (
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .B(_5457__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[1] [2]),
    .D(_5455__bF$buf2),
    .Y(_5591_)
);

AOI22X1 _15056_ (
    .A(_5460__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [2]),
    .C(_5462__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_5592_)
);

OAI22X1 _15057_ (
    .A(_4031_),
    .B(_5465__bF$buf2),
    .C(_5466__bF$buf2),
    .D(_4016_),
    .Y(_5593_)
);

OAI22X1 _15058_ (
    .A(_4019_),
    .B(_5471__bF$buf2),
    .C(_4054_),
    .D(_5472__bF$buf2),
    .Y(_5594_)
);

NOR2X1 _15059_ (
    .A(_5593_),
    .B(_5594_),
    .Y(_5595_)
);

NAND3X1 _15060_ (
    .A(_5592_),
    .B(_5591_),
    .C(_5595_),
    .Y(_5596_)
);

NOR2X1 _15061_ (
    .A(_5596_),
    .B(_5590_),
    .Y(_5597_)
);

NOR3X1 _15062_ (
    .A(_4033_),
    .B(_5558__bF$buf2),
    .C(_5555__bF$buf2),
    .Y(_5598_)
);

NAND2X1 _15063_ (
    .A(\datapath_1.regfile_1.regOut[22] [2]),
    .B(_5563__bF$buf2),
    .Y(_5599_)
);

NAND2X1 _15064_ (
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .B(_5565__bF$buf2),
    .Y(_5600_)
);

AOI22X1 _15065_ (
    .A(_5560__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [2]),
    .C(\datapath_1.regfile_1.regOut[24] [2]),
    .D(_5561__bF$buf2),
    .Y(_5601_)
);

NAND3X1 _15066_ (
    .A(_5599_),
    .B(_5601_),
    .C(_5600_),
    .Y(_5602_)
);

INVX1 _15067_ (
    .A(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_5603_)
);

OAI22X1 _15068_ (
    .A(_4026_),
    .B(_5506__bF$buf0),
    .C(_5603_),
    .D(_5511__bF$buf2),
    .Y(_5604_)
);

INVX1 _15069_ (
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_5605_)
);

INVX1 _15070_ (
    .A(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_5606_)
);

OAI22X1 _15071_ (
    .A(_5514__bF$buf2),
    .B(_5605_),
    .C(_5606_),
    .D(_5513__bF$buf2),
    .Y(_5607_)
);

NOR2X1 _15072_ (
    .A(_5607_),
    .B(_5604_),
    .Y(_5608_)
);

OAI22X1 _15073_ (
    .A(_5518__bF$buf2),
    .B(_4015_),
    .C(_4025_),
    .D(_5517__bF$buf2),
    .Y(_5609_)
);

OAI22X1 _15074_ (
    .A(_4022_),
    .B(_5520__bF$buf2),
    .C(_5521__bF$buf2),
    .D(_4030_),
    .Y(_5610_)
);

NOR2X1 _15075_ (
    .A(_5609_),
    .B(_5610_),
    .Y(_5611_)
);

NAND2X1 _15076_ (
    .A(_5608_),
    .B(_5611_),
    .Y(_5612_)
);

NOR3X1 _15077_ (
    .A(_5602_),
    .B(_5598_),
    .C(_5612_),
    .Y(_5613_)
);

AOI21X1 _15078_ (
    .A(_5597_),
    .B(_5613_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [2])
);

OAI22X1 _15079_ (
    .A(_4106_),
    .B(_5433__bF$buf1),
    .C(_5436__bF$buf1),
    .D(_4109_),
    .Y(_5614_)
);

NOR2X1 _15080_ (
    .A(_4083_),
    .B(_5428__bF$buf0),
    .Y(_5615_)
);

INVX1 _15081_ (
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_5616_)
);

NOR3X1 _15082_ (
    .A(_5421__bF$buf1),
    .B(_5616_),
    .C(_5423__bF$buf0),
    .Y(_5617_)
);

NOR3X1 _15083_ (
    .A(_5615_),
    .B(_5617_),
    .C(_5614_),
    .Y(_5618_)
);

INVX1 _15084_ (
    .A(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_5619_)
);

OAI22X1 _15085_ (
    .A(_4080_),
    .B(_5484__bF$buf1),
    .C(_5485__bF$buf1),
    .D(_5619_),
    .Y(_5620_)
);

AOI21X1 _15086_ (
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .B(_5482__bF$buf1),
    .C(_5620_),
    .Y(_5621_)
);

INVX1 _15087_ (
    .A(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_5622_)
);

INVX1 _15088_ (
    .A(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_5623_)
);

OAI22X1 _15089_ (
    .A(_5623_),
    .B(_5449_),
    .C(_5450_),
    .D(_5622_),
    .Y(_5624_)
);

INVX1 _15090_ (
    .A(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_5625_)
);

OAI22X1 _15091_ (
    .A(_5443_),
    .B(_4105_),
    .C(_5625_),
    .D(_5447_),
    .Y(_5626_)
);

NOR2X1 _15092_ (
    .A(_5624_),
    .B(_5626_),
    .Y(_5627_)
);

NAND3X1 _15093_ (
    .A(_5621_),
    .B(_5627_),
    .C(_5618_),
    .Y(_5628_)
);

AOI22X1 _15094_ (
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .B(_5457__bF$buf1),
    .C(\datapath_1.regfile_1.regOut[1] [3]),
    .D(_5455__bF$buf1),
    .Y(_5629_)
);

AOI22X1 _15095_ (
    .A(_5460__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [3]),
    .C(_5462__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_5630_)
);

INVX1 _15096_ (
    .A(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_5631_)
);

INVX1 _15097_ (
    .A(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_5632_)
);

OAI22X1 _15098_ (
    .A(_5632_),
    .B(_5465__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_5631_),
    .Y(_5633_)
);

INVX1 _15099_ (
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_5634_)
);

OAI22X1 _15100_ (
    .A(_5634_),
    .B(_5471__bF$buf1),
    .C(_4081_),
    .D(_5472__bF$buf1),
    .Y(_5635_)
);

NOR2X1 _15101_ (
    .A(_5633_),
    .B(_5635_),
    .Y(_5636_)
);

NAND3X1 _15102_ (
    .A(_5630_),
    .B(_5629_),
    .C(_5636_),
    .Y(_5637_)
);

NOR2X1 _15103_ (
    .A(_5637_),
    .B(_5628_),
    .Y(_5638_)
);

NOR3X1 _15104_ (
    .A(_4075_),
    .B(_5558__bF$buf1),
    .C(_5555__bF$buf1),
    .Y(_5639_)
);

NAND2X1 _15105_ (
    .A(\datapath_1.regfile_1.regOut[27] [3]),
    .B(_5478__bF$buf2),
    .Y(_5640_)
);

NOR3X1 _15106_ (
    .A(_5445_),
    .B(_5468_),
    .C(_5499_),
    .Y(_5641_)
);

AND2X2 _15107_ (
    .A(_5470_),
    .B(\datapath_1.PCJump_27_bF$buf1 ),
    .Y(_5642_)
);

AOI22X1 _15108_ (
    .A(\datapath_1.regfile_1.regOut[29] [3]),
    .B(_5641_),
    .C(\datapath_1.regfile_1.regOut[31] [3]),
    .D(_5642_),
    .Y(_5643_)
);

NAND2X1 _15109_ (
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .B(_5489_),
    .Y(_5644_)
);

NAND3X1 _15110_ (
    .A(_5644_),
    .B(_5643_),
    .C(_5640_),
    .Y(_5645_)
);

OAI22X1 _15111_ (
    .A(_4100_),
    .B(_5506__bF$buf4),
    .C(_4073_),
    .D(_5511__bF$buf1),
    .Y(_5646_)
);

INVX1 _15112_ (
    .A(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_5647_)
);

OAI22X1 _15113_ (
    .A(_5514__bF$buf1),
    .B(_4095_),
    .C(_5647_),
    .D(_5513__bF$buf1),
    .Y(_5648_)
);

NOR2X1 _15114_ (
    .A(_5648_),
    .B(_5646_),
    .Y(_5649_)
);

OAI22X1 _15115_ (
    .A(_5518__bF$buf1),
    .B(_4093_),
    .C(_4072_),
    .D(_5517__bF$buf1),
    .Y(_5650_)
);

INVX1 _15116_ (
    .A(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_5651_)
);

OAI22X1 _15117_ (
    .A(_5651_),
    .B(_5520__bF$buf1),
    .C(_5521__bF$buf1),
    .D(_4092_),
    .Y(_5652_)
);

NOR2X1 _15118_ (
    .A(_5650_),
    .B(_5652_),
    .Y(_5653_)
);

NAND2X1 _15119_ (
    .A(_5649_),
    .B(_5653_),
    .Y(_5654_)
);

NOR3X1 _15120_ (
    .A(_5645_),
    .B(_5639_),
    .C(_5654_),
    .Y(_5655_)
);

AOI21X1 _15121_ (
    .A(_5638_),
    .B(_5655_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [3])
);

AOI22X1 _15122_ (
    .A(_5563__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[22] [4]),
    .C(_5565__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_5656_)
);

INVX1 _15123_ (
    .A(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_5657_)
);

INVX1 _15124_ (
    .A(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_5658_)
);

OAI22X1 _15125_ (
    .A(_5658_),
    .B(_5433__bF$buf0),
    .C(_5436__bF$buf0),
    .D(_5657_),
    .Y(_5659_)
);

AOI21X1 _15126_ (
    .A(\datapath_1.regfile_1.regOut[20] [4]),
    .B(_5424_),
    .C(_5659_),
    .Y(_5660_)
);

AOI22X1 _15127_ (
    .A(_5429_),
    .B(\datapath_1.regfile_1.regOut[19] [4]),
    .C(\datapath_1.regfile_1.regOut[24] [4]),
    .D(_5561__bF$buf1),
    .Y(_5661_)
);

NAND3X1 _15128_ (
    .A(_5661_),
    .B(_5656_),
    .C(_5660_),
    .Y(_5662_)
);

AOI22X1 _15129_ (
    .A(\datapath_1.regfile_1.regOut[4] [4]),
    .B(_5457__bF$buf0),
    .C(\datapath_1.regfile_1.regOut[1] [4]),
    .D(_5455__bF$buf0),
    .Y(_5663_)
);

AOI22X1 _15130_ (
    .A(_5460__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [4]),
    .C(_5462__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_5664_)
);

OAI22X1 _15131_ (
    .A(_4118_),
    .B(_5465__bF$buf0),
    .C(_5466__bF$buf0),
    .D(_4117_),
    .Y(_5665_)
);

OAI22X1 _15132_ (
    .A(_4121_),
    .B(_5471__bF$buf0),
    .C(_4120_),
    .D(_5472__bF$buf0),
    .Y(_5666_)
);

NOR2X1 _15133_ (
    .A(_5665_),
    .B(_5666_),
    .Y(_5667_)
);

NAND3X1 _15134_ (
    .A(_5664_),
    .B(_5663_),
    .C(_5667_),
    .Y(_5668_)
);

NOR2X1 _15135_ (
    .A(_5662_),
    .B(_5668_),
    .Y(_5669_)
);

NAND2X1 _15136_ (
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .B(_5560__bF$buf1),
    .Y(_5670_)
);

INVX1 _15137_ (
    .A(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_5671_)
);

OAI22X1 _15138_ (
    .A(_5671_),
    .B(_5484__bF$buf0),
    .C(_5485__bF$buf0),
    .D(_4145_),
    .Y(_5672_)
);

AOI21X1 _15139_ (
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .B(_5482__bF$buf0),
    .C(_5672_),
    .Y(_5673_)
);

INVX1 _15140_ (
    .A(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_5674_)
);

OAI22X1 _15141_ (
    .A(_4154_),
    .B(_5477_),
    .C(_5488__bF$buf1),
    .D(_5674_),
    .Y(_5675_)
);

INVX1 _15142_ (
    .A(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_5676_)
);

NAND3X1 _15143_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(\datapath_1.regfile_1.regOut[31] [4]),
    .C(_5470_),
    .Y(_5677_)
);

OAI21X1 _15144_ (
    .A(_5676_),
    .B(_5492__bF$buf1),
    .C(_5677_),
    .Y(_5678_)
);

NOR2X1 _15145_ (
    .A(_5678_),
    .B(_5675_),
    .Y(_5679_)
);

NAND3X1 _15146_ (
    .A(_5670_),
    .B(_5679_),
    .C(_5673_),
    .Y(_5680_)
);

NAND3X1 _15147_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [4]),
    .C(_5509_),
    .Y(_5681_)
);

OAI22X1 _15148_ (
    .A(_4143_),
    .B(_5506__bF$buf3),
    .C(_4142_),
    .D(_5511__bF$buf0),
    .Y(_5682_)
);

INVX1 _15149_ (
    .A(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_5683_)
);

OAI22X1 _15150_ (
    .A(_5514__bF$buf0),
    .B(_4150_),
    .C(_5683_),
    .D(_5513__bF$buf0),
    .Y(_5684_)
);

NOR2X1 _15151_ (
    .A(_5684_),
    .B(_5682_),
    .Y(_5685_)
);

OAI22X1 _15152_ (
    .A(_5518__bF$buf0),
    .B(_4128_),
    .C(_4129_),
    .D(_5517__bF$buf0),
    .Y(_5686_)
);

OAI22X1 _15153_ (
    .A(_4132_),
    .B(_5520__bF$buf0),
    .C(_5521__bF$buf0),
    .D(_4131_),
    .Y(_5687_)
);

NOR2X1 _15154_ (
    .A(_5686_),
    .B(_5687_),
    .Y(_5688_)
);

NAND3X1 _15155_ (
    .A(_5685_),
    .B(_5688_),
    .C(_5681_),
    .Y(_5689_)
);

NOR2X1 _15156_ (
    .A(_5680_),
    .B(_5689_),
    .Y(_5690_)
);

AOI21X1 _15157_ (
    .A(_5690_),
    .B(_5669_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [4])
);

NOR2X1 _15158_ (
    .A(_4194_),
    .B(_5428__bF$buf3),
    .Y(_5691_)
);

INVX1 _15159_ (
    .A(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_5692_)
);

NOR3X1 _15160_ (
    .A(_5421__bF$buf0),
    .B(_5692_),
    .C(_5423__bF$buf3),
    .Y(_5693_)
);

OAI22X1 _15161_ (
    .A(_4176_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_4197_),
    .Y(_5694_)
);

NOR3X1 _15162_ (
    .A(_5693_),
    .B(_5691_),
    .C(_5694_),
    .Y(_5695_)
);

INVX1 _15163_ (
    .A(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_5696_)
);

OAI22X1 _15164_ (
    .A(_4167_),
    .B(_5484__bF$buf4),
    .C(_5485__bF$buf4),
    .D(_5696_),
    .Y(_5697_)
);

AOI21X1 _15165_ (
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .B(_5482__bF$buf3),
    .C(_5697_),
    .Y(_5698_)
);

INVX1 _15166_ (
    .A(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_5699_)
);

OAI22X1 _15167_ (
    .A(_5492__bF$buf0),
    .B(_4189_),
    .C(_5699_),
    .D(_5493__bF$buf0),
    .Y(_5700_)
);

INVX1 _15168_ (
    .A(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_5701_)
);

INVX1 _15169_ (
    .A(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_5702_)
);

OAI22X1 _15170_ (
    .A(_5702_),
    .B(_5477_),
    .C(_5488__bF$buf0),
    .D(_5701_),
    .Y(_5703_)
);

NOR2X1 _15171_ (
    .A(_5703_),
    .B(_5700_),
    .Y(_5704_)
);

NAND3X1 _15172_ (
    .A(_5698_),
    .B(_5704_),
    .C(_5695_),
    .Y(_5705_)
);

AOI22X1 _15173_ (
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [5]),
    .D(_5455__bF$buf4),
    .Y(_5706_)
);

AOI22X1 _15174_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [5]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_5707_)
);

INVX1 _15175_ (
    .A(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_5708_)
);

INVX1 _15176_ (
    .A(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_5709_)
);

OAI22X1 _15177_ (
    .A(_5709_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_5708_),
    .Y(_5710_)
);

OAI22X1 _15178_ (
    .A(_4174_),
    .B(_5471__bF$buf4),
    .C(_4198_),
    .D(_5472__bF$buf4),
    .Y(_5711_)
);

NOR2X1 _15179_ (
    .A(_5710_),
    .B(_5711_),
    .Y(_5712_)
);

NAND3X1 _15180_ (
    .A(_5707_),
    .B(_5706_),
    .C(_5712_),
    .Y(_5713_)
);

NOR2X1 _15181_ (
    .A(_5713_),
    .B(_5705_),
    .Y(_5714_)
);

INVX1 _15182_ (
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_5715_)
);

NOR3X1 _15183_ (
    .A(_5715_),
    .B(_5558__bF$buf0),
    .C(_5555__bF$buf0),
    .Y(_5716_)
);

NAND2X1 _15184_ (
    .A(\datapath_1.regfile_1.regOut[22] [5]),
    .B(_5563__bF$buf0),
    .Y(_5717_)
);

NAND2X1 _15185_ (
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .B(_5565__bF$buf0),
    .Y(_5718_)
);

AOI22X1 _15186_ (
    .A(_5560__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [5]),
    .C(\datapath_1.regfile_1.regOut[24] [5]),
    .D(_5561__bF$buf0),
    .Y(_5719_)
);

NAND3X1 _15187_ (
    .A(_5717_),
    .B(_5719_),
    .C(_5718_),
    .Y(_5720_)
);

OAI22X1 _15188_ (
    .A(_4183_),
    .B(_5506__bF$buf2),
    .C(_4177_),
    .D(_5511__bF$buf4),
    .Y(_5721_)
);

INVX1 _15189_ (
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_5722_)
);

INVX1 _15190_ (
    .A(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_5723_)
);

OAI22X1 _15191_ (
    .A(_5514__bF$buf4),
    .B(_5722_),
    .C(_5723_),
    .D(_5513__bF$buf4),
    .Y(_5724_)
);

NOR2X1 _15192_ (
    .A(_5724_),
    .B(_5721_),
    .Y(_5725_)
);

OAI22X1 _15193_ (
    .A(_5518__bF$buf4),
    .B(_4186_),
    .C(_4190_),
    .D(_5517__bF$buf4),
    .Y(_5726_)
);

OAI22X1 _15194_ (
    .A(_4187_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_4201_),
    .Y(_5727_)
);

NOR2X1 _15195_ (
    .A(_5726_),
    .B(_5727_),
    .Y(_5728_)
);

NAND2X1 _15196_ (
    .A(_5725_),
    .B(_5728_),
    .Y(_5729_)
);

NOR3X1 _15197_ (
    .A(_5720_),
    .B(_5716_),
    .C(_5729_),
    .Y(_5730_)
);

AOI21X1 _15198_ (
    .A(_5714_),
    .B(_5730_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [5])
);

NAND2X1 _15199_ (
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .B(_5489_),
    .Y(_5731_)
);

AOI22X1 _15200_ (
    .A(\datapath_1.regfile_1.regOut[29] [6]),
    .B(_5641_),
    .C(\datapath_1.regfile_1.regOut[31] [6]),
    .D(_5642_),
    .Y(_5732_)
);

INVX1 _15201_ (
    .A(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_5733_)
);

INVX1 _15202_ (
    .A(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_5734_)
);

OAI22X1 _15203_ (
    .A(_5734_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_5733_),
    .Y(_5735_)
);

INVX1 _15204_ (
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_5736_)
);

OAI22X1 _15205_ (
    .A(_5481_),
    .B(_5736_),
    .C(_4245_),
    .D(_5477_),
    .Y(_5737_)
);

NOR2X1 _15206_ (
    .A(_5737_),
    .B(_5735_),
    .Y(_5738_)
);

NAND3X1 _15207_ (
    .A(_5732_),
    .B(_5731_),
    .C(_5738_),
    .Y(_5739_)
);

AOI22X1 _15208_ (
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [6]),
    .D(_5455__bF$buf3),
    .Y(_5740_)
);

AOI22X1 _15209_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [6]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_5741_)
);

INVX1 _15210_ (
    .A(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_5742_)
);

INVX1 _15211_ (
    .A(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_5743_)
);

OAI22X1 _15212_ (
    .A(_5743_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_5742_),
    .Y(_5744_)
);

INVX1 _15213_ (
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_5745_)
);

OAI22X1 _15214_ (
    .A(_5745_),
    .B(_5471__bF$buf3),
    .C(_4238_),
    .D(_5472__bF$buf3),
    .Y(_5746_)
);

NOR2X1 _15215_ (
    .A(_5744_),
    .B(_5746_),
    .Y(_5747_)
);

NAND3X1 _15216_ (
    .A(_5741_),
    .B(_5740_),
    .C(_5747_),
    .Y(_5748_)
);

NOR2X1 _15217_ (
    .A(_5739_),
    .B(_5748_),
    .Y(_5749_)
);

NAND2X1 _15218_ (
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .B(_5424_),
    .Y(_5750_)
);

INVX1 _15219_ (
    .A(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_5751_)
);

OAI22X1 _15220_ (
    .A(_4219_),
    .B(_5433__bF$buf3),
    .C(_5436__bF$buf3),
    .D(_5751_),
    .Y(_5752_)
);

AOI21X1 _15221_ (
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .B(_5429_),
    .C(_5752_),
    .Y(_5753_)
);

INVX1 _15222_ (
    .A(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_5754_)
);

INVX1 _15223_ (
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_5755_)
);

OAI22X1 _15224_ (
    .A(_5443_),
    .B(_5755_),
    .C(_5754_),
    .D(_5447_),
    .Y(_5756_)
);

OAI22X1 _15225_ (
    .A(_4243_),
    .B(_5449_),
    .C(_5450_),
    .D(_4242_),
    .Y(_5757_)
);

NOR2X1 _15226_ (
    .A(_5757_),
    .B(_5756_),
    .Y(_5758_)
);

NAND3X1 _15227_ (
    .A(_5753_),
    .B(_5750_),
    .C(_5758_),
    .Y(_5759_)
);

NAND3X1 _15228_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [6]),
    .C(_5509_),
    .Y(_5760_)
);

INVX1 _15229_ (
    .A(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_5761_)
);

OAI22X1 _15230_ (
    .A(_4232_),
    .B(_5506__bF$buf1),
    .C(_5761_),
    .D(_5511__bF$buf3),
    .Y(_5762_)
);

INVX1 _15231_ (
    .A(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_5763_)
);

OAI22X1 _15232_ (
    .A(_5514__bF$buf3),
    .B(_4228_),
    .C(_5763_),
    .D(_5513__bF$buf3),
    .Y(_5764_)
);

NOR2X1 _15233_ (
    .A(_5764_),
    .B(_5762_),
    .Y(_5765_)
);

OAI22X1 _15234_ (
    .A(_5518__bF$buf3),
    .B(_4208_),
    .C(_4220_),
    .D(_5517__bF$buf3),
    .Y(_5766_)
);

INVX1 _15235_ (
    .A(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_5767_)
);

OAI22X1 _15236_ (
    .A(_5767_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_4211_),
    .Y(_5768_)
);

NOR2X1 _15237_ (
    .A(_5766_),
    .B(_5768_),
    .Y(_5769_)
);

NAND3X1 _15238_ (
    .A(_5765_),
    .B(_5769_),
    .C(_5760_),
    .Y(_5770_)
);

NOR2X1 _15239_ (
    .A(_5759_),
    .B(_5770_),
    .Y(_5771_)
);

AOI21X1 _15240_ (
    .A(_5771_),
    .B(_5749_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [6])
);

NAND2X1 _15241_ (
    .A(\datapath_1.regfile_1.regOut[20] [7]),
    .B(_5424_),
    .Y(_5772_)
);

INVX1 _15242_ (
    .A(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_5773_)
);

OAI22X1 _15243_ (
    .A(_4287_),
    .B(_5433__bF$buf2),
    .C(_5436__bF$buf2),
    .D(_5773_),
    .Y(_5774_)
);

AOI21X1 _15244_ (
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .B(_5429_),
    .C(_5774_),
    .Y(_5775_)
);

INVX1 _15245_ (
    .A(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_5776_)
);

INVX1 _15246_ (
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_5777_)
);

OAI22X1 _15247_ (
    .A(_5443_),
    .B(_5777_),
    .C(_5776_),
    .D(_5447_),
    .Y(_5778_)
);

OAI22X1 _15248_ (
    .A(_4278_),
    .B(_5449_),
    .C(_5450_),
    .D(_4277_),
    .Y(_5779_)
);

NOR2X1 _15249_ (
    .A(_5779_),
    .B(_5778_),
    .Y(_5780_)
);

NAND3X1 _15250_ (
    .A(_5775_),
    .B(_5772_),
    .C(_5780_),
    .Y(_5781_)
);

AOI22X1 _15251_ (
    .A(\datapath_1.regfile_1.regOut[4] [7]),
    .B(_5457__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[1] [7]),
    .D(_5455__bF$buf2),
    .Y(_5782_)
);

AOI22X1 _15252_ (
    .A(_5460__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [7]),
    .C(_5462__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_5783_)
);

INVX1 _15253_ (
    .A(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_5784_)
);

OAI22X1 _15254_ (
    .A(_5784_),
    .B(_5465__bF$buf2),
    .C(_5466__bF$buf2),
    .D(_4267_),
    .Y(_5785_)
);

OAI22X1 _15255_ (
    .A(_4257_),
    .B(_5471__bF$buf2),
    .C(_4266_),
    .D(_5472__bF$buf2),
    .Y(_5786_)
);

NOR2X1 _15256_ (
    .A(_5785_),
    .B(_5786_),
    .Y(_5787_)
);

NAND3X1 _15257_ (
    .A(_5783_),
    .B(_5782_),
    .C(_5787_),
    .Y(_5788_)
);

NOR2X1 _15258_ (
    .A(_5781_),
    .B(_5788_),
    .Y(_5789_)
);

AOI22X1 _15259_ (
    .A(_5641_),
    .B(\datapath_1.regfile_1.regOut[29] [7]),
    .C(\datapath_1.regfile_1.regOut[28] [7]),
    .D(_5482__bF$buf2),
    .Y(_5790_)
);

AOI22X1 _15260_ (
    .A(_5642_),
    .B(\datapath_1.regfile_1.regOut[31] [7]),
    .C(\datapath_1.regfile_1.regOut[30] [7]),
    .D(_5489_),
    .Y(_5791_)
);

INVX1 _15261_ (
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_5792_)
);

OAI22X1 _15262_ (
    .A(_5792_),
    .B(_5484__bF$buf2),
    .C(_5485__bF$buf2),
    .D(_4263_),
    .Y(_5793_)
);

AOI21X1 _15263_ (
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .B(_5478__bF$buf1),
    .C(_5793_),
    .Y(_5794_)
);

NAND3X1 _15264_ (
    .A(_5791_),
    .B(_5790_),
    .C(_5794_),
    .Y(_5795_)
);

NAND3X1 _15265_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [7]),
    .C(_5509_),
    .Y(_5796_)
);

OAI22X1 _15266_ (
    .A(_4275_),
    .B(_5506__bF$buf0),
    .C(_4274_),
    .D(_5511__bF$buf2),
    .Y(_5797_)
);

INVX1 _15267_ (
    .A(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_5798_)
);

INVX1 _15268_ (
    .A(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_5799_)
);

OAI22X1 _15269_ (
    .A(_5514__bF$buf2),
    .B(_5798_),
    .C(_5799_),
    .D(_5513__bF$buf2),
    .Y(_5800_)
);

NOR2X1 _15270_ (
    .A(_5800_),
    .B(_5797_),
    .Y(_5801_)
);

OAI22X1 _15271_ (
    .A(_5518__bF$buf2),
    .B(_4253_),
    .C(_4254_),
    .D(_5517__bF$buf2),
    .Y(_5802_)
);

OAI22X1 _15272_ (
    .A(_4284_),
    .B(_5520__bF$buf2),
    .C(_5521__bF$buf2),
    .D(_4288_),
    .Y(_5803_)
);

NOR2X1 _15273_ (
    .A(_5802_),
    .B(_5803_),
    .Y(_5804_)
);

NAND3X1 _15274_ (
    .A(_5801_),
    .B(_5804_),
    .C(_5796_),
    .Y(_5805_)
);

NOR2X1 _15275_ (
    .A(_5795_),
    .B(_5805_),
    .Y(_5806_)
);

AOI21X1 _15276_ (
    .A(_5806_),
    .B(_5789_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [7])
);

AOI22X1 _15277_ (
    .A(_5563__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [8]),
    .C(_5565__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_5807_)
);

OAI22X1 _15278_ (
    .A(_4322_),
    .B(_5433__bF$buf1),
    .C(_5436__bF$buf1),
    .D(_4331_),
    .Y(_5808_)
);

AOI21X1 _15279_ (
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .B(_5429_),
    .C(_5808_),
    .Y(_5809_)
);

AOI22X1 _15280_ (
    .A(_5424_),
    .B(\datapath_1.regfile_1.regOut[20] [8]),
    .C(\datapath_1.regfile_1.regOut[24] [8]),
    .D(_5561__bF$buf3),
    .Y(_5810_)
);

NAND3X1 _15281_ (
    .A(_5810_),
    .B(_5807_),
    .C(_5809_),
    .Y(_5811_)
);

AOI22X1 _15282_ (
    .A(\datapath_1.regfile_1.regOut[4] [8]),
    .B(_5457__bF$buf1),
    .C(\datapath_1.regfile_1.regOut[1] [8]),
    .D(_5455__bF$buf1),
    .Y(_5812_)
);

AOI22X1 _15283_ (
    .A(_5460__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [8]),
    .C(_5462__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_5813_)
);

INVX1 _15284_ (
    .A(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_5814_)
);

OAI22X1 _15285_ (
    .A(_4339_),
    .B(_5465__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_5814_),
    .Y(_5815_)
);

OAI22X1 _15286_ (
    .A(_4305_),
    .B(_5471__bF$buf1),
    .C(_4313_),
    .D(_5472__bF$buf1),
    .Y(_5816_)
);

NOR2X1 _15287_ (
    .A(_5815_),
    .B(_5816_),
    .Y(_5817_)
);

NAND3X1 _15288_ (
    .A(_5813_),
    .B(_5812_),
    .C(_5817_),
    .Y(_5818_)
);

NOR2X1 _15289_ (
    .A(_5811_),
    .B(_5818_),
    .Y(_5819_)
);

NAND2X1 _15290_ (
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .B(_5560__bF$buf3),
    .Y(_5820_)
);

NAND3X1 _15291_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(\datapath_1.regfile_1.regOut[31] [8]),
    .C(_5470_),
    .Y(_5821_)
);

OAI21X1 _15292_ (
    .A(_4334_),
    .B(_5492__bF$buf4),
    .C(_5821_),
    .Y(_5822_)
);

OAI22X1 _15293_ (
    .A(_4300_),
    .B(_5481_),
    .C(_4325_),
    .D(_5488__bF$buf3),
    .Y(_5823_)
);

NOR2X1 _15294_ (
    .A(_5822_),
    .B(_5823_),
    .Y(_5824_)
);

INVX1 _15295_ (
    .A(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_5825_)
);

INVX1 _15296_ (
    .A(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_5826_)
);

OAI22X1 _15297_ (
    .A(_5826_),
    .B(_5484__bF$buf1),
    .C(_5485__bF$buf1),
    .D(_5825_),
    .Y(_5827_)
);

AOI21X1 _15298_ (
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .B(_5478__bF$buf0),
    .C(_5827_),
    .Y(_5828_)
);

NAND3X1 _15299_ (
    .A(_5820_),
    .B(_5824_),
    .C(_5828_),
    .Y(_5829_)
);

NAND3X1 _15300_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [8]),
    .C(_5509_),
    .Y(_5830_)
);

OAI22X1 _15301_ (
    .A(_4293_),
    .B(_5506__bF$buf4),
    .C(_4309_),
    .D(_5511__bF$buf1),
    .Y(_5831_)
);

INVX1 _15302_ (
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_5832_)
);

INVX1 _15303_ (
    .A(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_5833_)
);

OAI22X1 _15304_ (
    .A(_5514__bF$buf1),
    .B(_5832_),
    .C(_5833_),
    .D(_5513__bF$buf1),
    .Y(_5834_)
);

NOR2X1 _15305_ (
    .A(_5834_),
    .B(_5831_),
    .Y(_5835_)
);

OAI22X1 _15306_ (
    .A(_5518__bF$buf1),
    .B(_4297_),
    .C(_4323_),
    .D(_5517__bF$buf1),
    .Y(_5836_)
);

INVX1 _15307_ (
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_5837_)
);

OAI22X1 _15308_ (
    .A(_5837_),
    .B(_5520__bF$buf1),
    .C(_5521__bF$buf1),
    .D(_4318_),
    .Y(_5838_)
);

NOR2X1 _15309_ (
    .A(_5836_),
    .B(_5838_),
    .Y(_5839_)
);

NAND3X1 _15310_ (
    .A(_5835_),
    .B(_5839_),
    .C(_5830_),
    .Y(_5840_)
);

NOR2X1 _15311_ (
    .A(_5829_),
    .B(_5840_),
    .Y(_5841_)
);

AOI21X1 _15312_ (
    .A(_5841_),
    .B(_5819_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [8])
);

NAND2X1 _15313_ (
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .B(_5429_),
    .Y(_5842_)
);

INVX1 _15314_ (
    .A(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_5843_)
);

INVX1 _15315_ (
    .A(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_5844_)
);

OAI22X1 _15316_ (
    .A(_5844_),
    .B(_5433__bF$buf0),
    .C(_5436__bF$buf0),
    .D(_5843_),
    .Y(_5845_)
);

AOI21X1 _15317_ (
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .B(_5424_),
    .C(_5845_),
    .Y(_5846_)
);

INVX1 _15318_ (
    .A(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_5847_)
);

INVX1 _15319_ (
    .A(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_5848_)
);

OAI22X1 _15320_ (
    .A(_5443_),
    .B(_5848_),
    .C(_5847_),
    .D(_5447_),
    .Y(_5849_)
);

OAI22X1 _15321_ (
    .A(_4372_),
    .B(_5449_),
    .C(_5450_),
    .D(_4371_),
    .Y(_5850_)
);

NOR2X1 _15322_ (
    .A(_5850_),
    .B(_5849_),
    .Y(_5851_)
);

NAND3X1 _15323_ (
    .A(_5846_),
    .B(_5842_),
    .C(_5851_),
    .Y(_5852_)
);

AOI22X1 _15324_ (
    .A(\datapath_1.regfile_1.regOut[4] [9]),
    .B(_5457__bF$buf0),
    .C(\datapath_1.regfile_1.regOut[1] [9]),
    .D(_5455__bF$buf0),
    .Y(_5853_)
);

AOI22X1 _15325_ (
    .A(_5460__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [9]),
    .C(_5462__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_5854_)
);

INVX1 _15326_ (
    .A(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_5855_)
);

OAI22X1 _15327_ (
    .A(_5855_),
    .B(_5465__bF$buf0),
    .C(_5466__bF$buf0),
    .D(_4364_),
    .Y(_5856_)
);

OAI22X1 _15328_ (
    .A(_4351_),
    .B(_5471__bF$buf0),
    .C(_4363_),
    .D(_5472__bF$buf0),
    .Y(_5857_)
);

NOR2X1 _15329_ (
    .A(_5856_),
    .B(_5857_),
    .Y(_5858_)
);

NAND3X1 _15330_ (
    .A(_5854_),
    .B(_5853_),
    .C(_5858_),
    .Y(_5859_)
);

NOR2X1 _15331_ (
    .A(_5852_),
    .B(_5859_),
    .Y(_5860_)
);

NAND2X1 _15332_ (
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .B(_5478__bF$buf3),
    .Y(_5861_)
);

INVX1 _15333_ (
    .A(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_5862_)
);

OAI22X1 _15334_ (
    .A(_4360_),
    .B(_5484__bF$buf0),
    .C(_5485__bF$buf0),
    .D(_5862_),
    .Y(_5863_)
);

AOI21X1 _15335_ (
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .B(_5482__bF$buf1),
    .C(_5863_),
    .Y(_5864_)
);

INVX1 _15336_ (
    .A(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_5865_)
);

INVX1 _15337_ (
    .A(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_5866_)
);

OAI22X1 _15338_ (
    .A(_5492__bF$buf3),
    .B(_5866_),
    .C(_5865_),
    .D(_5493__bF$buf3),
    .Y(_5867_)
);

AOI21X1 _15339_ (
    .A(\datapath_1.regfile_1.regOut[30] [9]),
    .B(_5489_),
    .C(_5867_),
    .Y(_5868_)
);

NAND3X1 _15340_ (
    .A(_5861_),
    .B(_5868_),
    .C(_5864_),
    .Y(_5869_)
);

NAND3X1 _15341_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [9]),
    .C(_5509_),
    .Y(_5870_)
);

INVX1 _15342_ (
    .A(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_5871_)
);

OAI22X1 _15343_ (
    .A(_4354_),
    .B(_5506__bF$buf3),
    .C(_5871_),
    .D(_5511__bF$buf0),
    .Y(_5872_)
);

OAI22X1 _15344_ (
    .A(_5514__bF$buf0),
    .B(_4361_),
    .C(_4374_),
    .D(_5513__bF$buf0),
    .Y(_5873_)
);

NOR2X1 _15345_ (
    .A(_5873_),
    .B(_5872_),
    .Y(_5874_)
);

OAI22X1 _15346_ (
    .A(_5518__bF$buf0),
    .B(_4384_),
    .C(_4353_),
    .D(_5517__bF$buf0),
    .Y(_5875_)
);

OAI22X1 _15347_ (
    .A(_4382_),
    .B(_5520__bF$buf0),
    .C(_5521__bF$buf0),
    .D(_4381_),
    .Y(_5876_)
);

NOR2X1 _15348_ (
    .A(_5875_),
    .B(_5876_),
    .Y(_5877_)
);

NAND3X1 _15349_ (
    .A(_5874_),
    .B(_5877_),
    .C(_5870_),
    .Y(_5878_)
);

NOR2X1 _15350_ (
    .A(_5869_),
    .B(_5878_),
    .Y(_5879_)
);

AOI21X1 _15351_ (
    .A(_5879_),
    .B(_5860_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [9])
);

NAND2X1 _15352_ (
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .B(_5429_),
    .Y(_5880_)
);

INVX1 _15353_ (
    .A(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_5881_)
);

OAI22X1 _15354_ (
    .A(_5881_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_4406_),
    .Y(_5882_)
);

AOI21X1 _15355_ (
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .B(_5424_),
    .C(_5882_),
    .Y(_5883_)
);

INVX1 _15356_ (
    .A(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_5884_)
);

OAI22X1 _15357_ (
    .A(_5443_),
    .B(_5884_),
    .C(_4405_),
    .D(_5447_),
    .Y(_5885_)
);

INVX1 _15358_ (
    .A(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_5886_)
);

INVX1 _15359_ (
    .A(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_5887_)
);

OAI22X1 _15360_ (
    .A(_5887_),
    .B(_5449_),
    .C(_5450_),
    .D(_5886_),
    .Y(_5888_)
);

NOR2X1 _15361_ (
    .A(_5888_),
    .B(_5885_),
    .Y(_5889_)
);

NAND3X1 _15362_ (
    .A(_5883_),
    .B(_5880_),
    .C(_5889_),
    .Y(_5890_)
);

AOI22X1 _15363_ (
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [10]),
    .D(_5455__bF$buf4),
    .Y(_5891_)
);

AOI22X1 _15364_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [10]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_5892_)
);

OAI22X1 _15365_ (
    .A(_4419_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_4422_),
    .Y(_5893_)
);

OAI22X1 _15366_ (
    .A(_4418_),
    .B(_5471__bF$buf4),
    .C(_4421_),
    .D(_5472__bF$buf4),
    .Y(_5894_)
);

NOR2X1 _15367_ (
    .A(_5893_),
    .B(_5894_),
    .Y(_5895_)
);

NAND3X1 _15368_ (
    .A(_5892_),
    .B(_5891_),
    .C(_5895_),
    .Y(_5896_)
);

NOR2X1 _15369_ (
    .A(_5890_),
    .B(_5896_),
    .Y(_5897_)
);

NAND2X1 _15370_ (
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .B(_5478__bF$buf2),
    .Y(_5898_)
);

OAI22X1 _15371_ (
    .A(_4412_),
    .B(_5484__bF$buf4),
    .C(_5485__bF$buf4),
    .D(_4394_),
    .Y(_5899_)
);

AOI21X1 _15372_ (
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .B(_5482__bF$buf0),
    .C(_5899_),
    .Y(_5900_)
);

OAI22X1 _15373_ (
    .A(_5492__bF$buf2),
    .B(_4402_),
    .C(_4438_),
    .D(_5493__bF$buf2),
    .Y(_5901_)
);

AOI21X1 _15374_ (
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .B(_5489_),
    .C(_5901_),
    .Y(_5902_)
);

NAND3X1 _15375_ (
    .A(_5898_),
    .B(_5902_),
    .C(_5900_),
    .Y(_5903_)
);

NAND3X1 _15376_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [10]),
    .C(_5509_),
    .Y(_5904_)
);

OAI22X1 _15377_ (
    .A(_4391_),
    .B(_5506__bF$buf2),
    .C(_4426_),
    .D(_5511__bF$buf4),
    .Y(_5905_)
);

INVX1 _15378_ (
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_5906_)
);

INVX1 _15379_ (
    .A(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_5907_)
);

OAI22X1 _15380_ (
    .A(_5514__bF$buf4),
    .B(_5906_),
    .C(_5907_),
    .D(_5513__bF$buf4),
    .Y(_5908_)
);

NOR2X1 _15381_ (
    .A(_5908_),
    .B(_5905_),
    .Y(_5909_)
);

OAI22X1 _15382_ (
    .A(_5518__bF$buf4),
    .B(_4428_),
    .C(_4390_),
    .D(_5517__bF$buf4),
    .Y(_5910_)
);

OAI22X1 _15383_ (
    .A(_4436_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_4435_),
    .Y(_5911_)
);

NOR2X1 _15384_ (
    .A(_5910_),
    .B(_5911_),
    .Y(_5912_)
);

NAND3X1 _15385_ (
    .A(_5909_),
    .B(_5912_),
    .C(_5904_),
    .Y(_5913_)
);

NOR2X1 _15386_ (
    .A(_5903_),
    .B(_5913_),
    .Y(_5914_)
);

AOI21X1 _15387_ (
    .A(_5914_),
    .B(_5897_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [10])
);

NOR2X1 _15388_ (
    .A(_4475_),
    .B(_5428__bF$buf2),
    .Y(_5915_)
);

INVX1 _15389_ (
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_5916_)
);

NOR3X1 _15390_ (
    .A(_5421__bF$buf3),
    .B(_5916_),
    .C(_5423__bF$buf2),
    .Y(_5917_)
);

INVX1 _15391_ (
    .A(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_5918_)
);

INVX1 _15392_ (
    .A(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_5919_)
);

OAI22X1 _15393_ (
    .A(_5919_),
    .B(_5433__bF$buf3),
    .C(_5436__bF$buf3),
    .D(_5918_),
    .Y(_5920_)
);

NOR3X1 _15394_ (
    .A(_5917_),
    .B(_5915_),
    .C(_5920_),
    .Y(_5921_)
);

INVX1 _15395_ (
    .A(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_5922_)
);

OAI22X1 _15396_ (
    .A(_4482_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_5922_),
    .Y(_5923_)
);

AOI21X1 _15397_ (
    .A(\datapath_1.regfile_1.regOut[28] [11]),
    .B(_5482__bF$buf3),
    .C(_5923_),
    .Y(_5924_)
);

INVX1 _15398_ (
    .A(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_5925_)
);

INVX1 _15399_ (
    .A(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_5926_)
);

OAI22X1 _15400_ (
    .A(_5492__bF$buf1),
    .B(_5926_),
    .C(_5925_),
    .D(_5493__bF$buf1),
    .Y(_5927_)
);

INVX1 _15401_ (
    .A(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_5928_)
);

INVX1 _15402_ (
    .A(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_5929_)
);

OAI22X1 _15403_ (
    .A(_5929_),
    .B(_5477_),
    .C(_5488__bF$buf2),
    .D(_5928_),
    .Y(_5930_)
);

NOR2X1 _15404_ (
    .A(_5930_),
    .B(_5927_),
    .Y(_5931_)
);

NAND3X1 _15405_ (
    .A(_5924_),
    .B(_5931_),
    .C(_5921_),
    .Y(_5932_)
);

AOI22X1 _15406_ (
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [11]),
    .D(_5455__bF$buf3),
    .Y(_5933_)
);

AOI22X1 _15407_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [11]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_5934_)
);

INVX1 _15408_ (
    .A(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_5935_)
);

OAI22X1 _15409_ (
    .A(_5935_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_4448_),
    .Y(_5936_)
);

OAI22X1 _15410_ (
    .A(_4447_),
    .B(_5471__bF$buf3),
    .C(_4463_),
    .D(_5472__bF$buf3),
    .Y(_5937_)
);

NOR2X1 _15411_ (
    .A(_5936_),
    .B(_5937_),
    .Y(_5938_)
);

NAND3X1 _15412_ (
    .A(_5934_),
    .B(_5933_),
    .C(_5938_),
    .Y(_5939_)
);

NOR2X1 _15413_ (
    .A(_5939_),
    .B(_5932_),
    .Y(_5940_)
);

INVX1 _15414_ (
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_5941_)
);

NOR3X1 _15415_ (
    .A(_5941_),
    .B(_5558__bF$buf3),
    .C(_5555__bF$buf3),
    .Y(_5942_)
);

NAND2X1 _15416_ (
    .A(\datapath_1.regfile_1.regOut[22] [11]),
    .B(_5563__bF$buf2),
    .Y(_5943_)
);

NAND2X1 _15417_ (
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .B(_5565__bF$buf2),
    .Y(_5944_)
);

AOI22X1 _15418_ (
    .A(_5560__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [11]),
    .C(\datapath_1.regfile_1.regOut[24] [11]),
    .D(_5561__bF$buf2),
    .Y(_5945_)
);

NAND3X1 _15419_ (
    .A(_5943_),
    .B(_5945_),
    .C(_5944_),
    .Y(_5946_)
);

OAI22X1 _15420_ (
    .A(_4460_),
    .B(_5506__bF$buf1),
    .C(_4445_),
    .D(_5511__bF$buf3),
    .Y(_5947_)
);

OAI22X1 _15421_ (
    .A(_5514__bF$buf3),
    .B(_4471_),
    .C(_4472_),
    .D(_5513__bF$buf3),
    .Y(_5948_)
);

NOR2X1 _15422_ (
    .A(_5948_),
    .B(_5947_),
    .Y(_5949_)
);

OAI22X1 _15423_ (
    .A(_5518__bF$buf3),
    .B(_4456_),
    .C(_4480_),
    .D(_5517__bF$buf3),
    .Y(_5950_)
);

OAI22X1 _15424_ (
    .A(_4479_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_4483_),
    .Y(_5951_)
);

NOR2X1 _15425_ (
    .A(_5950_),
    .B(_5951_),
    .Y(_5952_)
);

NAND2X1 _15426_ (
    .A(_5949_),
    .B(_5952_),
    .Y(_5953_)
);

NOR3X1 _15427_ (
    .A(_5946_),
    .B(_5942_),
    .C(_5953_),
    .Y(_5954_)
);

AOI21X1 _15428_ (
    .A(_5940_),
    .B(_5954_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [11])
);

NOR2X1 _15429_ (
    .A(_4516_),
    .B(_5428__bF$buf1),
    .Y(_5955_)
);

INVX1 _15430_ (
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_5956_)
);

NOR3X1 _15431_ (
    .A(_5421__bF$buf2),
    .B(_5956_),
    .C(_5423__bF$buf1),
    .Y(_5957_)
);

OAI22X1 _15432_ (
    .A(_4519_),
    .B(_5433__bF$buf2),
    .C(_5436__bF$buf2),
    .D(_4515_),
    .Y(_5958_)
);

NOR3X1 _15433_ (
    .A(_5957_),
    .B(_5955_),
    .C(_5958_),
    .Y(_5959_)
);

INVX1 _15434_ (
    .A(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_5960_)
);

OAI22X1 _15435_ (
    .A(_4493_),
    .B(_5484__bF$buf2),
    .C(_5485__bF$buf2),
    .D(_5960_),
    .Y(_5961_)
);

AOI21X1 _15436_ (
    .A(\datapath_1.regfile_1.regOut[27] [12]),
    .B(_5478__bF$buf1),
    .C(_5961_),
    .Y(_5962_)
);

INVX1 _15437_ (
    .A(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_5963_)
);

OAI22X1 _15438_ (
    .A(_5963_),
    .B(_5449_),
    .C(_5450_),
    .D(_4518_),
    .Y(_5964_)
);

INVX1 _15439_ (
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_5965_)
);

INVX1 _15440_ (
    .A(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_5966_)
);

OAI22X1 _15441_ (
    .A(_5443_),
    .B(_5966_),
    .C(_5965_),
    .D(_5447_),
    .Y(_5967_)
);

NOR2X1 _15442_ (
    .A(_5964_),
    .B(_5967_),
    .Y(_5968_)
);

NAND3X1 _15443_ (
    .A(_5962_),
    .B(_5968_),
    .C(_5959_),
    .Y(_5969_)
);

AOI22X1 _15444_ (
    .A(\datapath_1.regfile_1.regOut[4] [12]),
    .B(_5457__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[1] [12]),
    .D(_5455__bF$buf2),
    .Y(_5970_)
);

AOI22X1 _15445_ (
    .A(_5460__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [12]),
    .C(_5462__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_5971_)
);

INVX1 _15446_ (
    .A(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_5972_)
);

OAI22X1 _15447_ (
    .A(_4531_),
    .B(_5465__bF$buf2),
    .C(_5466__bF$buf2),
    .D(_5972_),
    .Y(_5973_)
);

OAI22X1 _15448_ (
    .A(_4528_),
    .B(_5471__bF$buf2),
    .C(_4527_),
    .D(_5472__bF$buf2),
    .Y(_5974_)
);

NOR2X1 _15449_ (
    .A(_5973_),
    .B(_5974_),
    .Y(_5975_)
);

NAND3X1 _15450_ (
    .A(_5971_),
    .B(_5970_),
    .C(_5975_),
    .Y(_5976_)
);

NOR2X1 _15451_ (
    .A(_5976_),
    .B(_5969_),
    .Y(_5977_)
);

INVX1 _15452_ (
    .A(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_5978_)
);

NOR3X1 _15453_ (
    .A(_5978_),
    .B(_5558__bF$buf2),
    .C(_5555__bF$buf2),
    .Y(_5979_)
);

AOI22X1 _15454_ (
    .A(_5641_),
    .B(\datapath_1.regfile_1.regOut[29] [12]),
    .C(\datapath_1.regfile_1.regOut[28] [12]),
    .D(_5482__bF$buf2),
    .Y(_5980_)
);

AOI22X1 _15455_ (
    .A(_5642_),
    .B(\datapath_1.regfile_1.regOut[31] [12]),
    .C(\datapath_1.regfile_1.regOut[30] [12]),
    .D(_5489_),
    .Y(_5981_)
);

NAND2X1 _15456_ (
    .A(_5980_),
    .B(_5981_),
    .Y(_5982_)
);

INVX1 _15457_ (
    .A(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_5983_)
);

OAI22X1 _15458_ (
    .A(_4508_),
    .B(_5506__bF$buf0),
    .C(_5983_),
    .D(_5511__bF$buf2),
    .Y(_5984_)
);

INVX1 _15459_ (
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_5985_)
);

INVX1 _15460_ (
    .A(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_5986_)
);

OAI22X1 _15461_ (
    .A(_5514__bF$buf2),
    .B(_5985_),
    .C(_5986_),
    .D(_5513__bF$buf2),
    .Y(_5987_)
);

NOR2X1 _15462_ (
    .A(_5987_),
    .B(_5984_),
    .Y(_5988_)
);

OAI22X1 _15463_ (
    .A(_5518__bF$buf2),
    .B(_4500_),
    .C(_4524_),
    .D(_5517__bF$buf2),
    .Y(_5989_)
);

OAI22X1 _15464_ (
    .A(_4504_),
    .B(_5520__bF$buf2),
    .C(_5521__bF$buf2),
    .D(_4494_),
    .Y(_5990_)
);

NOR2X1 _15465_ (
    .A(_5989_),
    .B(_5990_),
    .Y(_5991_)
);

NAND2X1 _15466_ (
    .A(_5988_),
    .B(_5991_),
    .Y(_5992_)
);

NOR3X1 _15467_ (
    .A(_5982_),
    .B(_5979_),
    .C(_5992_),
    .Y(_5993_)
);

AOI21X1 _15468_ (
    .A(_5977_),
    .B(_5993_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [12])
);

NOR2X1 _15469_ (
    .A(_4566_),
    .B(_5428__bF$buf0),
    .Y(_5994_)
);

INVX1 _15470_ (
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_5995_)
);

NOR3X1 _15471_ (
    .A(_5421__bF$buf1),
    .B(_5995_),
    .C(_5423__bF$buf0),
    .Y(_5996_)
);

INVX1 _15472_ (
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_5997_)
);

INVX1 _15473_ (
    .A(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_5998_)
);

OAI22X1 _15474_ (
    .A(_5998_),
    .B(_5433__bF$buf1),
    .C(_5436__bF$buf1),
    .D(_5997_),
    .Y(_5999_)
);

NOR3X1 _15475_ (
    .A(_5996_),
    .B(_5994_),
    .C(_5999_),
    .Y(_6000_)
);

INVX1 _15476_ (
    .A(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_6001_)
);

INVX1 _15477_ (
    .A(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_6002_)
);

OAI22X1 _15478_ (
    .A(_6002_),
    .B(_5484__bF$buf1),
    .C(_5485__bF$buf1),
    .D(_6001_),
    .Y(_6003_)
);

AOI21X1 _15479_ (
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .B(_5482__bF$buf1),
    .C(_6003_),
    .Y(_6004_)
);

INVX1 _15480_ (
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_6005_)
);

OAI22X1 _15481_ (
    .A(_5492__bF$buf0),
    .B(_4551_),
    .C(_6005_),
    .D(_5493__bF$buf0),
    .Y(_6006_)
);

INVX1 _15482_ (
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_6007_)
);

OAI22X1 _15483_ (
    .A(_4539_),
    .B(_5477_),
    .C(_5488__bF$buf1),
    .D(_6007_),
    .Y(_6008_)
);

NOR2X1 _15484_ (
    .A(_6008_),
    .B(_6006_),
    .Y(_6009_)
);

NAND3X1 _15485_ (
    .A(_6004_),
    .B(_6009_),
    .C(_6000_),
    .Y(_6010_)
);

AOI22X1 _15486_ (
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .B(_5457__bF$buf1),
    .C(\datapath_1.regfile_1.regOut[1] [13]),
    .D(_5455__bF$buf1),
    .Y(_6011_)
);

AOI22X1 _15487_ (
    .A(_5460__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [13]),
    .C(_5462__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_6012_)
);

INVX1 _15488_ (
    .A(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_6013_)
);

INVX1 _15489_ (
    .A(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_6014_)
);

OAI22X1 _15490_ (
    .A(_6014_),
    .B(_5465__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_6013_),
    .Y(_6015_)
);

INVX1 _15491_ (
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_6016_)
);

OAI22X1 _15492_ (
    .A(_6016_),
    .B(_5471__bF$buf1),
    .C(_4567_),
    .D(_5472__bF$buf1),
    .Y(_6017_)
);

NOR2X1 _15493_ (
    .A(_6015_),
    .B(_6017_),
    .Y(_6018_)
);

NAND3X1 _15494_ (
    .A(_6012_),
    .B(_6011_),
    .C(_6018_),
    .Y(_6019_)
);

NOR2X1 _15495_ (
    .A(_6019_),
    .B(_6010_),
    .Y(_6020_)
);

NOR3X1 _15496_ (
    .A(_4563_),
    .B(_5558__bF$buf1),
    .C(_5555__bF$buf1),
    .Y(_6021_)
);

NAND2X1 _15497_ (
    .A(\datapath_1.regfile_1.regOut[21] [13]),
    .B(_5565__bF$buf1),
    .Y(_6022_)
);

NAND2X1 _15498_ (
    .A(\datapath_1.regfile_1.regOut[22] [13]),
    .B(_5563__bF$buf1),
    .Y(_6023_)
);

AOI22X1 _15499_ (
    .A(_5560__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [13]),
    .C(\datapath_1.regfile_1.regOut[24] [13]),
    .D(_5561__bF$buf1),
    .Y(_6024_)
);

NAND3X1 _15500_ (
    .A(_6022_),
    .B(_6024_),
    .C(_6023_),
    .Y(_6025_)
);

OAI22X1 _15501_ (
    .A(_4549_),
    .B(_5506__bF$buf4),
    .C(_4540_),
    .D(_5511__bF$buf1),
    .Y(_6026_)
);

INVX1 _15502_ (
    .A(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_6027_)
);

OAI22X1 _15503_ (
    .A(_5514__bF$buf1),
    .B(_4564_),
    .C(_6027_),
    .D(_5513__bF$buf1),
    .Y(_6028_)
);

NOR2X1 _15504_ (
    .A(_6028_),
    .B(_6026_),
    .Y(_6029_)
);

OAI22X1 _15505_ (
    .A(_5518__bF$buf1),
    .B(_4537_),
    .C(_4552_),
    .D(_5517__bF$buf1),
    .Y(_6030_)
);

INVX1 _15506_ (
    .A(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_6031_)
);

OAI22X1 _15507_ (
    .A(_6031_),
    .B(_5520__bF$buf1),
    .C(_5521__bF$buf1),
    .D(_4536_),
    .Y(_6032_)
);

NOR2X1 _15508_ (
    .A(_6030_),
    .B(_6032_),
    .Y(_6033_)
);

NAND2X1 _15509_ (
    .A(_6029_),
    .B(_6033_),
    .Y(_6034_)
);

NOR3X1 _15510_ (
    .A(_6025_),
    .B(_6021_),
    .C(_6034_),
    .Y(_6035_)
);

AOI21X1 _15511_ (
    .A(_6020_),
    .B(_6035_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [13])
);

NOR2X1 _15512_ (
    .A(_4583_),
    .B(_5428__bF$buf3),
    .Y(_6036_)
);

INVX1 _15513_ (
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_6037_)
);

NOR3X1 _15514_ (
    .A(_5421__bF$buf0),
    .B(_6037_),
    .C(_5423__bF$buf3),
    .Y(_6038_)
);

INVX1 _15515_ (
    .A(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_6039_)
);

OAI22X1 _15516_ (
    .A(_4614_),
    .B(_5433__bF$buf0),
    .C(_5436__bF$buf0),
    .D(_6039_),
    .Y(_6040_)
);

NOR3X1 _15517_ (
    .A(_6038_),
    .B(_6036_),
    .C(_6040_),
    .Y(_6041_)
);

INVX1 _15518_ (
    .A(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_6042_)
);

INVX1 _15519_ (
    .A(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_6043_)
);

OAI22X1 _15520_ (
    .A(_5492__bF$buf4),
    .B(_6043_),
    .C(_6042_),
    .D(_5493__bF$buf3),
    .Y(_6044_)
);

INVX1 _15521_ (
    .A(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_6045_)
);

OAI22X1 _15522_ (
    .A(_4602_),
    .B(_5481_),
    .C(_6045_),
    .D(_5488__bF$buf0),
    .Y(_6046_)
);

NOR2X1 _15523_ (
    .A(_6046_),
    .B(_6044_),
    .Y(_6047_)
);

INVX1 _15524_ (
    .A(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_6048_)
);

INVX1 _15525_ (
    .A(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_6049_)
);

OAI22X1 _15526_ (
    .A(_6049_),
    .B(_5484__bF$buf0),
    .C(_5485__bF$buf0),
    .D(_6048_),
    .Y(_6050_)
);

AOI21X1 _15527_ (
    .A(\datapath_1.regfile_1.regOut[27] [14]),
    .B(_5478__bF$buf0),
    .C(_6050_),
    .Y(_6051_)
);

NAND3X1 _15528_ (
    .A(_6047_),
    .B(_6051_),
    .C(_6041_),
    .Y(_6052_)
);

AOI22X1 _15529_ (
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .B(_5457__bF$buf0),
    .C(\datapath_1.regfile_1.regOut[1] [14]),
    .D(_5455__bF$buf0),
    .Y(_6053_)
);

AOI22X1 _15530_ (
    .A(_5460__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [14]),
    .C(_5462__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_6054_)
);

INVX1 _15531_ (
    .A(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_6055_)
);

OAI22X1 _15532_ (
    .A(_6055_),
    .B(_5465__bF$buf0),
    .C(_5466__bF$buf0),
    .D(_4594_),
    .Y(_6056_)
);

OAI22X1 _15533_ (
    .A(_4593_),
    .B(_5471__bF$buf0),
    .C(_4584_),
    .D(_5472__bF$buf0),
    .Y(_6057_)
);

NOR2X1 _15534_ (
    .A(_6056_),
    .B(_6057_),
    .Y(_6058_)
);

NAND3X1 _15535_ (
    .A(_6054_),
    .B(_6053_),
    .C(_6058_),
    .Y(_6059_)
);

NOR2X1 _15536_ (
    .A(_6059_),
    .B(_6052_),
    .Y(_6060_)
);

INVX1 _15537_ (
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_6061_)
);

NOR3X1 _15538_ (
    .A(_6061_),
    .B(_5558__bF$buf0),
    .C(_5555__bF$buf0),
    .Y(_6062_)
);

NAND2X1 _15539_ (
    .A(\datapath_1.regfile_1.regOut[21] [14]),
    .B(_5565__bF$buf0),
    .Y(_6063_)
);

NAND2X1 _15540_ (
    .A(\datapath_1.regfile_1.regOut[22] [14]),
    .B(_5563__bF$buf0),
    .Y(_6064_)
);

AOI22X1 _15541_ (
    .A(_5560__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [14]),
    .C(\datapath_1.regfile_1.regOut[24] [14]),
    .D(_5561__bF$buf0),
    .Y(_6065_)
);

NAND3X1 _15542_ (
    .A(_6063_),
    .B(_6065_),
    .C(_6064_),
    .Y(_6066_)
);

INVX1 _15543_ (
    .A(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_6067_)
);

OAI22X1 _15544_ (
    .A(_4603_),
    .B(_5506__bF$buf3),
    .C(_6067_),
    .D(_5511__bF$buf0),
    .Y(_6068_)
);

OAI22X1 _15545_ (
    .A(_5514__bF$buf0),
    .B(_4590_),
    .C(_4600_),
    .D(_5513__bF$buf0),
    .Y(_6069_)
);

NOR2X1 _15546_ (
    .A(_6069_),
    .B(_6068_),
    .Y(_6070_)
);

OAI22X1 _15547_ (
    .A(_5518__bF$buf0),
    .B(_4580_),
    .C(_4581_),
    .D(_5517__bF$buf0),
    .Y(_6071_)
);

OAI22X1 _15548_ (
    .A(_4611_),
    .B(_5520__bF$buf0),
    .C(_5521__bF$buf0),
    .D(_4615_),
    .Y(_6072_)
);

NOR2X1 _15549_ (
    .A(_6071_),
    .B(_6072_),
    .Y(_6073_)
);

NAND2X1 _15550_ (
    .A(_6073_),
    .B(_6070_),
    .Y(_6074_)
);

NOR3X1 _15551_ (
    .A(_6066_),
    .B(_6062_),
    .C(_6074_),
    .Y(_6075_)
);

AOI21X1 _15552_ (
    .A(_6060_),
    .B(_6075_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [14])
);

AOI22X1 _15553_ (
    .A(_5563__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[22] [15]),
    .C(_5565__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_6076_)
);

INVX1 _15554_ (
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_6077_)
);

OAI22X1 _15555_ (
    .A(_4623_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_6077_),
    .Y(_6078_)
);

AOI21X1 _15556_ (
    .A(\datapath_1.regfile_1.regOut[20] [15]),
    .B(_5424_),
    .C(_6078_),
    .Y(_6079_)
);

AOI22X1 _15557_ (
    .A(_5429_),
    .B(\datapath_1.regfile_1.regOut[19] [15]),
    .C(\datapath_1.regfile_1.regOut[24] [15]),
    .D(_5561__bF$buf3),
    .Y(_6080_)
);

NAND3X1 _15558_ (
    .A(_6080_),
    .B(_6076_),
    .C(_6079_),
    .Y(_6081_)
);

AOI22X1 _15559_ (
    .A(\datapath_1.regfile_1.regOut[4] [15]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [15]),
    .D(_5455__bF$buf4),
    .Y(_6082_)
);

AOI22X1 _15560_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [15]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_6083_)
);

OAI22X1 _15561_ (
    .A(_4660_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_4642_),
    .Y(_6084_)
);

INVX1 _15562_ (
    .A(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_6085_)
);

OAI22X1 _15563_ (
    .A(_6085_),
    .B(_5471__bF$buf4),
    .C(_4641_),
    .D(_5472__bF$buf4),
    .Y(_6086_)
);

NOR2X1 _15564_ (
    .A(_6084_),
    .B(_6086_),
    .Y(_6087_)
);

NAND3X1 _15565_ (
    .A(_6083_),
    .B(_6082_),
    .C(_6087_),
    .Y(_6088_)
);

NOR2X1 _15566_ (
    .A(_6081_),
    .B(_6088_),
    .Y(_6089_)
);

NAND2X1 _15567_ (
    .A(\datapath_1.regfile_1.regOut[23] [15]),
    .B(_5560__bF$buf3),
    .Y(_6090_)
);

INVX1 _15568_ (
    .A(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_6091_)
);

NAND3X1 _15569_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(\datapath_1.regfile_1.regOut[31] [15]),
    .C(_5470_),
    .Y(_6092_)
);

OAI21X1 _15570_ (
    .A(_6091_),
    .B(_5492__bF$buf3),
    .C(_6092_),
    .Y(_6093_)
);

INVX1 _15571_ (
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_6094_)
);

OAI22X1 _15572_ (
    .A(_4621_),
    .B(_5481_),
    .C(_6094_),
    .D(_5488__bF$buf3),
    .Y(_6095_)
);

NOR2X1 _15573_ (
    .A(_6093_),
    .B(_6095_),
    .Y(_6096_)
);

INVX1 _15574_ (
    .A(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_6097_)
);

OAI22X1 _15575_ (
    .A(_6097_),
    .B(_5484__bF$buf4),
    .C(_5485__bF$buf4),
    .D(_4638_),
    .Y(_6098_)
);

AOI21X1 _15576_ (
    .A(\datapath_1.regfile_1.regOut[27] [15]),
    .B(_5478__bF$buf3),
    .C(_6098_),
    .Y(_6099_)
);

NAND3X1 _15577_ (
    .A(_6090_),
    .B(_6096_),
    .C(_6099_),
    .Y(_6100_)
);

NAND3X1 _15578_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [15]),
    .C(_5509_),
    .Y(_6101_)
);

OAI22X1 _15579_ (
    .A(_4650_),
    .B(_5506__bF$buf2),
    .C(_4649_),
    .D(_5511__bF$buf4),
    .Y(_6102_)
);

INVX1 _15580_ (
    .A(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_6103_)
);

OAI22X1 _15581_ (
    .A(_5514__bF$buf4),
    .B(_6103_),
    .C(_4661_),
    .D(_5513__bF$buf4),
    .Y(_6104_)
);

NOR2X1 _15582_ (
    .A(_6104_),
    .B(_6102_),
    .Y(_6105_)
);

OAI22X1 _15583_ (
    .A(_5518__bF$buf4),
    .B(_4635_),
    .C(_4624_),
    .D(_5517__bF$buf4),
    .Y(_6106_)
);

OAI22X1 _15584_ (
    .A(_4658_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_4657_),
    .Y(_6107_)
);

NOR2X1 _15585_ (
    .A(_6106_),
    .B(_6107_),
    .Y(_6108_)
);

NAND3X1 _15586_ (
    .A(_6105_),
    .B(_6108_),
    .C(_6101_),
    .Y(_6109_)
);

NOR2X1 _15587_ (
    .A(_6100_),
    .B(_6109_),
    .Y(_6110_)
);

AOI21X1 _15588_ (
    .A(_6110_),
    .B(_6089_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [15])
);

AOI22X1 _15589_ (
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [16]),
    .D(_5455__bF$buf3),
    .Y(_6111_)
);

AOI22X1 _15590_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [16]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_6112_)
);

OAI22X1 _15591_ (
    .A(_4705_),
    .B(_5471__bF$buf3),
    .C(_4672_),
    .D(_5472__bF$buf3),
    .Y(_6113_)
);

OAI22X1 _15592_ (
    .A(_4684_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_4669_),
    .Y(_6114_)
);

NOR2X1 _15593_ (
    .A(_6114_),
    .B(_6113_),
    .Y(_6115_)
);

NAND3X1 _15594_ (
    .A(_6112_),
    .B(_6111_),
    .C(_6115_),
    .Y(_6116_)
);

NAND3X1 _15595_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [16]),
    .C(_5509_),
    .Y(_6117_)
);

INVX1 _15596_ (
    .A(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_6118_)
);

OAI22X1 _15597_ (
    .A(_4679_),
    .B(_5506__bF$buf1),
    .C(_6118_),
    .D(_5511__bF$buf3),
    .Y(_6119_)
);

INVX1 _15598_ (
    .A(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_6120_)
);

INVX1 _15599_ (
    .A(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_6121_)
);

OAI22X1 _15600_ (
    .A(_5514__bF$buf3),
    .B(_6120_),
    .C(_6121_),
    .D(_5513__bF$buf3),
    .Y(_6122_)
);

NOR2X1 _15601_ (
    .A(_6122_),
    .B(_6119_),
    .Y(_6123_)
);

OAI22X1 _15602_ (
    .A(_5518__bF$buf3),
    .B(_4668_),
    .C(_4678_),
    .D(_5517__bF$buf3),
    .Y(_6124_)
);

OAI22X1 _15603_ (
    .A(_4675_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_4683_),
    .Y(_6125_)
);

NOR2X1 _15604_ (
    .A(_6124_),
    .B(_6125_),
    .Y(_6126_)
);

NAND3X1 _15605_ (
    .A(_6123_),
    .B(_6126_),
    .C(_6117_),
    .Y(_6127_)
);

NOR2X1 _15606_ (
    .A(_6116_),
    .B(_6127_),
    .Y(_6128_)
);

NAND2X1 _15607_ (
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .B(_5429_),
    .Y(_6129_)
);

INVX1 _15608_ (
    .A(_5436__bF$buf3),
    .Y(_6130_)
);

NOR2X1 _15609_ (
    .A(_4707_),
    .B(_5433__bF$buf3),
    .Y(_6131_)
);

AOI21X1 _15610_ (
    .A(_6130_),
    .B(\datapath_1.regfile_1.regOut[18] [16]),
    .C(_6131_),
    .Y(_6132_)
);

AOI22X1 _15611_ (
    .A(_5424_),
    .B(\datapath_1.regfile_1.regOut[20] [16]),
    .C(\datapath_1.regfile_1.regOut[24] [16]),
    .D(_5561__bF$buf2),
    .Y(_6133_)
);

NAND3X1 _15612_ (
    .A(_6129_),
    .B(_6133_),
    .C(_6132_),
    .Y(_6134_)
);

INVX1 _15613_ (
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_6135_)
);

INVX1 _15614_ (
    .A(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_6136_)
);

OAI22X1 _15615_ (
    .A(_5481_),
    .B(_6135_),
    .C(_6136_),
    .D(_5492__bF$buf2),
    .Y(_6137_)
);

INVX1 _15616_ (
    .A(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_6138_)
);

OAI22X1 _15617_ (
    .A(_5488__bF$buf2),
    .B(_4694_),
    .C(_6138_),
    .D(_5493__bF$buf2),
    .Y(_6139_)
);

NOR2X1 _15618_ (
    .A(_6137_),
    .B(_6139_),
    .Y(_6140_)
);

OAI22X1 _15619_ (
    .A(_4695_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_4704_),
    .Y(_6141_)
);

AOI21X1 _15620_ (
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .B(_5478__bF$buf2),
    .C(_6141_),
    .Y(_6142_)
);

INVX1 _15621_ (
    .A(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_6143_)
);

OAI22X1 _15622_ (
    .A(_4686_),
    .B(_5449_),
    .C(_5450_),
    .D(_6143_),
    .Y(_6144_)
);

AOI21X1 _15623_ (
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .B(_5560__bF$buf2),
    .C(_6144_),
    .Y(_6145_)
);

NAND3X1 _15624_ (
    .A(_6140_),
    .B(_6145_),
    .C(_6142_),
    .Y(_6146_)
);

NOR2X1 _15625_ (
    .A(_6134_),
    .B(_6146_),
    .Y(_6147_)
);

AOI21X1 _15626_ (
    .A(_6128_),
    .B(_6147_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [16])
);

INVX1 _15627_ (
    .A(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_6148_)
);

OAI22X1 _15628_ (
    .A(_4754_),
    .B(_5433__bF$buf2),
    .C(_5436__bF$buf2),
    .D(_6148_),
    .Y(_6149_)
);

NOR2X1 _15629_ (
    .A(_4744_),
    .B(_5428__bF$buf2),
    .Y(_6150_)
);

INVX1 _15630_ (
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_6151_)
);

NOR3X1 _15631_ (
    .A(_5421__bF$buf3),
    .B(_6151_),
    .C(_5423__bF$buf2),
    .Y(_6152_)
);

NOR3X1 _15632_ (
    .A(_6150_),
    .B(_6152_),
    .C(_6149_),
    .Y(_6153_)
);

INVX1 _15633_ (
    .A(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_6154_)
);

OAI22X1 _15634_ (
    .A(_5492__bF$buf1),
    .B(_6154_),
    .C(_4742_),
    .D(_5493__bF$buf1),
    .Y(_6155_)
);

INVX1 _15635_ (
    .A(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_6156_)
);

INVX1 _15636_ (
    .A(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_6157_)
);

OAI22X1 _15637_ (
    .A(_6157_),
    .B(_5481_),
    .C(_6156_),
    .D(_5488__bF$buf1),
    .Y(_6158_)
);

NOR2X1 _15638_ (
    .A(_6158_),
    .B(_6155_),
    .Y(_6159_)
);

INVX1 _15639_ (
    .A(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_6160_)
);

OAI22X1 _15640_ (
    .A(_4718_),
    .B(_5484__bF$buf2),
    .C(_5485__bF$buf2),
    .D(_6160_),
    .Y(_6161_)
);

AOI21X1 _15641_ (
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .B(_5478__bF$buf1),
    .C(_6161_),
    .Y(_6162_)
);

NAND3X1 _15642_ (
    .A(_6159_),
    .B(_6162_),
    .C(_6153_),
    .Y(_6163_)
);

AOI22X1 _15643_ (
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .B(_5457__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[1] [17]),
    .D(_5455__bF$buf2),
    .Y(_6164_)
);

AOI22X1 _15644_ (
    .A(_5460__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [17]),
    .C(_5462__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_6165_)
);

OAI22X1 _15645_ (
    .A(_4719_),
    .B(_5471__bF$buf2),
    .C(_4752_),
    .D(_5472__bF$buf2),
    .Y(_6166_)
);

OAI22X1 _15646_ (
    .A(_4731_),
    .B(_5465__bF$buf2),
    .C(_5466__bF$buf2),
    .D(_4716_),
    .Y(_6167_)
);

NOR2X1 _15647_ (
    .A(_6167_),
    .B(_6166_),
    .Y(_6168_)
);

NAND3X1 _15648_ (
    .A(_6165_),
    .B(_6164_),
    .C(_6168_),
    .Y(_6169_)
);

NOR2X1 _15649_ (
    .A(_6169_),
    .B(_6163_),
    .Y(_6170_)
);

NOR3X1 _15650_ (
    .A(_4741_),
    .B(_5558__bF$buf3),
    .C(_5555__bF$buf3),
    .Y(_6171_)
);

AOI22X1 _15651_ (
    .A(_5560__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [17]),
    .C(\datapath_1.regfile_1.regOut[24] [17]),
    .D(_5561__bF$buf1),
    .Y(_6172_)
);

NAND2X1 _15652_ (
    .A(\datapath_1.regfile_1.regOut[22] [17]),
    .B(_5563__bF$buf2),
    .Y(_6173_)
);

NAND2X1 _15653_ (
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .B(_5565__bF$buf2),
    .Y(_6174_)
);

NAND3X1 _15654_ (
    .A(_6173_),
    .B(_6172_),
    .C(_6174_),
    .Y(_6175_)
);

INVX1 _15655_ (
    .A(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_6176_)
);

OAI22X1 _15656_ (
    .A(_4726_),
    .B(_5506__bF$buf0),
    .C(_6176_),
    .D(_5511__bF$buf2),
    .Y(_6177_)
);

INVX1 _15657_ (
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_6178_)
);

INVX1 _15658_ (
    .A(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_6179_)
);

OAI22X1 _15659_ (
    .A(_5514__bF$buf2),
    .B(_6178_),
    .C(_6179_),
    .D(_5513__bF$buf2),
    .Y(_6180_)
);

NOR2X1 _15660_ (
    .A(_6180_),
    .B(_6177_),
    .Y(_6181_)
);

OAI22X1 _15661_ (
    .A(_5518__bF$buf2),
    .B(_4715_),
    .C(_4725_),
    .D(_5517__bF$buf2),
    .Y(_6182_)
);

OAI22X1 _15662_ (
    .A(_4722_),
    .B(_5520__bF$buf2),
    .C(_5521__bF$buf2),
    .D(_4730_),
    .Y(_6183_)
);

NOR2X1 _15663_ (
    .A(_6182_),
    .B(_6183_),
    .Y(_6184_)
);

NAND2X1 _15664_ (
    .A(_6181_),
    .B(_6184_),
    .Y(_6185_)
);

NOR3X1 _15665_ (
    .A(_6175_),
    .B(_6171_),
    .C(_6185_),
    .Y(_6186_)
);

AOI21X1 _15666_ (
    .A(_6170_),
    .B(_6186_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [17])
);

NOR2X1 _15667_ (
    .A(_4766_),
    .B(_5428__bF$buf1),
    .Y(_6187_)
);

INVX1 _15668_ (
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_6188_)
);

NOR3X1 _15669_ (
    .A(_5421__bF$buf2),
    .B(_6188_),
    .C(_5423__bF$buf1),
    .Y(_6189_)
);

INVX1 _15670_ (
    .A(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_6190_)
);

INVX1 _15671_ (
    .A(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_6191_)
);

OAI22X1 _15672_ (
    .A(_6191_),
    .B(_5433__bF$buf1),
    .C(_5436__bF$buf1),
    .D(_6190_),
    .Y(_6192_)
);

NOR3X1 _15673_ (
    .A(_6189_),
    .B(_6187_),
    .C(_6192_),
    .Y(_6193_)
);

OAI22X1 _15674_ (
    .A(_5492__bF$buf0),
    .B(_4774_),
    .C(_4777_),
    .D(_5493__bF$buf0),
    .Y(_6194_)
);

AOI21X1 _15675_ (
    .A(\datapath_1.regfile_1.regOut[30] [18]),
    .B(_5489_),
    .C(_6194_),
    .Y(_6195_)
);

INVX1 _15676_ (
    .A(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_6196_)
);

OAI22X1 _15677_ (
    .A(_6196_),
    .B(_5484__bF$buf1),
    .C(_5485__bF$buf1),
    .D(_4797_),
    .Y(_6197_)
);

INVX1 _15678_ (
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_6198_)
);

OAI22X1 _15679_ (
    .A(_5481_),
    .B(_6198_),
    .C(_4800_),
    .D(_5477_),
    .Y(_6199_)
);

NOR2X1 _15680_ (
    .A(_6199_),
    .B(_6197_),
    .Y(_6200_)
);

NAND3X1 _15681_ (
    .A(_6195_),
    .B(_6200_),
    .C(_6193_),
    .Y(_6201_)
);

AOI22X1 _15682_ (
    .A(\datapath_1.regfile_1.regOut[4] [18]),
    .B(_5457__bF$buf1),
    .C(\datapath_1.regfile_1.regOut[1] [18]),
    .D(_5455__bF$buf1),
    .Y(_6202_)
);

AOI22X1 _15683_ (
    .A(_5460__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [18]),
    .C(_5462__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_6203_)
);

INVX1 _15684_ (
    .A(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_6204_)
);

OAI22X1 _15685_ (
    .A(_6204_),
    .B(_5465__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_4769_),
    .Y(_6205_)
);

OAI22X1 _15686_ (
    .A(_4790_),
    .B(_5471__bF$buf1),
    .C(_4767_),
    .D(_5472__bF$buf1),
    .Y(_6206_)
);

NOR2X1 _15687_ (
    .A(_6205_),
    .B(_6206_),
    .Y(_6207_)
);

NAND3X1 _15688_ (
    .A(_6203_),
    .B(_6202_),
    .C(_6207_),
    .Y(_6208_)
);

NOR2X1 _15689_ (
    .A(_6208_),
    .B(_6201_),
    .Y(_6209_)
);

NOR3X1 _15690_ (
    .A(_4792_),
    .B(_5558__bF$buf2),
    .C(_5555__bF$buf2),
    .Y(_6210_)
);

NAND2X1 _15691_ (
    .A(\datapath_1.regfile_1.regOut[22] [18]),
    .B(_5563__bF$buf1),
    .Y(_6211_)
);

AOI22X1 _15692_ (
    .A(_5560__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [18]),
    .C(\datapath_1.regfile_1.regOut[24] [18]),
    .D(_5561__bF$buf0),
    .Y(_6212_)
);

NAND2X1 _15693_ (
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .B(_5565__bF$buf1),
    .Y(_6213_)
);

NAND3X1 _15694_ (
    .A(_6211_),
    .B(_6213_),
    .C(_6212_),
    .Y(_6214_)
);

OAI22X1 _15695_ (
    .A(_4801_),
    .B(_5506__bF$buf4),
    .C(_4793_),
    .D(_5511__bF$buf1),
    .Y(_6215_)
);

INVX1 _15696_ (
    .A(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_6216_)
);

OAI22X1 _15697_ (
    .A(_5514__bF$buf1),
    .B(_6216_),
    .C(_4770_),
    .D(_5513__bF$buf1),
    .Y(_6217_)
);

NOR2X1 _15698_ (
    .A(_6217_),
    .B(_6215_),
    .Y(_6218_)
);

OAI22X1 _15699_ (
    .A(_5518__bF$buf1),
    .B(_4778_),
    .C(_4775_),
    .D(_5517__bF$buf1),
    .Y(_6219_)
);

INVX1 _15700_ (
    .A(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_6220_)
);

OAI22X1 _15701_ (
    .A(_6220_),
    .B(_5520__bF$buf1),
    .C(_5521__bF$buf1),
    .D(_4762_),
    .Y(_6221_)
);

NOR2X1 _15702_ (
    .A(_6219_),
    .B(_6221_),
    .Y(_6222_)
);

NAND2X1 _15703_ (
    .A(_6218_),
    .B(_6222_),
    .Y(_6223_)
);

NOR3X1 _15704_ (
    .A(_6214_),
    .B(_6210_),
    .C(_6223_),
    .Y(_6224_)
);

AOI21X1 _15705_ (
    .A(_6209_),
    .B(_6224_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [18])
);

NOR2X1 _15706_ (
    .A(_4825_),
    .B(_5428__bF$buf0),
    .Y(_6225_)
);

NOR3X1 _15707_ (
    .A(_5421__bF$buf1),
    .B(_4829_),
    .C(_5423__bF$buf0),
    .Y(_6226_)
);

INVX1 _15708_ (
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_6227_)
);

INVX1 _15709_ (
    .A(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_6228_)
);

OAI22X1 _15710_ (
    .A(_6228_),
    .B(_5433__bF$buf0),
    .C(_5436__bF$buf0),
    .D(_6227_),
    .Y(_6229_)
);

NOR3X1 _15711_ (
    .A(_6226_),
    .B(_6225_),
    .C(_6229_),
    .Y(_6230_)
);

INVX1 _15712_ (
    .A(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_6231_)
);

INVX1 _15713_ (
    .A(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_6232_)
);

OAI22X1 _15714_ (
    .A(_5492__bF$buf4),
    .B(_6232_),
    .C(_6231_),
    .D(_5493__bF$buf3),
    .Y(_6233_)
);

INVX1 _15715_ (
    .A(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_6234_)
);

OAI22X1 _15716_ (
    .A(_6234_),
    .B(_5481_),
    .C(_4846_),
    .D(_5488__bF$buf0),
    .Y(_6235_)
);

NOR2X1 _15717_ (
    .A(_6235_),
    .B(_6233_),
    .Y(_6236_)
);

OAI22X1 _15718_ (
    .A(_4847_),
    .B(_5484__bF$buf0),
    .C(_5485__bF$buf0),
    .D(_4828_),
    .Y(_6237_)
);

AOI21X1 _15719_ (
    .A(\datapath_1.regfile_1.regOut[27] [19]),
    .B(_5478__bF$buf0),
    .C(_6237_),
    .Y(_6238_)
);

NAND3X1 _15720_ (
    .A(_6236_),
    .B(_6238_),
    .C(_6230_),
    .Y(_6239_)
);

AOI22X1 _15721_ (
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .B(_5457__bF$buf0),
    .C(\datapath_1.regfile_1.regOut[1] [19]),
    .D(_5455__bF$buf0),
    .Y(_6240_)
);

AOI22X1 _15722_ (
    .A(_5460__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [19]),
    .C(_5462__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_6241_)
);

OAI22X1 _15723_ (
    .A(_4835_),
    .B(_5465__bF$buf0),
    .C(_5466__bF$buf0),
    .D(_4838_),
    .Y(_6242_)
);

OAI22X1 _15724_ (
    .A(_4834_),
    .B(_5471__bF$buf0),
    .C(_4837_),
    .D(_5472__bF$buf0),
    .Y(_6243_)
);

NOR2X1 _15725_ (
    .A(_6242_),
    .B(_6243_),
    .Y(_6244_)
);

NAND3X1 _15726_ (
    .A(_6241_),
    .B(_6240_),
    .C(_6244_),
    .Y(_6245_)
);

NOR2X1 _15727_ (
    .A(_6245_),
    .B(_6239_),
    .Y(_6246_)
);

INVX1 _15728_ (
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_6247_)
);

NOR3X1 _15729_ (
    .A(_6247_),
    .B(_5558__bF$buf1),
    .C(_5555__bF$buf1),
    .Y(_6248_)
);

NAND2X1 _15730_ (
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .B(_5563__bF$buf0),
    .Y(_6249_)
);

NAND2X1 _15731_ (
    .A(\datapath_1.regfile_1.regOut[21] [19]),
    .B(_5565__bF$buf0),
    .Y(_6250_)
);

AOI22X1 _15732_ (
    .A(_5560__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .C(\datapath_1.regfile_1.regOut[24] [19]),
    .D(_5561__bF$buf3),
    .Y(_6251_)
);

NAND3X1 _15733_ (
    .A(_6249_),
    .B(_6251_),
    .C(_6250_),
    .Y(_6252_)
);

OAI22X1 _15734_ (
    .A(_4819_),
    .B(_5506__bF$buf3),
    .C(_4814_),
    .D(_5511__bF$buf0),
    .Y(_6253_)
);

INVX1 _15735_ (
    .A(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_6254_)
);

OAI22X1 _15736_ (
    .A(_5514__bF$buf0),
    .B(_4813_),
    .C(_6254_),
    .D(_5513__bF$buf0),
    .Y(_6255_)
);

NOR2X1 _15737_ (
    .A(_6255_),
    .B(_6253_),
    .Y(_6256_)
);

OAI22X1 _15738_ (
    .A(_5518__bF$buf0),
    .B(_4850_),
    .C(_4821_),
    .D(_5517__bF$buf0),
    .Y(_6257_)
);

OAI22X1 _15739_ (
    .A(_4818_),
    .B(_5520__bF$buf0),
    .C(_5521__bF$buf0),
    .D(_4849_),
    .Y(_6258_)
);

NOR2X1 _15740_ (
    .A(_6257_),
    .B(_6258_),
    .Y(_6259_)
);

NAND2X1 _15741_ (
    .A(_6259_),
    .B(_6256_),
    .Y(_6260_)
);

NOR3X1 _15742_ (
    .A(_6252_),
    .B(_6248_),
    .C(_6260_),
    .Y(_6261_)
);

AOI21X1 _15743_ (
    .A(_6246_),
    .B(_6261_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [19])
);

NOR2X1 _15744_ (
    .A(_4859_),
    .B(_5428__bF$buf3),
    .Y(_6262_)
);

INVX1 _15745_ (
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_6263_)
);

NOR3X1 _15746_ (
    .A(_5421__bF$buf0),
    .B(_6263_),
    .C(_5423__bF$buf3),
    .Y(_6264_)
);

INVX1 _15747_ (
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_6265_)
);

INVX1 _15748_ (
    .A(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_6266_)
);

OAI22X1 _15749_ (
    .A(_6266_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_6265_),
    .Y(_6267_)
);

NOR3X1 _15750_ (
    .A(_6264_),
    .B(_6262_),
    .C(_6267_),
    .Y(_6268_)
);

INVX1 _15751_ (
    .A(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_6269_)
);

INVX1 _15752_ (
    .A(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_6270_)
);

OAI22X1 _15753_ (
    .A(_5492__bF$buf3),
    .B(_6270_),
    .C(_6269_),
    .D(_5493__bF$buf2),
    .Y(_6271_)
);

AOI21X1 _15754_ (
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .B(_5489_),
    .C(_6271_),
    .Y(_6272_)
);

OAI22X1 _15755_ (
    .A(_4893_),
    .B(_5484__bF$buf4),
    .C(_5485__bF$buf4),
    .D(_4885_),
    .Y(_6273_)
);

OAI22X1 _15756_ (
    .A(_5481_),
    .B(_4890_),
    .C(_4867_),
    .D(_5477_),
    .Y(_6274_)
);

NOR2X1 _15757_ (
    .A(_6274_),
    .B(_6273_),
    .Y(_6275_)
);

NAND3X1 _15758_ (
    .A(_6272_),
    .B(_6275_),
    .C(_6268_),
    .Y(_6276_)
);

AOI22X1 _15759_ (
    .A(\datapath_1.regfile_1.regOut[4] [20]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [20]),
    .D(_5455__bF$buf4),
    .Y(_6277_)
);

AOI22X1 _15760_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [20]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_6278_)
);

OAI22X1 _15761_ (
    .A(_4883_),
    .B(_5471__bF$buf4),
    .C(_4860_),
    .D(_5472__bF$buf4),
    .Y(_6279_)
);

INVX1 _15762_ (
    .A(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_6280_)
);

OAI22X1 _15763_ (
    .A(_6280_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_4862_),
    .Y(_6281_)
);

NOR2X1 _15764_ (
    .A(_6281_),
    .B(_6279_),
    .Y(_6282_)
);

NAND3X1 _15765_ (
    .A(_6278_),
    .B(_6277_),
    .C(_6282_),
    .Y(_6283_)
);

NOR2X1 _15766_ (
    .A(_6283_),
    .B(_6276_),
    .Y(_6284_)
);

INVX1 _15767_ (
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_6285_)
);

NOR3X1 _15768_ (
    .A(_6285_),
    .B(_5558__bF$buf0),
    .C(_5555__bF$buf0),
    .Y(_6286_)
);

NAND2X1 _15769_ (
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .B(_5565__bF$buf3),
    .Y(_6287_)
);

NAND2X1 _15770_ (
    .A(\datapath_1.regfile_1.regOut[22] [20]),
    .B(_5563__bF$buf3),
    .Y(_6288_)
);

AOI22X1 _15771_ (
    .A(_5560__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [20]),
    .C(\datapath_1.regfile_1.regOut[24] [20]),
    .D(_5561__bF$buf2),
    .Y(_6289_)
);

NAND3X1 _15772_ (
    .A(_6287_),
    .B(_6289_),
    .C(_6288_),
    .Y(_6290_)
);

OAI22X1 _15773_ (
    .A(_4894_),
    .B(_5506__bF$buf2),
    .C(_4886_),
    .D(_5511__bF$buf4),
    .Y(_6291_)
);

INVX1 _15774_ (
    .A(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_6292_)
);

OAI22X1 _15775_ (
    .A(_5514__bF$buf4),
    .B(_6292_),
    .C(_4863_),
    .D(_5513__bF$buf4),
    .Y(_6293_)
);

NOR2X1 _15776_ (
    .A(_6293_),
    .B(_6291_),
    .Y(_6294_)
);

OAI22X1 _15777_ (
    .A(_5518__bF$buf4),
    .B(_4871_),
    .C(_4868_),
    .D(_5517__bF$buf4),
    .Y(_6295_)
);

INVX1 _15778_ (
    .A(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_6296_)
);

OAI22X1 _15779_ (
    .A(_6296_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_4855_),
    .Y(_6297_)
);

NOR2X1 _15780_ (
    .A(_6295_),
    .B(_6297_),
    .Y(_6298_)
);

NAND2X1 _15781_ (
    .A(_6294_),
    .B(_6298_),
    .Y(_6299_)
);

NOR3X1 _15782_ (
    .A(_6290_),
    .B(_6286_),
    .C(_6299_),
    .Y(_6300_)
);

AOI21X1 _15783_ (
    .A(_6284_),
    .B(_6300_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [20])
);

NAND2X1 _15784_ (
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .B(_5429_),
    .Y(_6301_)
);

INVX1 _15785_ (
    .A(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_6302_)
);

OAI22X1 _15786_ (
    .A(_6302_),
    .B(_5433__bF$buf3),
    .C(_5436__bF$buf3),
    .D(_4942_),
    .Y(_6303_)
);

AOI21X1 _15787_ (
    .A(\datapath_1.regfile_1.regOut[20] [21]),
    .B(_5424_),
    .C(_6303_),
    .Y(_6304_)
);

INVX1 _15788_ (
    .A(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_6305_)
);

INVX1 _15789_ (
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_6306_)
);

OAI22X1 _15790_ (
    .A(_5443_),
    .B(_6306_),
    .C(_6305_),
    .D(_5447_),
    .Y(_6307_)
);

OAI22X1 _15791_ (
    .A(_4939_),
    .B(_5449_),
    .C(_5450_),
    .D(_4938_),
    .Y(_6308_)
);

NOR2X1 _15792_ (
    .A(_6308_),
    .B(_6307_),
    .Y(_6309_)
);

NAND3X1 _15793_ (
    .A(_6304_),
    .B(_6301_),
    .C(_6309_),
    .Y(_6310_)
);

AOI22X1 _15794_ (
    .A(\datapath_1.regfile_1.regOut[4] [21]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [21]),
    .D(_5455__bF$buf3),
    .Y(_6311_)
);

AOI22X1 _15795_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [21]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_6312_)
);

INVX1 _15796_ (
    .A(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_6313_)
);

INVX1 _15797_ (
    .A(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_6314_)
);

OAI22X1 _15798_ (
    .A(_6314_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_6313_),
    .Y(_6315_)
);

INVX1 _15799_ (
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_6316_)
);

OAI22X1 _15800_ (
    .A(_6316_),
    .B(_5471__bF$buf3),
    .C(_4932_),
    .D(_5472__bF$buf3),
    .Y(_6317_)
);

NOR2X1 _15801_ (
    .A(_6315_),
    .B(_6317_),
    .Y(_6318_)
);

NAND3X1 _15802_ (
    .A(_6312_),
    .B(_6311_),
    .C(_6318_),
    .Y(_6319_)
);

NOR2X1 _15803_ (
    .A(_6310_),
    .B(_6319_),
    .Y(_6320_)
);

NAND2X1 _15804_ (
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .B(_5478__bF$buf3),
    .Y(_6321_)
);

OAI22X1 _15805_ (
    .A(_4913_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_4916_),
    .Y(_6322_)
);

AOI21X1 _15806_ (
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .B(_5482__bF$buf0),
    .C(_6322_),
    .Y(_6323_)
);

OAI22X1 _15807_ (
    .A(_5492__bF$buf2),
    .B(_4904_),
    .C(_4928_),
    .D(_5493__bF$buf1),
    .Y(_6324_)
);

AOI21X1 _15808_ (
    .A(\datapath_1.regfile_1.regOut[30] [21]),
    .B(_5489_),
    .C(_6324_),
    .Y(_6325_)
);

NAND3X1 _15809_ (
    .A(_6321_),
    .B(_6325_),
    .C(_6323_),
    .Y(_6326_)
);

NAND3X1 _15810_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [21]),
    .C(_5509_),
    .Y(_6327_)
);

INVX1 _15811_ (
    .A(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_6328_)
);

OAI22X1 _15812_ (
    .A(_4908_),
    .B(_5506__bF$buf1),
    .C(_6328_),
    .D(_5511__bF$buf3),
    .Y(_6329_)
);

INVX1 _15813_ (
    .A(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_6330_)
);

INVX1 _15814_ (
    .A(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_6331_)
);

OAI22X1 _15815_ (
    .A(_5514__bF$buf3),
    .B(_6330_),
    .C(_6331_),
    .D(_5513__bF$buf3),
    .Y(_6332_)
);

NOR2X1 _15816_ (
    .A(_6332_),
    .B(_6329_),
    .Y(_6333_)
);

OAI22X1 _15817_ (
    .A(_5518__bF$buf3),
    .B(_4917_),
    .C(_4914_),
    .D(_5517__bF$buf3),
    .Y(_6334_)
);

OAI22X1 _15818_ (
    .A(_4902_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_4901_),
    .Y(_6335_)
);

NOR2X1 _15819_ (
    .A(_6334_),
    .B(_6335_),
    .Y(_6336_)
);

NAND3X1 _15820_ (
    .A(_6333_),
    .B(_6336_),
    .C(_6327_),
    .Y(_6337_)
);

NOR2X1 _15821_ (
    .A(_6326_),
    .B(_6337_),
    .Y(_6338_)
);

AOI21X1 _15822_ (
    .A(_6338_),
    .B(_6320_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [21])
);

NOR2X1 _15823_ (
    .A(_4960_),
    .B(_5428__bF$buf2),
    .Y(_6339_)
);

NOR3X1 _15824_ (
    .A(_5421__bF$buf3),
    .B(_4988_),
    .C(_5423__bF$buf2),
    .Y(_6340_)
);

INVX1 _15825_ (
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_6341_)
);

OAI22X1 _15826_ (
    .A(_4971_),
    .B(_5433__bF$buf2),
    .C(_5436__bF$buf2),
    .D(_6341_),
    .Y(_6342_)
);

NOR3X1 _15827_ (
    .A(_6340_),
    .B(_6339_),
    .C(_6342_),
    .Y(_6343_)
);

INVX1 _15828_ (
    .A(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_6344_)
);

INVX1 _15829_ (
    .A(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_6345_)
);

OAI22X1 _15830_ (
    .A(_6345_),
    .B(_5484__bF$buf2),
    .C(_5485__bF$buf2),
    .D(_6344_),
    .Y(_6346_)
);

AOI21X1 _15831_ (
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .B(_5482__bF$buf3),
    .C(_6346_),
    .Y(_6347_)
);

INVX1 _15832_ (
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_6348_)
);

INVX1 _15833_ (
    .A(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_6349_)
);

OAI22X1 _15834_ (
    .A(_5492__bF$buf1),
    .B(_6349_),
    .C(_6348_),
    .D(_5493__bF$buf0),
    .Y(_6350_)
);

INVX1 _15835_ (
    .A(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_6351_)
);

OAI22X1 _15836_ (
    .A(_6351_),
    .B(_5477_),
    .C(_5488__bF$buf3),
    .D(_4950_),
    .Y(_6352_)
);

NOR2X1 _15837_ (
    .A(_6352_),
    .B(_6350_),
    .Y(_6353_)
);

NAND3X1 _15838_ (
    .A(_6347_),
    .B(_6353_),
    .C(_6343_),
    .Y(_6354_)
);

AOI22X1 _15839_ (
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .B(_5457__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[1] [22]),
    .D(_5455__bF$buf2),
    .Y(_6355_)
);

AOI22X1 _15840_ (
    .A(_5460__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [22]),
    .C(_5462__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_6356_)
);

INVX1 _15841_ (
    .A(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_6357_)
);

OAI22X1 _15842_ (
    .A(_4989_),
    .B(_5465__bF$buf2),
    .C(_5466__bF$buf2),
    .D(_6357_),
    .Y(_6358_)
);

INVX1 _15843_ (
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_6359_)
);

OAI22X1 _15844_ (
    .A(_6359_),
    .B(_5471__bF$buf2),
    .C(_4958_),
    .D(_5472__bF$buf2),
    .Y(_6360_)
);

NOR2X1 _15845_ (
    .A(_6358_),
    .B(_6360_),
    .Y(_6361_)
);

NAND3X1 _15846_ (
    .A(_6356_),
    .B(_6355_),
    .C(_6361_),
    .Y(_6362_)
);

NOR2X1 _15847_ (
    .A(_6362_),
    .B(_6354_),
    .Y(_6363_)
);

NOR3X1 _15848_ (
    .A(_4957_),
    .B(_5558__bF$buf3),
    .C(_5555__bF$buf3),
    .Y(_6364_)
);

NAND2X1 _15849_ (
    .A(\datapath_1.regfile_1.regOut[21] [22]),
    .B(_5565__bF$buf2),
    .Y(_6365_)
);

NAND2X1 _15850_ (
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .B(_5563__bF$buf2),
    .Y(_6366_)
);

AOI22X1 _15851_ (
    .A(_5560__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [22]),
    .C(\datapath_1.regfile_1.regOut[24] [22]),
    .D(_5561__bF$buf1),
    .Y(_6367_)
);

NAND3X1 _15852_ (
    .A(_6365_),
    .B(_6367_),
    .C(_6366_),
    .Y(_6368_)
);

OAI22X1 _15853_ (
    .A(_4974_),
    .B(_5506__bF$buf0),
    .C(_4979_),
    .D(_5511__bF$buf2),
    .Y(_6369_)
);

INVX1 _15854_ (
    .A(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_6370_)
);

OAI22X1 _15855_ (
    .A(_5514__bF$buf2),
    .B(_6370_),
    .C(_4948_),
    .D(_5513__bF$buf2),
    .Y(_6371_)
);

NOR2X1 _15856_ (
    .A(_6371_),
    .B(_6369_),
    .Y(_6372_)
);

OAI22X1 _15857_ (
    .A(_5518__bF$buf2),
    .B(_4981_),
    .C(_4973_),
    .D(_5517__bF$buf2),
    .Y(_6373_)
);

OAI22X1 _15858_ (
    .A(_4986_),
    .B(_5520__bF$buf2),
    .C(_5521__bF$buf2),
    .D(_4985_),
    .Y(_6374_)
);

NOR2X1 _15859_ (
    .A(_6373_),
    .B(_6374_),
    .Y(_6375_)
);

NAND2X1 _15860_ (
    .A(_6372_),
    .B(_6375_),
    .Y(_6376_)
);

NOR3X1 _15861_ (
    .A(_6368_),
    .B(_6364_),
    .C(_6376_),
    .Y(_6377_)
);

AOI21X1 _15862_ (
    .A(_6363_),
    .B(_6377_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [22])
);

NOR2X1 _15863_ (
    .A(_5001_),
    .B(_5428__bF$buf1),
    .Y(_6378_)
);

INVX1 _15864_ (
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_6379_)
);

NOR3X1 _15865_ (
    .A(_5421__bF$buf2),
    .B(_6379_),
    .C(_5423__bF$buf1),
    .Y(_6380_)
);

INVX1 _15866_ (
    .A(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_6381_)
);

OAI22X1 _15867_ (
    .A(_5034_),
    .B(_5433__bF$buf1),
    .C(_5436__bF$buf1),
    .D(_6381_),
    .Y(_6382_)
);

NOR3X1 _15868_ (
    .A(_6380_),
    .B(_6378_),
    .C(_6382_),
    .Y(_6383_)
);

INVX1 _15869_ (
    .A(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_6384_)
);

INVX1 _15870_ (
    .A(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_6385_)
);

OAI22X1 _15871_ (
    .A(_6385_),
    .B(_5484__bF$buf1),
    .C(_5485__bF$buf1),
    .D(_6384_),
    .Y(_6386_)
);

AOI21X1 _15872_ (
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .B(_5482__bF$buf2),
    .C(_6386_),
    .Y(_6387_)
);

OAI22X1 _15873_ (
    .A(_5022_),
    .B(_5449_),
    .C(_5450_),
    .D(_5021_),
    .Y(_6388_)
);

INVX1 _15874_ (
    .A(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_6389_)
);

INVX1 _15875_ (
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_6390_)
);

OAI22X1 _15876_ (
    .A(_5443_),
    .B(_6390_),
    .C(_6389_),
    .D(_5447_),
    .Y(_6391_)
);

NOR2X1 _15877_ (
    .A(_6388_),
    .B(_6391_),
    .Y(_6392_)
);

NAND3X1 _15878_ (
    .A(_6387_),
    .B(_6392_),
    .C(_6383_),
    .Y(_6393_)
);

AOI22X1 _15879_ (
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .B(_5457__bF$buf1),
    .C(\datapath_1.regfile_1.regOut[1] [23]),
    .D(_5455__bF$buf1),
    .Y(_6394_)
);

AOI22X1 _15880_ (
    .A(_5460__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [23]),
    .C(_5462__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_6395_)
);

INVX1 _15881_ (
    .A(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_6396_)
);

OAI22X1 _15882_ (
    .A(_6396_),
    .B(_5465__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_5012_),
    .Y(_6397_)
);

OAI22X1 _15883_ (
    .A(_5011_),
    .B(_5471__bF$buf1),
    .C(_5002_),
    .D(_5472__bF$buf1),
    .Y(_6398_)
);

NOR2X1 _15884_ (
    .A(_6397_),
    .B(_6398_),
    .Y(_6399_)
);

NAND3X1 _15885_ (
    .A(_6395_),
    .B(_6394_),
    .C(_6399_),
    .Y(_6400_)
);

NOR2X1 _15886_ (
    .A(_6400_),
    .B(_6393_),
    .Y(_6401_)
);

NOR3X1 _15887_ (
    .A(_5008_),
    .B(_5558__bF$buf2),
    .C(_5555__bF$buf2),
    .Y(_6402_)
);

NAND2X1 _15888_ (
    .A(\datapath_1.regfile_1.regOut[27] [23]),
    .B(_5478__bF$buf2),
    .Y(_6403_)
);

NAND2X1 _15889_ (
    .A(\datapath_1.regfile_1.regOut[30] [23]),
    .B(_5489_),
    .Y(_6404_)
);

AOI22X1 _15890_ (
    .A(\datapath_1.regfile_1.regOut[29] [23]),
    .B(_5641_),
    .C(\datapath_1.regfile_1.regOut[31] [23]),
    .D(_5642_),
    .Y(_6405_)
);

NAND3X1 _15891_ (
    .A(_6404_),
    .B(_6405_),
    .C(_6403_),
    .Y(_6406_)
);

OAI22X1 _15892_ (
    .A(_5018_),
    .B(_5506__bF$buf4),
    .C(_5025_),
    .D(_5511__bF$buf1),
    .Y(_6407_)
);

INVX1 _15893_ (
    .A(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_6408_)
);

OAI22X1 _15894_ (
    .A(_5514__bF$buf1),
    .B(_5009_),
    .C(_6408_),
    .D(_5513__bF$buf1),
    .Y(_6409_)
);

NOR2X1 _15895_ (
    .A(_6409_),
    .B(_6407_),
    .Y(_6410_)
);

OAI22X1 _15896_ (
    .A(_5518__bF$buf1),
    .B(_4998_),
    .C(_4999_),
    .D(_5517__bF$buf1),
    .Y(_6411_)
);

OAI22X1 _15897_ (
    .A(_5031_),
    .B(_5520__bF$buf1),
    .C(_5521__bF$buf1),
    .D(_5035_),
    .Y(_6412_)
);

NOR2X1 _15898_ (
    .A(_6411_),
    .B(_6412_),
    .Y(_6413_)
);

NAND2X1 _15899_ (
    .A(_6410_),
    .B(_6413_),
    .Y(_6414_)
);

NOR3X1 _15900_ (
    .A(_6406_),
    .B(_6402_),
    .C(_6414_),
    .Y(_6415_)
);

AOI21X1 _15901_ (
    .A(_6401_),
    .B(_6415_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [23])
);

NOR2X1 _15902_ (
    .A(_5074_),
    .B(_5428__bF$buf0),
    .Y(_6416_)
);

INVX1 _15903_ (
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_6417_)
);

NOR3X1 _15904_ (
    .A(_5421__bF$buf1),
    .B(_6417_),
    .C(_5423__bF$buf0),
    .Y(_6418_)
);

INVX1 _15905_ (
    .A(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_6419_)
);

OAI22X1 _15906_ (
    .A(_5083_),
    .B(_5433__bF$buf0),
    .C(_5436__bF$buf0),
    .D(_6419_),
    .Y(_6420_)
);

NOR3X1 _15907_ (
    .A(_6418_),
    .B(_6416_),
    .C(_6420_),
    .Y(_6421_)
);

INVX1 _15908_ (
    .A(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_6422_)
);

INVX1 _15909_ (
    .A(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_6423_)
);

OAI22X1 _15910_ (
    .A(_6423_),
    .B(_5484__bF$buf0),
    .C(_5485__bF$buf0),
    .D(_6422_),
    .Y(_6424_)
);

AOI21X1 _15911_ (
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .B(_5482__bF$buf1),
    .C(_6424_),
    .Y(_6425_)
);

INVX1 _15912_ (
    .A(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_6426_)
);

OAI22X1 _15913_ (
    .A(_5492__bF$buf0),
    .B(_5041_),
    .C(_6426_),
    .D(_5493__bF$buf3),
    .Y(_6427_)
);

INVX1 _15914_ (
    .A(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_6428_)
);

OAI22X1 _15915_ (
    .A(_6428_),
    .B(_5477_),
    .C(_5488__bF$buf2),
    .D(_5040_),
    .Y(_6429_)
);

NOR2X1 _15916_ (
    .A(_6429_),
    .B(_6427_),
    .Y(_6430_)
);

NAND3X1 _15917_ (
    .A(_6425_),
    .B(_6430_),
    .C(_6421_),
    .Y(_6431_)
);

AOI22X1 _15918_ (
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .B(_5457__bF$buf0),
    .C(\datapath_1.regfile_1.regOut[1] [24]),
    .D(_5455__bF$buf0),
    .Y(_6432_)
);

AOI22X1 _15919_ (
    .A(_5460__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [24]),
    .C(_5462__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_6433_)
);

INVX1 _15920_ (
    .A(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_6434_)
);

OAI22X1 _15921_ (
    .A(_6434_),
    .B(_5465__bF$buf0),
    .C(_5466__bF$buf0),
    .D(_5044_),
    .Y(_6435_)
);

OAI22X1 _15922_ (
    .A(_5063_),
    .B(_5471__bF$buf0),
    .C(_5043_),
    .D(_5472__bF$buf0),
    .Y(_6436_)
);

NOR2X1 _15923_ (
    .A(_6435_),
    .B(_6436_),
    .Y(_6437_)
);

NAND3X1 _15924_ (
    .A(_6433_),
    .B(_6432_),
    .C(_6437_),
    .Y(_6438_)
);

NOR2X1 _15925_ (
    .A(_6438_),
    .B(_6431_),
    .Y(_6439_)
);

NOR3X1 _15926_ (
    .A(_5059_),
    .B(_5558__bF$buf1),
    .C(_5555__bF$buf1),
    .Y(_6440_)
);

NAND2X1 _15927_ (
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .B(_5565__bF$buf1),
    .Y(_6441_)
);

NAND2X1 _15928_ (
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .B(_5563__bF$buf1),
    .Y(_6442_)
);

AOI22X1 _15929_ (
    .A(_5560__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [24]),
    .C(\datapath_1.regfile_1.regOut[24] [24]),
    .D(_5561__bF$buf0),
    .Y(_6443_)
);

NAND3X1 _15930_ (
    .A(_6441_),
    .B(_6443_),
    .C(_6442_),
    .Y(_6444_)
);

OAI22X1 _15931_ (
    .A(_5056_),
    .B(_5506__bF$buf3),
    .C(_5051_),
    .D(_5511__bF$buf0),
    .Y(_6445_)
);

INVX1 _15932_ (
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_6446_)
);

OAI22X1 _15933_ (
    .A(_5514__bF$buf0),
    .B(_5070_),
    .C(_6446_),
    .D(_5513__bF$buf0),
    .Y(_6447_)
);

NOR2X1 _15934_ (
    .A(_6447_),
    .B(_6445_),
    .Y(_6448_)
);

OAI22X1 _15935_ (
    .A(_5518__bF$buf0),
    .B(_5047_),
    .C(_5048_),
    .D(_5517__bF$buf0),
    .Y(_6449_)
);

OAI22X1 _15936_ (
    .A(_5080_),
    .B(_5520__bF$buf0),
    .C(_5521__bF$buf0),
    .D(_5084_),
    .Y(_6450_)
);

NOR2X1 _15937_ (
    .A(_6449_),
    .B(_6450_),
    .Y(_6451_)
);

NAND2X1 _15938_ (
    .A(_6448_),
    .B(_6451_),
    .Y(_6452_)
);

NOR3X1 _15939_ (
    .A(_6444_),
    .B(_6440_),
    .C(_6452_),
    .Y(_6453_)
);

AOI21X1 _15940_ (
    .A(_6439_),
    .B(_6453_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [24])
);

NAND2X1 _15941_ (
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .B(_5429_),
    .Y(_6454_)
);

INVX1 _15942_ (
    .A(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_6455_)
);

INVX1 _15943_ (
    .A(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_6456_)
);

OAI22X1 _15944_ (
    .A(_6456_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_6455_),
    .Y(_6457_)
);

AOI21X1 _15945_ (
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .B(_5424_),
    .C(_6457_),
    .Y(_6458_)
);

INVX1 _15946_ (
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_6459_)
);

OAI22X1 _15947_ (
    .A(_5443_),
    .B(_6459_),
    .C(_5100_),
    .D(_5447_),
    .Y(_6460_)
);

OAI22X1 _15948_ (
    .A(_5123_),
    .B(_5449_),
    .C(_5450_),
    .D(_5122_),
    .Y(_6461_)
);

NOR2X1 _15949_ (
    .A(_6461_),
    .B(_6460_),
    .Y(_6462_)
);

NAND3X1 _15950_ (
    .A(_6458_),
    .B(_6454_),
    .C(_6462_),
    .Y(_6463_)
);

AOI22X1 _15951_ (
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [25]),
    .D(_5455__bF$buf4),
    .Y(_6464_)
);

AOI22X1 _15952_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [25]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_6465_)
);

OAI22X1 _15953_ (
    .A(_5134_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_5115_),
    .Y(_6466_)
);

OAI22X1 _15954_ (
    .A(_5114_),
    .B(_5471__bF$buf4),
    .C(_5097_),
    .D(_5472__bF$buf4),
    .Y(_6467_)
);

NOR2X1 _15955_ (
    .A(_6466_),
    .B(_6467_),
    .Y(_6468_)
);

NAND3X1 _15956_ (
    .A(_6465_),
    .B(_6464_),
    .C(_6468_),
    .Y(_6469_)
);

NOR2X1 _15957_ (
    .A(_6463_),
    .B(_6469_),
    .Y(_6470_)
);

NAND2X1 _15958_ (
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .B(_5478__bF$buf1),
    .Y(_6471_)
);

OAI22X1 _15959_ (
    .A(_5111_),
    .B(_5484__bF$buf4),
    .C(_5485__bF$buf4),
    .D(_5093_),
    .Y(_6472_)
);

AOI21X1 _15960_ (
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .B(_5482__bF$buf0),
    .C(_6472_),
    .Y(_6473_)
);

INVX1 _15961_ (
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_6474_)
);

INVX1 _15962_ (
    .A(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_6475_)
);

OAI22X1 _15963_ (
    .A(_5492__bF$buf4),
    .B(_6475_),
    .C(_6474_),
    .D(_5493__bF$buf2),
    .Y(_6476_)
);

AOI21X1 _15964_ (
    .A(\datapath_1.regfile_1.regOut[30] [25]),
    .B(_5489_),
    .C(_6476_),
    .Y(_6477_)
);

NAND3X1 _15965_ (
    .A(_6471_),
    .B(_6477_),
    .C(_6473_),
    .Y(_6478_)
);

NAND3X1 _15966_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [25]),
    .C(_5509_),
    .Y(_6479_)
);

OAI22X1 _15967_ (
    .A(_5108_),
    .B(_5506__bF$buf2),
    .C(_5090_),
    .D(_5511__bF$buf4),
    .Y(_6480_)
);

OAI22X1 _15968_ (
    .A(_5514__bF$buf4),
    .B(_5112_),
    .C(_5125_),
    .D(_5513__bF$buf4),
    .Y(_6481_)
);

NOR2X1 _15969_ (
    .A(_6481_),
    .B(_6480_),
    .Y(_6482_)
);

OAI22X1 _15970_ (
    .A(_5518__bF$buf4),
    .B(_5105_),
    .C(_5131_),
    .D(_5517__bF$buf4),
    .Y(_6483_)
);

OAI22X1 _15971_ (
    .A(_5130_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_5133_),
    .Y(_6484_)
);

NOR2X1 _15972_ (
    .A(_6483_),
    .B(_6484_),
    .Y(_6485_)
);

NAND3X1 _15973_ (
    .A(_6482_),
    .B(_6485_),
    .C(_6479_),
    .Y(_6486_)
);

NOR2X1 _15974_ (
    .A(_6478_),
    .B(_6486_),
    .Y(_6487_)
);

AOI21X1 _15975_ (
    .A(_6487_),
    .B(_6470_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [25])
);

AOI22X1 _15976_ (
    .A(_5563__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[22] [26]),
    .C(_5565__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_6488_)
);

INVX1 _15977_ (
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_6489_)
);

INVX1 _15978_ (
    .A(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_6490_)
);

OAI22X1 _15979_ (
    .A(_6490_),
    .B(_5433__bF$buf3),
    .C(_5436__bF$buf3),
    .D(_6489_),
    .Y(_6491_)
);

AOI21X1 _15980_ (
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .B(_5429_),
    .C(_6491_),
    .Y(_6492_)
);

AOI22X1 _15981_ (
    .A(_5424_),
    .B(\datapath_1.regfile_1.regOut[20] [26]),
    .C(\datapath_1.regfile_1.regOut[24] [26]),
    .D(_5561__bF$buf3),
    .Y(_6493_)
);

NAND3X1 _15982_ (
    .A(_6493_),
    .B(_6488_),
    .C(_6492_),
    .Y(_6494_)
);

AOI22X1 _15983_ (
    .A(\datapath_1.regfile_1.regOut[4] [26]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [26]),
    .D(_5455__bF$buf3),
    .Y(_6495_)
);

AOI22X1 _15984_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_6496_)
);

INVX1 _15985_ (
    .A(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_6497_)
);

OAI22X1 _15986_ (
    .A(_6497_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_5148_),
    .Y(_6498_)
);

OAI22X1 _15987_ (
    .A(_5169_),
    .B(_5471__bF$buf3),
    .C(_5146_),
    .D(_5472__bF$buf3),
    .Y(_6499_)
);

NOR2X1 _15988_ (
    .A(_6498_),
    .B(_6499_),
    .Y(_6500_)
);

NAND3X1 _15989_ (
    .A(_6496_),
    .B(_6495_),
    .C(_6500_),
    .Y(_6501_)
);

NOR2X1 _15990_ (
    .A(_6494_),
    .B(_6501_),
    .Y(_6502_)
);

NAND2X1 _15991_ (
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .B(_5560__bF$buf3),
    .Y(_6503_)
);

OAI22X1 _15992_ (
    .A(_5179_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_5177_),
    .Y(_6504_)
);

AOI21X1 _15993_ (
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .B(_5482__bF$buf3),
    .C(_6504_),
    .Y(_6505_)
);

OAI22X1 _15994_ (
    .A(_5153_),
    .B(_5477_),
    .C(_5488__bF$buf1),
    .D(_5156_),
    .Y(_6506_)
);

INVX1 _15995_ (
    .A(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_6507_)
);

NAND3X1 _15996_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(\datapath_1.regfile_1.regOut[31] [26]),
    .C(_5470_),
    .Y(_6508_)
);

OAI21X1 _15997_ (
    .A(_6507_),
    .B(_5492__bF$buf3),
    .C(_6508_),
    .Y(_6509_)
);

NOR2X1 _15998_ (
    .A(_6509_),
    .B(_6506_),
    .Y(_6510_)
);

NAND3X1 _15999_ (
    .A(_6503_),
    .B(_6510_),
    .C(_6505_),
    .Y(_6511_)
);

NAND3X1 _16000_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [26]),
    .C(_5509_),
    .Y(_6512_)
);

OAI22X1 _16001_ (
    .A(_5180_),
    .B(_5506__bF$buf1),
    .C(_5172_),
    .D(_5511__bF$buf3),
    .Y(_6513_)
);

INVX1 _16002_ (
    .A(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_6514_)
);

OAI22X1 _16003_ (
    .A(_5514__bF$buf3),
    .B(_6514_),
    .C(_5149_),
    .D(_5513__bF$buf3),
    .Y(_6515_)
);

NOR2X1 _16004_ (
    .A(_6515_),
    .B(_6513_),
    .Y(_6516_)
);

OAI22X1 _16005_ (
    .A(_5518__bF$buf3),
    .B(_5157_),
    .C(_5154_),
    .D(_5517__bF$buf3),
    .Y(_6517_)
);

INVX1 _16006_ (
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_6518_)
);

OAI22X1 _16007_ (
    .A(_6518_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_5141_),
    .Y(_6519_)
);

NOR2X1 _16008_ (
    .A(_6517_),
    .B(_6519_),
    .Y(_6520_)
);

NAND3X1 _16009_ (
    .A(_6516_),
    .B(_6520_),
    .C(_6512_),
    .Y(_6521_)
);

NOR2X1 _16010_ (
    .A(_6511_),
    .B(_6521_),
    .Y(_6522_)
);

AOI21X1 _16011_ (
    .A(_6522_),
    .B(_6502_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [26])
);

NOR2X1 _16012_ (
    .A(_5194_),
    .B(_5428__bF$buf3),
    .Y(_6523_)
);

INVX1 _16013_ (
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_6524_)
);

NOR3X1 _16014_ (
    .A(_5421__bF$buf0),
    .B(_6524_),
    .C(_5423__bF$buf3),
    .Y(_6525_)
);

INVX1 _16015_ (
    .A(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_6526_)
);

INVX1 _16016_ (
    .A(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_6527_)
);

OAI22X1 _16017_ (
    .A(_6527_),
    .B(_5433__bF$buf2),
    .C(_5436__bF$buf2),
    .D(_6526_),
    .Y(_6528_)
);

NOR3X1 _16018_ (
    .A(_6525_),
    .B(_6523_),
    .C(_6528_),
    .Y(_6529_)
);

OAI22X1 _16019_ (
    .A(_5492__bF$buf2),
    .B(_5207_),
    .C(_5218_),
    .D(_5493__bF$buf1),
    .Y(_6530_)
);

AOI21X1 _16020_ (
    .A(\datapath_1.regfile_1.regOut[30] [27]),
    .B(_5489_),
    .C(_6530_),
    .Y(_6531_)
);

OAI22X1 _16021_ (
    .A(_5224_),
    .B(_5484__bF$buf2),
    .C(_5485__bF$buf2),
    .D(_5226_),
    .Y(_6532_)
);

OAI22X1 _16022_ (
    .A(_5481_),
    .B(_5190_),
    .C(_5197_),
    .D(_5477_),
    .Y(_6533_)
);

NOR2X1 _16023_ (
    .A(_6533_),
    .B(_6532_),
    .Y(_6534_)
);

NAND3X1 _16024_ (
    .A(_6531_),
    .B(_6534_),
    .C(_6529_),
    .Y(_6535_)
);

AOI22X1 _16025_ (
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .B(_5457__bF$buf2),
    .C(\datapath_1.regfile_1.regOut[1] [27]),
    .D(_5455__bF$buf2),
    .Y(_6536_)
);

AOI22X1 _16026_ (
    .A(_5460__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [27]),
    .C(_5462__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_6537_)
);

INVX1 _16027_ (
    .A(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_6538_)
);

OAI22X1 _16028_ (
    .A(_6538_),
    .B(_5465__bF$buf2),
    .C(_5466__bF$buf2),
    .D(_5198_),
    .Y(_6539_)
);

INVX1 _16029_ (
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_6540_)
);

OAI22X1 _16030_ (
    .A(_6540_),
    .B(_5471__bF$buf2),
    .C(_5195_),
    .D(_5472__bF$buf2),
    .Y(_6541_)
);

NOR2X1 _16031_ (
    .A(_6539_),
    .B(_6541_),
    .Y(_6542_)
);

NAND3X1 _16032_ (
    .A(_6537_),
    .B(_6536_),
    .C(_6542_),
    .Y(_6543_)
);

NOR2X1 _16033_ (
    .A(_6543_),
    .B(_6535_),
    .Y(_6544_)
);

NOR3X1 _16034_ (
    .A(_5223_),
    .B(_5558__bF$buf0),
    .C(_5555__bF$buf0),
    .Y(_6545_)
);

NAND2X1 _16035_ (
    .A(\datapath_1.regfile_1.regOut[22] [27]),
    .B(_5563__bF$buf3),
    .Y(_6546_)
);

NAND2X1 _16036_ (
    .A(\datapath_1.regfile_1.regOut[21] [27]),
    .B(_5565__bF$buf3),
    .Y(_6547_)
);

AOI22X1 _16037_ (
    .A(_5560__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .C(\datapath_1.regfile_1.regOut[24] [27]),
    .D(_5561__bF$buf2),
    .Y(_6548_)
);

NAND3X1 _16038_ (
    .A(_6546_),
    .B(_6548_),
    .C(_6547_),
    .Y(_6549_)
);

OAI22X1 _16039_ (
    .A(_5205_),
    .B(_5506__bF$buf0),
    .C(_5216_),
    .D(_5511__bF$buf2),
    .Y(_6550_)
);

INVX1 _16040_ (
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_6551_)
);

INVX1 _16041_ (
    .A(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_6552_)
);

OAI22X1 _16042_ (
    .A(_5514__bF$buf2),
    .B(_6551_),
    .C(_6552_),
    .D(_5513__bF$buf2),
    .Y(_6553_)
);

NOR2X1 _16043_ (
    .A(_6553_),
    .B(_6550_),
    .Y(_6554_)
);

OAI22X1 _16044_ (
    .A(_5518__bF$buf2),
    .B(_5219_),
    .C(_5187_),
    .D(_5517__bF$buf2),
    .Y(_6555_)
);

OAI22X1 _16045_ (
    .A(_5191_),
    .B(_5520__bF$buf2),
    .C(_5521__bF$buf2),
    .D(_5204_),
    .Y(_6556_)
);

NOR2X1 _16046_ (
    .A(_6555_),
    .B(_6556_),
    .Y(_6557_)
);

NAND2X1 _16047_ (
    .A(_6554_),
    .B(_6557_),
    .Y(_6558_)
);

NOR3X1 _16048_ (
    .A(_6549_),
    .B(_6545_),
    .C(_6558_),
    .Y(_6559_)
);

AOI21X1 _16049_ (
    .A(_6544_),
    .B(_6559_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [27])
);

NOR2X1 _16050_ (
    .A(_5241_),
    .B(_5428__bF$buf2),
    .Y(_6560_)
);

INVX1 _16051_ (
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_6561_)
);

NOR3X1 _16052_ (
    .A(_5421__bF$buf3),
    .B(_6561_),
    .C(_5423__bF$buf2),
    .Y(_6562_)
);

INVX1 _16053_ (
    .A(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_6563_)
);

OAI22X1 _16054_ (
    .A(_5251_),
    .B(_5433__bF$buf1),
    .C(_5436__bF$buf1),
    .D(_6563_),
    .Y(_6564_)
);

NOR3X1 _16055_ (
    .A(_6562_),
    .B(_6560_),
    .C(_6564_),
    .Y(_6565_)
);

OAI22X1 _16056_ (
    .A(_5492__bF$buf1),
    .B(_5265_),
    .C(_5237_),
    .D(_5493__bF$buf0),
    .Y(_6566_)
);

OAI22X1 _16057_ (
    .A(_5270_),
    .B(_5481_),
    .C(_5254_),
    .D(_5488__bF$buf0),
    .Y(_6567_)
);

NOR2X1 _16058_ (
    .A(_6567_),
    .B(_6566_),
    .Y(_6568_)
);

OAI22X1 _16059_ (
    .A(_5273_),
    .B(_5484__bF$buf1),
    .C(_5485__bF$buf1),
    .D(_5244_),
    .Y(_6569_)
);

AOI21X1 _16060_ (
    .A(\datapath_1.regfile_1.regOut[27] [28]),
    .B(_5478__bF$buf0),
    .C(_6569_),
    .Y(_6570_)
);

NAND3X1 _16061_ (
    .A(_6568_),
    .B(_6570_),
    .C(_6565_),
    .Y(_6571_)
);

AOI22X1 _16062_ (
    .A(\datapath_1.regfile_1.regOut[4] [28]),
    .B(_5457__bF$buf1),
    .C(\datapath_1.regfile_1.regOut[1] [28]),
    .D(_5455__bF$buf1),
    .Y(_6572_)
);

AOI22X1 _16063_ (
    .A(_5460__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [28]),
    .C(_5462__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_6573_)
);

INVX1 _16064_ (
    .A(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_6574_)
);

OAI22X1 _16065_ (
    .A(_6574_),
    .B(_5465__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_5245_),
    .Y(_6575_)
);

INVX1 _16066_ (
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_6576_)
);

OAI22X1 _16067_ (
    .A(_6576_),
    .B(_5471__bF$buf1),
    .C(_5242_),
    .D(_5472__bF$buf1),
    .Y(_6577_)
);

NOR2X1 _16068_ (
    .A(_6575_),
    .B(_6577_),
    .Y(_6578_)
);

NAND3X1 _16069_ (
    .A(_6573_),
    .B(_6572_),
    .C(_6578_),
    .Y(_6579_)
);

NOR2X1 _16070_ (
    .A(_6579_),
    .B(_6571_),
    .Y(_6580_)
);

INVX1 _16071_ (
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_6581_)
);

NOR3X1 _16072_ (
    .A(_6581_),
    .B(_5558__bF$buf3),
    .C(_5555__bF$buf3),
    .Y(_6582_)
);

NAND2X1 _16073_ (
    .A(\datapath_1.regfile_1.regOut[22] [28]),
    .B(_5563__bF$buf2),
    .Y(_6583_)
);

NAND2X1 _16074_ (
    .A(\datapath_1.regfile_1.regOut[21] [28]),
    .B(_5565__bF$buf2),
    .Y(_6584_)
);

AOI22X1 _16075_ (
    .A(_5560__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [28]),
    .C(\datapath_1.regfile_1.regOut[24] [28]),
    .D(_5561__bF$buf1),
    .Y(_6585_)
);

NAND3X1 _16076_ (
    .A(_6583_),
    .B(_6585_),
    .C(_6584_),
    .Y(_6586_)
);

OAI22X1 _16077_ (
    .A(_5274_),
    .B(_5506__bF$buf4),
    .C(_5235_),
    .D(_5511__bF$buf1),
    .Y(_6587_)
);

INVX1 _16078_ (
    .A(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_6588_)
);

OAI22X1 _16079_ (
    .A(_5514__bF$buf1),
    .B(_6588_),
    .C(_5263_),
    .D(_5513__bF$buf1),
    .Y(_6589_)
);

NOR2X1 _16080_ (
    .A(_6589_),
    .B(_6587_),
    .Y(_6590_)
);

OAI22X1 _16081_ (
    .A(_5518__bF$buf1),
    .B(_5234_),
    .C(_5252_),
    .D(_5517__bF$buf1),
    .Y(_6591_)
);

OAI22X1 _16082_ (
    .A(_5266_),
    .B(_5520__bF$buf1),
    .C(_5521__bF$buf1),
    .D(_5238_),
    .Y(_6592_)
);

NOR2X1 _16083_ (
    .A(_6591_),
    .B(_6592_),
    .Y(_6593_)
);

NAND2X1 _16084_ (
    .A(_6590_),
    .B(_6593_),
    .Y(_6594_)
);

NOR3X1 _16085_ (
    .A(_6586_),
    .B(_6582_),
    .C(_6594_),
    .Y(_6595_)
);

AOI21X1 _16086_ (
    .A(_6580_),
    .B(_6595_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [28])
);

INVX1 _16087_ (
    .A(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_6596_)
);

OAI22X1 _16088_ (
    .A(_5304_),
    .B(_5433__bF$buf0),
    .C(_5436__bF$buf0),
    .D(_6596_),
    .Y(_6597_)
);

NOR2X1 _16089_ (
    .A(_5299_),
    .B(_5428__bF$buf1),
    .Y(_6598_)
);

INVX1 _16090_ (
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_6599_)
);

NOR3X1 _16091_ (
    .A(_5421__bF$buf2),
    .B(_6599_),
    .C(_5423__bF$buf1),
    .Y(_6600_)
);

NOR3X1 _16092_ (
    .A(_6598_),
    .B(_6600_),
    .C(_6597_),
    .Y(_6601_)
);

INVX1 _16093_ (
    .A(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_6602_)
);

OAI22X1 _16094_ (
    .A(_5314_),
    .B(_5484__bF$buf0),
    .C(_5485__bF$buf0),
    .D(_6602_),
    .Y(_6603_)
);

AOI21X1 _16095_ (
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .B(_5482__bF$buf2),
    .C(_6603_),
    .Y(_6604_)
);

INVX1 _16096_ (
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_6605_)
);

INVX1 _16097_ (
    .A(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_6606_)
);

OAI22X1 _16098_ (
    .A(_5492__bF$buf0),
    .B(_6606_),
    .C(_6605_),
    .D(_5493__bF$buf3),
    .Y(_6607_)
);

INVX1 _16099_ (
    .A(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_6608_)
);

OAI22X1 _16100_ (
    .A(_5317_),
    .B(_5477_),
    .C(_5488__bF$buf3),
    .D(_6608_),
    .Y(_6609_)
);

NOR2X1 _16101_ (
    .A(_6609_),
    .B(_6607_),
    .Y(_6610_)
);

NAND3X1 _16102_ (
    .A(_6604_),
    .B(_6610_),
    .C(_6601_),
    .Y(_6611_)
);

AOI22X1 _16103_ (
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .B(_5457__bF$buf0),
    .C(\datapath_1.regfile_1.regOut[1] [29]),
    .D(_5455__bF$buf0),
    .Y(_6612_)
);

AOI22X1 _16104_ (
    .A(_5460__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [29]),
    .C(_5462__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_6613_)
);

INVX1 _16105_ (
    .A(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_6614_)
);

OAI22X1 _16106_ (
    .A(_6614_),
    .B(_5465__bF$buf0),
    .C(_5466__bF$buf0),
    .D(_5285_),
    .Y(_6615_)
);

OAI22X1 _16107_ (
    .A(_5284_),
    .B(_5471__bF$buf0),
    .C(_5296_),
    .D(_5472__bF$buf0),
    .Y(_6616_)
);

NOR2X1 _16108_ (
    .A(_6615_),
    .B(_6616_),
    .Y(_6617_)
);

NAND3X1 _16109_ (
    .A(_6613_),
    .B(_6612_),
    .C(_6617_),
    .Y(_6618_)
);

NOR2X1 _16110_ (
    .A(_6618_),
    .B(_6611_),
    .Y(_6619_)
);

NOR3X1 _16111_ (
    .A(_5298_),
    .B(_5558__bF$buf2),
    .C(_5555__bF$buf2),
    .Y(_6620_)
);

NAND2X1 _16112_ (
    .A(\datapath_1.regfile_1.regOut[21] [29]),
    .B(_5565__bF$buf1),
    .Y(_6621_)
);

NAND2X1 _16113_ (
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .B(_5563__bF$buf1),
    .Y(_6622_)
);

AOI22X1 _16114_ (
    .A(_5560__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [29]),
    .C(\datapath_1.regfile_1.regOut[24] [29]),
    .D(_5561__bF$buf0),
    .Y(_6623_)
);

NAND3X1 _16115_ (
    .A(_6621_),
    .B(_6623_),
    .C(_6622_),
    .Y(_6624_)
);

INVX1 _16116_ (
    .A(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_6625_)
);

OAI22X1 _16117_ (
    .A(_5282_),
    .B(_5506__bF$buf3),
    .C(_6625_),
    .D(_5511__bF$buf0),
    .Y(_6626_)
);

INVX1 _16118_ (
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_6627_)
);

OAI22X1 _16119_ (
    .A(_5514__bF$buf0),
    .B(_6627_),
    .C(_5315_),
    .D(_5513__bF$buf0),
    .Y(_6628_)
);

NOR2X1 _16120_ (
    .A(_6628_),
    .B(_6626_),
    .Y(_6629_)
);

OAI22X1 _16121_ (
    .A(_5518__bF$buf0),
    .B(_5307_),
    .C(_5321_),
    .D(_5517__bF$buf0),
    .Y(_6630_)
);

OAI22X1 _16122_ (
    .A(_5318_),
    .B(_5520__bF$buf0),
    .C(_5521__bF$buf0),
    .D(_5305_),
    .Y(_6631_)
);

NOR2X1 _16123_ (
    .A(_6630_),
    .B(_6631_),
    .Y(_6632_)
);

NAND2X1 _16124_ (
    .A(_6629_),
    .B(_6632_),
    .Y(_6633_)
);

NOR3X1 _16125_ (
    .A(_6624_),
    .B(_6620_),
    .C(_6633_),
    .Y(_6634_)
);

AOI21X1 _16126_ (
    .A(_6619_),
    .B(_6634_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [29])
);

NAND2X1 _16127_ (
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .B(_5478__bF$buf3),
    .Y(_6635_)
);

INVX1 _16128_ (
    .A(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_6636_)
);

INVX1 _16129_ (
    .A(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_6637_)
);

OAI22X1 _16130_ (
    .A(_5481_),
    .B(_6636_),
    .C(_6637_),
    .D(_5492__bF$buf4),
    .Y(_6638_)
);

INVX1 _16131_ (
    .A(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_6639_)
);

INVX1 _16132_ (
    .A(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_6640_)
);

OAI22X1 _16133_ (
    .A(_5488__bF$buf2),
    .B(_6639_),
    .C(_6640_),
    .D(_5493__bF$buf2),
    .Y(_6641_)
);

NOR2X1 _16134_ (
    .A(_6638_),
    .B(_6641_),
    .Y(_6642_)
);

INVX1 _16135_ (
    .A(_5484__bF$buf4),
    .Y(_6643_)
);

INVX1 _16136_ (
    .A(_5485__bF$buf4),
    .Y(_6644_)
);

AOI22X1 _16137_ (
    .A(_6644_),
    .B(\datapath_1.regfile_1.regOut[26] [30]),
    .C(_6643_),
    .D(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_6645_)
);

NAND3X1 _16138_ (
    .A(_6635_),
    .B(_6645_),
    .C(_6642_),
    .Y(_6646_)
);

AOI22X1 _16139_ (
    .A(\datapath_1.regfile_1.regOut[4] [30]),
    .B(_5457__bF$buf4),
    .C(\datapath_1.regfile_1.regOut[1] [30]),
    .D(_5455__bF$buf4),
    .Y(_6647_)
);

AOI22X1 _16140_ (
    .A(_5460__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[6] [30]),
    .C(_5462__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_6648_)
);

INVX1 _16141_ (
    .A(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_6649_)
);

OAI22X1 _16142_ (
    .A(_6649_),
    .B(_5465__bF$buf4),
    .C(_5466__bF$buf4),
    .D(_5343_),
    .Y(_6650_)
);

OAI22X1 _16143_ (
    .A(_5330_),
    .B(_5471__bF$buf4),
    .C(_5342_),
    .D(_5472__bF$buf4),
    .Y(_6651_)
);

NOR2X1 _16144_ (
    .A(_6650_),
    .B(_6651_),
    .Y(_6652_)
);

NAND3X1 _16145_ (
    .A(_6648_),
    .B(_6647_),
    .C(_6652_),
    .Y(_6653_)
);

NOR2X1 _16146_ (
    .A(_6646_),
    .B(_6653_),
    .Y(_6654_)
);

AOI22X1 _16147_ (
    .A(_5429_),
    .B(\datapath_1.regfile_1.regOut[19] [30]),
    .C(\datapath_1.regfile_1.regOut[24] [30]),
    .D(_5561__bF$buf3),
    .Y(_6655_)
);

OAI22X1 _16148_ (
    .A(_5351_),
    .B(_5449_),
    .C(_5450_),
    .D(_5350_),
    .Y(_6656_)
);

AOI21X1 _16149_ (
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .B(_5560__bF$buf3),
    .C(_6656_),
    .Y(_6657_)
);

INVX1 _16150_ (
    .A(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_6658_)
);

INVX1 _16151_ (
    .A(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_6659_)
);

OAI22X1 _16152_ (
    .A(_6659_),
    .B(_5433__bF$buf4),
    .C(_5436__bF$buf4),
    .D(_6658_),
    .Y(_6660_)
);

AOI21X1 _16153_ (
    .A(\datapath_1.regfile_1.regOut[20] [30]),
    .B(_5424_),
    .C(_6660_),
    .Y(_6661_)
);

NAND3X1 _16154_ (
    .A(_6655_),
    .B(_6661_),
    .C(_6657_),
    .Y(_6662_)
);

NAND3X1 _16155_ (
    .A(_5502_),
    .B(\datapath_1.regfile_1.regOut[0] [30]),
    .C(_5509_),
    .Y(_6663_)
);

INVX1 _16156_ (
    .A(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_6664_)
);

OAI22X1 _16157_ (
    .A(_5333_),
    .B(_5506__bF$buf2),
    .C(_6664_),
    .D(_5511__bF$buf4),
    .Y(_6665_)
);

OAI22X1 _16158_ (
    .A(_5514__bF$buf4),
    .B(_5340_),
    .C(_5353_),
    .D(_5513__bF$buf4),
    .Y(_6666_)
);

NOR2X1 _16159_ (
    .A(_6666_),
    .B(_6665_),
    .Y(_6667_)
);

OAI22X1 _16160_ (
    .A(_5518__bF$buf4),
    .B(_5363_),
    .C(_5332_),
    .D(_5517__bF$buf4),
    .Y(_6668_)
);

OAI22X1 _16161_ (
    .A(_5361_),
    .B(_5520__bF$buf4),
    .C(_5521__bF$buf4),
    .D(_5360_),
    .Y(_6669_)
);

NOR2X1 _16162_ (
    .A(_6668_),
    .B(_6669_),
    .Y(_6670_)
);

NAND3X1 _16163_ (
    .A(_6667_),
    .B(_6670_),
    .C(_6663_),
    .Y(_6671_)
);

NOR2X1 _16164_ (
    .A(_6662_),
    .B(_6671_),
    .Y(_6672_)
);

AOI21X1 _16165_ (
    .A(_6672_),
    .B(_6654_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [30])
);

NOR2X1 _16166_ (
    .A(_5402_),
    .B(_5428__bF$buf0),
    .Y(_6673_)
);

NOR3X1 _16167_ (
    .A(_5421__bF$buf1),
    .B(_5369_),
    .C(_5423__bF$buf0),
    .Y(_6674_)
);

INVX1 _16168_ (
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_6675_)
);

OAI22X1 _16169_ (
    .A(_6675_),
    .B(_5433__bF$buf3),
    .C(_5436__bF$buf3),
    .D(_5372_),
    .Y(_6676_)
);

NOR3X1 _16170_ (
    .A(_6674_),
    .B(_6673_),
    .C(_6676_),
    .Y(_6677_)
);

OAI22X1 _16171_ (
    .A(_5411_),
    .B(_5484__bF$buf3),
    .C(_5485__bF$buf3),
    .D(_5376_),
    .Y(_6678_)
);

AOI21X1 _16172_ (
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .B(_5482__bF$buf1),
    .C(_6678_),
    .Y(_6679_)
);

INVX1 _16173_ (
    .A(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_6680_)
);

INVX1 _16174_ (
    .A(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_6681_)
);

OAI22X1 _16175_ (
    .A(_5492__bF$buf3),
    .B(_6681_),
    .C(_6680_),
    .D(_5493__bF$buf1),
    .Y(_6682_)
);

INVX1 _16176_ (
    .A(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_6683_)
);

INVX1 _16177_ (
    .A(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_6684_)
);

OAI22X1 _16178_ (
    .A(_6684_),
    .B(_5477_),
    .C(_5488__bF$buf1),
    .D(_6683_),
    .Y(_6685_)
);

NOR2X1 _16179_ (
    .A(_6685_),
    .B(_6682_),
    .Y(_6686_)
);

NAND3X1 _16180_ (
    .A(_6679_),
    .B(_6686_),
    .C(_6677_),
    .Y(_6687_)
);

AOI22X1 _16181_ (
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .B(_5457__bF$buf3),
    .C(\datapath_1.regfile_1.regOut[1] [31]),
    .D(_5455__bF$buf3),
    .Y(_6688_)
);

AOI22X1 _16182_ (
    .A(_5460__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [31]),
    .C(_5462__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_6689_)
);

OAI22X1 _16183_ (
    .A(_5414_),
    .B(_5471__bF$buf3),
    .C(_5377_),
    .D(_5472__bF$buf3),
    .Y(_6690_)
);

INVX1 _16184_ (
    .A(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_6691_)
);

INVX1 _16185_ (
    .A(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_6692_)
);

OAI22X1 _16186_ (
    .A(_6692_),
    .B(_5465__bF$buf3),
    .C(_5466__bF$buf3),
    .D(_6691_),
    .Y(_6693_)
);

NOR2X1 _16187_ (
    .A(_6693_),
    .B(_6690_),
    .Y(_6694_)
);

NAND3X1 _16188_ (
    .A(_6689_),
    .B(_6688_),
    .C(_6694_),
    .Y(_6695_)
);

NOR2X1 _16189_ (
    .A(_6695_),
    .B(_6687_),
    .Y(_6696_)
);

INVX1 _16190_ (
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_6697_)
);

NOR3X1 _16191_ (
    .A(_6697_),
    .B(_5558__bF$buf1),
    .C(_5555__bF$buf1),
    .Y(_6698_)
);

NAND2X1 _16192_ (
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .B(_5565__bF$buf0),
    .Y(_6699_)
);

NAND2X1 _16193_ (
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .B(_5563__bF$buf0),
    .Y(_6700_)
);

AOI22X1 _16194_ (
    .A(_5560__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [31]),
    .C(\datapath_1.regfile_1.regOut[24] [31]),
    .D(_5561__bF$buf2),
    .Y(_6701_)
);

NAND3X1 _16195_ (
    .A(_6699_),
    .B(_6701_),
    .C(_6700_),
    .Y(_6702_)
);

OAI22X1 _16196_ (
    .A(_5415_),
    .B(_5506__bF$buf1),
    .C(_5388_),
    .D(_5511__bF$buf3),
    .Y(_6703_)
);

OAI22X1 _16197_ (
    .A(_5514__bF$buf3),
    .B(_5412_),
    .C(_5400_),
    .D(_5513__bF$buf3),
    .Y(_6704_)
);

NOR2X1 _16198_ (
    .A(_6704_),
    .B(_6703_),
    .Y(_6705_)
);

OAI22X1 _16199_ (
    .A(_5518__bF$buf3),
    .B(_5373_),
    .C(_5407_),
    .D(_5517__bF$buf3),
    .Y(_6706_)
);

OAI22X1 _16200_ (
    .A(_5370_),
    .B(_5520__bF$buf3),
    .C(_5521__bF$buf3),
    .D(_5395_),
    .Y(_6707_)
);

NOR2X1 _16201_ (
    .A(_6706_),
    .B(_6707_),
    .Y(_6708_)
);

NAND2X1 _16202_ (
    .A(_6705_),
    .B(_6708_),
    .Y(_6709_)
);

NOR3X1 _16203_ (
    .A(_6702_),
    .B(_6698_),
    .C(_6709_),
    .Y(_6710_)
);

AOI21X1 _16204_ (
    .A(_6696_),
    .B(_6710_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [31])
);

INVX1 _16205_ (
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_6774_)
);

NAND2X1 _16206_ (
    .A(gnd),
    .B(gnd),
    .Y(_6775_)
);

OAI21X1 _16207_ (
    .A(gnd),
    .B(_6774_),
    .C(_6775_),
    .Y(_6711_[0])
);

INVX1 _16208_ (
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_6712_)
);

NAND2X1 _16209_ (
    .A(gnd),
    .B(gnd),
    .Y(_6713_)
);

OAI21X1 _16210_ (
    .A(gnd),
    .B(_6712_),
    .C(_6713_),
    .Y(_6711_[1])
);

INVX1 _16211_ (
    .A(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_6714_)
);

NAND2X1 _16212_ (
    .A(gnd),
    .B(gnd),
    .Y(_6715_)
);

OAI21X1 _16213_ (
    .A(gnd),
    .B(_6714_),
    .C(_6715_),
    .Y(_6711_[2])
);

INVX1 _16214_ (
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_6716_)
);

NAND2X1 _16215_ (
    .A(gnd),
    .B(gnd),
    .Y(_6717_)
);

OAI21X1 _16216_ (
    .A(gnd),
    .B(_6716_),
    .C(_6717_),
    .Y(_6711_[3])
);

INVX1 _16217_ (
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .Y(_6718_)
);

NAND2X1 _16218_ (
    .A(gnd),
    .B(gnd),
    .Y(_6719_)
);

OAI21X1 _16219_ (
    .A(gnd),
    .B(_6718_),
    .C(_6719_),
    .Y(_6711_[4])
);

INVX1 _16220_ (
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_6720_)
);

NAND2X1 _16221_ (
    .A(gnd),
    .B(gnd),
    .Y(_6721_)
);

OAI21X1 _16222_ (
    .A(gnd),
    .B(_6720_),
    .C(_6721_),
    .Y(_6711_[5])
);

INVX1 _16223_ (
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_6722_)
);

NAND2X1 _16224_ (
    .A(gnd),
    .B(gnd),
    .Y(_6723_)
);

OAI21X1 _16225_ (
    .A(gnd),
    .B(_6722_),
    .C(_6723_),
    .Y(_6711_[6])
);

INVX1 _16226_ (
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .Y(_6724_)
);

NAND2X1 _16227_ (
    .A(gnd),
    .B(gnd),
    .Y(_6725_)
);

OAI21X1 _16228_ (
    .A(gnd),
    .B(_6724_),
    .C(_6725_),
    .Y(_6711_[7])
);

INVX1 _16229_ (
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_6726_)
);

NAND2X1 _16230_ (
    .A(gnd),
    .B(gnd),
    .Y(_6727_)
);

OAI21X1 _16231_ (
    .A(gnd),
    .B(_6726_),
    .C(_6727_),
    .Y(_6711_[8])
);

INVX1 _16232_ (
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .Y(_6728_)
);

NAND2X1 _16233_ (
    .A(gnd),
    .B(gnd),
    .Y(_6729_)
);

OAI21X1 _16234_ (
    .A(gnd),
    .B(_6728_),
    .C(_6729_),
    .Y(_6711_[9])
);

INVX1 _16235_ (
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_6730_)
);

NAND2X1 _16236_ (
    .A(gnd),
    .B(gnd),
    .Y(_6731_)
);

OAI21X1 _16237_ (
    .A(gnd),
    .B(_6730_),
    .C(_6731_),
    .Y(_6711_[10])
);

INVX1 _16238_ (
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_6732_)
);

NAND2X1 _16239_ (
    .A(gnd),
    .B(gnd),
    .Y(_6733_)
);

OAI21X1 _16240_ (
    .A(gnd),
    .B(_6732_),
    .C(_6733_),
    .Y(_6711_[11])
);

INVX1 _16241_ (
    .A(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_6734_)
);

NAND2X1 _16242_ (
    .A(gnd),
    .B(gnd),
    .Y(_6735_)
);

OAI21X1 _16243_ (
    .A(gnd),
    .B(_6734_),
    .C(_6735_),
    .Y(_6711_[12])
);

INVX1 _16244_ (
    .A(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_6736_)
);

NAND2X1 _16245_ (
    .A(gnd),
    .B(gnd),
    .Y(_6737_)
);

OAI21X1 _16246_ (
    .A(gnd),
    .B(_6736_),
    .C(_6737_),
    .Y(_6711_[13])
);

INVX1 _16247_ (
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_6738_)
);

NAND2X1 _16248_ (
    .A(gnd),
    .B(gnd),
    .Y(_6739_)
);

OAI21X1 _16249_ (
    .A(gnd),
    .B(_6738_),
    .C(_6739_),
    .Y(_6711_[14])
);

INVX1 _16250_ (
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_6740_)
);

NAND2X1 _16251_ (
    .A(gnd),
    .B(gnd),
    .Y(_6741_)
);

OAI21X1 _16252_ (
    .A(gnd),
    .B(_6740_),
    .C(_6741_),
    .Y(_6711_[15])
);

INVX1 _16253_ (
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_6742_)
);

NAND2X1 _16254_ (
    .A(gnd),
    .B(gnd),
    .Y(_6743_)
);

OAI21X1 _16255_ (
    .A(gnd),
    .B(_6742_),
    .C(_6743_),
    .Y(_6711_[16])
);

INVX1 _16256_ (
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_6744_)
);

NAND2X1 _16257_ (
    .A(gnd),
    .B(gnd),
    .Y(_6745_)
);

OAI21X1 _16258_ (
    .A(gnd),
    .B(_6744_),
    .C(_6745_),
    .Y(_6711_[17])
);

INVX1 _16259_ (
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_6746_)
);

NAND2X1 _16260_ (
    .A(gnd),
    .B(gnd),
    .Y(_6747_)
);

OAI21X1 _16261_ (
    .A(gnd),
    .B(_6746_),
    .C(_6747_),
    .Y(_6711_[18])
);

INVX1 _16262_ (
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_6748_)
);

NAND2X1 _16263_ (
    .A(gnd),
    .B(gnd),
    .Y(_6749_)
);

OAI21X1 _16264_ (
    .A(gnd),
    .B(_6748_),
    .C(_6749_),
    .Y(_6711_[19])
);

INVX1 _16265_ (
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_6750_)
);

NAND2X1 _16266_ (
    .A(gnd),
    .B(gnd),
    .Y(_6751_)
);

OAI21X1 _16267_ (
    .A(gnd),
    .B(_6750_),
    .C(_6751_),
    .Y(_6711_[20])
);

INVX1 _16268_ (
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .Y(_6752_)
);

NAND2X1 _16269_ (
    .A(gnd),
    .B(gnd),
    .Y(_6753_)
);

OAI21X1 _16270_ (
    .A(gnd),
    .B(_6752_),
    .C(_6753_),
    .Y(_6711_[21])
);

INVX1 _16271_ (
    .A(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_6754_)
);

NAND2X1 _16272_ (
    .A(gnd),
    .B(gnd),
    .Y(_6755_)
);

OAI21X1 _16273_ (
    .A(gnd),
    .B(_6754_),
    .C(_6755_),
    .Y(_6711_[22])
);

INVX1 _16274_ (
    .A(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_6756_)
);

NAND2X1 _16275_ (
    .A(gnd),
    .B(gnd),
    .Y(_6757_)
);

OAI21X1 _16276_ (
    .A(gnd),
    .B(_6756_),
    .C(_6757_),
    .Y(_6711_[23])
);

INVX1 _16277_ (
    .A(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_6758_)
);

NAND2X1 _16278_ (
    .A(gnd),
    .B(gnd),
    .Y(_6759_)
);

OAI21X1 _16279_ (
    .A(gnd),
    .B(_6758_),
    .C(_6759_),
    .Y(_6711_[24])
);

INVX1 _16280_ (
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .Y(_6760_)
);

NAND2X1 _16281_ (
    .A(gnd),
    .B(gnd),
    .Y(_6761_)
);

OAI21X1 _16282_ (
    .A(gnd),
    .B(_6760_),
    .C(_6761_),
    .Y(_6711_[25])
);

INVX1 _16283_ (
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .Y(_6762_)
);

NAND2X1 _16284_ (
    .A(gnd),
    .B(gnd),
    .Y(_6763_)
);

OAI21X1 _16285_ (
    .A(gnd),
    .B(_6762_),
    .C(_6763_),
    .Y(_6711_[26])
);

INVX1 _16286_ (
    .A(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_6764_)
);

NAND2X1 _16287_ (
    .A(gnd),
    .B(gnd),
    .Y(_6765_)
);

OAI21X1 _16288_ (
    .A(gnd),
    .B(_6764_),
    .C(_6765_),
    .Y(_6711_[27])
);

INVX1 _16289_ (
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_6766_)
);

NAND2X1 _16290_ (
    .A(gnd),
    .B(gnd),
    .Y(_6767_)
);

OAI21X1 _16291_ (
    .A(gnd),
    .B(_6766_),
    .C(_6767_),
    .Y(_6711_[28])
);

INVX1 _16292_ (
    .A(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_6768_)
);

NAND2X1 _16293_ (
    .A(gnd),
    .B(gnd),
    .Y(_6769_)
);

OAI21X1 _16294_ (
    .A(gnd),
    .B(_6768_),
    .C(_6769_),
    .Y(_6711_[29])
);

INVX1 _16295_ (
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_6770_)
);

NAND2X1 _16296_ (
    .A(gnd),
    .B(gnd),
    .Y(_6771_)
);

OAI21X1 _16297_ (
    .A(gnd),
    .B(_6770_),
    .C(_6771_),
    .Y(_6711_[30])
);

INVX1 _16298_ (
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_6772_)
);

NAND2X1 _16299_ (
    .A(gnd),
    .B(gnd),
    .Y(_6773_)
);

OAI21X1 _16300_ (
    .A(gnd),
    .B(_6772_),
    .C(_6773_),
    .Y(_6711_[31])
);

DFFSR _16301_ (
    .CLK(clk_bF$buf35),
    .D(_6711_[0]),
    .Q(\datapath_1.regfile_1.regOut[0] [0]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _16302_ (
    .CLK(clk_bF$buf34),
    .D(_6711_[1]),
    .Q(\datapath_1.regfile_1.regOut[0] [1]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _16303_ (
    .CLK(clk_bF$buf33),
    .D(_6711_[2]),
    .Q(\datapath_1.regfile_1.regOut[0] [2]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _16304_ (
    .CLK(clk_bF$buf32),
    .D(_6711_[3]),
    .Q(\datapath_1.regfile_1.regOut[0] [3]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _16305_ (
    .CLK(clk_bF$buf31),
    .D(_6711_[4]),
    .Q(\datapath_1.regfile_1.regOut[0] [4]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _16306_ (
    .CLK(clk_bF$buf30),
    .D(_6711_[5]),
    .Q(\datapath_1.regfile_1.regOut[0] [5]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _16307_ (
    .CLK(clk_bF$buf29),
    .D(_6711_[6]),
    .Q(\datapath_1.regfile_1.regOut[0] [6]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _16308_ (
    .CLK(clk_bF$buf28),
    .D(_6711_[7]),
    .Q(\datapath_1.regfile_1.regOut[0] [7]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _16309_ (
    .CLK(clk_bF$buf27),
    .D(_6711_[8]),
    .Q(\datapath_1.regfile_1.regOut[0] [8]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _16310_ (
    .CLK(clk_bF$buf26),
    .D(_6711_[9]),
    .Q(\datapath_1.regfile_1.regOut[0] [9]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _16311_ (
    .CLK(clk_bF$buf25),
    .D(_6711_[10]),
    .Q(\datapath_1.regfile_1.regOut[0] [10]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _16312_ (
    .CLK(clk_bF$buf24),
    .D(_6711_[11]),
    .Q(\datapath_1.regfile_1.regOut[0] [11]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _16313_ (
    .CLK(clk_bF$buf23),
    .D(_6711_[12]),
    .Q(\datapath_1.regfile_1.regOut[0] [12]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _16314_ (
    .CLK(clk_bF$buf22),
    .D(_6711_[13]),
    .Q(\datapath_1.regfile_1.regOut[0] [13]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _16315_ (
    .CLK(clk_bF$buf21),
    .D(_6711_[14]),
    .Q(\datapath_1.regfile_1.regOut[0] [14]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _16316_ (
    .CLK(clk_bF$buf20),
    .D(_6711_[15]),
    .Q(\datapath_1.regfile_1.regOut[0] [15]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _16317_ (
    .CLK(clk_bF$buf19),
    .D(_6711_[16]),
    .Q(\datapath_1.regfile_1.regOut[0] [16]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _16318_ (
    .CLK(clk_bF$buf18),
    .D(_6711_[17]),
    .Q(\datapath_1.regfile_1.regOut[0] [17]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _16319_ (
    .CLK(clk_bF$buf17),
    .D(_6711_[18]),
    .Q(\datapath_1.regfile_1.regOut[0] [18]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _16320_ (
    .CLK(clk_bF$buf16),
    .D(_6711_[19]),
    .Q(\datapath_1.regfile_1.regOut[0] [19]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _16321_ (
    .CLK(clk_bF$buf15),
    .D(_6711_[20]),
    .Q(\datapath_1.regfile_1.regOut[0] [20]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _16322_ (
    .CLK(clk_bF$buf14),
    .D(_6711_[21]),
    .Q(\datapath_1.regfile_1.regOut[0] [21]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _16323_ (
    .CLK(clk_bF$buf13),
    .D(_6711_[22]),
    .Q(\datapath_1.regfile_1.regOut[0] [22]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _16324_ (
    .CLK(clk_bF$buf12),
    .D(_6711_[23]),
    .Q(\datapath_1.regfile_1.regOut[0] [23]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _16325_ (
    .CLK(clk_bF$buf11),
    .D(_6711_[24]),
    .Q(\datapath_1.regfile_1.regOut[0] [24]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _16326_ (
    .CLK(clk_bF$buf10),
    .D(_6711_[25]),
    .Q(\datapath_1.regfile_1.regOut[0] [25]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _16327_ (
    .CLK(clk_bF$buf9),
    .D(_6711_[26]),
    .Q(\datapath_1.regfile_1.regOut[0] [26]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _16328_ (
    .CLK(clk_bF$buf8),
    .D(_6711_[27]),
    .Q(\datapath_1.regfile_1.regOut[0] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _16329_ (
    .CLK(clk_bF$buf7),
    .D(_6711_[28]),
    .Q(\datapath_1.regfile_1.regOut[0] [28]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _16330_ (
    .CLK(clk_bF$buf6),
    .D(_6711_[29]),
    .Q(\datapath_1.regfile_1.regOut[0] [29]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _16331_ (
    .CLK(clk_bF$buf5),
    .D(_6711_[30]),
    .Q(\datapath_1.regfile_1.regOut[0] [30]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _16332_ (
    .CLK(clk_bF$buf4),
    .D(_6711_[31]),
    .Q(\datapath_1.regfile_1.regOut[0] [31]),
    .R(rst_bF$buf4),
    .S(vdd)
);

INVX1 _16333_ (
    .A(BranchNe),
    .Y(_6776_)
);

AOI21X1 _16334_ (
    .A(Branch),
    .B(ALUZero),
    .C(PCWrite),
    .Y(_6777_)
);

OAI21X1 _16335_ (
    .A(_6776_),
    .B(ALUZero),
    .C(_6777_),
    .Y(PCEn)
);

BUFX2 _6778_ (
    .A(gnd),
    .Y(MemRead)
);

BUFX2 _6779_ (
    .A(_0_),
    .Y(MemWrite)
);

BUFX2 _6780_ (
    .A(_1_[0]),
    .Y(memoryAddress[0])
);

BUFX2 _6781_ (
    .A(_1_[1]),
    .Y(memoryAddress[1])
);

BUFX2 _6782_ (
    .A(_1_[2]),
    .Y(memoryAddress[2])
);

BUFX2 _6783_ (
    .A(_1_[3]),
    .Y(memoryAddress[3])
);

BUFX2 _6784_ (
    .A(_1_[4]),
    .Y(memoryAddress[4])
);

BUFX2 _6785_ (
    .A(_1_[5]),
    .Y(memoryAddress[5])
);

BUFX2 _6786_ (
    .A(_1_[6]),
    .Y(memoryAddress[6])
);

BUFX2 _6787_ (
    .A(_1_[7]),
    .Y(memoryAddress[7])
);

BUFX2 _6788_ (
    .A(_1_[8]),
    .Y(memoryAddress[8])
);

BUFX2 _6789_ (
    .A(_1_[9]),
    .Y(memoryAddress[9])
);

BUFX2 _6790_ (
    .A(_1_[10]),
    .Y(memoryAddress[10])
);

BUFX2 _6791_ (
    .A(_1_[11]),
    .Y(memoryAddress[11])
);

BUFX2 _6792_ (
    .A(_1_[12]),
    .Y(memoryAddress[12])
);

BUFX2 _6793_ (
    .A(_1_[13]),
    .Y(memoryAddress[13])
);

BUFX2 _6794_ (
    .A(_1_[14]),
    .Y(memoryAddress[14])
);

BUFX2 _6795_ (
    .A(_1_[15]),
    .Y(memoryAddress[15])
);

BUFX2 _6796_ (
    .A(_1_[16]),
    .Y(memoryAddress[16])
);

BUFX2 _6797_ (
    .A(_1_[17]),
    .Y(memoryAddress[17])
);

BUFX2 _6798_ (
    .A(_1_[18]),
    .Y(memoryAddress[18])
);

BUFX2 _6799_ (
    .A(_1_[19]),
    .Y(memoryAddress[19])
);

BUFX2 _6800_ (
    .A(_1_[20]),
    .Y(memoryAddress[20])
);

BUFX2 _6801_ (
    .A(_1_[21]),
    .Y(memoryAddress[21])
);

BUFX2 _6802_ (
    .A(_1_[22]),
    .Y(memoryAddress[22])
);

BUFX2 _6803_ (
    .A(_1_[23]),
    .Y(memoryAddress[23])
);

BUFX2 _6804_ (
    .A(_1_[24]),
    .Y(memoryAddress[24])
);

BUFX2 _6805_ (
    .A(_1_[25]),
    .Y(memoryAddress[25])
);

BUFX2 _6806_ (
    .A(_1_[26]),
    .Y(memoryAddress[26])
);

BUFX2 _6807_ (
    .A(_1_[27]),
    .Y(memoryAddress[27])
);

BUFX2 _6808_ (
    .A(_1_[28]),
    .Y(memoryAddress[28])
);

BUFX2 _6809_ (
    .A(_1_[29]),
    .Y(memoryAddress[29])
);

BUFX2 _6810_ (
    .A(_1_[30]),
    .Y(memoryAddress[30])
);

BUFX2 _6811_ (
    .A(_1_[31]),
    .Y(memoryAddress[31])
);

BUFX2 _6812_ (
    .A(_2_[0]),
    .Y(memoryWriteData[0])
);

BUFX2 _6813_ (
    .A(_2_[1]),
    .Y(memoryWriteData[1])
);

BUFX2 _6814_ (
    .A(_2_[2]),
    .Y(memoryWriteData[2])
);

BUFX2 _6815_ (
    .A(_2_[3]),
    .Y(memoryWriteData[3])
);

BUFX2 _6816_ (
    .A(_2_[4]),
    .Y(memoryWriteData[4])
);

BUFX2 _6817_ (
    .A(_2_[5]),
    .Y(memoryWriteData[5])
);

BUFX2 _6818_ (
    .A(_2_[6]),
    .Y(memoryWriteData[6])
);

BUFX2 _6819_ (
    .A(_2_[7]),
    .Y(memoryWriteData[7])
);

BUFX2 _6820_ (
    .A(_2_[8]),
    .Y(memoryWriteData[8])
);

BUFX2 _6821_ (
    .A(_2_[9]),
    .Y(memoryWriteData[9])
);

BUFX2 _6822_ (
    .A(_2_[10]),
    .Y(memoryWriteData[10])
);

BUFX2 _6823_ (
    .A(_2_[11]),
    .Y(memoryWriteData[11])
);

BUFX2 _6824_ (
    .A(_2_[12]),
    .Y(memoryWriteData[12])
);

BUFX2 _6825_ (
    .A(_2_[13]),
    .Y(memoryWriteData[13])
);

BUFX2 _6826_ (
    .A(_2_[14]),
    .Y(memoryWriteData[14])
);

BUFX2 _6827_ (
    .A(_2_[15]),
    .Y(memoryWriteData[15])
);

BUFX2 _6828_ (
    .A(_2_[16]),
    .Y(memoryWriteData[16])
);

BUFX2 _6829_ (
    .A(_2_[17]),
    .Y(memoryWriteData[17])
);

BUFX2 _6830_ (
    .A(_2_[18]),
    .Y(memoryWriteData[18])
);

BUFX2 _6831_ (
    .A(_2_[19]),
    .Y(memoryWriteData[19])
);

BUFX2 _6832_ (
    .A(_2_[20]),
    .Y(memoryWriteData[20])
);

BUFX2 _6833_ (
    .A(_2_[21]),
    .Y(memoryWriteData[21])
);

BUFX2 _6834_ (
    .A(_2_[22]),
    .Y(memoryWriteData[22])
);

BUFX2 _6835_ (
    .A(_2_[23]),
    .Y(memoryWriteData[23])
);

BUFX2 _6836_ (
    .A(_2_[24]),
    .Y(memoryWriteData[24])
);

BUFX2 _6837_ (
    .A(_2_[25]),
    .Y(memoryWriteData[25])
);

BUFX2 _6838_ (
    .A(_2_[26]),
    .Y(memoryWriteData[26])
);

BUFX2 _6839_ (
    .A(_2_[27]),
    .Y(memoryWriteData[27])
);

BUFX2 _6840_ (
    .A(_2_[28]),
    .Y(memoryWriteData[28])
);

BUFX2 _6841_ (
    .A(_2_[29]),
    .Y(memoryWriteData[29])
);

BUFX2 _6842_ (
    .A(_2_[30]),
    .Y(memoryWriteData[30])
);

BUFX2 _6843_ (
    .A(_2_[31]),
    .Y(memoryWriteData[31])
);

INVX1 _6844_ (
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_66_)
);

NAND2X1 _6845_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .Y(_67_)
);

OAI21X1 _6846_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_66_),
    .C(_67_),
    .Y(_3_[0])
);

INVX1 _6847_ (
    .A(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_4_)
);

NAND2X1 _6848_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_5_)
);

OAI21X1 _6849_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_4_),
    .C(_5_),
    .Y(_3_[1])
);

INVX1 _6850_ (
    .A(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_6_)
);

NAND2X1 _6851_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_7_)
);

OAI21X1 _6852_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_6_),
    .C(_7_),
    .Y(_3_[2])
);

INVX1 _6853_ (
    .A(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_8_)
);

NAND2X1 _6854_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_9_)
);

OAI21X1 _6855_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_8_),
    .C(_9_),
    .Y(_3_[3])
);

INVX1 _6856_ (
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_10_)
);

NAND2X1 _6857_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_11_)
);

OAI21X1 _6858_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_10_),
    .C(_11_),
    .Y(_3_[4])
);

INVX1 _6859_ (
    .A(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_12_)
);

NAND2X1 _6860_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_13_)
);

OAI21X1 _6861_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_12_),
    .C(_13_),
    .Y(_3_[5])
);

INVX1 _6862_ (
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_14_)
);

NAND2X1 _6863_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_15_)
);

OAI21X1 _6864_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_14_),
    .C(_15_),
    .Y(_3_[6])
);

INVX1 _6865_ (
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_16_)
);

NAND2X1 _6866_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_17_)
);

OAI21X1 _6867_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_16_),
    .C(_17_),
    .Y(_3_[7])
);

INVX1 _6868_ (
    .A(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_18_)
);

NAND2X1 _6869_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_19_)
);

OAI21X1 _6870_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_18_),
    .C(_19_),
    .Y(_3_[8])
);

INVX1 _6871_ (
    .A(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_20_)
);

NAND2X1 _6872_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_21_)
);

OAI21X1 _6873_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_20_),
    .C(_21_),
    .Y(_3_[9])
);

INVX1 _6874_ (
    .A(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_22_)
);

NAND2X1 _6875_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_23_)
);

OAI21X1 _6876_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_22_),
    .C(_23_),
    .Y(_3_[10])
);

INVX1 _6877_ (
    .A(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_24_)
);

NAND2X1 _6878_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_25_)
);

OAI21X1 _6879_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_24_),
    .C(_25_),
    .Y(_3_[11])
);

INVX1 _6880_ (
    .A(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_26_)
);

NAND2X1 _6881_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_27_)
);

OAI21X1 _6882_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_26_),
    .C(_27_),
    .Y(_3_[12])
);

INVX1 _6883_ (
    .A(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_28_)
);

NAND2X1 _6884_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_29_)
);

OAI21X1 _6885_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_28_),
    .C(_29_),
    .Y(_3_[13])
);

INVX1 _6886_ (
    .A(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_30_)
);

NAND2X1 _6887_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_31_)
);

OAI21X1 _6888_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_30_),
    .C(_31_),
    .Y(_3_[14])
);

INVX1 _6889_ (
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_32_)
);

NAND2X1 _6890_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_33_)
);

OAI21X1 _6891_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_32_),
    .C(_33_),
    .Y(_3_[15])
);

INVX1 _6892_ (
    .A(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_34_)
);

NAND2X1 _6893_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_35_)
);

OAI21X1 _6894_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_34_),
    .C(_35_),
    .Y(_3_[16])
);

INVX1 _6895_ (
    .A(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_36_)
);

NAND2X1 _6896_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_37_)
);

OAI21X1 _6897_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_36_),
    .C(_37_),
    .Y(_3_[17])
);

INVX1 _6898_ (
    .A(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_38_)
);

NAND2X1 _6899_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_39_)
);

OAI21X1 _6900_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_38_),
    .C(_39_),
    .Y(_3_[18])
);

INVX1 _6901_ (
    .A(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_40_)
);

NAND2X1 _6902_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_41_)
);

OAI21X1 _6903_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_40_),
    .C(_41_),
    .Y(_3_[19])
);

INVX1 _6904_ (
    .A(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_42_)
);

NAND2X1 _6905_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_43_)
);

OAI21X1 _6906_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_42_),
    .C(_43_),
    .Y(_3_[20])
);

INVX1 _6907_ (
    .A(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_44_)
);

NAND2X1 _6908_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_45_)
);

OAI21X1 _6909_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_44_),
    .C(_45_),
    .Y(_3_[21])
);

INVX1 _6910_ (
    .A(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_46_)
);

NAND2X1 _6911_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_47_)
);

OAI21X1 _6912_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_46_),
    .C(_47_),
    .Y(_3_[22])
);

INVX1 _6913_ (
    .A(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_48_)
);

NAND2X1 _6914_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_49_)
);

OAI21X1 _6915_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_48_),
    .C(_49_),
    .Y(_3_[23])
);

INVX1 _6916_ (
    .A(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_50_)
);

NAND2X1 _6917_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_51_)
);

OAI21X1 _6918_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_50_),
    .C(_51_),
    .Y(_3_[24])
);

INVX1 _6919_ (
    .A(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_52_)
);

NAND2X1 _6920_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_53_)
);

OAI21X1 _6921_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_52_),
    .C(_53_),
    .Y(_3_[25])
);

INVX1 _6922_ (
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_54_)
);

NAND2X1 _6923_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_55_)
);

OAI21X1 _6924_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_54_),
    .C(_55_),
    .Y(_3_[26])
);

INVX1 _6925_ (
    .A(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_56_)
);

NAND2X1 _6926_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_57_)
);

OAI21X1 _6927_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_56_),
    .C(_57_),
    .Y(_3_[27])
);

INVX1 _6928_ (
    .A(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_58_)
);

NAND2X1 _6929_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_59_)
);

OAI21X1 _6930_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(_58_),
    .C(_59_),
    .Y(_3_[28])
);

INVX1 _6931_ (
    .A(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_60_)
);

NAND2X1 _6932_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_61_)
);

OAI21X1 _6933_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(_60_),
    .C(_61_),
    .Y(_3_[29])
);

INVX1 _6934_ (
    .A(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_62_)
);

NAND2X1 _6935_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_63_)
);

OAI21X1 _6936_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(_62_),
    .C(_63_),
    .Y(_3_[30])
);

INVX1 _6937_ (
    .A(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_64_)
);

NAND2X1 _6938_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_65_)
);

OAI21X1 _6939_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(_64_),
    .C(_65_),
    .Y(_3_[31])
);

DFFSR _6940_ (
    .CLK(clk_bF$buf3),
    .D(_3_[0]),
    .Q(\datapath_1.regfile_1.regOut[1] [0]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _6941_ (
    .CLK(clk_bF$buf2),
    .D(_3_[1]),
    .Q(\datapath_1.regfile_1.regOut[1] [1]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _6942_ (
    .CLK(clk_bF$buf1),
    .D(_3_[2]),
    .Q(\datapath_1.regfile_1.regOut[1] [2]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _6943_ (
    .CLK(clk_bF$buf0),
    .D(_3_[3]),
    .Q(\datapath_1.regfile_1.regOut[1] [3]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _6944_ (
    .CLK(clk_bF$buf113),
    .D(_3_[4]),
    .Q(\datapath_1.regfile_1.regOut[1] [4]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _6945_ (
    .CLK(clk_bF$buf112),
    .D(_3_[5]),
    .Q(\datapath_1.regfile_1.regOut[1] [5]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _6946_ (
    .CLK(clk_bF$buf111),
    .D(_3_[6]),
    .Q(\datapath_1.regfile_1.regOut[1] [6]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _6947_ (
    .CLK(clk_bF$buf110),
    .D(_3_[7]),
    .Q(\datapath_1.regfile_1.regOut[1] [7]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _6948_ (
    .CLK(clk_bF$buf109),
    .D(_3_[8]),
    .Q(\datapath_1.regfile_1.regOut[1] [8]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _6949_ (
    .CLK(clk_bF$buf108),
    .D(_3_[9]),
    .Q(\datapath_1.regfile_1.regOut[1] [9]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _6950_ (
    .CLK(clk_bF$buf107),
    .D(_3_[10]),
    .Q(\datapath_1.regfile_1.regOut[1] [10]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _6951_ (
    .CLK(clk_bF$buf106),
    .D(_3_[11]),
    .Q(\datapath_1.regfile_1.regOut[1] [11]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _6952_ (
    .CLK(clk_bF$buf105),
    .D(_3_[12]),
    .Q(\datapath_1.regfile_1.regOut[1] [12]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _6953_ (
    .CLK(clk_bF$buf104),
    .D(_3_[13]),
    .Q(\datapath_1.regfile_1.regOut[1] [13]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _6954_ (
    .CLK(clk_bF$buf103),
    .D(_3_[14]),
    .Q(\datapath_1.regfile_1.regOut[1] [14]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _6955_ (
    .CLK(clk_bF$buf102),
    .D(_3_[15]),
    .Q(\datapath_1.regfile_1.regOut[1] [15]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _6956_ (
    .CLK(clk_bF$buf101),
    .D(_3_[16]),
    .Q(\datapath_1.regfile_1.regOut[1] [16]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _6957_ (
    .CLK(clk_bF$buf100),
    .D(_3_[17]),
    .Q(\datapath_1.regfile_1.regOut[1] [17]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _6958_ (
    .CLK(clk_bF$buf99),
    .D(_3_[18]),
    .Q(\datapath_1.regfile_1.regOut[1] [18]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _6959_ (
    .CLK(clk_bF$buf98),
    .D(_3_[19]),
    .Q(\datapath_1.regfile_1.regOut[1] [19]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _6960_ (
    .CLK(clk_bF$buf97),
    .D(_3_[20]),
    .Q(\datapath_1.regfile_1.regOut[1] [20]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _6961_ (
    .CLK(clk_bF$buf96),
    .D(_3_[21]),
    .Q(\datapath_1.regfile_1.regOut[1] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _6962_ (
    .CLK(clk_bF$buf95),
    .D(_3_[22]),
    .Q(\datapath_1.regfile_1.regOut[1] [22]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _6963_ (
    .CLK(clk_bF$buf94),
    .D(_3_[23]),
    .Q(\datapath_1.regfile_1.regOut[1] [23]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _6964_ (
    .CLK(clk_bF$buf93),
    .D(_3_[24]),
    .Q(\datapath_1.regfile_1.regOut[1] [24]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _6965_ (
    .CLK(clk_bF$buf92),
    .D(_3_[25]),
    .Q(\datapath_1.regfile_1.regOut[1] [25]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _6966_ (
    .CLK(clk_bF$buf91),
    .D(_3_[26]),
    .Q(\datapath_1.regfile_1.regOut[1] [26]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _6967_ (
    .CLK(clk_bF$buf90),
    .D(_3_[27]),
    .Q(\datapath_1.regfile_1.regOut[1] [27]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _6968_ (
    .CLK(clk_bF$buf89),
    .D(_3_[28]),
    .Q(\datapath_1.regfile_1.regOut[1] [28]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _6969_ (
    .CLK(clk_bF$buf88),
    .D(_3_[29]),
    .Q(\datapath_1.regfile_1.regOut[1] [29]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _6970_ (
    .CLK(clk_bF$buf87),
    .D(_3_[30]),
    .Q(\datapath_1.regfile_1.regOut[1] [30]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _6971_ (
    .CLK(clk_bF$buf86),
    .D(_3_[31]),
    .Q(\datapath_1.regfile_1.regOut[1] [31]),
    .R(rst_bF$buf86),
    .S(vdd)
);

INVX1 _6972_ (
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_131_)
);

NAND2X1 _6973_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .Y(_132_)
);

OAI21X1 _6974_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_131_),
    .C(_132_),
    .Y(_68_[0])
);

INVX1 _6975_ (
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_69_)
);

NAND2X1 _6976_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_70_)
);

OAI21X1 _6977_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_69_),
    .C(_70_),
    .Y(_68_[1])
);

INVX1 _6978_ (
    .A(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_71_)
);

NAND2X1 _6979_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_72_)
);

OAI21X1 _6980_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_71_),
    .C(_72_),
    .Y(_68_[2])
);

INVX1 _6981_ (
    .A(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_73_)
);

NAND2X1 _6982_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_74_)
);

OAI21X1 _6983_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_73_),
    .C(_74_),
    .Y(_68_[3])
);

INVX1 _6984_ (
    .A(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_75_)
);

NAND2X1 _6985_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_76_)
);

OAI21X1 _6986_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_75_),
    .C(_76_),
    .Y(_68_[4])
);

INVX1 _6987_ (
    .A(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_77_)
);

NAND2X1 _6988_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_78_)
);

OAI21X1 _6989_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_77_),
    .C(_78_),
    .Y(_68_[5])
);

INVX1 _6990_ (
    .A(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_79_)
);

NAND2X1 _6991_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_80_)
);

OAI21X1 _6992_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_79_),
    .C(_80_),
    .Y(_68_[6])
);

INVX1 _6993_ (
    .A(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_81_)
);

NAND2X1 _6994_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_82_)
);

OAI21X1 _6995_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_81_),
    .C(_82_),
    .Y(_68_[7])
);

INVX1 _6996_ (
    .A(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_83_)
);

NAND2X1 _6997_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_84_)
);

OAI21X1 _6998_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_83_),
    .C(_84_),
    .Y(_68_[8])
);

INVX1 _6999_ (
    .A(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_85_)
);

NAND2X1 _7000_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_86_)
);

OAI21X1 _7001_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_85_),
    .C(_86_),
    .Y(_68_[9])
);

INVX1 _7002_ (
    .A(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_87_)
);

NAND2X1 _7003_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_88_)
);

OAI21X1 _7004_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_87_),
    .C(_88_),
    .Y(_68_[10])
);

INVX1 _7005_ (
    .A(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_89_)
);

NAND2X1 _7006_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_90_)
);

OAI21X1 _7007_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_89_),
    .C(_90_),
    .Y(_68_[11])
);

INVX1 _7008_ (
    .A(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_91_)
);

NAND2X1 _7009_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_92_)
);

OAI21X1 _7010_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_91_),
    .C(_92_),
    .Y(_68_[12])
);

INVX1 _7011_ (
    .A(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_93_)
);

NAND2X1 _7012_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_94_)
);

OAI21X1 _7013_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_93_),
    .C(_94_),
    .Y(_68_[13])
);

INVX1 _7014_ (
    .A(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_95_)
);

NAND2X1 _7015_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_96_)
);

OAI21X1 _7016_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_95_),
    .C(_96_),
    .Y(_68_[14])
);

INVX1 _7017_ (
    .A(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_97_)
);

NAND2X1 _7018_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_98_)
);

OAI21X1 _7019_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_97_),
    .C(_98_),
    .Y(_68_[15])
);

INVX1 _7020_ (
    .A(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_99_)
);

NAND2X1 _7021_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_100_)
);

OAI21X1 _7022_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_99_),
    .C(_100_),
    .Y(_68_[16])
);

INVX1 _7023_ (
    .A(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_101_)
);

NAND2X1 _7024_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_102_)
);

OAI21X1 _7025_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_101_),
    .C(_102_),
    .Y(_68_[17])
);

INVX1 _7026_ (
    .A(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_103_)
);

NAND2X1 _7027_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_104_)
);

OAI21X1 _7028_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_103_),
    .C(_104_),
    .Y(_68_[18])
);

INVX1 _7029_ (
    .A(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_105_)
);

NAND2X1 _7030_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_106_)
);

OAI21X1 _7031_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_105_),
    .C(_106_),
    .Y(_68_[19])
);

INVX1 _7032_ (
    .A(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_107_)
);

NAND2X1 _7033_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_108_)
);

OAI21X1 _7034_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_107_),
    .C(_108_),
    .Y(_68_[20])
);

INVX1 _7035_ (
    .A(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_109_)
);

NAND2X1 _7036_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_110_)
);

OAI21X1 _7037_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_109_),
    .C(_110_),
    .Y(_68_[21])
);

INVX1 _7038_ (
    .A(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_111_)
);

NAND2X1 _7039_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_112_)
);

OAI21X1 _7040_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_111_),
    .C(_112_),
    .Y(_68_[22])
);

INVX1 _7041_ (
    .A(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_113_)
);

NAND2X1 _7042_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_114_)
);

OAI21X1 _7043_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_113_),
    .C(_114_),
    .Y(_68_[23])
);

INVX1 _7044_ (
    .A(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_115_)
);

NAND2X1 _7045_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_116_)
);

OAI21X1 _7046_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_115_),
    .C(_116_),
    .Y(_68_[24])
);

INVX1 _7047_ (
    .A(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_117_)
);

NAND2X1 _7048_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_118_)
);

OAI21X1 _7049_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_117_),
    .C(_118_),
    .Y(_68_[25])
);

INVX1 _7050_ (
    .A(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_119_)
);

NAND2X1 _7051_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_120_)
);

OAI21X1 _7052_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_119_),
    .C(_120_),
    .Y(_68_[26])
);

INVX1 _7053_ (
    .A(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_121_)
);

NAND2X1 _7054_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_122_)
);

OAI21X1 _7055_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_121_),
    .C(_122_),
    .Y(_68_[27])
);

INVX1 _7056_ (
    .A(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_123_)
);

NAND2X1 _7057_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_124_)
);

OAI21X1 _7058_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(_123_),
    .C(_124_),
    .Y(_68_[28])
);

INVX1 _7059_ (
    .A(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_125_)
);

NAND2X1 _7060_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_126_)
);

OAI21X1 _7061_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(_125_),
    .C(_126_),
    .Y(_68_[29])
);

INVX1 _7062_ (
    .A(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_127_)
);

NAND2X1 _7063_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_128_)
);

OAI21X1 _7064_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(_127_),
    .C(_128_),
    .Y(_68_[30])
);

INVX1 _7065_ (
    .A(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_129_)
);

NAND2X1 _7066_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_130_)
);

OAI21X1 _7067_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(_129_),
    .C(_130_),
    .Y(_68_[31])
);

DFFSR _7068_ (
    .CLK(clk_bF$buf85),
    .D(_68_[0]),
    .Q(\datapath_1.regfile_1.regOut[2] [0]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _7069_ (
    .CLK(clk_bF$buf84),
    .D(_68_[1]),
    .Q(\datapath_1.regfile_1.regOut[2] [1]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _7070_ (
    .CLK(clk_bF$buf83),
    .D(_68_[2]),
    .Q(\datapath_1.regfile_1.regOut[2] [2]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _7071_ (
    .CLK(clk_bF$buf82),
    .D(_68_[3]),
    .Q(\datapath_1.regfile_1.regOut[2] [3]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _7072_ (
    .CLK(clk_bF$buf81),
    .D(_68_[4]),
    .Q(\datapath_1.regfile_1.regOut[2] [4]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _7073_ (
    .CLK(clk_bF$buf80),
    .D(_68_[5]),
    .Q(\datapath_1.regfile_1.regOut[2] [5]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _7074_ (
    .CLK(clk_bF$buf79),
    .D(_68_[6]),
    .Q(\datapath_1.regfile_1.regOut[2] [6]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _7075_ (
    .CLK(clk_bF$buf78),
    .D(_68_[7]),
    .Q(\datapath_1.regfile_1.regOut[2] [7]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _7076_ (
    .CLK(clk_bF$buf77),
    .D(_68_[8]),
    .Q(\datapath_1.regfile_1.regOut[2] [8]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _7077_ (
    .CLK(clk_bF$buf76),
    .D(_68_[9]),
    .Q(\datapath_1.regfile_1.regOut[2] [9]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _7078_ (
    .CLK(clk_bF$buf75),
    .D(_68_[10]),
    .Q(\datapath_1.regfile_1.regOut[2] [10]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _7079_ (
    .CLK(clk_bF$buf74),
    .D(_68_[11]),
    .Q(\datapath_1.regfile_1.regOut[2] [11]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _7080_ (
    .CLK(clk_bF$buf73),
    .D(_68_[12]),
    .Q(\datapath_1.regfile_1.regOut[2] [12]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _7081_ (
    .CLK(clk_bF$buf72),
    .D(_68_[13]),
    .Q(\datapath_1.regfile_1.regOut[2] [13]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _7082_ (
    .CLK(clk_bF$buf71),
    .D(_68_[14]),
    .Q(\datapath_1.regfile_1.regOut[2] [14]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _7083_ (
    .CLK(clk_bF$buf70),
    .D(_68_[15]),
    .Q(\datapath_1.regfile_1.regOut[2] [15]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _7084_ (
    .CLK(clk_bF$buf69),
    .D(_68_[16]),
    .Q(\datapath_1.regfile_1.regOut[2] [16]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _7085_ (
    .CLK(clk_bF$buf68),
    .D(_68_[17]),
    .Q(\datapath_1.regfile_1.regOut[2] [17]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _7086_ (
    .CLK(clk_bF$buf67),
    .D(_68_[18]),
    .Q(\datapath_1.regfile_1.regOut[2] [18]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _7087_ (
    .CLK(clk_bF$buf66),
    .D(_68_[19]),
    .Q(\datapath_1.regfile_1.regOut[2] [19]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _7088_ (
    .CLK(clk_bF$buf65),
    .D(_68_[20]),
    .Q(\datapath_1.regfile_1.regOut[2] [20]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _7089_ (
    .CLK(clk_bF$buf64),
    .D(_68_[21]),
    .Q(\datapath_1.regfile_1.regOut[2] [21]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _7090_ (
    .CLK(clk_bF$buf63),
    .D(_68_[22]),
    .Q(\datapath_1.regfile_1.regOut[2] [22]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _7091_ (
    .CLK(clk_bF$buf62),
    .D(_68_[23]),
    .Q(\datapath_1.regfile_1.regOut[2] [23]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _7092_ (
    .CLK(clk_bF$buf61),
    .D(_68_[24]),
    .Q(\datapath_1.regfile_1.regOut[2] [24]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _7093_ (
    .CLK(clk_bF$buf60),
    .D(_68_[25]),
    .Q(\datapath_1.regfile_1.regOut[2] [25]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _7094_ (
    .CLK(clk_bF$buf59),
    .D(_68_[26]),
    .Q(\datapath_1.regfile_1.regOut[2] [26]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _7095_ (
    .CLK(clk_bF$buf58),
    .D(_68_[27]),
    .Q(\datapath_1.regfile_1.regOut[2] [27]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _7096_ (
    .CLK(clk_bF$buf57),
    .D(_68_[28]),
    .Q(\datapath_1.regfile_1.regOut[2] [28]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _7097_ (
    .CLK(clk_bF$buf56),
    .D(_68_[29]),
    .Q(\datapath_1.regfile_1.regOut[2] [29]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _7098_ (
    .CLK(clk_bF$buf55),
    .D(_68_[30]),
    .Q(\datapath_1.regfile_1.regOut[2] [30]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _7099_ (
    .CLK(clk_bF$buf54),
    .D(_68_[31]),
    .Q(\datapath_1.regfile_1.regOut[2] [31]),
    .R(rst_bF$buf54),
    .S(vdd)
);

INVX1 _7100_ (
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .Y(_196_)
);

NAND2X1 _7101_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .Y(_197_)
);

OAI21X1 _7102_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_196_),
    .C(_197_),
    .Y(_133_[0])
);

INVX1 _7103_ (
    .A(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_134_)
);

NAND2X1 _7104_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_135_)
);

OAI21X1 _7105_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_134_),
    .C(_135_),
    .Y(_133_[1])
);

INVX1 _7106_ (
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_136_)
);

NAND2X1 _7107_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_137_)
);

OAI21X1 _7108_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_136_),
    .C(_137_),
    .Y(_133_[2])
);

INVX1 _7109_ (
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_138_)
);

NAND2X1 _7110_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_139_)
);

OAI21X1 _7111_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_138_),
    .C(_139_),
    .Y(_133_[3])
);

INVX1 _7112_ (
    .A(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_140_)
);

NAND2X1 _7113_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_141_)
);

OAI21X1 _7114_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_140_),
    .C(_141_),
    .Y(_133_[4])
);

INVX1 _7115_ (
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_142_)
);

NAND2X1 _7116_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_143_)
);

OAI21X1 _7117_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_142_),
    .C(_143_),
    .Y(_133_[5])
);

INVX1 _7118_ (
    .A(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_144_)
);

NAND2X1 _7119_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_145_)
);

OAI21X1 _7120_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_144_),
    .C(_145_),
    .Y(_133_[6])
);

INVX1 _7121_ (
    .A(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_146_)
);

NAND2X1 _7122_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_147_)
);

OAI21X1 _7123_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_146_),
    .C(_147_),
    .Y(_133_[7])
);

INVX1 _7124_ (
    .A(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_148_)
);

NAND2X1 _7125_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_149_)
);

OAI21X1 _7126_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_148_),
    .C(_149_),
    .Y(_133_[8])
);

INVX1 _7127_ (
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_150_)
);

NAND2X1 _7128_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_151_)
);

OAI21X1 _7129_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_150_),
    .C(_151_),
    .Y(_133_[9])
);

INVX1 _7130_ (
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_152_)
);

NAND2X1 _7131_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_153_)
);

OAI21X1 _7132_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_152_),
    .C(_153_),
    .Y(_133_[10])
);

INVX1 _7133_ (
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_154_)
);

NAND2X1 _7134_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_155_)
);

OAI21X1 _7135_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_154_),
    .C(_155_),
    .Y(_133_[11])
);

INVX1 _7136_ (
    .A(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_156_)
);

NAND2X1 _7137_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_157_)
);

OAI21X1 _7138_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_156_),
    .C(_157_),
    .Y(_133_[12])
);

INVX1 _7139_ (
    .A(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_158_)
);

NAND2X1 _7140_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_159_)
);

OAI21X1 _7141_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_158_),
    .C(_159_),
    .Y(_133_[13])
);

INVX1 _7142_ (
    .A(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_160_)
);

NAND2X1 _7143_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_161_)
);

OAI21X1 _7144_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_160_),
    .C(_161_),
    .Y(_133_[14])
);

INVX1 _7145_ (
    .A(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_162_)
);

NAND2X1 _7146_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_163_)
);

OAI21X1 _7147_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_162_),
    .C(_163_),
    .Y(_133_[15])
);

INVX1 _7148_ (
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_164_)
);

NAND2X1 _7149_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_165_)
);

OAI21X1 _7150_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_164_),
    .C(_165_),
    .Y(_133_[16])
);

INVX1 _7151_ (
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_166_)
);

NAND2X1 _7152_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_167_)
);

OAI21X1 _7153_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_166_),
    .C(_167_),
    .Y(_133_[17])
);

INVX1 _7154_ (
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_168_)
);

NAND2X1 _7155_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_169_)
);

OAI21X1 _7156_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_168_),
    .C(_169_),
    .Y(_133_[18])
);

INVX1 _7157_ (
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_170_)
);

NAND2X1 _7158_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_171_)
);

OAI21X1 _7159_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_170_),
    .C(_171_),
    .Y(_133_[19])
);

INVX1 _7160_ (
    .A(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_172_)
);

NAND2X1 _7161_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_173_)
);

OAI21X1 _7162_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_172_),
    .C(_173_),
    .Y(_133_[20])
);

INVX1 _7163_ (
    .A(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_174_)
);

NAND2X1 _7164_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_175_)
);

OAI21X1 _7165_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_174_),
    .C(_175_),
    .Y(_133_[21])
);

INVX1 _7166_ (
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_176_)
);

NAND2X1 _7167_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_177_)
);

OAI21X1 _7168_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_176_),
    .C(_177_),
    .Y(_133_[22])
);

INVX1 _7169_ (
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_178_)
);

NAND2X1 _7170_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_179_)
);

OAI21X1 _7171_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_178_),
    .C(_179_),
    .Y(_133_[23])
);

INVX1 _7172_ (
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_180_)
);

NAND2X1 _7173_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_181_)
);

OAI21X1 _7174_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_180_),
    .C(_181_),
    .Y(_133_[24])
);

INVX1 _7175_ (
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_182_)
);

NAND2X1 _7176_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_183_)
);

OAI21X1 _7177_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_182_),
    .C(_183_),
    .Y(_133_[25])
);

INVX1 _7178_ (
    .A(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_184_)
);

NAND2X1 _7179_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_185_)
);

OAI21X1 _7180_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_184_),
    .C(_185_),
    .Y(_133_[26])
);

INVX1 _7181_ (
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_186_)
);

NAND2X1 _7182_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_187_)
);

OAI21X1 _7183_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_186_),
    .C(_187_),
    .Y(_133_[27])
);

INVX1 _7184_ (
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_188_)
);

NAND2X1 _7185_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_189_)
);

OAI21X1 _7186_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(_188_),
    .C(_189_),
    .Y(_133_[28])
);

INVX1 _7187_ (
    .A(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_190_)
);

NAND2X1 _7188_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_191_)
);

OAI21X1 _7189_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(_190_),
    .C(_191_),
    .Y(_133_[29])
);

INVX1 _7190_ (
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_192_)
);

NAND2X1 _7191_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_193_)
);

OAI21X1 _7192_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(_192_),
    .C(_193_),
    .Y(_133_[30])
);

INVX1 _7193_ (
    .A(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_194_)
);

NAND2X1 _7194_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_195_)
);

OAI21X1 _7195_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(_194_),
    .C(_195_),
    .Y(_133_[31])
);

DFFSR _7196_ (
    .CLK(clk_bF$buf53),
    .D(_133_[0]),
    .Q(\datapath_1.regfile_1.regOut[3] [0]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _7197_ (
    .CLK(clk_bF$buf52),
    .D(_133_[1]),
    .Q(\datapath_1.regfile_1.regOut[3] [1]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _7198_ (
    .CLK(clk_bF$buf51),
    .D(_133_[2]),
    .Q(\datapath_1.regfile_1.regOut[3] [2]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _7199_ (
    .CLK(clk_bF$buf50),
    .D(_133_[3]),
    .Q(\datapath_1.regfile_1.regOut[3] [3]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _7200_ (
    .CLK(clk_bF$buf49),
    .D(_133_[4]),
    .Q(\datapath_1.regfile_1.regOut[3] [4]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _7201_ (
    .CLK(clk_bF$buf48),
    .D(_133_[5]),
    .Q(\datapath_1.regfile_1.regOut[3] [5]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _7202_ (
    .CLK(clk_bF$buf47),
    .D(_133_[6]),
    .Q(\datapath_1.regfile_1.regOut[3] [6]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _7203_ (
    .CLK(clk_bF$buf46),
    .D(_133_[7]),
    .Q(\datapath_1.regfile_1.regOut[3] [7]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _7204_ (
    .CLK(clk_bF$buf45),
    .D(_133_[8]),
    .Q(\datapath_1.regfile_1.regOut[3] [8]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _7205_ (
    .CLK(clk_bF$buf44),
    .D(_133_[9]),
    .Q(\datapath_1.regfile_1.regOut[3] [9]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _7206_ (
    .CLK(clk_bF$buf43),
    .D(_133_[10]),
    .Q(\datapath_1.regfile_1.regOut[3] [10]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _7207_ (
    .CLK(clk_bF$buf42),
    .D(_133_[11]),
    .Q(\datapath_1.regfile_1.regOut[3] [11]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _7208_ (
    .CLK(clk_bF$buf41),
    .D(_133_[12]),
    .Q(\datapath_1.regfile_1.regOut[3] [12]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _7209_ (
    .CLK(clk_bF$buf40),
    .D(_133_[13]),
    .Q(\datapath_1.regfile_1.regOut[3] [13]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _7210_ (
    .CLK(clk_bF$buf39),
    .D(_133_[14]),
    .Q(\datapath_1.regfile_1.regOut[3] [14]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _7211_ (
    .CLK(clk_bF$buf38),
    .D(_133_[15]),
    .Q(\datapath_1.regfile_1.regOut[3] [15]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _7212_ (
    .CLK(clk_bF$buf37),
    .D(_133_[16]),
    .Q(\datapath_1.regfile_1.regOut[3] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _7213_ (
    .CLK(clk_bF$buf36),
    .D(_133_[17]),
    .Q(\datapath_1.regfile_1.regOut[3] [17]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _7214_ (
    .CLK(clk_bF$buf35),
    .D(_133_[18]),
    .Q(\datapath_1.regfile_1.regOut[3] [18]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _7215_ (
    .CLK(clk_bF$buf34),
    .D(_133_[19]),
    .Q(\datapath_1.regfile_1.regOut[3] [19]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _7216_ (
    .CLK(clk_bF$buf33),
    .D(_133_[20]),
    .Q(\datapath_1.regfile_1.regOut[3] [20]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _7217_ (
    .CLK(clk_bF$buf32),
    .D(_133_[21]),
    .Q(\datapath_1.regfile_1.regOut[3] [21]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _7218_ (
    .CLK(clk_bF$buf31),
    .D(_133_[22]),
    .Q(\datapath_1.regfile_1.regOut[3] [22]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _7219_ (
    .CLK(clk_bF$buf30),
    .D(_133_[23]),
    .Q(\datapath_1.regfile_1.regOut[3] [23]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _7220_ (
    .CLK(clk_bF$buf29),
    .D(_133_[24]),
    .Q(\datapath_1.regfile_1.regOut[3] [24]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _7221_ (
    .CLK(clk_bF$buf28),
    .D(_133_[25]),
    .Q(\datapath_1.regfile_1.regOut[3] [25]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _7222_ (
    .CLK(clk_bF$buf27),
    .D(_133_[26]),
    .Q(\datapath_1.regfile_1.regOut[3] [26]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _7223_ (
    .CLK(clk_bF$buf26),
    .D(_133_[27]),
    .Q(\datapath_1.regfile_1.regOut[3] [27]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _7224_ (
    .CLK(clk_bF$buf25),
    .D(_133_[28]),
    .Q(\datapath_1.regfile_1.regOut[3] [28]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _7225_ (
    .CLK(clk_bF$buf24),
    .D(_133_[29]),
    .Q(\datapath_1.regfile_1.regOut[3] [29]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _7226_ (
    .CLK(clk_bF$buf23),
    .D(_133_[30]),
    .Q(\datapath_1.regfile_1.regOut[3] [30]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _7227_ (
    .CLK(clk_bF$buf22),
    .D(_133_[31]),
    .Q(\datapath_1.regfile_1.regOut[3] [31]),
    .R(rst_bF$buf22),
    .S(vdd)
);

INVX1 _7228_ (
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_261_)
);

NAND2X1 _7229_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .Y(_262_)
);

OAI21X1 _7230_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_261_),
    .C(_262_),
    .Y(_198_[0])
);

INVX1 _7231_ (
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_199_)
);

NAND2X1 _7232_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_200_)
);

OAI21X1 _7233_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_199_),
    .C(_200_),
    .Y(_198_[1])
);

INVX1 _7234_ (
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_201_)
);

NAND2X1 _7235_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_202_)
);

OAI21X1 _7236_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_201_),
    .C(_202_),
    .Y(_198_[2])
);

INVX1 _7237_ (
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_203_)
);

NAND2X1 _7238_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_204_)
);

OAI21X1 _7239_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_203_),
    .C(_204_),
    .Y(_198_[3])
);

INVX1 _7240_ (
    .A(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_205_)
);

NAND2X1 _7241_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_206_)
);

OAI21X1 _7242_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_205_),
    .C(_206_),
    .Y(_198_[4])
);

INVX1 _7243_ (
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .Y(_207_)
);

NAND2X1 _7244_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_208_)
);

OAI21X1 _7245_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_207_),
    .C(_208_),
    .Y(_198_[5])
);

INVX1 _7246_ (
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_209_)
);

NAND2X1 _7247_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_210_)
);

OAI21X1 _7248_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_209_),
    .C(_210_),
    .Y(_198_[6])
);

INVX1 _7249_ (
    .A(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_211_)
);

NAND2X1 _7250_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_212_)
);

OAI21X1 _7251_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_211_),
    .C(_212_),
    .Y(_198_[7])
);

INVX1 _7252_ (
    .A(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_213_)
);

NAND2X1 _7253_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_214_)
);

OAI21X1 _7254_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_213_),
    .C(_214_),
    .Y(_198_[8])
);

INVX1 _7255_ (
    .A(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_215_)
);

NAND2X1 _7256_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_216_)
);

OAI21X1 _7257_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_215_),
    .C(_216_),
    .Y(_198_[9])
);

INVX1 _7258_ (
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_217_)
);

NAND2X1 _7259_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_218_)
);

OAI21X1 _7260_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_217_),
    .C(_218_),
    .Y(_198_[10])
);

INVX1 _7261_ (
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_219_)
);

NAND2X1 _7262_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_220_)
);

OAI21X1 _7263_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_219_),
    .C(_220_),
    .Y(_198_[11])
);

INVX1 _7264_ (
    .A(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_221_)
);

NAND2X1 _7265_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_222_)
);

OAI21X1 _7266_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_221_),
    .C(_222_),
    .Y(_198_[12])
);

INVX1 _7267_ (
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_223_)
);

NAND2X1 _7268_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_224_)
);

OAI21X1 _7269_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_223_),
    .C(_224_),
    .Y(_198_[13])
);

INVX1 _7270_ (
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_225_)
);

NAND2X1 _7271_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_226_)
);

OAI21X1 _7272_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_225_),
    .C(_226_),
    .Y(_198_[14])
);

INVX1 _7273_ (
    .A(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_227_)
);

NAND2X1 _7274_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_228_)
);

OAI21X1 _7275_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_227_),
    .C(_228_),
    .Y(_198_[15])
);

INVX1 _7276_ (
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_229_)
);

NAND2X1 _7277_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_230_)
);

OAI21X1 _7278_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_229_),
    .C(_230_),
    .Y(_198_[16])
);

INVX1 _7279_ (
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_231_)
);

NAND2X1 _7280_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_232_)
);

OAI21X1 _7281_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_231_),
    .C(_232_),
    .Y(_198_[17])
);

INVX1 _7282_ (
    .A(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_233_)
);

NAND2X1 _7283_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_234_)
);

OAI21X1 _7284_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_233_),
    .C(_234_),
    .Y(_198_[18])
);

INVX1 _7285_ (
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_235_)
);

NAND2X1 _7286_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_236_)
);

OAI21X1 _7287_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_235_),
    .C(_236_),
    .Y(_198_[19])
);

INVX1 _7288_ (
    .A(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_237_)
);

NAND2X1 _7289_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_238_)
);

OAI21X1 _7290_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_237_),
    .C(_238_),
    .Y(_198_[20])
);

INVX1 _7291_ (
    .A(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_239_)
);

NAND2X1 _7292_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_240_)
);

OAI21X1 _7293_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_239_),
    .C(_240_),
    .Y(_198_[21])
);

INVX1 _7294_ (
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_241_)
);

NAND2X1 _7295_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_242_)
);

OAI21X1 _7296_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_241_),
    .C(_242_),
    .Y(_198_[22])
);

INVX1 _7297_ (
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_243_)
);

NAND2X1 _7298_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_244_)
);

OAI21X1 _7299_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_243_),
    .C(_244_),
    .Y(_198_[23])
);

INVX1 _7300_ (
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_245_)
);

NAND2X1 _7301_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_246_)
);

OAI21X1 _7302_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_245_),
    .C(_246_),
    .Y(_198_[24])
);

INVX1 _7303_ (
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_247_)
);

NAND2X1 _7304_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_248_)
);

OAI21X1 _7305_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_247_),
    .C(_248_),
    .Y(_198_[25])
);

INVX1 _7306_ (
    .A(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_249_)
);

NAND2X1 _7307_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_250_)
);

OAI21X1 _7308_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_249_),
    .C(_250_),
    .Y(_198_[26])
);

INVX1 _7309_ (
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_251_)
);

NAND2X1 _7310_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_252_)
);

OAI21X1 _7311_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_251_),
    .C(_252_),
    .Y(_198_[27])
);

INVX1 _7312_ (
    .A(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_253_)
);

NAND2X1 _7313_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_254_)
);

OAI21X1 _7314_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(_253_),
    .C(_254_),
    .Y(_198_[28])
);

INVX1 _7315_ (
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_255_)
);

NAND2X1 _7316_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_256_)
);

OAI21X1 _7317_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(_255_),
    .C(_256_),
    .Y(_198_[29])
);

INVX1 _7318_ (
    .A(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_257_)
);

NAND2X1 _7319_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_258_)
);

OAI21X1 _7320_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(_257_),
    .C(_258_),
    .Y(_198_[30])
);

INVX1 _7321_ (
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_259_)
);

NAND2X1 _7322_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_260_)
);

OAI21X1 _7323_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(_259_),
    .C(_260_),
    .Y(_198_[31])
);

DFFSR _7324_ (
    .CLK(clk_bF$buf21),
    .D(_198_[0]),
    .Q(\datapath_1.regfile_1.regOut[4] [0]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _7325_ (
    .CLK(clk_bF$buf20),
    .D(_198_[1]),
    .Q(\datapath_1.regfile_1.regOut[4] [1]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _7326_ (
    .CLK(clk_bF$buf19),
    .D(_198_[2]),
    .Q(\datapath_1.regfile_1.regOut[4] [2]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _7327_ (
    .CLK(clk_bF$buf18),
    .D(_198_[3]),
    .Q(\datapath_1.regfile_1.regOut[4] [3]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _7328_ (
    .CLK(clk_bF$buf17),
    .D(_198_[4]),
    .Q(\datapath_1.regfile_1.regOut[4] [4]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _7329_ (
    .CLK(clk_bF$buf16),
    .D(_198_[5]),
    .Q(\datapath_1.regfile_1.regOut[4] [5]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _7330_ (
    .CLK(clk_bF$buf15),
    .D(_198_[6]),
    .Q(\datapath_1.regfile_1.regOut[4] [6]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _7331_ (
    .CLK(clk_bF$buf14),
    .D(_198_[7]),
    .Q(\datapath_1.regfile_1.regOut[4] [7]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _7332_ (
    .CLK(clk_bF$buf13),
    .D(_198_[8]),
    .Q(\datapath_1.regfile_1.regOut[4] [8]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _7333_ (
    .CLK(clk_bF$buf12),
    .D(_198_[9]),
    .Q(\datapath_1.regfile_1.regOut[4] [9]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _7334_ (
    .CLK(clk_bF$buf11),
    .D(_198_[10]),
    .Q(\datapath_1.regfile_1.regOut[4] [10]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _7335_ (
    .CLK(clk_bF$buf10),
    .D(_198_[11]),
    .Q(\datapath_1.regfile_1.regOut[4] [11]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _7336_ (
    .CLK(clk_bF$buf9),
    .D(_198_[12]),
    .Q(\datapath_1.regfile_1.regOut[4] [12]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _7337_ (
    .CLK(clk_bF$buf8),
    .D(_198_[13]),
    .Q(\datapath_1.regfile_1.regOut[4] [13]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _7338_ (
    .CLK(clk_bF$buf7),
    .D(_198_[14]),
    .Q(\datapath_1.regfile_1.regOut[4] [14]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _7339_ (
    .CLK(clk_bF$buf6),
    .D(_198_[15]),
    .Q(\datapath_1.regfile_1.regOut[4] [15]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _7340_ (
    .CLK(clk_bF$buf5),
    .D(_198_[16]),
    .Q(\datapath_1.regfile_1.regOut[4] [16]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _7341_ (
    .CLK(clk_bF$buf4),
    .D(_198_[17]),
    .Q(\datapath_1.regfile_1.regOut[4] [17]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _7342_ (
    .CLK(clk_bF$buf3),
    .D(_198_[18]),
    .Q(\datapath_1.regfile_1.regOut[4] [18]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _7343_ (
    .CLK(clk_bF$buf2),
    .D(_198_[19]),
    .Q(\datapath_1.regfile_1.regOut[4] [19]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _7344_ (
    .CLK(clk_bF$buf1),
    .D(_198_[20]),
    .Q(\datapath_1.regfile_1.regOut[4] [20]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _7345_ (
    .CLK(clk_bF$buf0),
    .D(_198_[21]),
    .Q(\datapath_1.regfile_1.regOut[4] [21]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _7346_ (
    .CLK(clk_bF$buf113),
    .D(_198_[22]),
    .Q(\datapath_1.regfile_1.regOut[4] [22]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _7347_ (
    .CLK(clk_bF$buf112),
    .D(_198_[23]),
    .Q(\datapath_1.regfile_1.regOut[4] [23]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _7348_ (
    .CLK(clk_bF$buf111),
    .D(_198_[24]),
    .Q(\datapath_1.regfile_1.regOut[4] [24]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _7349_ (
    .CLK(clk_bF$buf110),
    .D(_198_[25]),
    .Q(\datapath_1.regfile_1.regOut[4] [25]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _7350_ (
    .CLK(clk_bF$buf109),
    .D(_198_[26]),
    .Q(\datapath_1.regfile_1.regOut[4] [26]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _7351_ (
    .CLK(clk_bF$buf108),
    .D(_198_[27]),
    .Q(\datapath_1.regfile_1.regOut[4] [27]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _7352_ (
    .CLK(clk_bF$buf107),
    .D(_198_[28]),
    .Q(\datapath_1.regfile_1.regOut[4] [28]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _7353_ (
    .CLK(clk_bF$buf106),
    .D(_198_[29]),
    .Q(\datapath_1.regfile_1.regOut[4] [29]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _7354_ (
    .CLK(clk_bF$buf105),
    .D(_198_[30]),
    .Q(\datapath_1.regfile_1.regOut[4] [30]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _7355_ (
    .CLK(clk_bF$buf104),
    .D(_198_[31]),
    .Q(\datapath_1.regfile_1.regOut[4] [31]),
    .R(rst_bF$buf104),
    .S(vdd)
);

INVX1 _7356_ (
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_326_)
);

NAND2X1 _7357_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .Y(_327_)
);

OAI21X1 _7358_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_326_),
    .C(_327_),
    .Y(_263_[0])
);

INVX1 _7359_ (
    .A(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_264_)
);

NAND2X1 _7360_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_265_)
);

OAI21X1 _7361_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_264_),
    .C(_265_),
    .Y(_263_[1])
);

INVX1 _7362_ (
    .A(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_266_)
);

NAND2X1 _7363_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_267_)
);

OAI21X1 _7364_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_266_),
    .C(_267_),
    .Y(_263_[2])
);

INVX1 _7365_ (
    .A(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_268_)
);

NAND2X1 _7366_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_269_)
);

OAI21X1 _7367_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_268_),
    .C(_269_),
    .Y(_263_[3])
);

INVX1 _7368_ (
    .A(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_270_)
);

NAND2X1 _7369_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_271_)
);

OAI21X1 _7370_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_270_),
    .C(_271_),
    .Y(_263_[4])
);

INVX1 _7371_ (
    .A(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_272_)
);

NAND2X1 _7372_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_273_)
);

OAI21X1 _7373_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_272_),
    .C(_273_),
    .Y(_263_[5])
);

INVX1 _7374_ (
    .A(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_274_)
);

NAND2X1 _7375_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_275_)
);

OAI21X1 _7376_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_274_),
    .C(_275_),
    .Y(_263_[6])
);

INVX1 _7377_ (
    .A(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_276_)
);

NAND2X1 _7378_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_277_)
);

OAI21X1 _7379_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_276_),
    .C(_277_),
    .Y(_263_[7])
);

INVX1 _7380_ (
    .A(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_278_)
);

NAND2X1 _7381_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_279_)
);

OAI21X1 _7382_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_278_),
    .C(_279_),
    .Y(_263_[8])
);

INVX1 _7383_ (
    .A(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_280_)
);

NAND2X1 _7384_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_281_)
);

OAI21X1 _7385_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_280_),
    .C(_281_),
    .Y(_263_[9])
);

INVX1 _7386_ (
    .A(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_282_)
);

NAND2X1 _7387_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_283_)
);

OAI21X1 _7388_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_282_),
    .C(_283_),
    .Y(_263_[10])
);

INVX1 _7389_ (
    .A(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_284_)
);

NAND2X1 _7390_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_285_)
);

OAI21X1 _7391_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_284_),
    .C(_285_),
    .Y(_263_[11])
);

INVX1 _7392_ (
    .A(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_286_)
);

NAND2X1 _7393_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_287_)
);

OAI21X1 _7394_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_286_),
    .C(_287_),
    .Y(_263_[12])
);

INVX1 _7395_ (
    .A(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_288_)
);

NAND2X1 _7396_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_289_)
);

OAI21X1 _7397_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_288_),
    .C(_289_),
    .Y(_263_[13])
);

INVX1 _7398_ (
    .A(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_290_)
);

NAND2X1 _7399_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_291_)
);

OAI21X1 _7400_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_290_),
    .C(_291_),
    .Y(_263_[14])
);

INVX1 _7401_ (
    .A(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_292_)
);

NAND2X1 _7402_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_293_)
);

OAI21X1 _7403_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_292_),
    .C(_293_),
    .Y(_263_[15])
);

INVX1 _7404_ (
    .A(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_294_)
);

NAND2X1 _7405_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_295_)
);

OAI21X1 _7406_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_294_),
    .C(_295_),
    .Y(_263_[16])
);

INVX1 _7407_ (
    .A(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_296_)
);

NAND2X1 _7408_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_297_)
);

OAI21X1 _7409_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_296_),
    .C(_297_),
    .Y(_263_[17])
);

INVX1 _7410_ (
    .A(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_298_)
);

NAND2X1 _7411_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_299_)
);

OAI21X1 _7412_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_298_),
    .C(_299_),
    .Y(_263_[18])
);

INVX1 _7413_ (
    .A(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_300_)
);

NAND2X1 _7414_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_301_)
);

OAI21X1 _7415_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_300_),
    .C(_301_),
    .Y(_263_[19])
);

INVX1 _7416_ (
    .A(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_302_)
);

NAND2X1 _7417_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_303_)
);

OAI21X1 _7418_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_302_),
    .C(_303_),
    .Y(_263_[20])
);

INVX1 _7419_ (
    .A(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_304_)
);

NAND2X1 _7420_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_305_)
);

OAI21X1 _7421_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_304_),
    .C(_305_),
    .Y(_263_[21])
);

INVX1 _7422_ (
    .A(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_306_)
);

NAND2X1 _7423_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_307_)
);

OAI21X1 _7424_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_306_),
    .C(_307_),
    .Y(_263_[22])
);

INVX1 _7425_ (
    .A(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_308_)
);

NAND2X1 _7426_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_309_)
);

OAI21X1 _7427_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_308_),
    .C(_309_),
    .Y(_263_[23])
);

INVX1 _7428_ (
    .A(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_310_)
);

NAND2X1 _7429_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_311_)
);

OAI21X1 _7430_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_310_),
    .C(_311_),
    .Y(_263_[24])
);

INVX1 _7431_ (
    .A(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_312_)
);

NAND2X1 _7432_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_313_)
);

OAI21X1 _7433_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_312_),
    .C(_313_),
    .Y(_263_[25])
);

INVX1 _7434_ (
    .A(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_314_)
);

NAND2X1 _7435_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_315_)
);

OAI21X1 _7436_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_314_),
    .C(_315_),
    .Y(_263_[26])
);

INVX1 _7437_ (
    .A(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_316_)
);

NAND2X1 _7438_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_317_)
);

OAI21X1 _7439_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_316_),
    .C(_317_),
    .Y(_263_[27])
);

INVX1 _7440_ (
    .A(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_318_)
);

NAND2X1 _7441_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_319_)
);

OAI21X1 _7442_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(_318_),
    .C(_319_),
    .Y(_263_[28])
);

INVX1 _7443_ (
    .A(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_320_)
);

NAND2X1 _7444_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_321_)
);

OAI21X1 _7445_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(_320_),
    .C(_321_),
    .Y(_263_[29])
);

INVX1 _7446_ (
    .A(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_322_)
);

NAND2X1 _7447_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_323_)
);

OAI21X1 _7448_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(_322_),
    .C(_323_),
    .Y(_263_[30])
);

INVX1 _7449_ (
    .A(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_324_)
);

NAND2X1 _7450_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_325_)
);

OAI21X1 _7451_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(_324_),
    .C(_325_),
    .Y(_263_[31])
);

DFFSR _7452_ (
    .CLK(clk_bF$buf103),
    .D(_263_[0]),
    .Q(\datapath_1.regfile_1.regOut[5] [0]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _7453_ (
    .CLK(clk_bF$buf102),
    .D(_263_[1]),
    .Q(\datapath_1.regfile_1.regOut[5] [1]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _7454_ (
    .CLK(clk_bF$buf101),
    .D(_263_[2]),
    .Q(\datapath_1.regfile_1.regOut[5] [2]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _7455_ (
    .CLK(clk_bF$buf100),
    .D(_263_[3]),
    .Q(\datapath_1.regfile_1.regOut[5] [3]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _7456_ (
    .CLK(clk_bF$buf99),
    .D(_263_[4]),
    .Q(\datapath_1.regfile_1.regOut[5] [4]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _7457_ (
    .CLK(clk_bF$buf98),
    .D(_263_[5]),
    .Q(\datapath_1.regfile_1.regOut[5] [5]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _7458_ (
    .CLK(clk_bF$buf97),
    .D(_263_[6]),
    .Q(\datapath_1.regfile_1.regOut[5] [6]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _7459_ (
    .CLK(clk_bF$buf96),
    .D(_263_[7]),
    .Q(\datapath_1.regfile_1.regOut[5] [7]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _7460_ (
    .CLK(clk_bF$buf95),
    .D(_263_[8]),
    .Q(\datapath_1.regfile_1.regOut[5] [8]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _7461_ (
    .CLK(clk_bF$buf94),
    .D(_263_[9]),
    .Q(\datapath_1.regfile_1.regOut[5] [9]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _7462_ (
    .CLK(clk_bF$buf93),
    .D(_263_[10]),
    .Q(\datapath_1.regfile_1.regOut[5] [10]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _7463_ (
    .CLK(clk_bF$buf92),
    .D(_263_[11]),
    .Q(\datapath_1.regfile_1.regOut[5] [11]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _7464_ (
    .CLK(clk_bF$buf91),
    .D(_263_[12]),
    .Q(\datapath_1.regfile_1.regOut[5] [12]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _7465_ (
    .CLK(clk_bF$buf90),
    .D(_263_[13]),
    .Q(\datapath_1.regfile_1.regOut[5] [13]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _7466_ (
    .CLK(clk_bF$buf89),
    .D(_263_[14]),
    .Q(\datapath_1.regfile_1.regOut[5] [14]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _7467_ (
    .CLK(clk_bF$buf88),
    .D(_263_[15]),
    .Q(\datapath_1.regfile_1.regOut[5] [15]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _7468_ (
    .CLK(clk_bF$buf87),
    .D(_263_[16]),
    .Q(\datapath_1.regfile_1.regOut[5] [16]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _7469_ (
    .CLK(clk_bF$buf86),
    .D(_263_[17]),
    .Q(\datapath_1.regfile_1.regOut[5] [17]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _7470_ (
    .CLK(clk_bF$buf85),
    .D(_263_[18]),
    .Q(\datapath_1.regfile_1.regOut[5] [18]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _7471_ (
    .CLK(clk_bF$buf84),
    .D(_263_[19]),
    .Q(\datapath_1.regfile_1.regOut[5] [19]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _7472_ (
    .CLK(clk_bF$buf83),
    .D(_263_[20]),
    .Q(\datapath_1.regfile_1.regOut[5] [20]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _7473_ (
    .CLK(clk_bF$buf82),
    .D(_263_[21]),
    .Q(\datapath_1.regfile_1.regOut[5] [21]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _7474_ (
    .CLK(clk_bF$buf81),
    .D(_263_[22]),
    .Q(\datapath_1.regfile_1.regOut[5] [22]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _7475_ (
    .CLK(clk_bF$buf80),
    .D(_263_[23]),
    .Q(\datapath_1.regfile_1.regOut[5] [23]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _7476_ (
    .CLK(clk_bF$buf79),
    .D(_263_[24]),
    .Q(\datapath_1.regfile_1.regOut[5] [24]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _7477_ (
    .CLK(clk_bF$buf78),
    .D(_263_[25]),
    .Q(\datapath_1.regfile_1.regOut[5] [25]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _7478_ (
    .CLK(clk_bF$buf77),
    .D(_263_[26]),
    .Q(\datapath_1.regfile_1.regOut[5] [26]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _7479_ (
    .CLK(clk_bF$buf76),
    .D(_263_[27]),
    .Q(\datapath_1.regfile_1.regOut[5] [27]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _7480_ (
    .CLK(clk_bF$buf75),
    .D(_263_[28]),
    .Q(\datapath_1.regfile_1.regOut[5] [28]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _7481_ (
    .CLK(clk_bF$buf74),
    .D(_263_[29]),
    .Q(\datapath_1.regfile_1.regOut[5] [29]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _7482_ (
    .CLK(clk_bF$buf73),
    .D(_263_[30]),
    .Q(\datapath_1.regfile_1.regOut[5] [30]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _7483_ (
    .CLK(clk_bF$buf72),
    .D(_263_[31]),
    .Q(\datapath_1.regfile_1.regOut[5] [31]),
    .R(rst_bF$buf72),
    .S(vdd)
);

INVX1 _7484_ (
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_391_)
);

NAND2X1 _7485_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .Y(_392_)
);

OAI21X1 _7486_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_391_),
    .C(_392_),
    .Y(_328_[0])
);

INVX1 _7487_ (
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_329_)
);

NAND2X1 _7488_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_330_)
);

OAI21X1 _7489_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_329_),
    .C(_330_),
    .Y(_328_[1])
);

INVX1 _7490_ (
    .A(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_331_)
);

NAND2X1 _7491_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_332_)
);

OAI21X1 _7492_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_331_),
    .C(_332_),
    .Y(_328_[2])
);

INVX1 _7493_ (
    .A(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_333_)
);

NAND2X1 _7494_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_334_)
);

OAI21X1 _7495_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_333_),
    .C(_334_),
    .Y(_328_[3])
);

INVX1 _7496_ (
    .A(\datapath_1.regfile_1.regOut[6] [4]),
    .Y(_335_)
);

NAND2X1 _7497_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_336_)
);

OAI21X1 _7498_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_335_),
    .C(_336_),
    .Y(_328_[4])
);

INVX1 _7499_ (
    .A(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_337_)
);

NAND2X1 _7500_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_338_)
);

OAI21X1 _7501_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_337_),
    .C(_338_),
    .Y(_328_[5])
);

INVX1 _7502_ (
    .A(\datapath_1.regfile_1.regOut[6] [6]),
    .Y(_339_)
);

NAND2X1 _7503_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_340_)
);

OAI21X1 _7504_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_339_),
    .C(_340_),
    .Y(_328_[6])
);

INVX1 _7505_ (
    .A(\datapath_1.regfile_1.regOut[6] [7]),
    .Y(_341_)
);

NAND2X1 _7506_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_342_)
);

OAI21X1 _7507_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_341_),
    .C(_342_),
    .Y(_328_[7])
);

INVX1 _7508_ (
    .A(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_343_)
);

NAND2X1 _7509_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_344_)
);

OAI21X1 _7510_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_343_),
    .C(_344_),
    .Y(_328_[8])
);

INVX1 _7511_ (
    .A(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_345_)
);

NAND2X1 _7512_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_346_)
);

OAI21X1 _7513_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_345_),
    .C(_346_),
    .Y(_328_[9])
);

INVX1 _7514_ (
    .A(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_347_)
);

NAND2X1 _7515_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_348_)
);

OAI21X1 _7516_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_347_),
    .C(_348_),
    .Y(_328_[10])
);

INVX1 _7517_ (
    .A(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_349_)
);

NAND2X1 _7518_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_350_)
);

OAI21X1 _7519_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_349_),
    .C(_350_),
    .Y(_328_[11])
);

INVX1 _7520_ (
    .A(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_351_)
);

NAND2X1 _7521_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_352_)
);

OAI21X1 _7522_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_351_),
    .C(_352_),
    .Y(_328_[12])
);

INVX1 _7523_ (
    .A(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_353_)
);

NAND2X1 _7524_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_354_)
);

OAI21X1 _7525_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_353_),
    .C(_354_),
    .Y(_328_[13])
);

INVX1 _7526_ (
    .A(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_355_)
);

NAND2X1 _7527_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_356_)
);

OAI21X1 _7528_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_355_),
    .C(_356_),
    .Y(_328_[14])
);

INVX1 _7529_ (
    .A(\datapath_1.regfile_1.regOut[6] [15]),
    .Y(_357_)
);

NAND2X1 _7530_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_358_)
);

OAI21X1 _7531_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_357_),
    .C(_358_),
    .Y(_328_[15])
);

INVX1 _7532_ (
    .A(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_359_)
);

NAND2X1 _7533_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_360_)
);

OAI21X1 _7534_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_359_),
    .C(_360_),
    .Y(_328_[16])
);

INVX1 _7535_ (
    .A(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_361_)
);

NAND2X1 _7536_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_362_)
);

OAI21X1 _7537_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_361_),
    .C(_362_),
    .Y(_328_[17])
);

INVX1 _7538_ (
    .A(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_363_)
);

NAND2X1 _7539_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_364_)
);

OAI21X1 _7540_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_363_),
    .C(_364_),
    .Y(_328_[18])
);

INVX1 _7541_ (
    .A(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_365_)
);

NAND2X1 _7542_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_366_)
);

OAI21X1 _7543_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_365_),
    .C(_366_),
    .Y(_328_[19])
);

INVX1 _7544_ (
    .A(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_367_)
);

NAND2X1 _7545_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_368_)
);

OAI21X1 _7546_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_367_),
    .C(_368_),
    .Y(_328_[20])
);

INVX1 _7547_ (
    .A(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_369_)
);

NAND2X1 _7548_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_370_)
);

OAI21X1 _7549_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_369_),
    .C(_370_),
    .Y(_328_[21])
);

INVX1 _7550_ (
    .A(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_371_)
);

NAND2X1 _7551_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_372_)
);

OAI21X1 _7552_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_371_),
    .C(_372_),
    .Y(_328_[22])
);

INVX1 _7553_ (
    .A(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_373_)
);

NAND2X1 _7554_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_374_)
);

OAI21X1 _7555_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_373_),
    .C(_374_),
    .Y(_328_[23])
);

INVX1 _7556_ (
    .A(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_375_)
);

NAND2X1 _7557_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_376_)
);

OAI21X1 _7558_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_375_),
    .C(_376_),
    .Y(_328_[24])
);

INVX1 _7559_ (
    .A(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_377_)
);

NAND2X1 _7560_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_378_)
);

OAI21X1 _7561_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_377_),
    .C(_378_),
    .Y(_328_[25])
);

INVX1 _7562_ (
    .A(\datapath_1.regfile_1.regOut[6] [26]),
    .Y(_379_)
);

NAND2X1 _7563_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_380_)
);

OAI21X1 _7564_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_379_),
    .C(_380_),
    .Y(_328_[26])
);

INVX1 _7565_ (
    .A(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_381_)
);

NAND2X1 _7566_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_382_)
);

OAI21X1 _7567_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_381_),
    .C(_382_),
    .Y(_328_[27])
);

INVX1 _7568_ (
    .A(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_383_)
);

NAND2X1 _7569_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_384_)
);

OAI21X1 _7570_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(_383_),
    .C(_384_),
    .Y(_328_[28])
);

INVX1 _7571_ (
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_385_)
);

NAND2X1 _7572_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_386_)
);

OAI21X1 _7573_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(_385_),
    .C(_386_),
    .Y(_328_[29])
);

INVX1 _7574_ (
    .A(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_387_)
);

NAND2X1 _7575_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_388_)
);

OAI21X1 _7576_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(_387_),
    .C(_388_),
    .Y(_328_[30])
);

INVX1 _7577_ (
    .A(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_389_)
);

NAND2X1 _7578_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_390_)
);

OAI21X1 _7579_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(_389_),
    .C(_390_),
    .Y(_328_[31])
);

DFFSR _7580_ (
    .CLK(clk_bF$buf71),
    .D(_328_[0]),
    .Q(\datapath_1.regfile_1.regOut[6] [0]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _7581_ (
    .CLK(clk_bF$buf70),
    .D(_328_[1]),
    .Q(\datapath_1.regfile_1.regOut[6] [1]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _7582_ (
    .CLK(clk_bF$buf69),
    .D(_328_[2]),
    .Q(\datapath_1.regfile_1.regOut[6] [2]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _7583_ (
    .CLK(clk_bF$buf68),
    .D(_328_[3]),
    .Q(\datapath_1.regfile_1.regOut[6] [3]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _7584_ (
    .CLK(clk_bF$buf67),
    .D(_328_[4]),
    .Q(\datapath_1.regfile_1.regOut[6] [4]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _7585_ (
    .CLK(clk_bF$buf66),
    .D(_328_[5]),
    .Q(\datapath_1.regfile_1.regOut[6] [5]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _7586_ (
    .CLK(clk_bF$buf65),
    .D(_328_[6]),
    .Q(\datapath_1.regfile_1.regOut[6] [6]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _7587_ (
    .CLK(clk_bF$buf64),
    .D(_328_[7]),
    .Q(\datapath_1.regfile_1.regOut[6] [7]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _7588_ (
    .CLK(clk_bF$buf63),
    .D(_328_[8]),
    .Q(\datapath_1.regfile_1.regOut[6] [8]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _7589_ (
    .CLK(clk_bF$buf62),
    .D(_328_[9]),
    .Q(\datapath_1.regfile_1.regOut[6] [9]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _7590_ (
    .CLK(clk_bF$buf61),
    .D(_328_[10]),
    .Q(\datapath_1.regfile_1.regOut[6] [10]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _7591_ (
    .CLK(clk_bF$buf60),
    .D(_328_[11]),
    .Q(\datapath_1.regfile_1.regOut[6] [11]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _7592_ (
    .CLK(clk_bF$buf59),
    .D(_328_[12]),
    .Q(\datapath_1.regfile_1.regOut[6] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _7593_ (
    .CLK(clk_bF$buf58),
    .D(_328_[13]),
    .Q(\datapath_1.regfile_1.regOut[6] [13]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _7594_ (
    .CLK(clk_bF$buf57),
    .D(_328_[14]),
    .Q(\datapath_1.regfile_1.regOut[6] [14]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _7595_ (
    .CLK(clk_bF$buf56),
    .D(_328_[15]),
    .Q(\datapath_1.regfile_1.regOut[6] [15]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _7596_ (
    .CLK(clk_bF$buf55),
    .D(_328_[16]),
    .Q(\datapath_1.regfile_1.regOut[6] [16]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _7597_ (
    .CLK(clk_bF$buf54),
    .D(_328_[17]),
    .Q(\datapath_1.regfile_1.regOut[6] [17]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _7598_ (
    .CLK(clk_bF$buf53),
    .D(_328_[18]),
    .Q(\datapath_1.regfile_1.regOut[6] [18]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _7599_ (
    .CLK(clk_bF$buf52),
    .D(_328_[19]),
    .Q(\datapath_1.regfile_1.regOut[6] [19]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _7600_ (
    .CLK(clk_bF$buf51),
    .D(_328_[20]),
    .Q(\datapath_1.regfile_1.regOut[6] [20]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _7601_ (
    .CLK(clk_bF$buf50),
    .D(_328_[21]),
    .Q(\datapath_1.regfile_1.regOut[6] [21]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _7602_ (
    .CLK(clk_bF$buf49),
    .D(_328_[22]),
    .Q(\datapath_1.regfile_1.regOut[6] [22]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _7603_ (
    .CLK(clk_bF$buf48),
    .D(_328_[23]),
    .Q(\datapath_1.regfile_1.regOut[6] [23]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _7604_ (
    .CLK(clk_bF$buf47),
    .D(_328_[24]),
    .Q(\datapath_1.regfile_1.regOut[6] [24]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _7605_ (
    .CLK(clk_bF$buf46),
    .D(_328_[25]),
    .Q(\datapath_1.regfile_1.regOut[6] [25]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _7606_ (
    .CLK(clk_bF$buf45),
    .D(_328_[26]),
    .Q(\datapath_1.regfile_1.regOut[6] [26]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _7607_ (
    .CLK(clk_bF$buf44),
    .D(_328_[27]),
    .Q(\datapath_1.regfile_1.regOut[6] [27]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _7608_ (
    .CLK(clk_bF$buf43),
    .D(_328_[28]),
    .Q(\datapath_1.regfile_1.regOut[6] [28]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _7609_ (
    .CLK(clk_bF$buf42),
    .D(_328_[29]),
    .Q(\datapath_1.regfile_1.regOut[6] [29]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _7610_ (
    .CLK(clk_bF$buf41),
    .D(_328_[30]),
    .Q(\datapath_1.regfile_1.regOut[6] [30]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _7611_ (
    .CLK(clk_bF$buf40),
    .D(_328_[31]),
    .Q(\datapath_1.regfile_1.regOut[6] [31]),
    .R(rst_bF$buf40),
    .S(vdd)
);

INVX1 _7612_ (
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .Y(_456_)
);

NAND2X1 _7613_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .Y(_457_)
);

OAI21X1 _7614_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_456_),
    .C(_457_),
    .Y(_393_[0])
);

INVX1 _7615_ (
    .A(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_394_)
);

NAND2X1 _7616_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_395_)
);

OAI21X1 _7617_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_394_),
    .C(_395_),
    .Y(_393_[1])
);

INVX1 _7618_ (
    .A(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_396_)
);

NAND2X1 _7619_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_397_)
);

OAI21X1 _7620_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_396_),
    .C(_397_),
    .Y(_393_[2])
);

INVX1 _7621_ (
    .A(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_398_)
);

NAND2X1 _7622_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_399_)
);

OAI21X1 _7623_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_398_),
    .C(_399_),
    .Y(_393_[3])
);

INVX1 _7624_ (
    .A(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_400_)
);

NAND2X1 _7625_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_401_)
);

OAI21X1 _7626_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_400_),
    .C(_401_),
    .Y(_393_[4])
);

INVX1 _7627_ (
    .A(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_402_)
);

NAND2X1 _7628_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_403_)
);

OAI21X1 _7629_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_402_),
    .C(_403_),
    .Y(_393_[5])
);

INVX1 _7630_ (
    .A(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_404_)
);

NAND2X1 _7631_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_405_)
);

OAI21X1 _7632_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_404_),
    .C(_405_),
    .Y(_393_[6])
);

INVX1 _7633_ (
    .A(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_406_)
);

NAND2X1 _7634_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_407_)
);

OAI21X1 _7635_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_406_),
    .C(_407_),
    .Y(_393_[7])
);

INVX1 _7636_ (
    .A(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_408_)
);

NAND2X1 _7637_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_409_)
);

OAI21X1 _7638_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_408_),
    .C(_409_),
    .Y(_393_[8])
);

INVX1 _7639_ (
    .A(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_410_)
);

NAND2X1 _7640_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_411_)
);

OAI21X1 _7641_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_410_),
    .C(_411_),
    .Y(_393_[9])
);

INVX1 _7642_ (
    .A(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_412_)
);

NAND2X1 _7643_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_413_)
);

OAI21X1 _7644_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_412_),
    .C(_413_),
    .Y(_393_[10])
);

INVX1 _7645_ (
    .A(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_414_)
);

NAND2X1 _7646_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_415_)
);

OAI21X1 _7647_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_414_),
    .C(_415_),
    .Y(_393_[11])
);

INVX1 _7648_ (
    .A(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_416_)
);

NAND2X1 _7649_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_417_)
);

OAI21X1 _7650_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_416_),
    .C(_417_),
    .Y(_393_[12])
);

INVX1 _7651_ (
    .A(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_418_)
);

NAND2X1 _7652_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_419_)
);

OAI21X1 _7653_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_418_),
    .C(_419_),
    .Y(_393_[13])
);

INVX1 _7654_ (
    .A(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_420_)
);

NAND2X1 _7655_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_421_)
);

OAI21X1 _7656_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_420_),
    .C(_421_),
    .Y(_393_[14])
);

INVX1 _7657_ (
    .A(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_422_)
);

NAND2X1 _7658_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_423_)
);

OAI21X1 _7659_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_422_),
    .C(_423_),
    .Y(_393_[15])
);

INVX1 _7660_ (
    .A(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_424_)
);

NAND2X1 _7661_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_425_)
);

OAI21X1 _7662_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_424_),
    .C(_425_),
    .Y(_393_[16])
);

INVX1 _7663_ (
    .A(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_426_)
);

NAND2X1 _7664_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_427_)
);

OAI21X1 _7665_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_426_),
    .C(_427_),
    .Y(_393_[17])
);

INVX1 _7666_ (
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_428_)
);

NAND2X1 _7667_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_429_)
);

OAI21X1 _7668_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_428_),
    .C(_429_),
    .Y(_393_[18])
);

INVX1 _7669_ (
    .A(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_430_)
);

NAND2X1 _7670_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_431_)
);

OAI21X1 _7671_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_430_),
    .C(_431_),
    .Y(_393_[19])
);

INVX1 _7672_ (
    .A(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_432_)
);

NAND2X1 _7673_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_433_)
);

OAI21X1 _7674_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_432_),
    .C(_433_),
    .Y(_393_[20])
);

INVX1 _7675_ (
    .A(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_434_)
);

NAND2X1 _7676_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_435_)
);

OAI21X1 _7677_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_434_),
    .C(_435_),
    .Y(_393_[21])
);

INVX1 _7678_ (
    .A(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_436_)
);

NAND2X1 _7679_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_437_)
);

OAI21X1 _7680_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_436_),
    .C(_437_),
    .Y(_393_[22])
);

INVX1 _7681_ (
    .A(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_438_)
);

NAND2X1 _7682_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_439_)
);

OAI21X1 _7683_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_438_),
    .C(_439_),
    .Y(_393_[23])
);

INVX1 _7684_ (
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_440_)
);

NAND2X1 _7685_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_441_)
);

OAI21X1 _7686_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_440_),
    .C(_441_),
    .Y(_393_[24])
);

INVX1 _7687_ (
    .A(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_442_)
);

NAND2X1 _7688_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_443_)
);

OAI21X1 _7689_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_442_),
    .C(_443_),
    .Y(_393_[25])
);

INVX1 _7690_ (
    .A(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_444_)
);

NAND2X1 _7691_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_445_)
);

OAI21X1 _7692_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_444_),
    .C(_445_),
    .Y(_393_[26])
);

INVX1 _7693_ (
    .A(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_446_)
);

NAND2X1 _7694_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_447_)
);

OAI21X1 _7695_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_446_),
    .C(_447_),
    .Y(_393_[27])
);

INVX1 _7696_ (
    .A(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_448_)
);

NAND2X1 _7697_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_449_)
);

OAI21X1 _7698_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(_448_),
    .C(_449_),
    .Y(_393_[28])
);

INVX1 _7699_ (
    .A(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_450_)
);

NAND2X1 _7700_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_451_)
);

OAI21X1 _7701_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(_450_),
    .C(_451_),
    .Y(_393_[29])
);

INVX1 _7702_ (
    .A(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_452_)
);

NAND2X1 _7703_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_453_)
);

OAI21X1 _7704_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(_452_),
    .C(_453_),
    .Y(_393_[30])
);

INVX1 _7705_ (
    .A(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_454_)
);

NAND2X1 _7706_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_455_)
);

OAI21X1 _7707_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(_454_),
    .C(_455_),
    .Y(_393_[31])
);

DFFSR _7708_ (
    .CLK(clk_bF$buf39),
    .D(_393_[0]),
    .Q(\datapath_1.regfile_1.regOut[7] [0]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _7709_ (
    .CLK(clk_bF$buf38),
    .D(_393_[1]),
    .Q(\datapath_1.regfile_1.regOut[7] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _7710_ (
    .CLK(clk_bF$buf37),
    .D(_393_[2]),
    .Q(\datapath_1.regfile_1.regOut[7] [2]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _7711_ (
    .CLK(clk_bF$buf36),
    .D(_393_[3]),
    .Q(\datapath_1.regfile_1.regOut[7] [3]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _7712_ (
    .CLK(clk_bF$buf35),
    .D(_393_[4]),
    .Q(\datapath_1.regfile_1.regOut[7] [4]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _7713_ (
    .CLK(clk_bF$buf34),
    .D(_393_[5]),
    .Q(\datapath_1.regfile_1.regOut[7] [5]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _7714_ (
    .CLK(clk_bF$buf33),
    .D(_393_[6]),
    .Q(\datapath_1.regfile_1.regOut[7] [6]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _7715_ (
    .CLK(clk_bF$buf32),
    .D(_393_[7]),
    .Q(\datapath_1.regfile_1.regOut[7] [7]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _7716_ (
    .CLK(clk_bF$buf31),
    .D(_393_[8]),
    .Q(\datapath_1.regfile_1.regOut[7] [8]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _7717_ (
    .CLK(clk_bF$buf30),
    .D(_393_[9]),
    .Q(\datapath_1.regfile_1.regOut[7] [9]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _7718_ (
    .CLK(clk_bF$buf29),
    .D(_393_[10]),
    .Q(\datapath_1.regfile_1.regOut[7] [10]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _7719_ (
    .CLK(clk_bF$buf28),
    .D(_393_[11]),
    .Q(\datapath_1.regfile_1.regOut[7] [11]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _7720_ (
    .CLK(clk_bF$buf27),
    .D(_393_[12]),
    .Q(\datapath_1.regfile_1.regOut[7] [12]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _7721_ (
    .CLK(clk_bF$buf26),
    .D(_393_[13]),
    .Q(\datapath_1.regfile_1.regOut[7] [13]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _7722_ (
    .CLK(clk_bF$buf25),
    .D(_393_[14]),
    .Q(\datapath_1.regfile_1.regOut[7] [14]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _7723_ (
    .CLK(clk_bF$buf24),
    .D(_393_[15]),
    .Q(\datapath_1.regfile_1.regOut[7] [15]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _7724_ (
    .CLK(clk_bF$buf23),
    .D(_393_[16]),
    .Q(\datapath_1.regfile_1.regOut[7] [16]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _7725_ (
    .CLK(clk_bF$buf22),
    .D(_393_[17]),
    .Q(\datapath_1.regfile_1.regOut[7] [17]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _7726_ (
    .CLK(clk_bF$buf21),
    .D(_393_[18]),
    .Q(\datapath_1.regfile_1.regOut[7] [18]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _7727_ (
    .CLK(clk_bF$buf20),
    .D(_393_[19]),
    .Q(\datapath_1.regfile_1.regOut[7] [19]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _7728_ (
    .CLK(clk_bF$buf19),
    .D(_393_[20]),
    .Q(\datapath_1.regfile_1.regOut[7] [20]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _7729_ (
    .CLK(clk_bF$buf18),
    .D(_393_[21]),
    .Q(\datapath_1.regfile_1.regOut[7] [21]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _7730_ (
    .CLK(clk_bF$buf17),
    .D(_393_[22]),
    .Q(\datapath_1.regfile_1.regOut[7] [22]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _7731_ (
    .CLK(clk_bF$buf16),
    .D(_393_[23]),
    .Q(\datapath_1.regfile_1.regOut[7] [23]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _7732_ (
    .CLK(clk_bF$buf15),
    .D(_393_[24]),
    .Q(\datapath_1.regfile_1.regOut[7] [24]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _7733_ (
    .CLK(clk_bF$buf14),
    .D(_393_[25]),
    .Q(\datapath_1.regfile_1.regOut[7] [25]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _7734_ (
    .CLK(clk_bF$buf13),
    .D(_393_[26]),
    .Q(\datapath_1.regfile_1.regOut[7] [26]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _7735_ (
    .CLK(clk_bF$buf12),
    .D(_393_[27]),
    .Q(\datapath_1.regfile_1.regOut[7] [27]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _7736_ (
    .CLK(clk_bF$buf11),
    .D(_393_[28]),
    .Q(\datapath_1.regfile_1.regOut[7] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _7737_ (
    .CLK(clk_bF$buf10),
    .D(_393_[29]),
    .Q(\datapath_1.regfile_1.regOut[7] [29]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _7738_ (
    .CLK(clk_bF$buf9),
    .D(_393_[30]),
    .Q(\datapath_1.regfile_1.regOut[7] [30]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _7739_ (
    .CLK(clk_bF$buf8),
    .D(_393_[31]),
    .Q(\datapath_1.regfile_1.regOut[7] [31]),
    .R(rst_bF$buf8),
    .S(vdd)
);

INVX1 _7740_ (
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_521_)
);

NAND2X1 _7741_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .Y(_522_)
);

OAI21X1 _7742_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_521_),
    .C(_522_),
    .Y(_458_[0])
);

INVX1 _7743_ (
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_459_)
);

NAND2X1 _7744_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_460_)
);

OAI21X1 _7745_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_459_),
    .C(_460_),
    .Y(_458_[1])
);

INVX1 _7746_ (
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_461_)
);

NAND2X1 _7747_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_462_)
);

OAI21X1 _7748_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_461_),
    .C(_462_),
    .Y(_458_[2])
);

INVX1 _7749_ (
    .A(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_463_)
);

NAND2X1 _7750_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_464_)
);

OAI21X1 _7751_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_463_),
    .C(_464_),
    .Y(_458_[3])
);

INVX1 _7752_ (
    .A(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_465_)
);

NAND2X1 _7753_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_466_)
);

OAI21X1 _7754_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_465_),
    .C(_466_),
    .Y(_458_[4])
);

INVX1 _7755_ (
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_467_)
);

NAND2X1 _7756_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_468_)
);

OAI21X1 _7757_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_467_),
    .C(_468_),
    .Y(_458_[5])
);

INVX1 _7758_ (
    .A(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_469_)
);

NAND2X1 _7759_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_470_)
);

OAI21X1 _7760_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_469_),
    .C(_470_),
    .Y(_458_[6])
);

INVX1 _7761_ (
    .A(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_471_)
);

NAND2X1 _7762_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_472_)
);

OAI21X1 _7763_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_471_),
    .C(_472_),
    .Y(_458_[7])
);

INVX1 _7764_ (
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_473_)
);

NAND2X1 _7765_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_474_)
);

OAI21X1 _7766_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_473_),
    .C(_474_),
    .Y(_458_[8])
);

INVX1 _7767_ (
    .A(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_475_)
);

NAND2X1 _7768_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_476_)
);

OAI21X1 _7769_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_475_),
    .C(_476_),
    .Y(_458_[9])
);

INVX1 _7770_ (
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_477_)
);

NAND2X1 _7771_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_478_)
);

OAI21X1 _7772_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_477_),
    .C(_478_),
    .Y(_458_[10])
);

INVX1 _7773_ (
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_479_)
);

NAND2X1 _7774_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_480_)
);

OAI21X1 _7775_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_479_),
    .C(_480_),
    .Y(_458_[11])
);

INVX1 _7776_ (
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_481_)
);

NAND2X1 _7777_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_482_)
);

OAI21X1 _7778_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_481_),
    .C(_482_),
    .Y(_458_[12])
);

INVX1 _7779_ (
    .A(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_483_)
);

NAND2X1 _7780_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_484_)
);

OAI21X1 _7781_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_483_),
    .C(_484_),
    .Y(_458_[13])
);

INVX1 _7782_ (
    .A(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_485_)
);

NAND2X1 _7783_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_486_)
);

OAI21X1 _7784_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_485_),
    .C(_486_),
    .Y(_458_[14])
);

INVX1 _7785_ (
    .A(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_487_)
);

NAND2X1 _7786_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_488_)
);

OAI21X1 _7787_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_487_),
    .C(_488_),
    .Y(_458_[15])
);

INVX1 _7788_ (
    .A(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_489_)
);

NAND2X1 _7789_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_490_)
);

OAI21X1 _7790_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_489_),
    .C(_490_),
    .Y(_458_[16])
);

INVX1 _7791_ (
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_491_)
);

NAND2X1 _7792_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_492_)
);

OAI21X1 _7793_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_491_),
    .C(_492_),
    .Y(_458_[17])
);

INVX1 _7794_ (
    .A(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_493_)
);

NAND2X1 _7795_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_494_)
);

OAI21X1 _7796_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_493_),
    .C(_494_),
    .Y(_458_[18])
);

INVX1 _7797_ (
    .A(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_495_)
);

NAND2X1 _7798_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_496_)
);

OAI21X1 _7799_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_495_),
    .C(_496_),
    .Y(_458_[19])
);

INVX1 _7800_ (
    .A(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_497_)
);

NAND2X1 _7801_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_498_)
);

OAI21X1 _7802_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_497_),
    .C(_498_),
    .Y(_458_[20])
);

INVX1 _7803_ (
    .A(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_499_)
);

NAND2X1 _7804_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_500_)
);

OAI21X1 _7805_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_499_),
    .C(_500_),
    .Y(_458_[21])
);

INVX1 _7806_ (
    .A(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_501_)
);

NAND2X1 _7807_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_502_)
);

OAI21X1 _7808_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_501_),
    .C(_502_),
    .Y(_458_[22])
);

INVX1 _7809_ (
    .A(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_503_)
);

NAND2X1 _7810_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_504_)
);

OAI21X1 _7811_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_503_),
    .C(_504_),
    .Y(_458_[23])
);

INVX1 _7812_ (
    .A(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_505_)
);

NAND2X1 _7813_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_506_)
);

OAI21X1 _7814_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_505_),
    .C(_506_),
    .Y(_458_[24])
);

INVX1 _7815_ (
    .A(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_507_)
);

NAND2X1 _7816_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_508_)
);

OAI21X1 _7817_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_507_),
    .C(_508_),
    .Y(_458_[25])
);

INVX1 _7818_ (
    .A(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_509_)
);

NAND2X1 _7819_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_510_)
);

OAI21X1 _7820_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_509_),
    .C(_510_),
    .Y(_458_[26])
);

INVX1 _7821_ (
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_511_)
);

NAND2X1 _7822_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_512_)
);

OAI21X1 _7823_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_511_),
    .C(_512_),
    .Y(_458_[27])
);

INVX1 _7824_ (
    .A(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_513_)
);

NAND2X1 _7825_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_514_)
);

OAI21X1 _7826_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(_513_),
    .C(_514_),
    .Y(_458_[28])
);

INVX1 _7827_ (
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_515_)
);

NAND2X1 _7828_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_516_)
);

OAI21X1 _7829_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(_515_),
    .C(_516_),
    .Y(_458_[29])
);

INVX1 _7830_ (
    .A(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_517_)
);

NAND2X1 _7831_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_518_)
);

OAI21X1 _7832_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(_517_),
    .C(_518_),
    .Y(_458_[30])
);

INVX1 _7833_ (
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_519_)
);

NAND2X1 _7834_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_520_)
);

OAI21X1 _7835_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(_519_),
    .C(_520_),
    .Y(_458_[31])
);

DFFSR _7836_ (
    .CLK(clk_bF$buf7),
    .D(_458_[0]),
    .Q(\datapath_1.regfile_1.regOut[8] [0]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _7837_ (
    .CLK(clk_bF$buf6),
    .D(_458_[1]),
    .Q(\datapath_1.regfile_1.regOut[8] [1]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _7838_ (
    .CLK(clk_bF$buf5),
    .D(_458_[2]),
    .Q(\datapath_1.regfile_1.regOut[8] [2]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _7839_ (
    .CLK(clk_bF$buf4),
    .D(_458_[3]),
    .Q(\datapath_1.regfile_1.regOut[8] [3]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _7840_ (
    .CLK(clk_bF$buf3),
    .D(_458_[4]),
    .Q(\datapath_1.regfile_1.regOut[8] [4]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _7841_ (
    .CLK(clk_bF$buf2),
    .D(_458_[5]),
    .Q(\datapath_1.regfile_1.regOut[8] [5]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _7842_ (
    .CLK(clk_bF$buf1),
    .D(_458_[6]),
    .Q(\datapath_1.regfile_1.regOut[8] [6]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _7843_ (
    .CLK(clk_bF$buf0),
    .D(_458_[7]),
    .Q(\datapath_1.regfile_1.regOut[8] [7]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _7844_ (
    .CLK(clk_bF$buf113),
    .D(_458_[8]),
    .Q(\datapath_1.regfile_1.regOut[8] [8]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _7845_ (
    .CLK(clk_bF$buf112),
    .D(_458_[9]),
    .Q(\datapath_1.regfile_1.regOut[8] [9]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _7846_ (
    .CLK(clk_bF$buf111),
    .D(_458_[10]),
    .Q(\datapath_1.regfile_1.regOut[8] [10]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _7847_ (
    .CLK(clk_bF$buf110),
    .D(_458_[11]),
    .Q(\datapath_1.regfile_1.regOut[8] [11]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _7848_ (
    .CLK(clk_bF$buf109),
    .D(_458_[12]),
    .Q(\datapath_1.regfile_1.regOut[8] [12]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _7849_ (
    .CLK(clk_bF$buf108),
    .D(_458_[13]),
    .Q(\datapath_1.regfile_1.regOut[8] [13]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _7850_ (
    .CLK(clk_bF$buf107),
    .D(_458_[14]),
    .Q(\datapath_1.regfile_1.regOut[8] [14]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _7851_ (
    .CLK(clk_bF$buf106),
    .D(_458_[15]),
    .Q(\datapath_1.regfile_1.regOut[8] [15]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _7852_ (
    .CLK(clk_bF$buf105),
    .D(_458_[16]),
    .Q(\datapath_1.regfile_1.regOut[8] [16]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _7853_ (
    .CLK(clk_bF$buf104),
    .D(_458_[17]),
    .Q(\datapath_1.regfile_1.regOut[8] [17]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _7854_ (
    .CLK(clk_bF$buf103),
    .D(_458_[18]),
    .Q(\datapath_1.regfile_1.regOut[8] [18]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _7855_ (
    .CLK(clk_bF$buf102),
    .D(_458_[19]),
    .Q(\datapath_1.regfile_1.regOut[8] [19]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _7856_ (
    .CLK(clk_bF$buf101),
    .D(_458_[20]),
    .Q(\datapath_1.regfile_1.regOut[8] [20]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _7857_ (
    .CLK(clk_bF$buf100),
    .D(_458_[21]),
    .Q(\datapath_1.regfile_1.regOut[8] [21]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _7858_ (
    .CLK(clk_bF$buf99),
    .D(_458_[22]),
    .Q(\datapath_1.regfile_1.regOut[8] [22]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _7859_ (
    .CLK(clk_bF$buf98),
    .D(_458_[23]),
    .Q(\datapath_1.regfile_1.regOut[8] [23]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _7860_ (
    .CLK(clk_bF$buf97),
    .D(_458_[24]),
    .Q(\datapath_1.regfile_1.regOut[8] [24]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _7861_ (
    .CLK(clk_bF$buf96),
    .D(_458_[25]),
    .Q(\datapath_1.regfile_1.regOut[8] [25]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _7862_ (
    .CLK(clk_bF$buf95),
    .D(_458_[26]),
    .Q(\datapath_1.regfile_1.regOut[8] [26]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _7863_ (
    .CLK(clk_bF$buf94),
    .D(_458_[27]),
    .Q(\datapath_1.regfile_1.regOut[8] [27]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _7864_ (
    .CLK(clk_bF$buf93),
    .D(_458_[28]),
    .Q(\datapath_1.regfile_1.regOut[8] [28]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _7865_ (
    .CLK(clk_bF$buf92),
    .D(_458_[29]),
    .Q(\datapath_1.regfile_1.regOut[8] [29]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _7866_ (
    .CLK(clk_bF$buf91),
    .D(_458_[30]),
    .Q(\datapath_1.regfile_1.regOut[8] [30]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _7867_ (
    .CLK(clk_bF$buf90),
    .D(_458_[31]),
    .Q(\datapath_1.regfile_1.regOut[8] [31]),
    .R(rst_bF$buf90),
    .S(vdd)
);

INVX1 _7868_ (
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_586_)
);

NAND2X1 _7869_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .Y(_587_)
);

OAI21X1 _7870_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_586_),
    .C(_587_),
    .Y(_523_[0])
);

INVX1 _7871_ (
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_524_)
);

NAND2X1 _7872_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_525_)
);

OAI21X1 _7873_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_524_),
    .C(_525_),
    .Y(_523_[1])
);

INVX1 _7874_ (
    .A(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_526_)
);

NAND2X1 _7875_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_527_)
);

OAI21X1 _7876_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_526_),
    .C(_527_),
    .Y(_523_[2])
);

INVX1 _7877_ (
    .A(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_528_)
);

NAND2X1 _7878_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_529_)
);

OAI21X1 _7879_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_528_),
    .C(_529_),
    .Y(_523_[3])
);

INVX1 _7880_ (
    .A(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_530_)
);

NAND2X1 _7881_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_531_)
);

OAI21X1 _7882_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_530_),
    .C(_531_),
    .Y(_523_[4])
);

INVX1 _7883_ (
    .A(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_532_)
);

NAND2X1 _7884_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_533_)
);

OAI21X1 _7885_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_532_),
    .C(_533_),
    .Y(_523_[5])
);

INVX1 _7886_ (
    .A(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_534_)
);

NAND2X1 _7887_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_535_)
);

OAI21X1 _7888_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_534_),
    .C(_535_),
    .Y(_523_[6])
);

INVX1 _7889_ (
    .A(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_536_)
);

NAND2X1 _7890_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_537_)
);

OAI21X1 _7891_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_536_),
    .C(_537_),
    .Y(_523_[7])
);

INVX1 _7892_ (
    .A(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_538_)
);

NAND2X1 _7893_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_539_)
);

OAI21X1 _7894_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_538_),
    .C(_539_),
    .Y(_523_[8])
);

INVX1 _7895_ (
    .A(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_540_)
);

NAND2X1 _7896_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_541_)
);

OAI21X1 _7897_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_540_),
    .C(_541_),
    .Y(_523_[9])
);

INVX1 _7898_ (
    .A(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_542_)
);

NAND2X1 _7899_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_543_)
);

OAI21X1 _7900_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_542_),
    .C(_543_),
    .Y(_523_[10])
);

INVX1 _7901_ (
    .A(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_544_)
);

NAND2X1 _7902_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_545_)
);

OAI21X1 _7903_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_544_),
    .C(_545_),
    .Y(_523_[11])
);

INVX1 _7904_ (
    .A(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_546_)
);

NAND2X1 _7905_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_547_)
);

OAI21X1 _7906_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_546_),
    .C(_547_),
    .Y(_523_[12])
);

INVX1 _7907_ (
    .A(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_548_)
);

NAND2X1 _7908_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_549_)
);

OAI21X1 _7909_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_548_),
    .C(_549_),
    .Y(_523_[13])
);

INVX1 _7910_ (
    .A(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_550_)
);

NAND2X1 _7911_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_551_)
);

OAI21X1 _7912_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_550_),
    .C(_551_),
    .Y(_523_[14])
);

INVX1 _7913_ (
    .A(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_552_)
);

NAND2X1 _7914_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_553_)
);

OAI21X1 _7915_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_552_),
    .C(_553_),
    .Y(_523_[15])
);

INVX1 _7916_ (
    .A(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_554_)
);

NAND2X1 _7917_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_555_)
);

OAI21X1 _7918_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_554_),
    .C(_555_),
    .Y(_523_[16])
);

INVX1 _7919_ (
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_556_)
);

NAND2X1 _7920_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_557_)
);

OAI21X1 _7921_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_556_),
    .C(_557_),
    .Y(_523_[17])
);

INVX1 _7922_ (
    .A(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_558_)
);

NAND2X1 _7923_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_559_)
);

OAI21X1 _7924_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_558_),
    .C(_559_),
    .Y(_523_[18])
);

INVX1 _7925_ (
    .A(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_560_)
);

NAND2X1 _7926_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_561_)
);

OAI21X1 _7927_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_560_),
    .C(_561_),
    .Y(_523_[19])
);

INVX1 _7928_ (
    .A(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_562_)
);

NAND2X1 _7929_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_563_)
);

OAI21X1 _7930_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_562_),
    .C(_563_),
    .Y(_523_[20])
);

INVX1 _7931_ (
    .A(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_564_)
);

NAND2X1 _7932_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_565_)
);

OAI21X1 _7933_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_564_),
    .C(_565_),
    .Y(_523_[21])
);

INVX1 _7934_ (
    .A(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_566_)
);

NAND2X1 _7935_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_567_)
);

OAI21X1 _7936_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_566_),
    .C(_567_),
    .Y(_523_[22])
);

INVX1 _7937_ (
    .A(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_568_)
);

NAND2X1 _7938_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_569_)
);

OAI21X1 _7939_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_568_),
    .C(_569_),
    .Y(_523_[23])
);

INVX1 _7940_ (
    .A(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_570_)
);

NAND2X1 _7941_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_571_)
);

OAI21X1 _7942_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_570_),
    .C(_571_),
    .Y(_523_[24])
);

INVX1 _7943_ (
    .A(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_572_)
);

NAND2X1 _7944_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_573_)
);

OAI21X1 _7945_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_572_),
    .C(_573_),
    .Y(_523_[25])
);

INVX1 _7946_ (
    .A(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_574_)
);

NAND2X1 _7947_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_575_)
);

OAI21X1 _7948_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_574_),
    .C(_575_),
    .Y(_523_[26])
);

INVX1 _7949_ (
    .A(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_576_)
);

NAND2X1 _7950_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_577_)
);

OAI21X1 _7951_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_576_),
    .C(_577_),
    .Y(_523_[27])
);

INVX1 _7952_ (
    .A(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_578_)
);

NAND2X1 _7953_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_579_)
);

OAI21X1 _7954_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(_578_),
    .C(_579_),
    .Y(_523_[28])
);

INVX1 _7955_ (
    .A(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_580_)
);

NAND2X1 _7956_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_581_)
);

OAI21X1 _7957_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(_580_),
    .C(_581_),
    .Y(_523_[29])
);

INVX1 _7958_ (
    .A(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_582_)
);

NAND2X1 _7959_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_583_)
);

OAI21X1 _7960_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(_582_),
    .C(_583_),
    .Y(_523_[30])
);

INVX1 _7961_ (
    .A(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_584_)
);

NAND2X1 _7962_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_585_)
);

OAI21X1 _7963_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(_584_),
    .C(_585_),
    .Y(_523_[31])
);

DFFSR _7964_ (
    .CLK(clk_bF$buf89),
    .D(_523_[0]),
    .Q(\datapath_1.regfile_1.regOut[9] [0]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _7965_ (
    .CLK(clk_bF$buf88),
    .D(_523_[1]),
    .Q(\datapath_1.regfile_1.regOut[9] [1]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _7966_ (
    .CLK(clk_bF$buf87),
    .D(_523_[2]),
    .Q(\datapath_1.regfile_1.regOut[9] [2]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _7967_ (
    .CLK(clk_bF$buf86),
    .D(_523_[3]),
    .Q(\datapath_1.regfile_1.regOut[9] [3]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _7968_ (
    .CLK(clk_bF$buf85),
    .D(_523_[4]),
    .Q(\datapath_1.regfile_1.regOut[9] [4]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _7969_ (
    .CLK(clk_bF$buf84),
    .D(_523_[5]),
    .Q(\datapath_1.regfile_1.regOut[9] [5]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _7970_ (
    .CLK(clk_bF$buf83),
    .D(_523_[6]),
    .Q(\datapath_1.regfile_1.regOut[9] [6]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _7971_ (
    .CLK(clk_bF$buf82),
    .D(_523_[7]),
    .Q(\datapath_1.regfile_1.regOut[9] [7]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _7972_ (
    .CLK(clk_bF$buf81),
    .D(_523_[8]),
    .Q(\datapath_1.regfile_1.regOut[9] [8]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _7973_ (
    .CLK(clk_bF$buf80),
    .D(_523_[9]),
    .Q(\datapath_1.regfile_1.regOut[9] [9]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _7974_ (
    .CLK(clk_bF$buf79),
    .D(_523_[10]),
    .Q(\datapath_1.regfile_1.regOut[9] [10]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _7975_ (
    .CLK(clk_bF$buf78),
    .D(_523_[11]),
    .Q(\datapath_1.regfile_1.regOut[9] [11]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _7976_ (
    .CLK(clk_bF$buf77),
    .D(_523_[12]),
    .Q(\datapath_1.regfile_1.regOut[9] [12]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _7977_ (
    .CLK(clk_bF$buf76),
    .D(_523_[13]),
    .Q(\datapath_1.regfile_1.regOut[9] [13]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _7978_ (
    .CLK(clk_bF$buf75),
    .D(_523_[14]),
    .Q(\datapath_1.regfile_1.regOut[9] [14]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _7979_ (
    .CLK(clk_bF$buf74),
    .D(_523_[15]),
    .Q(\datapath_1.regfile_1.regOut[9] [15]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _7980_ (
    .CLK(clk_bF$buf73),
    .D(_523_[16]),
    .Q(\datapath_1.regfile_1.regOut[9] [16]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _7981_ (
    .CLK(clk_bF$buf72),
    .D(_523_[17]),
    .Q(\datapath_1.regfile_1.regOut[9] [17]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _7982_ (
    .CLK(clk_bF$buf71),
    .D(_523_[18]),
    .Q(\datapath_1.regfile_1.regOut[9] [18]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _7983_ (
    .CLK(clk_bF$buf70),
    .D(_523_[19]),
    .Q(\datapath_1.regfile_1.regOut[9] [19]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _7984_ (
    .CLK(clk_bF$buf69),
    .D(_523_[20]),
    .Q(\datapath_1.regfile_1.regOut[9] [20]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _7985_ (
    .CLK(clk_bF$buf68),
    .D(_523_[21]),
    .Q(\datapath_1.regfile_1.regOut[9] [21]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _7986_ (
    .CLK(clk_bF$buf67),
    .D(_523_[22]),
    .Q(\datapath_1.regfile_1.regOut[9] [22]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _7987_ (
    .CLK(clk_bF$buf66),
    .D(_523_[23]),
    .Q(\datapath_1.regfile_1.regOut[9] [23]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _7988_ (
    .CLK(clk_bF$buf65),
    .D(_523_[24]),
    .Q(\datapath_1.regfile_1.regOut[9] [24]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _7989_ (
    .CLK(clk_bF$buf64),
    .D(_523_[25]),
    .Q(\datapath_1.regfile_1.regOut[9] [25]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _7990_ (
    .CLK(clk_bF$buf63),
    .D(_523_[26]),
    .Q(\datapath_1.regfile_1.regOut[9] [26]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _7991_ (
    .CLK(clk_bF$buf62),
    .D(_523_[27]),
    .Q(\datapath_1.regfile_1.regOut[9] [27]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _7992_ (
    .CLK(clk_bF$buf61),
    .D(_523_[28]),
    .Q(\datapath_1.regfile_1.regOut[9] [28]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _7993_ (
    .CLK(clk_bF$buf60),
    .D(_523_[29]),
    .Q(\datapath_1.regfile_1.regOut[9] [29]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _7994_ (
    .CLK(clk_bF$buf59),
    .D(_523_[30]),
    .Q(\datapath_1.regfile_1.regOut[9] [30]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _7995_ (
    .CLK(clk_bF$buf58),
    .D(_523_[31]),
    .Q(\datapath_1.regfile_1.regOut[9] [31]),
    .R(rst_bF$buf58),
    .S(vdd)
);

INVX1 _7996_ (
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_651_)
);

NAND2X1 _7997_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .Y(_652_)
);

OAI21X1 _7998_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_651_),
    .C(_652_),
    .Y(_588_[0])
);

INVX1 _7999_ (
    .A(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_589_)
);

NAND2X1 _8000_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_590_)
);

OAI21X1 _8001_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_589_),
    .C(_590_),
    .Y(_588_[1])
);

INVX1 _8002_ (
    .A(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_591_)
);

NAND2X1 _8003_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_592_)
);

OAI21X1 _8004_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_591_),
    .C(_592_),
    .Y(_588_[2])
);

INVX1 _8005_ (
    .A(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_593_)
);

NAND2X1 _8006_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_594_)
);

OAI21X1 _8007_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_593_),
    .C(_594_),
    .Y(_588_[3])
);

INVX1 _8008_ (
    .A(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_595_)
);

NAND2X1 _8009_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_596_)
);

OAI21X1 _8010_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_595_),
    .C(_596_),
    .Y(_588_[4])
);

INVX1 _8011_ (
    .A(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_597_)
);

NAND2X1 _8012_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_598_)
);

OAI21X1 _8013_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_597_),
    .C(_598_),
    .Y(_588_[5])
);

INVX1 _8014_ (
    .A(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_599_)
);

NAND2X1 _8015_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_600_)
);

OAI21X1 _8016_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_599_),
    .C(_600_),
    .Y(_588_[6])
);

INVX1 _8017_ (
    .A(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_601_)
);

NAND2X1 _8018_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_602_)
);

OAI21X1 _8019_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_601_),
    .C(_602_),
    .Y(_588_[7])
);

INVX1 _8020_ (
    .A(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_603_)
);

NAND2X1 _8021_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_604_)
);

OAI21X1 _8022_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_603_),
    .C(_604_),
    .Y(_588_[8])
);

INVX1 _8023_ (
    .A(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_605_)
);

NAND2X1 _8024_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_606_)
);

OAI21X1 _8025_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_605_),
    .C(_606_),
    .Y(_588_[9])
);

INVX1 _8026_ (
    .A(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_607_)
);

NAND2X1 _8027_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_608_)
);

OAI21X1 _8028_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_607_),
    .C(_608_),
    .Y(_588_[10])
);

INVX1 _8029_ (
    .A(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_609_)
);

NAND2X1 _8030_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_610_)
);

OAI21X1 _8031_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_609_),
    .C(_610_),
    .Y(_588_[11])
);

INVX1 _8032_ (
    .A(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_611_)
);

NAND2X1 _8033_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_612_)
);

OAI21X1 _8034_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_611_),
    .C(_612_),
    .Y(_588_[12])
);

INVX1 _8035_ (
    .A(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_613_)
);

NAND2X1 _8036_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_614_)
);

OAI21X1 _8037_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_613_),
    .C(_614_),
    .Y(_588_[13])
);

INVX1 _8038_ (
    .A(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_615_)
);

NAND2X1 _8039_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_616_)
);

OAI21X1 _8040_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_615_),
    .C(_616_),
    .Y(_588_[14])
);

INVX1 _8041_ (
    .A(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_617_)
);

NAND2X1 _8042_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_618_)
);

OAI21X1 _8043_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_617_),
    .C(_618_),
    .Y(_588_[15])
);

INVX1 _8044_ (
    .A(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_619_)
);

NAND2X1 _8045_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_620_)
);

OAI21X1 _8046_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_619_),
    .C(_620_),
    .Y(_588_[16])
);

INVX1 _8047_ (
    .A(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_621_)
);

NAND2X1 _8048_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_622_)
);

OAI21X1 _8049_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_621_),
    .C(_622_),
    .Y(_588_[17])
);

INVX1 _8050_ (
    .A(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_623_)
);

NAND2X1 _8051_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_624_)
);

OAI21X1 _8052_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_623_),
    .C(_624_),
    .Y(_588_[18])
);

INVX1 _8053_ (
    .A(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_625_)
);

NAND2X1 _8054_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_626_)
);

OAI21X1 _8055_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_625_),
    .C(_626_),
    .Y(_588_[19])
);

INVX1 _8056_ (
    .A(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_627_)
);

NAND2X1 _8057_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_628_)
);

OAI21X1 _8058_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_627_),
    .C(_628_),
    .Y(_588_[20])
);

INVX1 _8059_ (
    .A(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_629_)
);

NAND2X1 _8060_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_630_)
);

OAI21X1 _8061_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_629_),
    .C(_630_),
    .Y(_588_[21])
);

INVX1 _8062_ (
    .A(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_631_)
);

NAND2X1 _8063_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_632_)
);

OAI21X1 _8064_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_631_),
    .C(_632_),
    .Y(_588_[22])
);

INVX1 _8065_ (
    .A(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_633_)
);

NAND2X1 _8066_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_634_)
);

OAI21X1 _8067_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_633_),
    .C(_634_),
    .Y(_588_[23])
);

INVX1 _8068_ (
    .A(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_635_)
);

NAND2X1 _8069_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_636_)
);

OAI21X1 _8070_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_635_),
    .C(_636_),
    .Y(_588_[24])
);

INVX1 _8071_ (
    .A(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_637_)
);

NAND2X1 _8072_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_638_)
);

OAI21X1 _8073_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_637_),
    .C(_638_),
    .Y(_588_[25])
);

INVX1 _8074_ (
    .A(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_639_)
);

NAND2X1 _8075_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_640_)
);

OAI21X1 _8076_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_639_),
    .C(_640_),
    .Y(_588_[26])
);

INVX1 _8077_ (
    .A(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_641_)
);

NAND2X1 _8078_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_642_)
);

OAI21X1 _8079_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_641_),
    .C(_642_),
    .Y(_588_[27])
);

INVX1 _8080_ (
    .A(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_643_)
);

NAND2X1 _8081_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_644_)
);

OAI21X1 _8082_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(_643_),
    .C(_644_),
    .Y(_588_[28])
);

INVX1 _8083_ (
    .A(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_645_)
);

NAND2X1 _8084_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_646_)
);

OAI21X1 _8085_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(_645_),
    .C(_646_),
    .Y(_588_[29])
);

INVX1 _8086_ (
    .A(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_647_)
);

NAND2X1 _8087_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_648_)
);

OAI21X1 _8088_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(_647_),
    .C(_648_),
    .Y(_588_[30])
);

INVX1 _8089_ (
    .A(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_649_)
);

NAND2X1 _8090_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_650_)
);

OAI21X1 _8091_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(_649_),
    .C(_650_),
    .Y(_588_[31])
);

DFFSR _8092_ (
    .CLK(clk_bF$buf57),
    .D(_588_[0]),
    .Q(\datapath_1.regfile_1.regOut[10] [0]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _8093_ (
    .CLK(clk_bF$buf56),
    .D(_588_[1]),
    .Q(\datapath_1.regfile_1.regOut[10] [1]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _8094_ (
    .CLK(clk_bF$buf55),
    .D(_588_[2]),
    .Q(\datapath_1.regfile_1.regOut[10] [2]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _8095_ (
    .CLK(clk_bF$buf54),
    .D(_588_[3]),
    .Q(\datapath_1.regfile_1.regOut[10] [3]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _8096_ (
    .CLK(clk_bF$buf53),
    .D(_588_[4]),
    .Q(\datapath_1.regfile_1.regOut[10] [4]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _8097_ (
    .CLK(clk_bF$buf52),
    .D(_588_[5]),
    .Q(\datapath_1.regfile_1.regOut[10] [5]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _8098_ (
    .CLK(clk_bF$buf51),
    .D(_588_[6]),
    .Q(\datapath_1.regfile_1.regOut[10] [6]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _8099_ (
    .CLK(clk_bF$buf50),
    .D(_588_[7]),
    .Q(\datapath_1.regfile_1.regOut[10] [7]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _8100_ (
    .CLK(clk_bF$buf49),
    .D(_588_[8]),
    .Q(\datapath_1.regfile_1.regOut[10] [8]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _8101_ (
    .CLK(clk_bF$buf48),
    .D(_588_[9]),
    .Q(\datapath_1.regfile_1.regOut[10] [9]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _8102_ (
    .CLK(clk_bF$buf47),
    .D(_588_[10]),
    .Q(\datapath_1.regfile_1.regOut[10] [10]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _8103_ (
    .CLK(clk_bF$buf46),
    .D(_588_[11]),
    .Q(\datapath_1.regfile_1.regOut[10] [11]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _8104_ (
    .CLK(clk_bF$buf45),
    .D(_588_[12]),
    .Q(\datapath_1.regfile_1.regOut[10] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _8105_ (
    .CLK(clk_bF$buf44),
    .D(_588_[13]),
    .Q(\datapath_1.regfile_1.regOut[10] [13]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _8106_ (
    .CLK(clk_bF$buf43),
    .D(_588_[14]),
    .Q(\datapath_1.regfile_1.regOut[10] [14]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _8107_ (
    .CLK(clk_bF$buf42),
    .D(_588_[15]),
    .Q(\datapath_1.regfile_1.regOut[10] [15]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _8108_ (
    .CLK(clk_bF$buf41),
    .D(_588_[16]),
    .Q(\datapath_1.regfile_1.regOut[10] [16]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _8109_ (
    .CLK(clk_bF$buf40),
    .D(_588_[17]),
    .Q(\datapath_1.regfile_1.regOut[10] [17]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _8110_ (
    .CLK(clk_bF$buf39),
    .D(_588_[18]),
    .Q(\datapath_1.regfile_1.regOut[10] [18]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _8111_ (
    .CLK(clk_bF$buf38),
    .D(_588_[19]),
    .Q(\datapath_1.regfile_1.regOut[10] [19]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _8112_ (
    .CLK(clk_bF$buf37),
    .D(_588_[20]),
    .Q(\datapath_1.regfile_1.regOut[10] [20]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _8113_ (
    .CLK(clk_bF$buf36),
    .D(_588_[21]),
    .Q(\datapath_1.regfile_1.regOut[10] [21]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _8114_ (
    .CLK(clk_bF$buf35),
    .D(_588_[22]),
    .Q(\datapath_1.regfile_1.regOut[10] [22]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _8115_ (
    .CLK(clk_bF$buf34),
    .D(_588_[23]),
    .Q(\datapath_1.regfile_1.regOut[10] [23]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _8116_ (
    .CLK(clk_bF$buf33),
    .D(_588_[24]),
    .Q(\datapath_1.regfile_1.regOut[10] [24]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _8117_ (
    .CLK(clk_bF$buf32),
    .D(_588_[25]),
    .Q(\datapath_1.regfile_1.regOut[10] [25]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _8118_ (
    .CLK(clk_bF$buf31),
    .D(_588_[26]),
    .Q(\datapath_1.regfile_1.regOut[10] [26]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _8119_ (
    .CLK(clk_bF$buf30),
    .D(_588_[27]),
    .Q(\datapath_1.regfile_1.regOut[10] [27]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _8120_ (
    .CLK(clk_bF$buf29),
    .D(_588_[28]),
    .Q(\datapath_1.regfile_1.regOut[10] [28]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _8121_ (
    .CLK(clk_bF$buf28),
    .D(_588_[29]),
    .Q(\datapath_1.regfile_1.regOut[10] [29]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _8122_ (
    .CLK(clk_bF$buf27),
    .D(_588_[30]),
    .Q(\datapath_1.regfile_1.regOut[10] [30]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _8123_ (
    .CLK(clk_bF$buf26),
    .D(_588_[31]),
    .Q(\datapath_1.regfile_1.regOut[10] [31]),
    .R(rst_bF$buf26),
    .S(vdd)
);

INVX1 _8124_ (
    .A(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_716_)
);

NAND2X1 _8125_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .Y(_717_)
);

OAI21X1 _8126_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_716_),
    .C(_717_),
    .Y(_653_[0])
);

INVX1 _8127_ (
    .A(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_654_)
);

NAND2X1 _8128_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_655_)
);

OAI21X1 _8129_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_654_),
    .C(_655_),
    .Y(_653_[1])
);

INVX1 _8130_ (
    .A(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_656_)
);

NAND2X1 _8131_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_657_)
);

OAI21X1 _8132_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_656_),
    .C(_657_),
    .Y(_653_[2])
);

INVX1 _8133_ (
    .A(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_658_)
);

NAND2X1 _8134_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_659_)
);

OAI21X1 _8135_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_658_),
    .C(_659_),
    .Y(_653_[3])
);

INVX1 _8136_ (
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_660_)
);

NAND2X1 _8137_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_661_)
);

OAI21X1 _8138_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_660_),
    .C(_661_),
    .Y(_653_[4])
);

INVX1 _8139_ (
    .A(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_662_)
);

NAND2X1 _8140_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_663_)
);

OAI21X1 _8141_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_662_),
    .C(_663_),
    .Y(_653_[5])
);

INVX1 _8142_ (
    .A(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_664_)
);

NAND2X1 _8143_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_665_)
);

OAI21X1 _8144_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_664_),
    .C(_665_),
    .Y(_653_[6])
);

INVX1 _8145_ (
    .A(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_666_)
);

NAND2X1 _8146_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_667_)
);

OAI21X1 _8147_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_666_),
    .C(_667_),
    .Y(_653_[7])
);

INVX1 _8148_ (
    .A(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_668_)
);

NAND2X1 _8149_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_669_)
);

OAI21X1 _8150_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_668_),
    .C(_669_),
    .Y(_653_[8])
);

INVX1 _8151_ (
    .A(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_670_)
);

NAND2X1 _8152_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_671_)
);

OAI21X1 _8153_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_670_),
    .C(_671_),
    .Y(_653_[9])
);

INVX1 _8154_ (
    .A(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_672_)
);

NAND2X1 _8155_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_673_)
);

OAI21X1 _8156_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_672_),
    .C(_673_),
    .Y(_653_[10])
);

INVX1 _8157_ (
    .A(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_674_)
);

NAND2X1 _8158_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_675_)
);

OAI21X1 _8159_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_674_),
    .C(_675_),
    .Y(_653_[11])
);

INVX1 _8160_ (
    .A(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_676_)
);

NAND2X1 _8161_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_677_)
);

OAI21X1 _8162_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_676_),
    .C(_677_),
    .Y(_653_[12])
);

INVX1 _8163_ (
    .A(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_678_)
);

NAND2X1 _8164_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_679_)
);

OAI21X1 _8165_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_678_),
    .C(_679_),
    .Y(_653_[13])
);

INVX1 _8166_ (
    .A(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_680_)
);

NAND2X1 _8167_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_681_)
);

OAI21X1 _8168_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_680_),
    .C(_681_),
    .Y(_653_[14])
);

INVX1 _8169_ (
    .A(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_682_)
);

NAND2X1 _8170_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_683_)
);

OAI21X1 _8171_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_682_),
    .C(_683_),
    .Y(_653_[15])
);

INVX1 _8172_ (
    .A(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_684_)
);

NAND2X1 _8173_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_685_)
);

OAI21X1 _8174_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_684_),
    .C(_685_),
    .Y(_653_[16])
);

INVX1 _8175_ (
    .A(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_686_)
);

NAND2X1 _8176_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_687_)
);

OAI21X1 _8177_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_686_),
    .C(_687_),
    .Y(_653_[17])
);

INVX1 _8178_ (
    .A(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_688_)
);

NAND2X1 _8179_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_689_)
);

OAI21X1 _8180_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_688_),
    .C(_689_),
    .Y(_653_[18])
);

INVX1 _8181_ (
    .A(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_690_)
);

NAND2X1 _8182_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_691_)
);

OAI21X1 _8183_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_690_),
    .C(_691_),
    .Y(_653_[19])
);

INVX1 _8184_ (
    .A(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_692_)
);

NAND2X1 _8185_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_693_)
);

OAI21X1 _8186_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_692_),
    .C(_693_),
    .Y(_653_[20])
);

INVX1 _8187_ (
    .A(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_694_)
);

NAND2X1 _8188_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_695_)
);

OAI21X1 _8189_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_694_),
    .C(_695_),
    .Y(_653_[21])
);

INVX1 _8190_ (
    .A(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_696_)
);

NAND2X1 _8191_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_697_)
);

OAI21X1 _8192_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_696_),
    .C(_697_),
    .Y(_653_[22])
);

INVX1 _8193_ (
    .A(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_698_)
);

NAND2X1 _8194_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_699_)
);

OAI21X1 _8195_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_698_),
    .C(_699_),
    .Y(_653_[23])
);

INVX1 _8196_ (
    .A(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_700_)
);

NAND2X1 _8197_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_701_)
);

OAI21X1 _8198_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_700_),
    .C(_701_),
    .Y(_653_[24])
);

INVX1 _8199_ (
    .A(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_702_)
);

NAND2X1 _8200_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_703_)
);

OAI21X1 _8201_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_702_),
    .C(_703_),
    .Y(_653_[25])
);

INVX1 _8202_ (
    .A(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_704_)
);

NAND2X1 _8203_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_705_)
);

OAI21X1 _8204_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_704_),
    .C(_705_),
    .Y(_653_[26])
);

INVX1 _8205_ (
    .A(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_706_)
);

NAND2X1 _8206_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_707_)
);

OAI21X1 _8207_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_706_),
    .C(_707_),
    .Y(_653_[27])
);

INVX1 _8208_ (
    .A(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_708_)
);

NAND2X1 _8209_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_709_)
);

OAI21X1 _8210_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(_708_),
    .C(_709_),
    .Y(_653_[28])
);

INVX1 _8211_ (
    .A(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_710_)
);

NAND2X1 _8212_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_711_)
);

OAI21X1 _8213_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(_710_),
    .C(_711_),
    .Y(_653_[29])
);

INVX1 _8214_ (
    .A(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_712_)
);

NAND2X1 _8215_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_713_)
);

OAI21X1 _8216_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(_712_),
    .C(_713_),
    .Y(_653_[30])
);

INVX1 _8217_ (
    .A(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_714_)
);

NAND2X1 _8218_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_715_)
);

OAI21X1 _8219_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(_714_),
    .C(_715_),
    .Y(_653_[31])
);

DFFSR _8220_ (
    .CLK(clk_bF$buf25),
    .D(_653_[0]),
    .Q(\datapath_1.regfile_1.regOut[11] [0]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _8221_ (
    .CLK(clk_bF$buf24),
    .D(_653_[1]),
    .Q(\datapath_1.regfile_1.regOut[11] [1]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _8222_ (
    .CLK(clk_bF$buf23),
    .D(_653_[2]),
    .Q(\datapath_1.regfile_1.regOut[11] [2]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _8223_ (
    .CLK(clk_bF$buf22),
    .D(_653_[3]),
    .Q(\datapath_1.regfile_1.regOut[11] [3]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _8224_ (
    .CLK(clk_bF$buf21),
    .D(_653_[4]),
    .Q(\datapath_1.regfile_1.regOut[11] [4]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _8225_ (
    .CLK(clk_bF$buf20),
    .D(_653_[5]),
    .Q(\datapath_1.regfile_1.regOut[11] [5]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _8226_ (
    .CLK(clk_bF$buf19),
    .D(_653_[6]),
    .Q(\datapath_1.regfile_1.regOut[11] [6]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _8227_ (
    .CLK(clk_bF$buf18),
    .D(_653_[7]),
    .Q(\datapath_1.regfile_1.regOut[11] [7]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _8228_ (
    .CLK(clk_bF$buf17),
    .D(_653_[8]),
    .Q(\datapath_1.regfile_1.regOut[11] [8]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _8229_ (
    .CLK(clk_bF$buf16),
    .D(_653_[9]),
    .Q(\datapath_1.regfile_1.regOut[11] [9]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _8230_ (
    .CLK(clk_bF$buf15),
    .D(_653_[10]),
    .Q(\datapath_1.regfile_1.regOut[11] [10]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _8231_ (
    .CLK(clk_bF$buf14),
    .D(_653_[11]),
    .Q(\datapath_1.regfile_1.regOut[11] [11]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _8232_ (
    .CLK(clk_bF$buf13),
    .D(_653_[12]),
    .Q(\datapath_1.regfile_1.regOut[11] [12]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _8233_ (
    .CLK(clk_bF$buf12),
    .D(_653_[13]),
    .Q(\datapath_1.regfile_1.regOut[11] [13]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _8234_ (
    .CLK(clk_bF$buf11),
    .D(_653_[14]),
    .Q(\datapath_1.regfile_1.regOut[11] [14]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _8235_ (
    .CLK(clk_bF$buf10),
    .D(_653_[15]),
    .Q(\datapath_1.regfile_1.regOut[11] [15]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _8236_ (
    .CLK(clk_bF$buf9),
    .D(_653_[16]),
    .Q(\datapath_1.regfile_1.regOut[11] [16]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _8237_ (
    .CLK(clk_bF$buf8),
    .D(_653_[17]),
    .Q(\datapath_1.regfile_1.regOut[11] [17]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _8238_ (
    .CLK(clk_bF$buf7),
    .D(_653_[18]),
    .Q(\datapath_1.regfile_1.regOut[11] [18]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _8239_ (
    .CLK(clk_bF$buf6),
    .D(_653_[19]),
    .Q(\datapath_1.regfile_1.regOut[11] [19]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _8240_ (
    .CLK(clk_bF$buf5),
    .D(_653_[20]),
    .Q(\datapath_1.regfile_1.regOut[11] [20]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _8241_ (
    .CLK(clk_bF$buf4),
    .D(_653_[21]),
    .Q(\datapath_1.regfile_1.regOut[11] [21]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _8242_ (
    .CLK(clk_bF$buf3),
    .D(_653_[22]),
    .Q(\datapath_1.regfile_1.regOut[11] [22]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _8243_ (
    .CLK(clk_bF$buf2),
    .D(_653_[23]),
    .Q(\datapath_1.regfile_1.regOut[11] [23]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _8244_ (
    .CLK(clk_bF$buf1),
    .D(_653_[24]),
    .Q(\datapath_1.regfile_1.regOut[11] [24]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _8245_ (
    .CLK(clk_bF$buf0),
    .D(_653_[25]),
    .Q(\datapath_1.regfile_1.regOut[11] [25]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _8246_ (
    .CLK(clk_bF$buf113),
    .D(_653_[26]),
    .Q(\datapath_1.regfile_1.regOut[11] [26]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _8247_ (
    .CLK(clk_bF$buf112),
    .D(_653_[27]),
    .Q(\datapath_1.regfile_1.regOut[11] [27]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _8248_ (
    .CLK(clk_bF$buf111),
    .D(_653_[28]),
    .Q(\datapath_1.regfile_1.regOut[11] [28]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _8249_ (
    .CLK(clk_bF$buf110),
    .D(_653_[29]),
    .Q(\datapath_1.regfile_1.regOut[11] [29]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _8250_ (
    .CLK(clk_bF$buf109),
    .D(_653_[30]),
    .Q(\datapath_1.regfile_1.regOut[11] [30]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _8251_ (
    .CLK(clk_bF$buf108),
    .D(_653_[31]),
    .Q(\datapath_1.regfile_1.regOut[11] [31]),
    .R(rst_bF$buf108),
    .S(vdd)
);

INVX1 _8252_ (
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_781_)
);

NAND2X1 _8253_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .Y(_782_)
);

OAI21X1 _8254_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_781_),
    .C(_782_),
    .Y(_718_[0])
);

INVX1 _8255_ (
    .A(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_719_)
);

NAND2X1 _8256_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_720_)
);

OAI21X1 _8257_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_719_),
    .C(_720_),
    .Y(_718_[1])
);

INVX1 _8258_ (
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_721_)
);

NAND2X1 _8259_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_722_)
);

OAI21X1 _8260_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_721_),
    .C(_722_),
    .Y(_718_[2])
);

INVX1 _8261_ (
    .A(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_723_)
);

NAND2X1 _8262_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_724_)
);

OAI21X1 _8263_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_723_),
    .C(_724_),
    .Y(_718_[3])
);

INVX1 _8264_ (
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_725_)
);

NAND2X1 _8265_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_726_)
);

OAI21X1 _8266_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_725_),
    .C(_726_),
    .Y(_718_[4])
);

INVX1 _8267_ (
    .A(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_727_)
);

NAND2X1 _8268_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_728_)
);

OAI21X1 _8269_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_727_),
    .C(_728_),
    .Y(_718_[5])
);

INVX1 _8270_ (
    .A(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_729_)
);

NAND2X1 _8271_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_730_)
);

OAI21X1 _8272_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_729_),
    .C(_730_),
    .Y(_718_[6])
);

INVX1 _8273_ (
    .A(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_731_)
);

NAND2X1 _8274_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_732_)
);

OAI21X1 _8275_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_731_),
    .C(_732_),
    .Y(_718_[7])
);

INVX1 _8276_ (
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_733_)
);

NAND2X1 _8277_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_734_)
);

OAI21X1 _8278_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_733_),
    .C(_734_),
    .Y(_718_[8])
);

INVX1 _8279_ (
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_735_)
);

NAND2X1 _8280_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_736_)
);

OAI21X1 _8281_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_735_),
    .C(_736_),
    .Y(_718_[9])
);

INVX1 _8282_ (
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_737_)
);

NAND2X1 _8283_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_738_)
);

OAI21X1 _8284_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_737_),
    .C(_738_),
    .Y(_718_[10])
);

INVX1 _8285_ (
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_739_)
);

NAND2X1 _8286_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_740_)
);

OAI21X1 _8287_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_739_),
    .C(_740_),
    .Y(_718_[11])
);

INVX1 _8288_ (
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_741_)
);

NAND2X1 _8289_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_742_)
);

OAI21X1 _8290_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_741_),
    .C(_742_),
    .Y(_718_[12])
);

INVX1 _8291_ (
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_743_)
);

NAND2X1 _8292_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_744_)
);

OAI21X1 _8293_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_743_),
    .C(_744_),
    .Y(_718_[13])
);

INVX1 _8294_ (
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_745_)
);

NAND2X1 _8295_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_746_)
);

OAI21X1 _8296_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_745_),
    .C(_746_),
    .Y(_718_[14])
);

INVX1 _8297_ (
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_747_)
);

NAND2X1 _8298_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_748_)
);

OAI21X1 _8299_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_747_),
    .C(_748_),
    .Y(_718_[15])
);

INVX1 _8300_ (
    .A(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_749_)
);

NAND2X1 _8301_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_750_)
);

OAI21X1 _8302_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_749_),
    .C(_750_),
    .Y(_718_[16])
);

INVX1 _8303_ (
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_751_)
);

NAND2X1 _8304_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_752_)
);

OAI21X1 _8305_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_751_),
    .C(_752_),
    .Y(_718_[17])
);

INVX1 _8306_ (
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_753_)
);

NAND2X1 _8307_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_754_)
);

OAI21X1 _8308_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_753_),
    .C(_754_),
    .Y(_718_[18])
);

INVX1 _8309_ (
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_755_)
);

NAND2X1 _8310_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_756_)
);

OAI21X1 _8311_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_755_),
    .C(_756_),
    .Y(_718_[19])
);

INVX1 _8312_ (
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_757_)
);

NAND2X1 _8313_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_758_)
);

OAI21X1 _8314_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_757_),
    .C(_758_),
    .Y(_718_[20])
);

INVX1 _8315_ (
    .A(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_759_)
);

NAND2X1 _8316_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_760_)
);

OAI21X1 _8317_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_759_),
    .C(_760_),
    .Y(_718_[21])
);

INVX1 _8318_ (
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_761_)
);

NAND2X1 _8319_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_762_)
);

OAI21X1 _8320_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_761_),
    .C(_762_),
    .Y(_718_[22])
);

INVX1 _8321_ (
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_763_)
);

NAND2X1 _8322_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_764_)
);

OAI21X1 _8323_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_763_),
    .C(_764_),
    .Y(_718_[23])
);

INVX1 _8324_ (
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_765_)
);

NAND2X1 _8325_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_766_)
);

OAI21X1 _8326_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_765_),
    .C(_766_),
    .Y(_718_[24])
);

INVX1 _8327_ (
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_767_)
);

NAND2X1 _8328_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_768_)
);

OAI21X1 _8329_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_767_),
    .C(_768_),
    .Y(_718_[25])
);

INVX1 _8330_ (
    .A(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_769_)
);

NAND2X1 _8331_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_770_)
);

OAI21X1 _8332_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_769_),
    .C(_770_),
    .Y(_718_[26])
);

INVX1 _8333_ (
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_771_)
);

NAND2X1 _8334_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_772_)
);

OAI21X1 _8335_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_771_),
    .C(_772_),
    .Y(_718_[27])
);

INVX1 _8336_ (
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_773_)
);

NAND2X1 _8337_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_774_)
);

OAI21X1 _8338_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(_773_),
    .C(_774_),
    .Y(_718_[28])
);

INVX1 _8339_ (
    .A(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_775_)
);

NAND2X1 _8340_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_776_)
);

OAI21X1 _8341_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(_775_),
    .C(_776_),
    .Y(_718_[29])
);

INVX1 _8342_ (
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_777_)
);

NAND2X1 _8343_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_778_)
);

OAI21X1 _8344_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(_777_),
    .C(_778_),
    .Y(_718_[30])
);

INVX1 _8345_ (
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_779_)
);

NAND2X1 _8346_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_780_)
);

OAI21X1 _8347_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(_779_),
    .C(_780_),
    .Y(_718_[31])
);

DFFSR _8348_ (
    .CLK(clk_bF$buf107),
    .D(_718_[0]),
    .Q(\datapath_1.regfile_1.regOut[12] [0]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _8349_ (
    .CLK(clk_bF$buf106),
    .D(_718_[1]),
    .Q(\datapath_1.regfile_1.regOut[12] [1]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _8350_ (
    .CLK(clk_bF$buf105),
    .D(_718_[2]),
    .Q(\datapath_1.regfile_1.regOut[12] [2]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _8351_ (
    .CLK(clk_bF$buf104),
    .D(_718_[3]),
    .Q(\datapath_1.regfile_1.regOut[12] [3]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _8352_ (
    .CLK(clk_bF$buf103),
    .D(_718_[4]),
    .Q(\datapath_1.regfile_1.regOut[12] [4]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _8353_ (
    .CLK(clk_bF$buf102),
    .D(_718_[5]),
    .Q(\datapath_1.regfile_1.regOut[12] [5]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _8354_ (
    .CLK(clk_bF$buf101),
    .D(_718_[6]),
    .Q(\datapath_1.regfile_1.regOut[12] [6]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _8355_ (
    .CLK(clk_bF$buf100),
    .D(_718_[7]),
    .Q(\datapath_1.regfile_1.regOut[12] [7]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _8356_ (
    .CLK(clk_bF$buf99),
    .D(_718_[8]),
    .Q(\datapath_1.regfile_1.regOut[12] [8]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _8357_ (
    .CLK(clk_bF$buf98),
    .D(_718_[9]),
    .Q(\datapath_1.regfile_1.regOut[12] [9]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _8358_ (
    .CLK(clk_bF$buf97),
    .D(_718_[10]),
    .Q(\datapath_1.regfile_1.regOut[12] [10]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _8359_ (
    .CLK(clk_bF$buf96),
    .D(_718_[11]),
    .Q(\datapath_1.regfile_1.regOut[12] [11]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _8360_ (
    .CLK(clk_bF$buf95),
    .D(_718_[12]),
    .Q(\datapath_1.regfile_1.regOut[12] [12]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _8361_ (
    .CLK(clk_bF$buf94),
    .D(_718_[13]),
    .Q(\datapath_1.regfile_1.regOut[12] [13]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _8362_ (
    .CLK(clk_bF$buf93),
    .D(_718_[14]),
    .Q(\datapath_1.regfile_1.regOut[12] [14]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _8363_ (
    .CLK(clk_bF$buf92),
    .D(_718_[15]),
    .Q(\datapath_1.regfile_1.regOut[12] [15]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _8364_ (
    .CLK(clk_bF$buf91),
    .D(_718_[16]),
    .Q(\datapath_1.regfile_1.regOut[12] [16]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _8365_ (
    .CLK(clk_bF$buf90),
    .D(_718_[17]),
    .Q(\datapath_1.regfile_1.regOut[12] [17]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _8366_ (
    .CLK(clk_bF$buf89),
    .D(_718_[18]),
    .Q(\datapath_1.regfile_1.regOut[12] [18]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _8367_ (
    .CLK(clk_bF$buf88),
    .D(_718_[19]),
    .Q(\datapath_1.regfile_1.regOut[12] [19]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _8368_ (
    .CLK(clk_bF$buf87),
    .D(_718_[20]),
    .Q(\datapath_1.regfile_1.regOut[12] [20]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _8369_ (
    .CLK(clk_bF$buf86),
    .D(_718_[21]),
    .Q(\datapath_1.regfile_1.regOut[12] [21]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _8370_ (
    .CLK(clk_bF$buf85),
    .D(_718_[22]),
    .Q(\datapath_1.regfile_1.regOut[12] [22]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _8371_ (
    .CLK(clk_bF$buf84),
    .D(_718_[23]),
    .Q(\datapath_1.regfile_1.regOut[12] [23]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _8372_ (
    .CLK(clk_bF$buf83),
    .D(_718_[24]),
    .Q(\datapath_1.regfile_1.regOut[12] [24]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _8373_ (
    .CLK(clk_bF$buf82),
    .D(_718_[25]),
    .Q(\datapath_1.regfile_1.regOut[12] [25]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _8374_ (
    .CLK(clk_bF$buf81),
    .D(_718_[26]),
    .Q(\datapath_1.regfile_1.regOut[12] [26]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _8375_ (
    .CLK(clk_bF$buf80),
    .D(_718_[27]),
    .Q(\datapath_1.regfile_1.regOut[12] [27]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _8376_ (
    .CLK(clk_bF$buf79),
    .D(_718_[28]),
    .Q(\datapath_1.regfile_1.regOut[12] [28]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _8377_ (
    .CLK(clk_bF$buf78),
    .D(_718_[29]),
    .Q(\datapath_1.regfile_1.regOut[12] [29]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _8378_ (
    .CLK(clk_bF$buf77),
    .D(_718_[30]),
    .Q(\datapath_1.regfile_1.regOut[12] [30]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _8379_ (
    .CLK(clk_bF$buf76),
    .D(_718_[31]),
    .Q(\datapath_1.regfile_1.regOut[12] [31]),
    .R(rst_bF$buf76),
    .S(vdd)
);

INVX1 _8380_ (
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_846_)
);

NAND2X1 _8381_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .Y(_847_)
);

OAI21X1 _8382_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_846_),
    .C(_847_),
    .Y(_783_[0])
);

INVX1 _8383_ (
    .A(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_784_)
);

NAND2X1 _8384_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_785_)
);

OAI21X1 _8385_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_784_),
    .C(_785_),
    .Y(_783_[1])
);

INVX1 _8386_ (
    .A(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_786_)
);

NAND2X1 _8387_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_787_)
);

OAI21X1 _8388_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_786_),
    .C(_787_),
    .Y(_783_[2])
);

INVX1 _8389_ (
    .A(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_788_)
);

NAND2X1 _8390_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_789_)
);

OAI21X1 _8391_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_788_),
    .C(_789_),
    .Y(_783_[3])
);

INVX1 _8392_ (
    .A(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_790_)
);

NAND2X1 _8393_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_791_)
);

OAI21X1 _8394_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_790_),
    .C(_791_),
    .Y(_783_[4])
);

INVX1 _8395_ (
    .A(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_792_)
);

NAND2X1 _8396_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_793_)
);

OAI21X1 _8397_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_792_),
    .C(_793_),
    .Y(_783_[5])
);

INVX1 _8398_ (
    .A(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_794_)
);

NAND2X1 _8399_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_795_)
);

OAI21X1 _8400_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_794_),
    .C(_795_),
    .Y(_783_[6])
);

INVX1 _8401_ (
    .A(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_796_)
);

NAND2X1 _8402_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_797_)
);

OAI21X1 _8403_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_796_),
    .C(_797_),
    .Y(_783_[7])
);

INVX1 _8404_ (
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_798_)
);

NAND2X1 _8405_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_799_)
);

OAI21X1 _8406_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_798_),
    .C(_799_),
    .Y(_783_[8])
);

INVX1 _8407_ (
    .A(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_800_)
);

NAND2X1 _8408_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_801_)
);

OAI21X1 _8409_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_800_),
    .C(_801_),
    .Y(_783_[9])
);

INVX1 _8410_ (
    .A(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_802_)
);

NAND2X1 _8411_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_803_)
);

OAI21X1 _8412_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_802_),
    .C(_803_),
    .Y(_783_[10])
);

INVX1 _8413_ (
    .A(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_804_)
);

NAND2X1 _8414_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_805_)
);

OAI21X1 _8415_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_804_),
    .C(_805_),
    .Y(_783_[11])
);

INVX1 _8416_ (
    .A(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_806_)
);

NAND2X1 _8417_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_807_)
);

OAI21X1 _8418_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_806_),
    .C(_807_),
    .Y(_783_[12])
);

INVX1 _8419_ (
    .A(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_808_)
);

NAND2X1 _8420_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_809_)
);

OAI21X1 _8421_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_808_),
    .C(_809_),
    .Y(_783_[13])
);

INVX1 _8422_ (
    .A(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_810_)
);

NAND2X1 _8423_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_811_)
);

OAI21X1 _8424_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_810_),
    .C(_811_),
    .Y(_783_[14])
);

INVX1 _8425_ (
    .A(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_812_)
);

NAND2X1 _8426_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_813_)
);

OAI21X1 _8427_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_812_),
    .C(_813_),
    .Y(_783_[15])
);

INVX1 _8428_ (
    .A(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_814_)
);

NAND2X1 _8429_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_815_)
);

OAI21X1 _8430_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_814_),
    .C(_815_),
    .Y(_783_[16])
);

INVX1 _8431_ (
    .A(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_816_)
);

NAND2X1 _8432_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_817_)
);

OAI21X1 _8433_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_816_),
    .C(_817_),
    .Y(_783_[17])
);

INVX1 _8434_ (
    .A(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_818_)
);

NAND2X1 _8435_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_819_)
);

OAI21X1 _8436_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_818_),
    .C(_819_),
    .Y(_783_[18])
);

INVX1 _8437_ (
    .A(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_820_)
);

NAND2X1 _8438_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_821_)
);

OAI21X1 _8439_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_820_),
    .C(_821_),
    .Y(_783_[19])
);

INVX1 _8440_ (
    .A(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_822_)
);

NAND2X1 _8441_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_823_)
);

OAI21X1 _8442_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_822_),
    .C(_823_),
    .Y(_783_[20])
);

INVX1 _8443_ (
    .A(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_824_)
);

NAND2X1 _8444_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_825_)
);

OAI21X1 _8445_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_824_),
    .C(_825_),
    .Y(_783_[21])
);

INVX1 _8446_ (
    .A(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_826_)
);

NAND2X1 _8447_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_827_)
);

OAI21X1 _8448_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_826_),
    .C(_827_),
    .Y(_783_[22])
);

INVX1 _8449_ (
    .A(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_828_)
);

NAND2X1 _8450_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_829_)
);

OAI21X1 _8451_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_828_),
    .C(_829_),
    .Y(_783_[23])
);

INVX1 _8452_ (
    .A(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_830_)
);

NAND2X1 _8453_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_831_)
);

OAI21X1 _8454_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_830_),
    .C(_831_),
    .Y(_783_[24])
);

INVX1 _8455_ (
    .A(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_832_)
);

NAND2X1 _8456_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_833_)
);

OAI21X1 _8457_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_832_),
    .C(_833_),
    .Y(_783_[25])
);

INVX1 _8458_ (
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_834_)
);

NAND2X1 _8459_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_835_)
);

OAI21X1 _8460_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_834_),
    .C(_835_),
    .Y(_783_[26])
);

INVX1 _8461_ (
    .A(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_836_)
);

NAND2X1 _8462_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_837_)
);

OAI21X1 _8463_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_836_),
    .C(_837_),
    .Y(_783_[27])
);

INVX1 _8464_ (
    .A(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_838_)
);

NAND2X1 _8465_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_839_)
);

OAI21X1 _8466_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(_838_),
    .C(_839_),
    .Y(_783_[28])
);

INVX1 _8467_ (
    .A(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_840_)
);

NAND2X1 _8468_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_841_)
);

OAI21X1 _8469_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(_840_),
    .C(_841_),
    .Y(_783_[29])
);

INVX1 _8470_ (
    .A(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_842_)
);

NAND2X1 _8471_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_843_)
);

OAI21X1 _8472_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(_842_),
    .C(_843_),
    .Y(_783_[30])
);

INVX1 _8473_ (
    .A(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_844_)
);

NAND2X1 _8474_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_845_)
);

OAI21X1 _8475_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(_844_),
    .C(_845_),
    .Y(_783_[31])
);

DFFSR _8476_ (
    .CLK(clk_bF$buf75),
    .D(_783_[0]),
    .Q(\datapath_1.regfile_1.regOut[13] [0]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _8477_ (
    .CLK(clk_bF$buf74),
    .D(_783_[1]),
    .Q(\datapath_1.regfile_1.regOut[13] [1]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _8478_ (
    .CLK(clk_bF$buf73),
    .D(_783_[2]),
    .Q(\datapath_1.regfile_1.regOut[13] [2]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _8479_ (
    .CLK(clk_bF$buf72),
    .D(_783_[3]),
    .Q(\datapath_1.regfile_1.regOut[13] [3]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _8480_ (
    .CLK(clk_bF$buf71),
    .D(_783_[4]),
    .Q(\datapath_1.regfile_1.regOut[13] [4]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _8481_ (
    .CLK(clk_bF$buf70),
    .D(_783_[5]),
    .Q(\datapath_1.regfile_1.regOut[13] [5]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _8482_ (
    .CLK(clk_bF$buf69),
    .D(_783_[6]),
    .Q(\datapath_1.regfile_1.regOut[13] [6]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _8483_ (
    .CLK(clk_bF$buf68),
    .D(_783_[7]),
    .Q(\datapath_1.regfile_1.regOut[13] [7]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _8484_ (
    .CLK(clk_bF$buf67),
    .D(_783_[8]),
    .Q(\datapath_1.regfile_1.regOut[13] [8]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _8485_ (
    .CLK(clk_bF$buf66),
    .D(_783_[9]),
    .Q(\datapath_1.regfile_1.regOut[13] [9]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _8486_ (
    .CLK(clk_bF$buf65),
    .D(_783_[10]),
    .Q(\datapath_1.regfile_1.regOut[13] [10]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _8487_ (
    .CLK(clk_bF$buf64),
    .D(_783_[11]),
    .Q(\datapath_1.regfile_1.regOut[13] [11]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _8488_ (
    .CLK(clk_bF$buf63),
    .D(_783_[12]),
    .Q(\datapath_1.regfile_1.regOut[13] [12]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _8489_ (
    .CLK(clk_bF$buf62),
    .D(_783_[13]),
    .Q(\datapath_1.regfile_1.regOut[13] [13]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _8490_ (
    .CLK(clk_bF$buf61),
    .D(_783_[14]),
    .Q(\datapath_1.regfile_1.regOut[13] [14]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _8491_ (
    .CLK(clk_bF$buf60),
    .D(_783_[15]),
    .Q(\datapath_1.regfile_1.regOut[13] [15]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _8492_ (
    .CLK(clk_bF$buf59),
    .D(_783_[16]),
    .Q(\datapath_1.regfile_1.regOut[13] [16]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _8493_ (
    .CLK(clk_bF$buf58),
    .D(_783_[17]),
    .Q(\datapath_1.regfile_1.regOut[13] [17]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _8494_ (
    .CLK(clk_bF$buf57),
    .D(_783_[18]),
    .Q(\datapath_1.regfile_1.regOut[13] [18]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _8495_ (
    .CLK(clk_bF$buf56),
    .D(_783_[19]),
    .Q(\datapath_1.regfile_1.regOut[13] [19]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _8496_ (
    .CLK(clk_bF$buf55),
    .D(_783_[20]),
    .Q(\datapath_1.regfile_1.regOut[13] [20]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _8497_ (
    .CLK(clk_bF$buf54),
    .D(_783_[21]),
    .Q(\datapath_1.regfile_1.regOut[13] [21]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _8498_ (
    .CLK(clk_bF$buf53),
    .D(_783_[22]),
    .Q(\datapath_1.regfile_1.regOut[13] [22]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _8499_ (
    .CLK(clk_bF$buf52),
    .D(_783_[23]),
    .Q(\datapath_1.regfile_1.regOut[13] [23]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _8500_ (
    .CLK(clk_bF$buf51),
    .D(_783_[24]),
    .Q(\datapath_1.regfile_1.regOut[13] [24]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _8501_ (
    .CLK(clk_bF$buf50),
    .D(_783_[25]),
    .Q(\datapath_1.regfile_1.regOut[13] [25]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _8502_ (
    .CLK(clk_bF$buf49),
    .D(_783_[26]),
    .Q(\datapath_1.regfile_1.regOut[13] [26]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _8503_ (
    .CLK(clk_bF$buf48),
    .D(_783_[27]),
    .Q(\datapath_1.regfile_1.regOut[13] [27]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _8504_ (
    .CLK(clk_bF$buf47),
    .D(_783_[28]),
    .Q(\datapath_1.regfile_1.regOut[13] [28]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _8505_ (
    .CLK(clk_bF$buf46),
    .D(_783_[29]),
    .Q(\datapath_1.regfile_1.regOut[13] [29]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _8506_ (
    .CLK(clk_bF$buf45),
    .D(_783_[30]),
    .Q(\datapath_1.regfile_1.regOut[13] [30]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _8507_ (
    .CLK(clk_bF$buf44),
    .D(_783_[31]),
    .Q(\datapath_1.regfile_1.regOut[13] [31]),
    .R(rst_bF$buf44),
    .S(vdd)
);

INVX1 _8508_ (
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_911_)
);

NAND2X1 _8509_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .Y(_912_)
);

OAI21X1 _8510_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_911_),
    .C(_912_),
    .Y(_848_[0])
);

INVX1 _8511_ (
    .A(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_849_)
);

NAND2X1 _8512_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_850_)
);

OAI21X1 _8513_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_849_),
    .C(_850_),
    .Y(_848_[1])
);

INVX1 _8514_ (
    .A(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_851_)
);

NAND2X1 _8515_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_852_)
);

OAI21X1 _8516_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_851_),
    .C(_852_),
    .Y(_848_[2])
);

INVX1 _8517_ (
    .A(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_853_)
);

NAND2X1 _8518_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_854_)
);

OAI21X1 _8519_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_853_),
    .C(_854_),
    .Y(_848_[3])
);

INVX1 _8520_ (
    .A(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_855_)
);

NAND2X1 _8521_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_856_)
);

OAI21X1 _8522_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_855_),
    .C(_856_),
    .Y(_848_[4])
);

INVX1 _8523_ (
    .A(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_857_)
);

NAND2X1 _8524_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_858_)
);

OAI21X1 _8525_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_857_),
    .C(_858_),
    .Y(_848_[5])
);

INVX1 _8526_ (
    .A(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_859_)
);

NAND2X1 _8527_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_860_)
);

OAI21X1 _8528_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_859_),
    .C(_860_),
    .Y(_848_[6])
);

INVX1 _8529_ (
    .A(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_861_)
);

NAND2X1 _8530_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_862_)
);

OAI21X1 _8531_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_861_),
    .C(_862_),
    .Y(_848_[7])
);

INVX1 _8532_ (
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_863_)
);

NAND2X1 _8533_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_864_)
);

OAI21X1 _8534_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_863_),
    .C(_864_),
    .Y(_848_[8])
);

INVX1 _8535_ (
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_865_)
);

NAND2X1 _8536_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_866_)
);

OAI21X1 _8537_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_865_),
    .C(_866_),
    .Y(_848_[9])
);

INVX1 _8538_ (
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_867_)
);

NAND2X1 _8539_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_868_)
);

OAI21X1 _8540_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_867_),
    .C(_868_),
    .Y(_848_[10])
);

INVX1 _8541_ (
    .A(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_869_)
);

NAND2X1 _8542_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_870_)
);

OAI21X1 _8543_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_869_),
    .C(_870_),
    .Y(_848_[11])
);

INVX1 _8544_ (
    .A(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_871_)
);

NAND2X1 _8545_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_872_)
);

OAI21X1 _8546_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_871_),
    .C(_872_),
    .Y(_848_[12])
);

INVX1 _8547_ (
    .A(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_873_)
);

NAND2X1 _8548_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_874_)
);

OAI21X1 _8549_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_873_),
    .C(_874_),
    .Y(_848_[13])
);

INVX1 _8550_ (
    .A(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_875_)
);

NAND2X1 _8551_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_876_)
);

OAI21X1 _8552_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_875_),
    .C(_876_),
    .Y(_848_[14])
);

INVX1 _8553_ (
    .A(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_877_)
);

NAND2X1 _8554_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_878_)
);

OAI21X1 _8555_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_877_),
    .C(_878_),
    .Y(_848_[15])
);

INVX1 _8556_ (
    .A(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_879_)
);

NAND2X1 _8557_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_880_)
);

OAI21X1 _8558_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_879_),
    .C(_880_),
    .Y(_848_[16])
);

INVX1 _8559_ (
    .A(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_881_)
);

NAND2X1 _8560_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_882_)
);

OAI21X1 _8561_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_881_),
    .C(_882_),
    .Y(_848_[17])
);

INVX1 _8562_ (
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_883_)
);

NAND2X1 _8563_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_884_)
);

OAI21X1 _8564_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_883_),
    .C(_884_),
    .Y(_848_[18])
);

INVX1 _8565_ (
    .A(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_885_)
);

NAND2X1 _8566_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_886_)
);

OAI21X1 _8567_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_885_),
    .C(_886_),
    .Y(_848_[19])
);

INVX1 _8568_ (
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_887_)
);

NAND2X1 _8569_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_888_)
);

OAI21X1 _8570_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_887_),
    .C(_888_),
    .Y(_848_[20])
);

INVX1 _8571_ (
    .A(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_889_)
);

NAND2X1 _8572_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_890_)
);

OAI21X1 _8573_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_889_),
    .C(_890_),
    .Y(_848_[21])
);

INVX1 _8574_ (
    .A(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_891_)
);

NAND2X1 _8575_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_892_)
);

OAI21X1 _8576_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_891_),
    .C(_892_),
    .Y(_848_[22])
);

INVX1 _8577_ (
    .A(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_893_)
);

NAND2X1 _8578_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_894_)
);

OAI21X1 _8579_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_893_),
    .C(_894_),
    .Y(_848_[23])
);

INVX1 _8580_ (
    .A(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_895_)
);

NAND2X1 _8581_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_896_)
);

OAI21X1 _8582_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_895_),
    .C(_896_),
    .Y(_848_[24])
);

INVX1 _8583_ (
    .A(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_897_)
);

NAND2X1 _8584_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_898_)
);

OAI21X1 _8585_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_897_),
    .C(_898_),
    .Y(_848_[25])
);

INVX1 _8586_ (
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_899_)
);

NAND2X1 _8587_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_900_)
);

OAI21X1 _8588_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_899_),
    .C(_900_),
    .Y(_848_[26])
);

INVX1 _8589_ (
    .A(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_901_)
);

NAND2X1 _8590_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_902_)
);

OAI21X1 _8591_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_901_),
    .C(_902_),
    .Y(_848_[27])
);

INVX1 _8592_ (
    .A(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_903_)
);

NAND2X1 _8593_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_904_)
);

OAI21X1 _8594_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(_903_),
    .C(_904_),
    .Y(_848_[28])
);

INVX1 _8595_ (
    .A(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_905_)
);

NAND2X1 _8596_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_906_)
);

OAI21X1 _8597_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(_905_),
    .C(_906_),
    .Y(_848_[29])
);

INVX1 _8598_ (
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_907_)
);

NAND2X1 _8599_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_908_)
);

OAI21X1 _8600_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(_907_),
    .C(_908_),
    .Y(_848_[30])
);

INVX1 _8601_ (
    .A(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_909_)
);

NAND2X1 _8602_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_910_)
);

OAI21X1 _8603_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(_909_),
    .C(_910_),
    .Y(_848_[31])
);

DFFSR _8604_ (
    .CLK(clk_bF$buf43),
    .D(_848_[0]),
    .Q(\datapath_1.regfile_1.regOut[14] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _8605_ (
    .CLK(clk_bF$buf42),
    .D(_848_[1]),
    .Q(\datapath_1.regfile_1.regOut[14] [1]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _8606_ (
    .CLK(clk_bF$buf41),
    .D(_848_[2]),
    .Q(\datapath_1.regfile_1.regOut[14] [2]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _8607_ (
    .CLK(clk_bF$buf40),
    .D(_848_[3]),
    .Q(\datapath_1.regfile_1.regOut[14] [3]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _8608_ (
    .CLK(clk_bF$buf39),
    .D(_848_[4]),
    .Q(\datapath_1.regfile_1.regOut[14] [4]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _8609_ (
    .CLK(clk_bF$buf38),
    .D(_848_[5]),
    .Q(\datapath_1.regfile_1.regOut[14] [5]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _8610_ (
    .CLK(clk_bF$buf37),
    .D(_848_[6]),
    .Q(\datapath_1.regfile_1.regOut[14] [6]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _8611_ (
    .CLK(clk_bF$buf36),
    .D(_848_[7]),
    .Q(\datapath_1.regfile_1.regOut[14] [7]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _8612_ (
    .CLK(clk_bF$buf35),
    .D(_848_[8]),
    .Q(\datapath_1.regfile_1.regOut[14] [8]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _8613_ (
    .CLK(clk_bF$buf34),
    .D(_848_[9]),
    .Q(\datapath_1.regfile_1.regOut[14] [9]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _8614_ (
    .CLK(clk_bF$buf33),
    .D(_848_[10]),
    .Q(\datapath_1.regfile_1.regOut[14] [10]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _8615_ (
    .CLK(clk_bF$buf32),
    .D(_848_[11]),
    .Q(\datapath_1.regfile_1.regOut[14] [11]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _8616_ (
    .CLK(clk_bF$buf31),
    .D(_848_[12]),
    .Q(\datapath_1.regfile_1.regOut[14] [12]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _8617_ (
    .CLK(clk_bF$buf30),
    .D(_848_[13]),
    .Q(\datapath_1.regfile_1.regOut[14] [13]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _8618_ (
    .CLK(clk_bF$buf29),
    .D(_848_[14]),
    .Q(\datapath_1.regfile_1.regOut[14] [14]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _8619_ (
    .CLK(clk_bF$buf28),
    .D(_848_[15]),
    .Q(\datapath_1.regfile_1.regOut[14] [15]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _8620_ (
    .CLK(clk_bF$buf27),
    .D(_848_[16]),
    .Q(\datapath_1.regfile_1.regOut[14] [16]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _8621_ (
    .CLK(clk_bF$buf26),
    .D(_848_[17]),
    .Q(\datapath_1.regfile_1.regOut[14] [17]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _8622_ (
    .CLK(clk_bF$buf25),
    .D(_848_[18]),
    .Q(\datapath_1.regfile_1.regOut[14] [18]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _8623_ (
    .CLK(clk_bF$buf24),
    .D(_848_[19]),
    .Q(\datapath_1.regfile_1.regOut[14] [19]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _8624_ (
    .CLK(clk_bF$buf23),
    .D(_848_[20]),
    .Q(\datapath_1.regfile_1.regOut[14] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _8625_ (
    .CLK(clk_bF$buf22),
    .D(_848_[21]),
    .Q(\datapath_1.regfile_1.regOut[14] [21]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _8626_ (
    .CLK(clk_bF$buf21),
    .D(_848_[22]),
    .Q(\datapath_1.regfile_1.regOut[14] [22]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _8627_ (
    .CLK(clk_bF$buf20),
    .D(_848_[23]),
    .Q(\datapath_1.regfile_1.regOut[14] [23]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _8628_ (
    .CLK(clk_bF$buf19),
    .D(_848_[24]),
    .Q(\datapath_1.regfile_1.regOut[14] [24]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _8629_ (
    .CLK(clk_bF$buf18),
    .D(_848_[25]),
    .Q(\datapath_1.regfile_1.regOut[14] [25]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _8630_ (
    .CLK(clk_bF$buf17),
    .D(_848_[26]),
    .Q(\datapath_1.regfile_1.regOut[14] [26]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _8631_ (
    .CLK(clk_bF$buf16),
    .D(_848_[27]),
    .Q(\datapath_1.regfile_1.regOut[14] [27]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _8632_ (
    .CLK(clk_bF$buf15),
    .D(_848_[28]),
    .Q(\datapath_1.regfile_1.regOut[14] [28]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _8633_ (
    .CLK(clk_bF$buf14),
    .D(_848_[29]),
    .Q(\datapath_1.regfile_1.regOut[14] [29]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _8634_ (
    .CLK(clk_bF$buf13),
    .D(_848_[30]),
    .Q(\datapath_1.regfile_1.regOut[14] [30]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _8635_ (
    .CLK(clk_bF$buf12),
    .D(_848_[31]),
    .Q(\datapath_1.regfile_1.regOut[14] [31]),
    .R(rst_bF$buf12),
    .S(vdd)
);

INVX1 _8636_ (
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_976_)
);

NAND2X1 _8637_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .Y(_977_)
);

OAI21X1 _8638_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_976_),
    .C(_977_),
    .Y(_913_[0])
);

INVX1 _8639_ (
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_914_)
);

NAND2X1 _8640_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_915_)
);

OAI21X1 _8641_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_914_),
    .C(_915_),
    .Y(_913_[1])
);

INVX1 _8642_ (
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_916_)
);

NAND2X1 _8643_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_917_)
);

OAI21X1 _8644_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_916_),
    .C(_917_),
    .Y(_913_[2])
);

INVX1 _8645_ (
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_918_)
);

NAND2X1 _8646_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_919_)
);

OAI21X1 _8647_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_918_),
    .C(_919_),
    .Y(_913_[3])
);

INVX1 _8648_ (
    .A(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_920_)
);

NAND2X1 _8649_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_921_)
);

OAI21X1 _8650_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_920_),
    .C(_921_),
    .Y(_913_[4])
);

INVX1 _8651_ (
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_922_)
);

NAND2X1 _8652_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_923_)
);

OAI21X1 _8653_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_922_),
    .C(_923_),
    .Y(_913_[5])
);

INVX1 _8654_ (
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_924_)
);

NAND2X1 _8655_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_925_)
);

OAI21X1 _8656_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_924_),
    .C(_925_),
    .Y(_913_[6])
);

INVX1 _8657_ (
    .A(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_926_)
);

NAND2X1 _8658_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_927_)
);

OAI21X1 _8659_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_926_),
    .C(_927_),
    .Y(_913_[7])
);

INVX1 _8660_ (
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_928_)
);

NAND2X1 _8661_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_929_)
);

OAI21X1 _8662_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_928_),
    .C(_929_),
    .Y(_913_[8])
);

INVX1 _8663_ (
    .A(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_930_)
);

NAND2X1 _8664_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_931_)
);

OAI21X1 _8665_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_930_),
    .C(_931_),
    .Y(_913_[9])
);

INVX1 _8666_ (
    .A(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_932_)
);

NAND2X1 _8667_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_933_)
);

OAI21X1 _8668_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_932_),
    .C(_933_),
    .Y(_913_[10])
);

INVX1 _8669_ (
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_934_)
);

NAND2X1 _8670_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_935_)
);

OAI21X1 _8671_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_934_),
    .C(_935_),
    .Y(_913_[11])
);

INVX1 _8672_ (
    .A(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_936_)
);

NAND2X1 _8673_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_937_)
);

OAI21X1 _8674_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_936_),
    .C(_937_),
    .Y(_913_[12])
);

INVX1 _8675_ (
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_938_)
);

NAND2X1 _8676_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_939_)
);

OAI21X1 _8677_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_938_),
    .C(_939_),
    .Y(_913_[13])
);

INVX1 _8678_ (
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_940_)
);

NAND2X1 _8679_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_941_)
);

OAI21X1 _8680_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_940_),
    .C(_941_),
    .Y(_913_[14])
);

INVX1 _8681_ (
    .A(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_942_)
);

NAND2X1 _8682_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_943_)
);

OAI21X1 _8683_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_942_),
    .C(_943_),
    .Y(_913_[15])
);

INVX1 _8684_ (
    .A(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_944_)
);

NAND2X1 _8685_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_945_)
);

OAI21X1 _8686_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_944_),
    .C(_945_),
    .Y(_913_[16])
);

INVX1 _8687_ (
    .A(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_946_)
);

NAND2X1 _8688_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_947_)
);

OAI21X1 _8689_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_946_),
    .C(_947_),
    .Y(_913_[17])
);

INVX1 _8690_ (
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_948_)
);

NAND2X1 _8691_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_949_)
);

OAI21X1 _8692_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_948_),
    .C(_949_),
    .Y(_913_[18])
);

INVX1 _8693_ (
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_950_)
);

NAND2X1 _8694_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_951_)
);

OAI21X1 _8695_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_950_),
    .C(_951_),
    .Y(_913_[19])
);

INVX1 _8696_ (
    .A(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_952_)
);

NAND2X1 _8697_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_953_)
);

OAI21X1 _8698_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_952_),
    .C(_953_),
    .Y(_913_[20])
);

INVX1 _8699_ (
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_954_)
);

NAND2X1 _8700_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_955_)
);

OAI21X1 _8701_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_954_),
    .C(_955_),
    .Y(_913_[21])
);

INVX1 _8702_ (
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_956_)
);

NAND2X1 _8703_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_957_)
);

OAI21X1 _8704_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_956_),
    .C(_957_),
    .Y(_913_[22])
);

INVX1 _8705_ (
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_958_)
);

NAND2X1 _8706_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_959_)
);

OAI21X1 _8707_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_958_),
    .C(_959_),
    .Y(_913_[23])
);

INVX1 _8708_ (
    .A(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_960_)
);

NAND2X1 _8709_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_961_)
);

OAI21X1 _8710_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_960_),
    .C(_961_),
    .Y(_913_[24])
);

INVX1 _8711_ (
    .A(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_962_)
);

NAND2X1 _8712_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_963_)
);

OAI21X1 _8713_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_962_),
    .C(_963_),
    .Y(_913_[25])
);

INVX1 _8714_ (
    .A(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_964_)
);

NAND2X1 _8715_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_965_)
);

OAI21X1 _8716_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_964_),
    .C(_965_),
    .Y(_913_[26])
);

INVX1 _8717_ (
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_966_)
);

NAND2X1 _8718_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_967_)
);

OAI21X1 _8719_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_966_),
    .C(_967_),
    .Y(_913_[27])
);

INVX1 _8720_ (
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_968_)
);

NAND2X1 _8721_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_969_)
);

OAI21X1 _8722_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(_968_),
    .C(_969_),
    .Y(_913_[28])
);

INVX1 _8723_ (
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_970_)
);

NAND2X1 _8724_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_971_)
);

OAI21X1 _8725_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(_970_),
    .C(_971_),
    .Y(_913_[29])
);

INVX1 _8726_ (
    .A(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_972_)
);

NAND2X1 _8727_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_973_)
);

OAI21X1 _8728_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(_972_),
    .C(_973_),
    .Y(_913_[30])
);

INVX1 _8729_ (
    .A(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_974_)
);

NAND2X1 _8730_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_975_)
);

OAI21X1 _8731_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(_974_),
    .C(_975_),
    .Y(_913_[31])
);

DFFSR _8732_ (
    .CLK(clk_bF$buf11),
    .D(_913_[0]),
    .Q(\datapath_1.regfile_1.regOut[15] [0]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _8733_ (
    .CLK(clk_bF$buf10),
    .D(_913_[1]),
    .Q(\datapath_1.regfile_1.regOut[15] [1]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _8734_ (
    .CLK(clk_bF$buf9),
    .D(_913_[2]),
    .Q(\datapath_1.regfile_1.regOut[15] [2]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _8735_ (
    .CLK(clk_bF$buf8),
    .D(_913_[3]),
    .Q(\datapath_1.regfile_1.regOut[15] [3]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _8736_ (
    .CLK(clk_bF$buf7),
    .D(_913_[4]),
    .Q(\datapath_1.regfile_1.regOut[15] [4]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _8737_ (
    .CLK(clk_bF$buf6),
    .D(_913_[5]),
    .Q(\datapath_1.regfile_1.regOut[15] [5]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _8738_ (
    .CLK(clk_bF$buf5),
    .D(_913_[6]),
    .Q(\datapath_1.regfile_1.regOut[15] [6]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _8739_ (
    .CLK(clk_bF$buf4),
    .D(_913_[7]),
    .Q(\datapath_1.regfile_1.regOut[15] [7]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _8740_ (
    .CLK(clk_bF$buf3),
    .D(_913_[8]),
    .Q(\datapath_1.regfile_1.regOut[15] [8]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _8741_ (
    .CLK(clk_bF$buf2),
    .D(_913_[9]),
    .Q(\datapath_1.regfile_1.regOut[15] [9]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _8742_ (
    .CLK(clk_bF$buf1),
    .D(_913_[10]),
    .Q(\datapath_1.regfile_1.regOut[15] [10]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _8743_ (
    .CLK(clk_bF$buf0),
    .D(_913_[11]),
    .Q(\datapath_1.regfile_1.regOut[15] [11]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _8744_ (
    .CLK(clk_bF$buf113),
    .D(_913_[12]),
    .Q(\datapath_1.regfile_1.regOut[15] [12]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _8745_ (
    .CLK(clk_bF$buf112),
    .D(_913_[13]),
    .Q(\datapath_1.regfile_1.regOut[15] [13]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _8746_ (
    .CLK(clk_bF$buf111),
    .D(_913_[14]),
    .Q(\datapath_1.regfile_1.regOut[15] [14]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _8747_ (
    .CLK(clk_bF$buf110),
    .D(_913_[15]),
    .Q(\datapath_1.regfile_1.regOut[15] [15]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _8748_ (
    .CLK(clk_bF$buf109),
    .D(_913_[16]),
    .Q(\datapath_1.regfile_1.regOut[15] [16]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _8749_ (
    .CLK(clk_bF$buf108),
    .D(_913_[17]),
    .Q(\datapath_1.regfile_1.regOut[15] [17]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _8750_ (
    .CLK(clk_bF$buf107),
    .D(_913_[18]),
    .Q(\datapath_1.regfile_1.regOut[15] [18]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _8751_ (
    .CLK(clk_bF$buf106),
    .D(_913_[19]),
    .Q(\datapath_1.regfile_1.regOut[15] [19]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _8752_ (
    .CLK(clk_bF$buf105),
    .D(_913_[20]),
    .Q(\datapath_1.regfile_1.regOut[15] [20]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _8753_ (
    .CLK(clk_bF$buf104),
    .D(_913_[21]),
    .Q(\datapath_1.regfile_1.regOut[15] [21]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _8754_ (
    .CLK(clk_bF$buf103),
    .D(_913_[22]),
    .Q(\datapath_1.regfile_1.regOut[15] [22]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _8755_ (
    .CLK(clk_bF$buf102),
    .D(_913_[23]),
    .Q(\datapath_1.regfile_1.regOut[15] [23]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _8756_ (
    .CLK(clk_bF$buf101),
    .D(_913_[24]),
    .Q(\datapath_1.regfile_1.regOut[15] [24]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _8757_ (
    .CLK(clk_bF$buf100),
    .D(_913_[25]),
    .Q(\datapath_1.regfile_1.regOut[15] [25]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _8758_ (
    .CLK(clk_bF$buf99),
    .D(_913_[26]),
    .Q(\datapath_1.regfile_1.regOut[15] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _8759_ (
    .CLK(clk_bF$buf98),
    .D(_913_[27]),
    .Q(\datapath_1.regfile_1.regOut[15] [27]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _8760_ (
    .CLK(clk_bF$buf97),
    .D(_913_[28]),
    .Q(\datapath_1.regfile_1.regOut[15] [28]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _8761_ (
    .CLK(clk_bF$buf96),
    .D(_913_[29]),
    .Q(\datapath_1.regfile_1.regOut[15] [29]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _8762_ (
    .CLK(clk_bF$buf95),
    .D(_913_[30]),
    .Q(\datapath_1.regfile_1.regOut[15] [30]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _8763_ (
    .CLK(clk_bF$buf94),
    .D(_913_[31]),
    .Q(\datapath_1.regfile_1.regOut[15] [31]),
    .R(rst_bF$buf94),
    .S(vdd)
);

INVX1 _8764_ (
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_1041_)
);

NAND2X1 _8765_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .Y(_1042_)
);

OAI21X1 _8766_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_1041_),
    .C(_1042_),
    .Y(_978_[0])
);

INVX1 _8767_ (
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_979_)
);

NAND2X1 _8768_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_980_)
);

OAI21X1 _8769_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_979_),
    .C(_980_),
    .Y(_978_[1])
);

INVX1 _8770_ (
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_981_)
);

NAND2X1 _8771_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_982_)
);

OAI21X1 _8772_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_981_),
    .C(_982_),
    .Y(_978_[2])
);

INVX1 _8773_ (
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_983_)
);

NAND2X1 _8774_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_984_)
);

OAI21X1 _8775_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_983_),
    .C(_984_),
    .Y(_978_[3])
);

INVX1 _8776_ (
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_985_)
);

NAND2X1 _8777_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_986_)
);

OAI21X1 _8778_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_985_),
    .C(_986_),
    .Y(_978_[4])
);

INVX1 _8779_ (
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_987_)
);

NAND2X1 _8780_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_988_)
);

OAI21X1 _8781_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_987_),
    .C(_988_),
    .Y(_978_[5])
);

INVX1 _8782_ (
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_989_)
);

NAND2X1 _8783_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_990_)
);

OAI21X1 _8784_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_989_),
    .C(_990_),
    .Y(_978_[6])
);

INVX1 _8785_ (
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_991_)
);

NAND2X1 _8786_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_992_)
);

OAI21X1 _8787_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_991_),
    .C(_992_),
    .Y(_978_[7])
);

INVX1 _8788_ (
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_993_)
);

NAND2X1 _8789_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_994_)
);

OAI21X1 _8790_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_993_),
    .C(_994_),
    .Y(_978_[8])
);

INVX1 _8791_ (
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_995_)
);

NAND2X1 _8792_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_996_)
);

OAI21X1 _8793_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_995_),
    .C(_996_),
    .Y(_978_[9])
);

INVX1 _8794_ (
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_997_)
);

NAND2X1 _8795_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_998_)
);

OAI21X1 _8796_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_997_),
    .C(_998_),
    .Y(_978_[10])
);

INVX1 _8797_ (
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_999_)
);

NAND2X1 _8798_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1000_)
);

OAI21X1 _8799_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_999_),
    .C(_1000_),
    .Y(_978_[11])
);

INVX1 _8800_ (
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_1001_)
);

NAND2X1 _8801_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1002_)
);

OAI21X1 _8802_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_1001_),
    .C(_1002_),
    .Y(_978_[12])
);

INVX1 _8803_ (
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_1003_)
);

NAND2X1 _8804_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1004_)
);

OAI21X1 _8805_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_1003_),
    .C(_1004_),
    .Y(_978_[13])
);

INVX1 _8806_ (
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_1005_)
);

NAND2X1 _8807_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1006_)
);

OAI21X1 _8808_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_1005_),
    .C(_1006_),
    .Y(_978_[14])
);

INVX1 _8809_ (
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_1007_)
);

NAND2X1 _8810_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1008_)
);

OAI21X1 _8811_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_1007_),
    .C(_1008_),
    .Y(_978_[15])
);

INVX1 _8812_ (
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_1009_)
);

NAND2X1 _8813_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1010_)
);

OAI21X1 _8814_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_1009_),
    .C(_1010_),
    .Y(_978_[16])
);

INVX1 _8815_ (
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_1011_)
);

NAND2X1 _8816_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1012_)
);

OAI21X1 _8817_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_1011_),
    .C(_1012_),
    .Y(_978_[17])
);

INVX1 _8818_ (
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_1013_)
);

NAND2X1 _8819_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1014_)
);

OAI21X1 _8820_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_1013_),
    .C(_1014_),
    .Y(_978_[18])
);

INVX1 _8821_ (
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_1015_)
);

NAND2X1 _8822_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1016_)
);

OAI21X1 _8823_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_1015_),
    .C(_1016_),
    .Y(_978_[19])
);

INVX1 _8824_ (
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_1017_)
);

NAND2X1 _8825_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1018_)
);

OAI21X1 _8826_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_1017_),
    .C(_1018_),
    .Y(_978_[20])
);

INVX1 _8827_ (
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_1019_)
);

NAND2X1 _8828_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1020_)
);

OAI21X1 _8829_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_1019_),
    .C(_1020_),
    .Y(_978_[21])
);

INVX1 _8830_ (
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_1021_)
);

NAND2X1 _8831_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1022_)
);

OAI21X1 _8832_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_1021_),
    .C(_1022_),
    .Y(_978_[22])
);

INVX1 _8833_ (
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_1023_)
);

NAND2X1 _8834_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1024_)
);

OAI21X1 _8835_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_1023_),
    .C(_1024_),
    .Y(_978_[23])
);

INVX1 _8836_ (
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_1025_)
);

NAND2X1 _8837_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1026_)
);

OAI21X1 _8838_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_1025_),
    .C(_1026_),
    .Y(_978_[24])
);

INVX1 _8839_ (
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_1027_)
);

NAND2X1 _8840_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_1028_)
);

OAI21X1 _8841_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_1027_),
    .C(_1028_),
    .Y(_978_[25])
);

INVX1 _8842_ (
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_1029_)
);

NAND2X1 _8843_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1030_)
);

OAI21X1 _8844_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_1029_),
    .C(_1030_),
    .Y(_978_[26])
);

INVX1 _8845_ (
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_1031_)
);

NAND2X1 _8846_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1032_)
);

OAI21X1 _8847_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_1031_),
    .C(_1032_),
    .Y(_978_[27])
);

INVX1 _8848_ (
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_1033_)
);

NAND2X1 _8849_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1034_)
);

OAI21X1 _8850_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(_1033_),
    .C(_1034_),
    .Y(_978_[28])
);

INVX1 _8851_ (
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_1035_)
);

NAND2X1 _8852_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1036_)
);

OAI21X1 _8853_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(_1035_),
    .C(_1036_),
    .Y(_978_[29])
);

INVX1 _8854_ (
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_1037_)
);

NAND2X1 _8855_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1038_)
);

OAI21X1 _8856_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(_1037_),
    .C(_1038_),
    .Y(_978_[30])
);

INVX1 _8857_ (
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_1039_)
);

NAND2X1 _8858_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1040_)
);

OAI21X1 _8859_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(_1039_),
    .C(_1040_),
    .Y(_978_[31])
);

DFFSR _8860_ (
    .CLK(clk_bF$buf93),
    .D(_978_[0]),
    .Q(\datapath_1.regfile_1.regOut[16] [0]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _8861_ (
    .CLK(clk_bF$buf92),
    .D(_978_[1]),
    .Q(\datapath_1.regfile_1.regOut[16] [1]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _8862_ (
    .CLK(clk_bF$buf91),
    .D(_978_[2]),
    .Q(\datapath_1.regfile_1.regOut[16] [2]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _8863_ (
    .CLK(clk_bF$buf90),
    .D(_978_[3]),
    .Q(\datapath_1.regfile_1.regOut[16] [3]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _8864_ (
    .CLK(clk_bF$buf89),
    .D(_978_[4]),
    .Q(\datapath_1.regfile_1.regOut[16] [4]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _8865_ (
    .CLK(clk_bF$buf88),
    .D(_978_[5]),
    .Q(\datapath_1.regfile_1.regOut[16] [5]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _8866_ (
    .CLK(clk_bF$buf87),
    .D(_978_[6]),
    .Q(\datapath_1.regfile_1.regOut[16] [6]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _8867_ (
    .CLK(clk_bF$buf86),
    .D(_978_[7]),
    .Q(\datapath_1.regfile_1.regOut[16] [7]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _8868_ (
    .CLK(clk_bF$buf85),
    .D(_978_[8]),
    .Q(\datapath_1.regfile_1.regOut[16] [8]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _8869_ (
    .CLK(clk_bF$buf84),
    .D(_978_[9]),
    .Q(\datapath_1.regfile_1.regOut[16] [9]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _8870_ (
    .CLK(clk_bF$buf83),
    .D(_978_[10]),
    .Q(\datapath_1.regfile_1.regOut[16] [10]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _8871_ (
    .CLK(clk_bF$buf82),
    .D(_978_[11]),
    .Q(\datapath_1.regfile_1.regOut[16] [11]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _8872_ (
    .CLK(clk_bF$buf81),
    .D(_978_[12]),
    .Q(\datapath_1.regfile_1.regOut[16] [12]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _8873_ (
    .CLK(clk_bF$buf80),
    .D(_978_[13]),
    .Q(\datapath_1.regfile_1.regOut[16] [13]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _8874_ (
    .CLK(clk_bF$buf79),
    .D(_978_[14]),
    .Q(\datapath_1.regfile_1.regOut[16] [14]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _8875_ (
    .CLK(clk_bF$buf78),
    .D(_978_[15]),
    .Q(\datapath_1.regfile_1.regOut[16] [15]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _8876_ (
    .CLK(clk_bF$buf77),
    .D(_978_[16]),
    .Q(\datapath_1.regfile_1.regOut[16] [16]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _8877_ (
    .CLK(clk_bF$buf76),
    .D(_978_[17]),
    .Q(\datapath_1.regfile_1.regOut[16] [17]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _8878_ (
    .CLK(clk_bF$buf75),
    .D(_978_[18]),
    .Q(\datapath_1.regfile_1.regOut[16] [18]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _8879_ (
    .CLK(clk_bF$buf74),
    .D(_978_[19]),
    .Q(\datapath_1.regfile_1.regOut[16] [19]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _8880_ (
    .CLK(clk_bF$buf73),
    .D(_978_[20]),
    .Q(\datapath_1.regfile_1.regOut[16] [20]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _8881_ (
    .CLK(clk_bF$buf72),
    .D(_978_[21]),
    .Q(\datapath_1.regfile_1.regOut[16] [21]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _8882_ (
    .CLK(clk_bF$buf71),
    .D(_978_[22]),
    .Q(\datapath_1.regfile_1.regOut[16] [22]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _8883_ (
    .CLK(clk_bF$buf70),
    .D(_978_[23]),
    .Q(\datapath_1.regfile_1.regOut[16] [23]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _8884_ (
    .CLK(clk_bF$buf69),
    .D(_978_[24]),
    .Q(\datapath_1.regfile_1.regOut[16] [24]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _8885_ (
    .CLK(clk_bF$buf68),
    .D(_978_[25]),
    .Q(\datapath_1.regfile_1.regOut[16] [25]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _8886_ (
    .CLK(clk_bF$buf67),
    .D(_978_[26]),
    .Q(\datapath_1.regfile_1.regOut[16] [26]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _8887_ (
    .CLK(clk_bF$buf66),
    .D(_978_[27]),
    .Q(\datapath_1.regfile_1.regOut[16] [27]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _8888_ (
    .CLK(clk_bF$buf65),
    .D(_978_[28]),
    .Q(\datapath_1.regfile_1.regOut[16] [28]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _8889_ (
    .CLK(clk_bF$buf64),
    .D(_978_[29]),
    .Q(\datapath_1.regfile_1.regOut[16] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _8890_ (
    .CLK(clk_bF$buf63),
    .D(_978_[30]),
    .Q(\datapath_1.regfile_1.regOut[16] [30]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _8891_ (
    .CLK(clk_bF$buf62),
    .D(_978_[31]),
    .Q(\datapath_1.regfile_1.regOut[16] [31]),
    .R(rst_bF$buf62),
    .S(vdd)
);

INVX1 _8892_ (
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_1106_)
);

NAND2X1 _8893_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .Y(_1107_)
);

OAI21X1 _8894_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1106_),
    .C(_1107_),
    .Y(_1043_[0])
);

INVX1 _8895_ (
    .A(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_1044_)
);

NAND2X1 _8896_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1045_)
);

OAI21X1 _8897_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1044_),
    .C(_1045_),
    .Y(_1043_[1])
);

INVX1 _8898_ (
    .A(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_1046_)
);

NAND2X1 _8899_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1047_)
);

OAI21X1 _8900_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1046_),
    .C(_1047_),
    .Y(_1043_[2])
);

INVX1 _8901_ (
    .A(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_1048_)
);

NAND2X1 _8902_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1049_)
);

OAI21X1 _8903_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1048_),
    .C(_1049_),
    .Y(_1043_[3])
);

INVX1 _8904_ (
    .A(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_1050_)
);

NAND2X1 _8905_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1051_)
);

OAI21X1 _8906_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1050_),
    .C(_1051_),
    .Y(_1043_[4])
);

INVX1 _8907_ (
    .A(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_1052_)
);

NAND2X1 _8908_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1053_)
);

OAI21X1 _8909_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1052_),
    .C(_1053_),
    .Y(_1043_[5])
);

INVX1 _8910_ (
    .A(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_1054_)
);

NAND2X1 _8911_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1055_)
);

OAI21X1 _8912_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1054_),
    .C(_1055_),
    .Y(_1043_[6])
);

INVX1 _8913_ (
    .A(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_1056_)
);

NAND2X1 _8914_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1057_)
);

OAI21X1 _8915_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1056_),
    .C(_1057_),
    .Y(_1043_[7])
);

INVX1 _8916_ (
    .A(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_1058_)
);

NAND2X1 _8917_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1059_)
);

OAI21X1 _8918_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1058_),
    .C(_1059_),
    .Y(_1043_[8])
);

INVX1 _8919_ (
    .A(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_1060_)
);

NAND2X1 _8920_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1061_)
);

OAI21X1 _8921_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1060_),
    .C(_1061_),
    .Y(_1043_[9])
);

INVX1 _8922_ (
    .A(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_1062_)
);

NAND2X1 _8923_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1063_)
);

OAI21X1 _8924_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1062_),
    .C(_1063_),
    .Y(_1043_[10])
);

INVX1 _8925_ (
    .A(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_1064_)
);

NAND2X1 _8926_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1065_)
);

OAI21X1 _8927_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1064_),
    .C(_1065_),
    .Y(_1043_[11])
);

INVX1 _8928_ (
    .A(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_1066_)
);

NAND2X1 _8929_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1067_)
);

OAI21X1 _8930_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1066_),
    .C(_1067_),
    .Y(_1043_[12])
);

INVX1 _8931_ (
    .A(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_1068_)
);

NAND2X1 _8932_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1069_)
);

OAI21X1 _8933_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1068_),
    .C(_1069_),
    .Y(_1043_[13])
);

INVX1 _8934_ (
    .A(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_1070_)
);

NAND2X1 _8935_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1071_)
);

OAI21X1 _8936_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1070_),
    .C(_1071_),
    .Y(_1043_[14])
);

INVX1 _8937_ (
    .A(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_1072_)
);

NAND2X1 _8938_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1073_)
);

OAI21X1 _8939_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1072_),
    .C(_1073_),
    .Y(_1043_[15])
);

INVX1 _8940_ (
    .A(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_1074_)
);

NAND2X1 _8941_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1075_)
);

OAI21X1 _8942_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1074_),
    .C(_1075_),
    .Y(_1043_[16])
);

INVX1 _8943_ (
    .A(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_1076_)
);

NAND2X1 _8944_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1077_)
);

OAI21X1 _8945_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1076_),
    .C(_1077_),
    .Y(_1043_[17])
);

INVX1 _8946_ (
    .A(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_1078_)
);

NAND2X1 _8947_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1079_)
);

OAI21X1 _8948_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1078_),
    .C(_1079_),
    .Y(_1043_[18])
);

INVX1 _8949_ (
    .A(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_1080_)
);

NAND2X1 _8950_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1081_)
);

OAI21X1 _8951_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1080_),
    .C(_1081_),
    .Y(_1043_[19])
);

INVX1 _8952_ (
    .A(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_1082_)
);

NAND2X1 _8953_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1083_)
);

OAI21X1 _8954_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1082_),
    .C(_1083_),
    .Y(_1043_[20])
);

INVX1 _8955_ (
    .A(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_1084_)
);

NAND2X1 _8956_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1085_)
);

OAI21X1 _8957_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1084_),
    .C(_1085_),
    .Y(_1043_[21])
);

INVX1 _8958_ (
    .A(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_1086_)
);

NAND2X1 _8959_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1087_)
);

OAI21X1 _8960_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1086_),
    .C(_1087_),
    .Y(_1043_[22])
);

INVX1 _8961_ (
    .A(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_1088_)
);

NAND2X1 _8962_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1089_)
);

OAI21X1 _8963_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1088_),
    .C(_1089_),
    .Y(_1043_[23])
);

INVX1 _8964_ (
    .A(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_1090_)
);

NAND2X1 _8965_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1091_)
);

OAI21X1 _8966_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1090_),
    .C(_1091_),
    .Y(_1043_[24])
);

INVX1 _8967_ (
    .A(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_1092_)
);

NAND2X1 _8968_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1093_)
);

OAI21X1 _8969_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1092_),
    .C(_1093_),
    .Y(_1043_[25])
);

INVX1 _8970_ (
    .A(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_1094_)
);

NAND2X1 _8971_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1095_)
);

OAI21X1 _8972_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1094_),
    .C(_1095_),
    .Y(_1043_[26])
);

INVX1 _8973_ (
    .A(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_1096_)
);

NAND2X1 _8974_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1097_)
);

OAI21X1 _8975_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1096_),
    .C(_1097_),
    .Y(_1043_[27])
);

INVX1 _8976_ (
    .A(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_1098_)
);

NAND2X1 _8977_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1099_)
);

OAI21X1 _8978_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(_1098_),
    .C(_1099_),
    .Y(_1043_[28])
);

INVX1 _8979_ (
    .A(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_1100_)
);

NAND2X1 _8980_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1101_)
);

OAI21X1 _8981_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(_1100_),
    .C(_1101_),
    .Y(_1043_[29])
);

INVX1 _8982_ (
    .A(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_1102_)
);

NAND2X1 _8983_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1103_)
);

OAI21X1 _8984_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(_1102_),
    .C(_1103_),
    .Y(_1043_[30])
);

INVX1 _8985_ (
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_1104_)
);

NAND2X1 _8986_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1105_)
);

OAI21X1 _8987_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(_1104_),
    .C(_1105_),
    .Y(_1043_[31])
);

DFFSR _8988_ (
    .CLK(clk_bF$buf61),
    .D(_1043_[0]),
    .Q(\datapath_1.regfile_1.regOut[17] [0]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _8989_ (
    .CLK(clk_bF$buf60),
    .D(_1043_[1]),
    .Q(\datapath_1.regfile_1.regOut[17] [1]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _8990_ (
    .CLK(clk_bF$buf59),
    .D(_1043_[2]),
    .Q(\datapath_1.regfile_1.regOut[17] [2]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _8991_ (
    .CLK(clk_bF$buf58),
    .D(_1043_[3]),
    .Q(\datapath_1.regfile_1.regOut[17] [3]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _8992_ (
    .CLK(clk_bF$buf57),
    .D(_1043_[4]),
    .Q(\datapath_1.regfile_1.regOut[17] [4]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _8993_ (
    .CLK(clk_bF$buf56),
    .D(_1043_[5]),
    .Q(\datapath_1.regfile_1.regOut[17] [5]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _8994_ (
    .CLK(clk_bF$buf55),
    .D(_1043_[6]),
    .Q(\datapath_1.regfile_1.regOut[17] [6]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _8995_ (
    .CLK(clk_bF$buf54),
    .D(_1043_[7]),
    .Q(\datapath_1.regfile_1.regOut[17] [7]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _8996_ (
    .CLK(clk_bF$buf53),
    .D(_1043_[8]),
    .Q(\datapath_1.regfile_1.regOut[17] [8]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _8997_ (
    .CLK(clk_bF$buf52),
    .D(_1043_[9]),
    .Q(\datapath_1.regfile_1.regOut[17] [9]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _8998_ (
    .CLK(clk_bF$buf51),
    .D(_1043_[10]),
    .Q(\datapath_1.regfile_1.regOut[17] [10]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _8999_ (
    .CLK(clk_bF$buf50),
    .D(_1043_[11]),
    .Q(\datapath_1.regfile_1.regOut[17] [11]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _9000_ (
    .CLK(clk_bF$buf49),
    .D(_1043_[12]),
    .Q(\datapath_1.regfile_1.regOut[17] [12]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _9001_ (
    .CLK(clk_bF$buf48),
    .D(_1043_[13]),
    .Q(\datapath_1.regfile_1.regOut[17] [13]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _9002_ (
    .CLK(clk_bF$buf47),
    .D(_1043_[14]),
    .Q(\datapath_1.regfile_1.regOut[17] [14]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _9003_ (
    .CLK(clk_bF$buf46),
    .D(_1043_[15]),
    .Q(\datapath_1.regfile_1.regOut[17] [15]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _9004_ (
    .CLK(clk_bF$buf45),
    .D(_1043_[16]),
    .Q(\datapath_1.regfile_1.regOut[17] [16]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _9005_ (
    .CLK(clk_bF$buf44),
    .D(_1043_[17]),
    .Q(\datapath_1.regfile_1.regOut[17] [17]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _9006_ (
    .CLK(clk_bF$buf43),
    .D(_1043_[18]),
    .Q(\datapath_1.regfile_1.regOut[17] [18]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _9007_ (
    .CLK(clk_bF$buf42),
    .D(_1043_[19]),
    .Q(\datapath_1.regfile_1.regOut[17] [19]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _9008_ (
    .CLK(clk_bF$buf41),
    .D(_1043_[20]),
    .Q(\datapath_1.regfile_1.regOut[17] [20]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _9009_ (
    .CLK(clk_bF$buf40),
    .D(_1043_[21]),
    .Q(\datapath_1.regfile_1.regOut[17] [21]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _9010_ (
    .CLK(clk_bF$buf39),
    .D(_1043_[22]),
    .Q(\datapath_1.regfile_1.regOut[17] [22]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _9011_ (
    .CLK(clk_bF$buf38),
    .D(_1043_[23]),
    .Q(\datapath_1.regfile_1.regOut[17] [23]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _9012_ (
    .CLK(clk_bF$buf37),
    .D(_1043_[24]),
    .Q(\datapath_1.regfile_1.regOut[17] [24]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _9013_ (
    .CLK(clk_bF$buf36),
    .D(_1043_[25]),
    .Q(\datapath_1.regfile_1.regOut[17] [25]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _9014_ (
    .CLK(clk_bF$buf35),
    .D(_1043_[26]),
    .Q(\datapath_1.regfile_1.regOut[17] [26]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _9015_ (
    .CLK(clk_bF$buf34),
    .D(_1043_[27]),
    .Q(\datapath_1.regfile_1.regOut[17] [27]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _9016_ (
    .CLK(clk_bF$buf33),
    .D(_1043_[28]),
    .Q(\datapath_1.regfile_1.regOut[17] [28]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _9017_ (
    .CLK(clk_bF$buf32),
    .D(_1043_[29]),
    .Q(\datapath_1.regfile_1.regOut[17] [29]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _9018_ (
    .CLK(clk_bF$buf31),
    .D(_1043_[30]),
    .Q(\datapath_1.regfile_1.regOut[17] [30]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _9019_ (
    .CLK(clk_bF$buf30),
    .D(_1043_[31]),
    .Q(\datapath_1.regfile_1.regOut[17] [31]),
    .R(rst_bF$buf30),
    .S(vdd)
);

INVX1 _9020_ (
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_1171_)
);

NAND2X1 _9021_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .Y(_1172_)
);

OAI21X1 _9022_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1171_),
    .C(_1172_),
    .Y(_1108_[0])
);

INVX1 _9023_ (
    .A(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_1109_)
);

NAND2X1 _9024_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1110_)
);

OAI21X1 _9025_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1109_),
    .C(_1110_),
    .Y(_1108_[1])
);

INVX1 _9026_ (
    .A(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_1111_)
);

NAND2X1 _9027_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1112_)
);

OAI21X1 _9028_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1111_),
    .C(_1112_),
    .Y(_1108_[2])
);

INVX1 _9029_ (
    .A(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_1113_)
);

NAND2X1 _9030_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1114_)
);

OAI21X1 _9031_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1113_),
    .C(_1114_),
    .Y(_1108_[3])
);

INVX1 _9032_ (
    .A(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_1115_)
);

NAND2X1 _9033_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1116_)
);

OAI21X1 _9034_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1115_),
    .C(_1116_),
    .Y(_1108_[4])
);

INVX1 _9035_ (
    .A(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_1117_)
);

NAND2X1 _9036_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1118_)
);

OAI21X1 _9037_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1117_),
    .C(_1118_),
    .Y(_1108_[5])
);

INVX1 _9038_ (
    .A(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_1119_)
);

NAND2X1 _9039_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1120_)
);

OAI21X1 _9040_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1119_),
    .C(_1120_),
    .Y(_1108_[6])
);

INVX1 _9041_ (
    .A(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_1121_)
);

NAND2X1 _9042_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1122_)
);

OAI21X1 _9043_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1121_),
    .C(_1122_),
    .Y(_1108_[7])
);

INVX1 _9044_ (
    .A(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_1123_)
);

NAND2X1 _9045_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1124_)
);

OAI21X1 _9046_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1123_),
    .C(_1124_),
    .Y(_1108_[8])
);

INVX1 _9047_ (
    .A(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_1125_)
);

NAND2X1 _9048_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1126_)
);

OAI21X1 _9049_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1125_),
    .C(_1126_),
    .Y(_1108_[9])
);

INVX1 _9050_ (
    .A(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_1127_)
);

NAND2X1 _9051_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1128_)
);

OAI21X1 _9052_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1127_),
    .C(_1128_),
    .Y(_1108_[10])
);

INVX1 _9053_ (
    .A(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_1129_)
);

NAND2X1 _9054_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1130_)
);

OAI21X1 _9055_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1129_),
    .C(_1130_),
    .Y(_1108_[11])
);

INVX1 _9056_ (
    .A(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_1131_)
);

NAND2X1 _9057_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1132_)
);

OAI21X1 _9058_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1131_),
    .C(_1132_),
    .Y(_1108_[12])
);

INVX1 _9059_ (
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_1133_)
);

NAND2X1 _9060_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1134_)
);

OAI21X1 _9061_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1133_),
    .C(_1134_),
    .Y(_1108_[13])
);

INVX1 _9062_ (
    .A(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_1135_)
);

NAND2X1 _9063_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1136_)
);

OAI21X1 _9064_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1135_),
    .C(_1136_),
    .Y(_1108_[14])
);

INVX1 _9065_ (
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_1137_)
);

NAND2X1 _9066_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1138_)
);

OAI21X1 _9067_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1137_),
    .C(_1138_),
    .Y(_1108_[15])
);

INVX1 _9068_ (
    .A(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_1139_)
);

NAND2X1 _9069_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1140_)
);

OAI21X1 _9070_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1139_),
    .C(_1140_),
    .Y(_1108_[16])
);

INVX1 _9071_ (
    .A(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_1141_)
);

NAND2X1 _9072_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1142_)
);

OAI21X1 _9073_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1141_),
    .C(_1142_),
    .Y(_1108_[17])
);

INVX1 _9074_ (
    .A(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_1143_)
);

NAND2X1 _9075_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1144_)
);

OAI21X1 _9076_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1143_),
    .C(_1144_),
    .Y(_1108_[18])
);

INVX1 _9077_ (
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_1145_)
);

NAND2X1 _9078_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1146_)
);

OAI21X1 _9079_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1145_),
    .C(_1146_),
    .Y(_1108_[19])
);

INVX1 _9080_ (
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_1147_)
);

NAND2X1 _9081_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1148_)
);

OAI21X1 _9082_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1147_),
    .C(_1148_),
    .Y(_1108_[20])
);

INVX1 _9083_ (
    .A(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_1149_)
);

NAND2X1 _9084_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1150_)
);

OAI21X1 _9085_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1149_),
    .C(_1150_),
    .Y(_1108_[21])
);

INVX1 _9086_ (
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_1151_)
);

NAND2X1 _9087_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_1152_)
);

OAI21X1 _9088_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1151_),
    .C(_1152_),
    .Y(_1108_[22])
);

INVX1 _9089_ (
    .A(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_1153_)
);

NAND2X1 _9090_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1154_)
);

OAI21X1 _9091_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1153_),
    .C(_1154_),
    .Y(_1108_[23])
);

INVX1 _9092_ (
    .A(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_1155_)
);

NAND2X1 _9093_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1156_)
);

OAI21X1 _9094_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1155_),
    .C(_1156_),
    .Y(_1108_[24])
);

INVX1 _9095_ (
    .A(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_1157_)
);

NAND2X1 _9096_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1158_)
);

OAI21X1 _9097_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1157_),
    .C(_1158_),
    .Y(_1108_[25])
);

INVX1 _9098_ (
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_1159_)
);

NAND2X1 _9099_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1160_)
);

OAI21X1 _9100_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1159_),
    .C(_1160_),
    .Y(_1108_[26])
);

INVX1 _9101_ (
    .A(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_1161_)
);

NAND2X1 _9102_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1162_)
);

OAI21X1 _9103_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1161_),
    .C(_1162_),
    .Y(_1108_[27])
);

INVX1 _9104_ (
    .A(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_1163_)
);

NAND2X1 _9105_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1164_)
);

OAI21X1 _9106_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(_1163_),
    .C(_1164_),
    .Y(_1108_[28])
);

INVX1 _9107_ (
    .A(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_1165_)
);

NAND2X1 _9108_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1166_)
);

OAI21X1 _9109_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(_1165_),
    .C(_1166_),
    .Y(_1108_[29])
);

INVX1 _9110_ (
    .A(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_1167_)
);

NAND2X1 _9111_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1168_)
);

OAI21X1 _9112_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(_1167_),
    .C(_1168_),
    .Y(_1108_[30])
);

INVX1 _9113_ (
    .A(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_1169_)
);

NAND2X1 _9114_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1170_)
);

OAI21X1 _9115_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(_1169_),
    .C(_1170_),
    .Y(_1108_[31])
);

DFFSR _9116_ (
    .CLK(clk_bF$buf29),
    .D(_1108_[0]),
    .Q(\datapath_1.regfile_1.regOut[18] [0]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _9117_ (
    .CLK(clk_bF$buf28),
    .D(_1108_[1]),
    .Q(\datapath_1.regfile_1.regOut[18] [1]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _9118_ (
    .CLK(clk_bF$buf27),
    .D(_1108_[2]),
    .Q(\datapath_1.regfile_1.regOut[18] [2]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _9119_ (
    .CLK(clk_bF$buf26),
    .D(_1108_[3]),
    .Q(\datapath_1.regfile_1.regOut[18] [3]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _9120_ (
    .CLK(clk_bF$buf25),
    .D(_1108_[4]),
    .Q(\datapath_1.regfile_1.regOut[18] [4]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _9121_ (
    .CLK(clk_bF$buf24),
    .D(_1108_[5]),
    .Q(\datapath_1.regfile_1.regOut[18] [5]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _9122_ (
    .CLK(clk_bF$buf23),
    .D(_1108_[6]),
    .Q(\datapath_1.regfile_1.regOut[18] [6]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _9123_ (
    .CLK(clk_bF$buf22),
    .D(_1108_[7]),
    .Q(\datapath_1.regfile_1.regOut[18] [7]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _9124_ (
    .CLK(clk_bF$buf21),
    .D(_1108_[8]),
    .Q(\datapath_1.regfile_1.regOut[18] [8]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _9125_ (
    .CLK(clk_bF$buf20),
    .D(_1108_[9]),
    .Q(\datapath_1.regfile_1.regOut[18] [9]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _9126_ (
    .CLK(clk_bF$buf19),
    .D(_1108_[10]),
    .Q(\datapath_1.regfile_1.regOut[18] [10]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _9127_ (
    .CLK(clk_bF$buf18),
    .D(_1108_[11]),
    .Q(\datapath_1.regfile_1.regOut[18] [11]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _9128_ (
    .CLK(clk_bF$buf17),
    .D(_1108_[12]),
    .Q(\datapath_1.regfile_1.regOut[18] [12]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _9129_ (
    .CLK(clk_bF$buf16),
    .D(_1108_[13]),
    .Q(\datapath_1.regfile_1.regOut[18] [13]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _9130_ (
    .CLK(clk_bF$buf15),
    .D(_1108_[14]),
    .Q(\datapath_1.regfile_1.regOut[18] [14]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _9131_ (
    .CLK(clk_bF$buf14),
    .D(_1108_[15]),
    .Q(\datapath_1.regfile_1.regOut[18] [15]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _9132_ (
    .CLK(clk_bF$buf13),
    .D(_1108_[16]),
    .Q(\datapath_1.regfile_1.regOut[18] [16]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _9133_ (
    .CLK(clk_bF$buf12),
    .D(_1108_[17]),
    .Q(\datapath_1.regfile_1.regOut[18] [17]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _9134_ (
    .CLK(clk_bF$buf11),
    .D(_1108_[18]),
    .Q(\datapath_1.regfile_1.regOut[18] [18]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _9135_ (
    .CLK(clk_bF$buf10),
    .D(_1108_[19]),
    .Q(\datapath_1.regfile_1.regOut[18] [19]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _9136_ (
    .CLK(clk_bF$buf9),
    .D(_1108_[20]),
    .Q(\datapath_1.regfile_1.regOut[18] [20]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _9137_ (
    .CLK(clk_bF$buf8),
    .D(_1108_[21]),
    .Q(\datapath_1.regfile_1.regOut[18] [21]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _9138_ (
    .CLK(clk_bF$buf7),
    .D(_1108_[22]),
    .Q(\datapath_1.regfile_1.regOut[18] [22]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _9139_ (
    .CLK(clk_bF$buf6),
    .D(_1108_[23]),
    .Q(\datapath_1.regfile_1.regOut[18] [23]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _9140_ (
    .CLK(clk_bF$buf5),
    .D(_1108_[24]),
    .Q(\datapath_1.regfile_1.regOut[18] [24]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _9141_ (
    .CLK(clk_bF$buf4),
    .D(_1108_[25]),
    .Q(\datapath_1.regfile_1.regOut[18] [25]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _9142_ (
    .CLK(clk_bF$buf3),
    .D(_1108_[26]),
    .Q(\datapath_1.regfile_1.regOut[18] [26]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _9143_ (
    .CLK(clk_bF$buf2),
    .D(_1108_[27]),
    .Q(\datapath_1.regfile_1.regOut[18] [27]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _9144_ (
    .CLK(clk_bF$buf1),
    .D(_1108_[28]),
    .Q(\datapath_1.regfile_1.regOut[18] [28]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _9145_ (
    .CLK(clk_bF$buf0),
    .D(_1108_[29]),
    .Q(\datapath_1.regfile_1.regOut[18] [29]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _9146_ (
    .CLK(clk_bF$buf113),
    .D(_1108_[30]),
    .Q(\datapath_1.regfile_1.regOut[18] [30]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _9147_ (
    .CLK(clk_bF$buf112),
    .D(_1108_[31]),
    .Q(\datapath_1.regfile_1.regOut[18] [31]),
    .R(rst_bF$buf112),
    .S(vdd)
);

INVX1 _9148_ (
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_1236_)
);

NAND2X1 _9149_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .Y(_1237_)
);

OAI21X1 _9150_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1236_),
    .C(_1237_),
    .Y(_1173_[0])
);

INVX1 _9151_ (
    .A(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_1174_)
);

NAND2X1 _9152_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1175_)
);

OAI21X1 _9153_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1174_),
    .C(_1175_),
    .Y(_1173_[1])
);

INVX1 _9154_ (
    .A(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_1176_)
);

NAND2X1 _9155_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1177_)
);

OAI21X1 _9156_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1176_),
    .C(_1177_),
    .Y(_1173_[2])
);

INVX1 _9157_ (
    .A(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_1178_)
);

NAND2X1 _9158_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1179_)
);

OAI21X1 _9159_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1178_),
    .C(_1179_),
    .Y(_1173_[3])
);

INVX1 _9160_ (
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_1180_)
);

NAND2X1 _9161_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1181_)
);

OAI21X1 _9162_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1180_),
    .C(_1181_),
    .Y(_1173_[4])
);

INVX1 _9163_ (
    .A(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_1182_)
);

NAND2X1 _9164_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1183_)
);

OAI21X1 _9165_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1182_),
    .C(_1183_),
    .Y(_1173_[5])
);

INVX1 _9166_ (
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_1184_)
);

NAND2X1 _9167_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1185_)
);

OAI21X1 _9168_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1184_),
    .C(_1185_),
    .Y(_1173_[6])
);

INVX1 _9169_ (
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_1186_)
);

NAND2X1 _9170_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1187_)
);

OAI21X1 _9171_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1186_),
    .C(_1187_),
    .Y(_1173_[7])
);

INVX1 _9172_ (
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_1188_)
);

NAND2X1 _9173_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1189_)
);

OAI21X1 _9174_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1188_),
    .C(_1189_),
    .Y(_1173_[8])
);

INVX1 _9175_ (
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_1190_)
);

NAND2X1 _9176_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1191_)
);

OAI21X1 _9177_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1190_),
    .C(_1191_),
    .Y(_1173_[9])
);

INVX1 _9178_ (
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_1192_)
);

NAND2X1 _9179_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1193_)
);

OAI21X1 _9180_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1192_),
    .C(_1193_),
    .Y(_1173_[10])
);

INVX1 _9181_ (
    .A(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_1194_)
);

NAND2X1 _9182_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1195_)
);

OAI21X1 _9183_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1194_),
    .C(_1195_),
    .Y(_1173_[11])
);

INVX1 _9184_ (
    .A(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_1196_)
);

NAND2X1 _9185_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1197_)
);

OAI21X1 _9186_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1196_),
    .C(_1197_),
    .Y(_1173_[12])
);

INVX1 _9187_ (
    .A(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_1198_)
);

NAND2X1 _9188_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1199_)
);

OAI21X1 _9189_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1198_),
    .C(_1199_),
    .Y(_1173_[13])
);

INVX1 _9190_ (
    .A(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_1200_)
);

NAND2X1 _9191_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1201_)
);

OAI21X1 _9192_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1200_),
    .C(_1201_),
    .Y(_1173_[14])
);

INVX1 _9193_ (
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_1202_)
);

NAND2X1 _9194_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1203_)
);

OAI21X1 _9195_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1202_),
    .C(_1203_),
    .Y(_1173_[15])
);

INVX1 _9196_ (
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_1204_)
);

NAND2X1 _9197_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1205_)
);

OAI21X1 _9198_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1204_),
    .C(_1205_),
    .Y(_1173_[16])
);

INVX1 _9199_ (
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_1206_)
);

NAND2X1 _9200_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1207_)
);

OAI21X1 _9201_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1206_),
    .C(_1207_),
    .Y(_1173_[17])
);

INVX1 _9202_ (
    .A(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_1208_)
);

NAND2X1 _9203_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1209_)
);

OAI21X1 _9204_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1208_),
    .C(_1209_),
    .Y(_1173_[18])
);

INVX1 _9205_ (
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_1210_)
);

NAND2X1 _9206_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1211_)
);

OAI21X1 _9207_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1210_),
    .C(_1211_),
    .Y(_1173_[19])
);

INVX1 _9208_ (
    .A(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_1212_)
);

NAND2X1 _9209_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1213_)
);

OAI21X1 _9210_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1212_),
    .C(_1213_),
    .Y(_1173_[20])
);

INVX1 _9211_ (
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_1214_)
);

NAND2X1 _9212_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1215_)
);

OAI21X1 _9213_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1214_),
    .C(_1215_),
    .Y(_1173_[21])
);

INVX1 _9214_ (
    .A(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_1216_)
);

NAND2X1 _9215_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1217_)
);

OAI21X1 _9216_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1216_),
    .C(_1217_),
    .Y(_1173_[22])
);

INVX1 _9217_ (
    .A(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_1218_)
);

NAND2X1 _9218_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1219_)
);

OAI21X1 _9219_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1218_),
    .C(_1219_),
    .Y(_1173_[23])
);

INVX1 _9220_ (
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_1220_)
);

NAND2X1 _9221_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1221_)
);

OAI21X1 _9222_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1220_),
    .C(_1221_),
    .Y(_1173_[24])
);

INVX1 _9223_ (
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_1222_)
);

NAND2X1 _9224_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1223_)
);

OAI21X1 _9225_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1222_),
    .C(_1223_),
    .Y(_1173_[25])
);

INVX1 _9226_ (
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_1224_)
);

NAND2X1 _9227_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1225_)
);

OAI21X1 _9228_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1224_),
    .C(_1225_),
    .Y(_1173_[26])
);

INVX1 _9229_ (
    .A(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_1226_)
);

NAND2X1 _9230_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1227_)
);

OAI21X1 _9231_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1226_),
    .C(_1227_),
    .Y(_1173_[27])
);

INVX1 _9232_ (
    .A(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_1228_)
);

NAND2X1 _9233_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1229_)
);

OAI21X1 _9234_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(_1228_),
    .C(_1229_),
    .Y(_1173_[28])
);

INVX1 _9235_ (
    .A(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_1230_)
);

NAND2X1 _9236_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1231_)
);

OAI21X1 _9237_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(_1230_),
    .C(_1231_),
    .Y(_1173_[29])
);

INVX1 _9238_ (
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_1232_)
);

NAND2X1 _9239_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1233_)
);

OAI21X1 _9240_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(_1232_),
    .C(_1233_),
    .Y(_1173_[30])
);

INVX1 _9241_ (
    .A(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_1234_)
);

NAND2X1 _9242_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1235_)
);

OAI21X1 _9243_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(_1234_),
    .C(_1235_),
    .Y(_1173_[31])
);

DFFSR _9244_ (
    .CLK(clk_bF$buf111),
    .D(_1173_[0]),
    .Q(\datapath_1.regfile_1.regOut[19] [0]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _9245_ (
    .CLK(clk_bF$buf110),
    .D(_1173_[1]),
    .Q(\datapath_1.regfile_1.regOut[19] [1]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _9246_ (
    .CLK(clk_bF$buf109),
    .D(_1173_[2]),
    .Q(\datapath_1.regfile_1.regOut[19] [2]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _9247_ (
    .CLK(clk_bF$buf108),
    .D(_1173_[3]),
    .Q(\datapath_1.regfile_1.regOut[19] [3]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _9248_ (
    .CLK(clk_bF$buf107),
    .D(_1173_[4]),
    .Q(\datapath_1.regfile_1.regOut[19] [4]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _9249_ (
    .CLK(clk_bF$buf106),
    .D(_1173_[5]),
    .Q(\datapath_1.regfile_1.regOut[19] [5]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _9250_ (
    .CLK(clk_bF$buf105),
    .D(_1173_[6]),
    .Q(\datapath_1.regfile_1.regOut[19] [6]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _9251_ (
    .CLK(clk_bF$buf104),
    .D(_1173_[7]),
    .Q(\datapath_1.regfile_1.regOut[19] [7]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _9252_ (
    .CLK(clk_bF$buf103),
    .D(_1173_[8]),
    .Q(\datapath_1.regfile_1.regOut[19] [8]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _9253_ (
    .CLK(clk_bF$buf102),
    .D(_1173_[9]),
    .Q(\datapath_1.regfile_1.regOut[19] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _9254_ (
    .CLK(clk_bF$buf101),
    .D(_1173_[10]),
    .Q(\datapath_1.regfile_1.regOut[19] [10]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _9255_ (
    .CLK(clk_bF$buf100),
    .D(_1173_[11]),
    .Q(\datapath_1.regfile_1.regOut[19] [11]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _9256_ (
    .CLK(clk_bF$buf99),
    .D(_1173_[12]),
    .Q(\datapath_1.regfile_1.regOut[19] [12]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _9257_ (
    .CLK(clk_bF$buf98),
    .D(_1173_[13]),
    .Q(\datapath_1.regfile_1.regOut[19] [13]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _9258_ (
    .CLK(clk_bF$buf97),
    .D(_1173_[14]),
    .Q(\datapath_1.regfile_1.regOut[19] [14]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _9259_ (
    .CLK(clk_bF$buf96),
    .D(_1173_[15]),
    .Q(\datapath_1.regfile_1.regOut[19] [15]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _9260_ (
    .CLK(clk_bF$buf95),
    .D(_1173_[16]),
    .Q(\datapath_1.regfile_1.regOut[19] [16]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _9261_ (
    .CLK(clk_bF$buf94),
    .D(_1173_[17]),
    .Q(\datapath_1.regfile_1.regOut[19] [17]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _9262_ (
    .CLK(clk_bF$buf93),
    .D(_1173_[18]),
    .Q(\datapath_1.regfile_1.regOut[19] [18]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _9263_ (
    .CLK(clk_bF$buf92),
    .D(_1173_[19]),
    .Q(\datapath_1.regfile_1.regOut[19] [19]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _9264_ (
    .CLK(clk_bF$buf91),
    .D(_1173_[20]),
    .Q(\datapath_1.regfile_1.regOut[19] [20]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _9265_ (
    .CLK(clk_bF$buf90),
    .D(_1173_[21]),
    .Q(\datapath_1.regfile_1.regOut[19] [21]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _9266_ (
    .CLK(clk_bF$buf89),
    .D(_1173_[22]),
    .Q(\datapath_1.regfile_1.regOut[19] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _9267_ (
    .CLK(clk_bF$buf88),
    .D(_1173_[23]),
    .Q(\datapath_1.regfile_1.regOut[19] [23]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _9268_ (
    .CLK(clk_bF$buf87),
    .D(_1173_[24]),
    .Q(\datapath_1.regfile_1.regOut[19] [24]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _9269_ (
    .CLK(clk_bF$buf86),
    .D(_1173_[25]),
    .Q(\datapath_1.regfile_1.regOut[19] [25]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _9270_ (
    .CLK(clk_bF$buf85),
    .D(_1173_[26]),
    .Q(\datapath_1.regfile_1.regOut[19] [26]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _9271_ (
    .CLK(clk_bF$buf84),
    .D(_1173_[27]),
    .Q(\datapath_1.regfile_1.regOut[19] [27]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _9272_ (
    .CLK(clk_bF$buf83),
    .D(_1173_[28]),
    .Q(\datapath_1.regfile_1.regOut[19] [28]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _9273_ (
    .CLK(clk_bF$buf82),
    .D(_1173_[29]),
    .Q(\datapath_1.regfile_1.regOut[19] [29]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _9274_ (
    .CLK(clk_bF$buf81),
    .D(_1173_[30]),
    .Q(\datapath_1.regfile_1.regOut[19] [30]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _9275_ (
    .CLK(clk_bF$buf80),
    .D(_1173_[31]),
    .Q(\datapath_1.regfile_1.regOut[19] [31]),
    .R(rst_bF$buf80),
    .S(vdd)
);

INVX1 _9276_ (
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_1301_)
);

NAND2X1 _9277_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .Y(_1302_)
);

OAI21X1 _9278_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1301_),
    .C(_1302_),
    .Y(_1238_[0])
);

INVX1 _9279_ (
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_1239_)
);

NAND2X1 _9280_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1240_)
);

OAI21X1 _9281_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1239_),
    .C(_1240_),
    .Y(_1238_[1])
);

INVX1 _9282_ (
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_1241_)
);

NAND2X1 _9283_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1242_)
);

OAI21X1 _9284_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1241_),
    .C(_1242_),
    .Y(_1238_[2])
);

INVX1 _9285_ (
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_1243_)
);

NAND2X1 _9286_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1244_)
);

OAI21X1 _9287_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1243_),
    .C(_1244_),
    .Y(_1238_[3])
);

INVX1 _9288_ (
    .A(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_1245_)
);

NAND2X1 _9289_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1246_)
);

OAI21X1 _9290_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1245_),
    .C(_1246_),
    .Y(_1238_[4])
);

INVX1 _9291_ (
    .A(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_1247_)
);

NAND2X1 _9292_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1248_)
);

OAI21X1 _9293_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1247_),
    .C(_1248_),
    .Y(_1238_[5])
);

INVX1 _9294_ (
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_1249_)
);

NAND2X1 _9295_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1250_)
);

OAI21X1 _9296_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1249_),
    .C(_1250_),
    .Y(_1238_[6])
);

INVX1 _9297_ (
    .A(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_1251_)
);

NAND2X1 _9298_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1252_)
);

OAI21X1 _9299_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1251_),
    .C(_1252_),
    .Y(_1238_[7])
);

INVX1 _9300_ (
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_1253_)
);

NAND2X1 _9301_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1254_)
);

OAI21X1 _9302_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1253_),
    .C(_1254_),
    .Y(_1238_[8])
);

INVX1 _9303_ (
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_1255_)
);

NAND2X1 _9304_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1256_)
);

OAI21X1 _9305_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1255_),
    .C(_1256_),
    .Y(_1238_[9])
);

INVX1 _9306_ (
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_1257_)
);

NAND2X1 _9307_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1258_)
);

OAI21X1 _9308_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1257_),
    .C(_1258_),
    .Y(_1238_[10])
);

INVX1 _9309_ (
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_1259_)
);

NAND2X1 _9310_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1260_)
);

OAI21X1 _9311_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1259_),
    .C(_1260_),
    .Y(_1238_[11])
);

INVX1 _9312_ (
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_1261_)
);

NAND2X1 _9313_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1262_)
);

OAI21X1 _9314_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1261_),
    .C(_1262_),
    .Y(_1238_[12])
);

INVX1 _9315_ (
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_1263_)
);

NAND2X1 _9316_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1264_)
);

OAI21X1 _9317_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1263_),
    .C(_1264_),
    .Y(_1238_[13])
);

INVX1 _9318_ (
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_1265_)
);

NAND2X1 _9319_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1266_)
);

OAI21X1 _9320_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1265_),
    .C(_1266_),
    .Y(_1238_[14])
);

INVX1 _9321_ (
    .A(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_1267_)
);

NAND2X1 _9322_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1268_)
);

OAI21X1 _9323_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1267_),
    .C(_1268_),
    .Y(_1238_[15])
);

INVX1 _9324_ (
    .A(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_1269_)
);

NAND2X1 _9325_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1270_)
);

OAI21X1 _9326_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1269_),
    .C(_1270_),
    .Y(_1238_[16])
);

INVX1 _9327_ (
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_1271_)
);

NAND2X1 _9328_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1272_)
);

OAI21X1 _9329_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1271_),
    .C(_1272_),
    .Y(_1238_[17])
);

INVX1 _9330_ (
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_1273_)
);

NAND2X1 _9331_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1274_)
);

OAI21X1 _9332_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1273_),
    .C(_1274_),
    .Y(_1238_[18])
);

INVX1 _9333_ (
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_1275_)
);

NAND2X1 _9334_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1276_)
);

OAI21X1 _9335_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1275_),
    .C(_1276_),
    .Y(_1238_[19])
);

INVX1 _9336_ (
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_1277_)
);

NAND2X1 _9337_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1278_)
);

OAI21X1 _9338_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1277_),
    .C(_1278_),
    .Y(_1238_[20])
);

INVX1 _9339_ (
    .A(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_1279_)
);

NAND2X1 _9340_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1280_)
);

OAI21X1 _9341_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1279_),
    .C(_1280_),
    .Y(_1238_[21])
);

INVX1 _9342_ (
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_1281_)
);

NAND2X1 _9343_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1282_)
);

OAI21X1 _9344_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1281_),
    .C(_1282_),
    .Y(_1238_[22])
);

INVX1 _9345_ (
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_1283_)
);

NAND2X1 _9346_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1284_)
);

OAI21X1 _9347_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1283_),
    .C(_1284_),
    .Y(_1238_[23])
);

INVX1 _9348_ (
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_1285_)
);

NAND2X1 _9349_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1286_)
);

OAI21X1 _9350_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1285_),
    .C(_1286_),
    .Y(_1238_[24])
);

INVX1 _9351_ (
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_1287_)
);

NAND2X1 _9352_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1288_)
);

OAI21X1 _9353_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1287_),
    .C(_1288_),
    .Y(_1238_[25])
);

INVX1 _9354_ (
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_1289_)
);

NAND2X1 _9355_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1290_)
);

OAI21X1 _9356_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1289_),
    .C(_1290_),
    .Y(_1238_[26])
);

INVX1 _9357_ (
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_1291_)
);

NAND2X1 _9358_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1292_)
);

OAI21X1 _9359_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1291_),
    .C(_1292_),
    .Y(_1238_[27])
);

INVX1 _9360_ (
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_1293_)
);

NAND2X1 _9361_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1294_)
);

OAI21X1 _9362_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(_1293_),
    .C(_1294_),
    .Y(_1238_[28])
);

INVX1 _9363_ (
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_1295_)
);

NAND2X1 _9364_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_1296_)
);

OAI21X1 _9365_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(_1295_),
    .C(_1296_),
    .Y(_1238_[29])
);

INVX1 _9366_ (
    .A(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_1297_)
);

NAND2X1 _9367_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1298_)
);

OAI21X1 _9368_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(_1297_),
    .C(_1298_),
    .Y(_1238_[30])
);

INVX1 _9369_ (
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_1299_)
);

NAND2X1 _9370_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_1300_)
);

OAI21X1 _9371_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(_1299_),
    .C(_1300_),
    .Y(_1238_[31])
);

DFFSR _9372_ (
    .CLK(clk_bF$buf79),
    .D(_1238_[0]),
    .Q(\datapath_1.regfile_1.regOut[20] [0]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _9373_ (
    .CLK(clk_bF$buf78),
    .D(_1238_[1]),
    .Q(\datapath_1.regfile_1.regOut[20] [1]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _9374_ (
    .CLK(clk_bF$buf77),
    .D(_1238_[2]),
    .Q(\datapath_1.regfile_1.regOut[20] [2]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _9375_ (
    .CLK(clk_bF$buf76),
    .D(_1238_[3]),
    .Q(\datapath_1.regfile_1.regOut[20] [3]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _9376_ (
    .CLK(clk_bF$buf75),
    .D(_1238_[4]),
    .Q(\datapath_1.regfile_1.regOut[20] [4]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _9377_ (
    .CLK(clk_bF$buf74),
    .D(_1238_[5]),
    .Q(\datapath_1.regfile_1.regOut[20] [5]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _9378_ (
    .CLK(clk_bF$buf73),
    .D(_1238_[6]),
    .Q(\datapath_1.regfile_1.regOut[20] [6]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _9379_ (
    .CLK(clk_bF$buf72),
    .D(_1238_[7]),
    .Q(\datapath_1.regfile_1.regOut[20] [7]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _9380_ (
    .CLK(clk_bF$buf71),
    .D(_1238_[8]),
    .Q(\datapath_1.regfile_1.regOut[20] [8]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _9381_ (
    .CLK(clk_bF$buf70),
    .D(_1238_[9]),
    .Q(\datapath_1.regfile_1.regOut[20] [9]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _9382_ (
    .CLK(clk_bF$buf69),
    .D(_1238_[10]),
    .Q(\datapath_1.regfile_1.regOut[20] [10]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _9383_ (
    .CLK(clk_bF$buf68),
    .D(_1238_[11]),
    .Q(\datapath_1.regfile_1.regOut[20] [11]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _9384_ (
    .CLK(clk_bF$buf67),
    .D(_1238_[12]),
    .Q(\datapath_1.regfile_1.regOut[20] [12]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _9385_ (
    .CLK(clk_bF$buf66),
    .D(_1238_[13]),
    .Q(\datapath_1.regfile_1.regOut[20] [13]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _9386_ (
    .CLK(clk_bF$buf65),
    .D(_1238_[14]),
    .Q(\datapath_1.regfile_1.regOut[20] [14]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _9387_ (
    .CLK(clk_bF$buf64),
    .D(_1238_[15]),
    .Q(\datapath_1.regfile_1.regOut[20] [15]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _9388_ (
    .CLK(clk_bF$buf63),
    .D(_1238_[16]),
    .Q(\datapath_1.regfile_1.regOut[20] [16]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _9389_ (
    .CLK(clk_bF$buf62),
    .D(_1238_[17]),
    .Q(\datapath_1.regfile_1.regOut[20] [17]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _9390_ (
    .CLK(clk_bF$buf61),
    .D(_1238_[18]),
    .Q(\datapath_1.regfile_1.regOut[20] [18]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _9391_ (
    .CLK(clk_bF$buf60),
    .D(_1238_[19]),
    .Q(\datapath_1.regfile_1.regOut[20] [19]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _9392_ (
    .CLK(clk_bF$buf59),
    .D(_1238_[20]),
    .Q(\datapath_1.regfile_1.regOut[20] [20]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _9393_ (
    .CLK(clk_bF$buf58),
    .D(_1238_[21]),
    .Q(\datapath_1.regfile_1.regOut[20] [21]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _9394_ (
    .CLK(clk_bF$buf57),
    .D(_1238_[22]),
    .Q(\datapath_1.regfile_1.regOut[20] [22]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _9395_ (
    .CLK(clk_bF$buf56),
    .D(_1238_[23]),
    .Q(\datapath_1.regfile_1.regOut[20] [23]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _9396_ (
    .CLK(clk_bF$buf55),
    .D(_1238_[24]),
    .Q(\datapath_1.regfile_1.regOut[20] [24]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _9397_ (
    .CLK(clk_bF$buf54),
    .D(_1238_[25]),
    .Q(\datapath_1.regfile_1.regOut[20] [25]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _9398_ (
    .CLK(clk_bF$buf53),
    .D(_1238_[26]),
    .Q(\datapath_1.regfile_1.regOut[20] [26]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _9399_ (
    .CLK(clk_bF$buf52),
    .D(_1238_[27]),
    .Q(\datapath_1.regfile_1.regOut[20] [27]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _9400_ (
    .CLK(clk_bF$buf51),
    .D(_1238_[28]),
    .Q(\datapath_1.regfile_1.regOut[20] [28]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _9401_ (
    .CLK(clk_bF$buf50),
    .D(_1238_[29]),
    .Q(\datapath_1.regfile_1.regOut[20] [29]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _9402_ (
    .CLK(clk_bF$buf49),
    .D(_1238_[30]),
    .Q(\datapath_1.regfile_1.regOut[20] [30]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _9403_ (
    .CLK(clk_bF$buf48),
    .D(_1238_[31]),
    .Q(\datapath_1.regfile_1.regOut[20] [31]),
    .R(rst_bF$buf48),
    .S(vdd)
);

INVX1 _9404_ (
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_1366_)
);

NAND2X1 _9405_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .Y(_1367_)
);

OAI21X1 _9406_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1366_),
    .C(_1367_),
    .Y(_1303_[0])
);

INVX1 _9407_ (
    .A(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_1304_)
);

NAND2X1 _9408_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1305_)
);

OAI21X1 _9409_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1304_),
    .C(_1305_),
    .Y(_1303_[1])
);

INVX1 _9410_ (
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_1306_)
);

NAND2X1 _9411_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1307_)
);

OAI21X1 _9412_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1306_),
    .C(_1307_),
    .Y(_1303_[2])
);

INVX1 _9413_ (
    .A(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_1308_)
);

NAND2X1 _9414_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_1309_)
);

OAI21X1 _9415_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1308_),
    .C(_1309_),
    .Y(_1303_[3])
);

INVX1 _9416_ (
    .A(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_1310_)
);

NAND2X1 _9417_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1311_)
);

OAI21X1 _9418_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1310_),
    .C(_1311_),
    .Y(_1303_[4])
);

INVX1 _9419_ (
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_1312_)
);

NAND2X1 _9420_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1313_)
);

OAI21X1 _9421_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1312_),
    .C(_1313_),
    .Y(_1303_[5])
);

INVX1 _9422_ (
    .A(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_1314_)
);

NAND2X1 _9423_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1315_)
);

OAI21X1 _9424_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1314_),
    .C(_1315_),
    .Y(_1303_[6])
);

INVX1 _9425_ (
    .A(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_1316_)
);

NAND2X1 _9426_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1317_)
);

OAI21X1 _9427_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1316_),
    .C(_1317_),
    .Y(_1303_[7])
);

INVX1 _9428_ (
    .A(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_1318_)
);

NAND2X1 _9429_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1319_)
);

OAI21X1 _9430_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1318_),
    .C(_1319_),
    .Y(_1303_[8])
);

INVX1 _9431_ (
    .A(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_1320_)
);

NAND2X1 _9432_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1321_)
);

OAI21X1 _9433_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1320_),
    .C(_1321_),
    .Y(_1303_[9])
);

INVX1 _9434_ (
    .A(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_1322_)
);

NAND2X1 _9435_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1323_)
);

OAI21X1 _9436_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1322_),
    .C(_1323_),
    .Y(_1303_[10])
);

INVX1 _9437_ (
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_1324_)
);

NAND2X1 _9438_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1325_)
);

OAI21X1 _9439_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1324_),
    .C(_1325_),
    .Y(_1303_[11])
);

INVX1 _9440_ (
    .A(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_1326_)
);

NAND2X1 _9441_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1327_)
);

OAI21X1 _9442_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1326_),
    .C(_1327_),
    .Y(_1303_[12])
);

INVX1 _9443_ (
    .A(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_1328_)
);

NAND2X1 _9444_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1329_)
);

OAI21X1 _9445_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1328_),
    .C(_1329_),
    .Y(_1303_[13])
);

INVX1 _9446_ (
    .A(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_1330_)
);

NAND2X1 _9447_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1331_)
);

OAI21X1 _9448_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1330_),
    .C(_1331_),
    .Y(_1303_[14])
);

INVX1 _9449_ (
    .A(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_1332_)
);

NAND2X1 _9450_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1333_)
);

OAI21X1 _9451_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1332_),
    .C(_1333_),
    .Y(_1303_[15])
);

INVX1 _9452_ (
    .A(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_1334_)
);

NAND2X1 _9453_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1335_)
);

OAI21X1 _9454_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1334_),
    .C(_1335_),
    .Y(_1303_[16])
);

INVX1 _9455_ (
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_1336_)
);

NAND2X1 _9456_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1337_)
);

OAI21X1 _9457_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1336_),
    .C(_1337_),
    .Y(_1303_[17])
);

INVX1 _9458_ (
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_1338_)
);

NAND2X1 _9459_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1339_)
);

OAI21X1 _9460_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1338_),
    .C(_1339_),
    .Y(_1303_[18])
);

INVX1 _9461_ (
    .A(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_1340_)
);

NAND2X1 _9462_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1341_)
);

OAI21X1 _9463_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1340_),
    .C(_1341_),
    .Y(_1303_[19])
);

INVX1 _9464_ (
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_1342_)
);

NAND2X1 _9465_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1343_)
);

OAI21X1 _9466_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1342_),
    .C(_1343_),
    .Y(_1303_[20])
);

INVX1 _9467_ (
    .A(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_1344_)
);

NAND2X1 _9468_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1345_)
);

OAI21X1 _9469_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1344_),
    .C(_1345_),
    .Y(_1303_[21])
);

INVX1 _9470_ (
    .A(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_1346_)
);

NAND2X1 _9471_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1347_)
);

OAI21X1 _9472_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1346_),
    .C(_1347_),
    .Y(_1303_[22])
);

INVX1 _9473_ (
    .A(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_1348_)
);

NAND2X1 _9474_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1349_)
);

OAI21X1 _9475_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1348_),
    .C(_1349_),
    .Y(_1303_[23])
);

INVX1 _9476_ (
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_1350_)
);

NAND2X1 _9477_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1351_)
);

OAI21X1 _9478_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1350_),
    .C(_1351_),
    .Y(_1303_[24])
);

INVX1 _9479_ (
    .A(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_1352_)
);

NAND2X1 _9480_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_1353_)
);

OAI21X1 _9481_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1352_),
    .C(_1353_),
    .Y(_1303_[25])
);

INVX1 _9482_ (
    .A(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_1354_)
);

NAND2X1 _9483_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1355_)
);

OAI21X1 _9484_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1354_),
    .C(_1355_),
    .Y(_1303_[26])
);

INVX1 _9485_ (
    .A(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_1356_)
);

NAND2X1 _9486_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1357_)
);

OAI21X1 _9487_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1356_),
    .C(_1357_),
    .Y(_1303_[27])
);

INVX1 _9488_ (
    .A(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_1358_)
);

NAND2X1 _9489_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1359_)
);

OAI21X1 _9490_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(_1358_),
    .C(_1359_),
    .Y(_1303_[28])
);

INVX1 _9491_ (
    .A(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_1360_)
);

NAND2X1 _9492_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1361_)
);

OAI21X1 _9493_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(_1360_),
    .C(_1361_),
    .Y(_1303_[29])
);

INVX1 _9494_ (
    .A(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_1362_)
);

NAND2X1 _9495_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1363_)
);

OAI21X1 _9496_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(_1362_),
    .C(_1363_),
    .Y(_1303_[30])
);

INVX1 _9497_ (
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_1364_)
);

NAND2X1 _9498_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1365_)
);

OAI21X1 _9499_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(_1364_),
    .C(_1365_),
    .Y(_1303_[31])
);

DFFSR _9500_ (
    .CLK(clk_bF$buf47),
    .D(_1303_[0]),
    .Q(\datapath_1.regfile_1.regOut[21] [0]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _9501_ (
    .CLK(clk_bF$buf46),
    .D(_1303_[1]),
    .Q(\datapath_1.regfile_1.regOut[21] [1]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _9502_ (
    .CLK(clk_bF$buf45),
    .D(_1303_[2]),
    .Q(\datapath_1.regfile_1.regOut[21] [2]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _9503_ (
    .CLK(clk_bF$buf44),
    .D(_1303_[3]),
    .Q(\datapath_1.regfile_1.regOut[21] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _9504_ (
    .CLK(clk_bF$buf43),
    .D(_1303_[4]),
    .Q(\datapath_1.regfile_1.regOut[21] [4]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _9505_ (
    .CLK(clk_bF$buf42),
    .D(_1303_[5]),
    .Q(\datapath_1.regfile_1.regOut[21] [5]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _9506_ (
    .CLK(clk_bF$buf41),
    .D(_1303_[6]),
    .Q(\datapath_1.regfile_1.regOut[21] [6]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _9507_ (
    .CLK(clk_bF$buf40),
    .D(_1303_[7]),
    .Q(\datapath_1.regfile_1.regOut[21] [7]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _9508_ (
    .CLK(clk_bF$buf39),
    .D(_1303_[8]),
    .Q(\datapath_1.regfile_1.regOut[21] [8]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _9509_ (
    .CLK(clk_bF$buf38),
    .D(_1303_[9]),
    .Q(\datapath_1.regfile_1.regOut[21] [9]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _9510_ (
    .CLK(clk_bF$buf37),
    .D(_1303_[10]),
    .Q(\datapath_1.regfile_1.regOut[21] [10]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _9511_ (
    .CLK(clk_bF$buf36),
    .D(_1303_[11]),
    .Q(\datapath_1.regfile_1.regOut[21] [11]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _9512_ (
    .CLK(clk_bF$buf35),
    .D(_1303_[12]),
    .Q(\datapath_1.regfile_1.regOut[21] [12]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _9513_ (
    .CLK(clk_bF$buf34),
    .D(_1303_[13]),
    .Q(\datapath_1.regfile_1.regOut[21] [13]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _9514_ (
    .CLK(clk_bF$buf33),
    .D(_1303_[14]),
    .Q(\datapath_1.regfile_1.regOut[21] [14]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _9515_ (
    .CLK(clk_bF$buf32),
    .D(_1303_[15]),
    .Q(\datapath_1.regfile_1.regOut[21] [15]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _9516_ (
    .CLK(clk_bF$buf31),
    .D(_1303_[16]),
    .Q(\datapath_1.regfile_1.regOut[21] [16]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _9517_ (
    .CLK(clk_bF$buf30),
    .D(_1303_[17]),
    .Q(\datapath_1.regfile_1.regOut[21] [17]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _9518_ (
    .CLK(clk_bF$buf29),
    .D(_1303_[18]),
    .Q(\datapath_1.regfile_1.regOut[21] [18]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _9519_ (
    .CLK(clk_bF$buf28),
    .D(_1303_[19]),
    .Q(\datapath_1.regfile_1.regOut[21] [19]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _9520_ (
    .CLK(clk_bF$buf27),
    .D(_1303_[20]),
    .Q(\datapath_1.regfile_1.regOut[21] [20]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _9521_ (
    .CLK(clk_bF$buf26),
    .D(_1303_[21]),
    .Q(\datapath_1.regfile_1.regOut[21] [21]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _9522_ (
    .CLK(clk_bF$buf25),
    .D(_1303_[22]),
    .Q(\datapath_1.regfile_1.regOut[21] [22]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _9523_ (
    .CLK(clk_bF$buf24),
    .D(_1303_[23]),
    .Q(\datapath_1.regfile_1.regOut[21] [23]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _9524_ (
    .CLK(clk_bF$buf23),
    .D(_1303_[24]),
    .Q(\datapath_1.regfile_1.regOut[21] [24]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _9525_ (
    .CLK(clk_bF$buf22),
    .D(_1303_[25]),
    .Q(\datapath_1.regfile_1.regOut[21] [25]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _9526_ (
    .CLK(clk_bF$buf21),
    .D(_1303_[26]),
    .Q(\datapath_1.regfile_1.regOut[21] [26]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _9527_ (
    .CLK(clk_bF$buf20),
    .D(_1303_[27]),
    .Q(\datapath_1.regfile_1.regOut[21] [27]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _9528_ (
    .CLK(clk_bF$buf19),
    .D(_1303_[28]),
    .Q(\datapath_1.regfile_1.regOut[21] [28]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _9529_ (
    .CLK(clk_bF$buf18),
    .D(_1303_[29]),
    .Q(\datapath_1.regfile_1.regOut[21] [29]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _9530_ (
    .CLK(clk_bF$buf17),
    .D(_1303_[30]),
    .Q(\datapath_1.regfile_1.regOut[21] [30]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _9531_ (
    .CLK(clk_bF$buf16),
    .D(_1303_[31]),
    .Q(\datapath_1.regfile_1.regOut[21] [31]),
    .R(rst_bF$buf16),
    .S(vdd)
);

INVX1 _9532_ (
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_1431_)
);

NAND2X1 _9533_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .Y(_1432_)
);

OAI21X1 _9534_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1431_),
    .C(_1432_),
    .Y(_1368_[0])
);

INVX1 _9535_ (
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_1369_)
);

NAND2X1 _9536_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1370_)
);

OAI21X1 _9537_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1369_),
    .C(_1370_),
    .Y(_1368_[1])
);

INVX1 _9538_ (
    .A(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_1371_)
);

NAND2X1 _9539_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1372_)
);

OAI21X1 _9540_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1371_),
    .C(_1372_),
    .Y(_1368_[2])
);

INVX1 _9541_ (
    .A(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_1373_)
);

NAND2X1 _9542_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1374_)
);

OAI21X1 _9543_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1373_),
    .C(_1374_),
    .Y(_1368_[3])
);

INVX1 _9544_ (
    .A(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_1375_)
);

NAND2X1 _9545_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1376_)
);

OAI21X1 _9546_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1375_),
    .C(_1376_),
    .Y(_1368_[4])
);

INVX1 _9547_ (
    .A(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_1377_)
);

NAND2X1 _9548_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1378_)
);

OAI21X1 _9549_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1377_),
    .C(_1378_),
    .Y(_1368_[5])
);

INVX1 _9550_ (
    .A(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_1379_)
);

NAND2X1 _9551_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1380_)
);

OAI21X1 _9552_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1379_),
    .C(_1380_),
    .Y(_1368_[6])
);

INVX1 _9553_ (
    .A(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_1381_)
);

NAND2X1 _9554_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1382_)
);

OAI21X1 _9555_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1381_),
    .C(_1382_),
    .Y(_1368_[7])
);

INVX1 _9556_ (
    .A(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_1383_)
);

NAND2X1 _9557_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1384_)
);

OAI21X1 _9558_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1383_),
    .C(_1384_),
    .Y(_1368_[8])
);

INVX1 _9559_ (
    .A(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_1385_)
);

NAND2X1 _9560_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1386_)
);

OAI21X1 _9561_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1385_),
    .C(_1386_),
    .Y(_1368_[9])
);

INVX1 _9562_ (
    .A(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_1387_)
);

NAND2X1 _9563_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1388_)
);

OAI21X1 _9564_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1387_),
    .C(_1388_),
    .Y(_1368_[10])
);

INVX1 _9565_ (
    .A(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_1389_)
);

NAND2X1 _9566_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1390_)
);

OAI21X1 _9567_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1389_),
    .C(_1390_),
    .Y(_1368_[11])
);

INVX1 _9568_ (
    .A(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_1391_)
);

NAND2X1 _9569_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1392_)
);

OAI21X1 _9570_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1391_),
    .C(_1392_),
    .Y(_1368_[12])
);

INVX1 _9571_ (
    .A(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_1393_)
);

NAND2X1 _9572_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1394_)
);

OAI21X1 _9573_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1393_),
    .C(_1394_),
    .Y(_1368_[13])
);

INVX1 _9574_ (
    .A(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_1395_)
);

NAND2X1 _9575_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1396_)
);

OAI21X1 _9576_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1395_),
    .C(_1396_),
    .Y(_1368_[14])
);

INVX1 _9577_ (
    .A(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_1397_)
);

NAND2X1 _9578_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1398_)
);

OAI21X1 _9579_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1397_),
    .C(_1398_),
    .Y(_1368_[15])
);

INVX1 _9580_ (
    .A(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_1399_)
);

NAND2X1 _9581_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1400_)
);

OAI21X1 _9582_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1399_),
    .C(_1400_),
    .Y(_1368_[16])
);

INVX1 _9583_ (
    .A(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_1401_)
);

NAND2X1 _9584_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1402_)
);

OAI21X1 _9585_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1401_),
    .C(_1402_),
    .Y(_1368_[17])
);

INVX1 _9586_ (
    .A(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_1403_)
);

NAND2X1 _9587_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1404_)
);

OAI21X1 _9588_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1403_),
    .C(_1404_),
    .Y(_1368_[18])
);

INVX1 _9589_ (
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_1405_)
);

NAND2X1 _9590_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1406_)
);

OAI21X1 _9591_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1405_),
    .C(_1406_),
    .Y(_1368_[19])
);

INVX1 _9592_ (
    .A(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_1407_)
);

NAND2X1 _9593_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1408_)
);

OAI21X1 _9594_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1407_),
    .C(_1408_),
    .Y(_1368_[20])
);

INVX1 _9595_ (
    .A(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_1409_)
);

NAND2X1 _9596_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1410_)
);

OAI21X1 _9597_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1409_),
    .C(_1410_),
    .Y(_1368_[21])
);

INVX1 _9598_ (
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_1411_)
);

NAND2X1 _9599_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1412_)
);

OAI21X1 _9600_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1411_),
    .C(_1412_),
    .Y(_1368_[22])
);

INVX1 _9601_ (
    .A(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_1413_)
);

NAND2X1 _9602_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1414_)
);

OAI21X1 _9603_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1413_),
    .C(_1414_),
    .Y(_1368_[23])
);

INVX1 _9604_ (
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_1415_)
);

NAND2X1 _9605_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1416_)
);

OAI21X1 _9606_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1415_),
    .C(_1416_),
    .Y(_1368_[24])
);

INVX1 _9607_ (
    .A(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_1417_)
);

NAND2X1 _9608_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1418_)
);

OAI21X1 _9609_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1417_),
    .C(_1418_),
    .Y(_1368_[25])
);

INVX1 _9610_ (
    .A(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_1419_)
);

NAND2X1 _9611_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1420_)
);

OAI21X1 _9612_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1419_),
    .C(_1420_),
    .Y(_1368_[26])
);

INVX1 _9613_ (
    .A(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_1421_)
);

NAND2X1 _9614_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1422_)
);

OAI21X1 _9615_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1421_),
    .C(_1422_),
    .Y(_1368_[27])
);

INVX1 _9616_ (
    .A(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_1423_)
);

NAND2X1 _9617_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1424_)
);

OAI21X1 _9618_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(_1423_),
    .C(_1424_),
    .Y(_1368_[28])
);

INVX1 _9619_ (
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_1425_)
);

NAND2X1 _9620_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1426_)
);

OAI21X1 _9621_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(_1425_),
    .C(_1426_),
    .Y(_1368_[29])
);

INVX1 _9622_ (
    .A(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_1427_)
);

NAND2X1 _9623_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1428_)
);

OAI21X1 _9624_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(_1427_),
    .C(_1428_),
    .Y(_1368_[30])
);

INVX1 _9625_ (
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_1429_)
);

NAND2X1 _9626_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1430_)
);

OAI21X1 _9627_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(_1429_),
    .C(_1430_),
    .Y(_1368_[31])
);

DFFSR _9628_ (
    .CLK(clk_bF$buf15),
    .D(_1368_[0]),
    .Q(\datapath_1.regfile_1.regOut[22] [0]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _9629_ (
    .CLK(clk_bF$buf14),
    .D(_1368_[1]),
    .Q(\datapath_1.regfile_1.regOut[22] [1]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _9630_ (
    .CLK(clk_bF$buf13),
    .D(_1368_[2]),
    .Q(\datapath_1.regfile_1.regOut[22] [2]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _9631_ (
    .CLK(clk_bF$buf12),
    .D(_1368_[3]),
    .Q(\datapath_1.regfile_1.regOut[22] [3]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _9632_ (
    .CLK(clk_bF$buf11),
    .D(_1368_[4]),
    .Q(\datapath_1.regfile_1.regOut[22] [4]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _9633_ (
    .CLK(clk_bF$buf10),
    .D(_1368_[5]),
    .Q(\datapath_1.regfile_1.regOut[22] [5]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _9634_ (
    .CLK(clk_bF$buf9),
    .D(_1368_[6]),
    .Q(\datapath_1.regfile_1.regOut[22] [6]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _9635_ (
    .CLK(clk_bF$buf8),
    .D(_1368_[7]),
    .Q(\datapath_1.regfile_1.regOut[22] [7]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _9636_ (
    .CLK(clk_bF$buf7),
    .D(_1368_[8]),
    .Q(\datapath_1.regfile_1.regOut[22] [8]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _9637_ (
    .CLK(clk_bF$buf6),
    .D(_1368_[9]),
    .Q(\datapath_1.regfile_1.regOut[22] [9]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _9638_ (
    .CLK(clk_bF$buf5),
    .D(_1368_[10]),
    .Q(\datapath_1.regfile_1.regOut[22] [10]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _9639_ (
    .CLK(clk_bF$buf4),
    .D(_1368_[11]),
    .Q(\datapath_1.regfile_1.regOut[22] [11]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _9640_ (
    .CLK(clk_bF$buf3),
    .D(_1368_[12]),
    .Q(\datapath_1.regfile_1.regOut[22] [12]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _9641_ (
    .CLK(clk_bF$buf2),
    .D(_1368_[13]),
    .Q(\datapath_1.regfile_1.regOut[22] [13]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _9642_ (
    .CLK(clk_bF$buf1),
    .D(_1368_[14]),
    .Q(\datapath_1.regfile_1.regOut[22] [14]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _9643_ (
    .CLK(clk_bF$buf0),
    .D(_1368_[15]),
    .Q(\datapath_1.regfile_1.regOut[22] [15]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _9644_ (
    .CLK(clk_bF$buf113),
    .D(_1368_[16]),
    .Q(\datapath_1.regfile_1.regOut[22] [16]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _9645_ (
    .CLK(clk_bF$buf112),
    .D(_1368_[17]),
    .Q(\datapath_1.regfile_1.regOut[22] [17]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _9646_ (
    .CLK(clk_bF$buf111),
    .D(_1368_[18]),
    .Q(\datapath_1.regfile_1.regOut[22] [18]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _9647_ (
    .CLK(clk_bF$buf110),
    .D(_1368_[19]),
    .Q(\datapath_1.regfile_1.regOut[22] [19]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _9648_ (
    .CLK(clk_bF$buf109),
    .D(_1368_[20]),
    .Q(\datapath_1.regfile_1.regOut[22] [20]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _9649_ (
    .CLK(clk_bF$buf108),
    .D(_1368_[21]),
    .Q(\datapath_1.regfile_1.regOut[22] [21]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _9650_ (
    .CLK(clk_bF$buf107),
    .D(_1368_[22]),
    .Q(\datapath_1.regfile_1.regOut[22] [22]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _9651_ (
    .CLK(clk_bF$buf106),
    .D(_1368_[23]),
    .Q(\datapath_1.regfile_1.regOut[22] [23]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _9652_ (
    .CLK(clk_bF$buf105),
    .D(_1368_[24]),
    .Q(\datapath_1.regfile_1.regOut[22] [24]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _9653_ (
    .CLK(clk_bF$buf104),
    .D(_1368_[25]),
    .Q(\datapath_1.regfile_1.regOut[22] [25]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _9654_ (
    .CLK(clk_bF$buf103),
    .D(_1368_[26]),
    .Q(\datapath_1.regfile_1.regOut[22] [26]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _9655_ (
    .CLK(clk_bF$buf102),
    .D(_1368_[27]),
    .Q(\datapath_1.regfile_1.regOut[22] [27]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _9656_ (
    .CLK(clk_bF$buf101),
    .D(_1368_[28]),
    .Q(\datapath_1.regfile_1.regOut[22] [28]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _9657_ (
    .CLK(clk_bF$buf100),
    .D(_1368_[29]),
    .Q(\datapath_1.regfile_1.regOut[22] [29]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _9658_ (
    .CLK(clk_bF$buf99),
    .D(_1368_[30]),
    .Q(\datapath_1.regfile_1.regOut[22] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _9659_ (
    .CLK(clk_bF$buf98),
    .D(_1368_[31]),
    .Q(\datapath_1.regfile_1.regOut[22] [31]),
    .R(rst_bF$buf98),
    .S(vdd)
);

INVX1 _9660_ (
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_1496_)
);

NAND2X1 _9661_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .Y(_1497_)
);

OAI21X1 _9662_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1496_),
    .C(_1497_),
    .Y(_1433_[0])
);

INVX1 _9663_ (
    .A(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_1434_)
);

NAND2X1 _9664_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1435_)
);

OAI21X1 _9665_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1434_),
    .C(_1435_),
    .Y(_1433_[1])
);

INVX1 _9666_ (
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_1436_)
);

NAND2X1 _9667_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1437_)
);

OAI21X1 _9668_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1436_),
    .C(_1437_),
    .Y(_1433_[2])
);

INVX1 _9669_ (
    .A(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_1438_)
);

NAND2X1 _9670_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1439_)
);

OAI21X1 _9671_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1438_),
    .C(_1439_),
    .Y(_1433_[3])
);

INVX1 _9672_ (
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_1440_)
);

NAND2X1 _9673_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1441_)
);

OAI21X1 _9674_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1440_),
    .C(_1441_),
    .Y(_1433_[4])
);

INVX1 _9675_ (
    .A(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_1442_)
);

NAND2X1 _9676_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1443_)
);

OAI21X1 _9677_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1442_),
    .C(_1443_),
    .Y(_1433_[5])
);

INVX1 _9678_ (
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_1444_)
);

NAND2X1 _9679_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1445_)
);

OAI21X1 _9680_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1444_),
    .C(_1445_),
    .Y(_1433_[6])
);

INVX1 _9681_ (
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_1446_)
);

NAND2X1 _9682_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1447_)
);

OAI21X1 _9683_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1446_),
    .C(_1447_),
    .Y(_1433_[7])
);

INVX1 _9684_ (
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_1448_)
);

NAND2X1 _9685_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1449_)
);

OAI21X1 _9686_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1448_),
    .C(_1449_),
    .Y(_1433_[8])
);

INVX1 _9687_ (
    .A(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_1450_)
);

NAND2X1 _9688_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1451_)
);

OAI21X1 _9689_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1450_),
    .C(_1451_),
    .Y(_1433_[9])
);

INVX1 _9690_ (
    .A(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_1452_)
);

NAND2X1 _9691_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1453_)
);

OAI21X1 _9692_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1452_),
    .C(_1453_),
    .Y(_1433_[10])
);

INVX1 _9693_ (
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_1454_)
);

NAND2X1 _9694_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1455_)
);

OAI21X1 _9695_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1454_),
    .C(_1455_),
    .Y(_1433_[11])
);

INVX1 _9696_ (
    .A(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_1456_)
);

NAND2X1 _9697_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1457_)
);

OAI21X1 _9698_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1456_),
    .C(_1457_),
    .Y(_1433_[12])
);

INVX1 _9699_ (
    .A(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_1458_)
);

NAND2X1 _9700_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1459_)
);

OAI21X1 _9701_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1458_),
    .C(_1459_),
    .Y(_1433_[13])
);

INVX1 _9702_ (
    .A(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_1460_)
);

NAND2X1 _9703_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1461_)
);

OAI21X1 _9704_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1460_),
    .C(_1461_),
    .Y(_1433_[14])
);

INVX1 _9705_ (
    .A(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_1462_)
);

NAND2X1 _9706_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1463_)
);

OAI21X1 _9707_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1462_),
    .C(_1463_),
    .Y(_1433_[15])
);

INVX1 _9708_ (
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_1464_)
);

NAND2X1 _9709_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1465_)
);

OAI21X1 _9710_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1464_),
    .C(_1465_),
    .Y(_1433_[16])
);

INVX1 _9711_ (
    .A(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_1466_)
);

NAND2X1 _9712_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1467_)
);

OAI21X1 _9713_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1466_),
    .C(_1467_),
    .Y(_1433_[17])
);

INVX1 _9714_ (
    .A(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_1468_)
);

NAND2X1 _9715_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1469_)
);

OAI21X1 _9716_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1468_),
    .C(_1469_),
    .Y(_1433_[18])
);

INVX1 _9717_ (
    .A(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_1470_)
);

NAND2X1 _9718_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1471_)
);

OAI21X1 _9719_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1470_),
    .C(_1471_),
    .Y(_1433_[19])
);

INVX1 _9720_ (
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_1472_)
);

NAND2X1 _9721_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1473_)
);

OAI21X1 _9722_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1472_),
    .C(_1473_),
    .Y(_1433_[20])
);

INVX1 _9723_ (
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_1474_)
);

NAND2X1 _9724_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1475_)
);

OAI21X1 _9725_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1474_),
    .C(_1475_),
    .Y(_1433_[21])
);

INVX1 _9726_ (
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_1476_)
);

NAND2X1 _9727_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_1477_)
);

OAI21X1 _9728_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1476_),
    .C(_1477_),
    .Y(_1433_[22])
);

INVX1 _9729_ (
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_1478_)
);

NAND2X1 _9730_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1479_)
);

OAI21X1 _9731_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1478_),
    .C(_1479_),
    .Y(_1433_[23])
);

INVX1 _9732_ (
    .A(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_1480_)
);

NAND2X1 _9733_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1481_)
);

OAI21X1 _9734_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1480_),
    .C(_1481_),
    .Y(_1433_[24])
);

INVX1 _9735_ (
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_1482_)
);

NAND2X1 _9736_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1483_)
);

OAI21X1 _9737_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1482_),
    .C(_1483_),
    .Y(_1433_[25])
);

INVX1 _9738_ (
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .Y(_1484_)
);

NAND2X1 _9739_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1485_)
);

OAI21X1 _9740_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1484_),
    .C(_1485_),
    .Y(_1433_[26])
);

INVX1 _9741_ (
    .A(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_1486_)
);

NAND2X1 _9742_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1487_)
);

OAI21X1 _9743_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1486_),
    .C(_1487_),
    .Y(_1433_[27])
);

INVX1 _9744_ (
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_1488_)
);

NAND2X1 _9745_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1489_)
);

OAI21X1 _9746_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(_1488_),
    .C(_1489_),
    .Y(_1433_[28])
);

INVX1 _9747_ (
    .A(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_1490_)
);

NAND2X1 _9748_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1491_)
);

OAI21X1 _9749_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(_1490_),
    .C(_1491_),
    .Y(_1433_[29])
);

INVX1 _9750_ (
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_1492_)
);

NAND2X1 _9751_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1493_)
);

OAI21X1 _9752_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(_1492_),
    .C(_1493_),
    .Y(_1433_[30])
);

INVX1 _9753_ (
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_1494_)
);

NAND2X1 _9754_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1495_)
);

OAI21X1 _9755_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(_1494_),
    .C(_1495_),
    .Y(_1433_[31])
);

DFFSR _9756_ (
    .CLK(clk_bF$buf97),
    .D(_1433_[0]),
    .Q(\datapath_1.regfile_1.regOut[23] [0]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _9757_ (
    .CLK(clk_bF$buf96),
    .D(_1433_[1]),
    .Q(\datapath_1.regfile_1.regOut[23] [1]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _9758_ (
    .CLK(clk_bF$buf95),
    .D(_1433_[2]),
    .Q(\datapath_1.regfile_1.regOut[23] [2]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _9759_ (
    .CLK(clk_bF$buf94),
    .D(_1433_[3]),
    .Q(\datapath_1.regfile_1.regOut[23] [3]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _9760_ (
    .CLK(clk_bF$buf93),
    .D(_1433_[4]),
    .Q(\datapath_1.regfile_1.regOut[23] [4]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _9761_ (
    .CLK(clk_bF$buf92),
    .D(_1433_[5]),
    .Q(\datapath_1.regfile_1.regOut[23] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _9762_ (
    .CLK(clk_bF$buf91),
    .D(_1433_[6]),
    .Q(\datapath_1.regfile_1.regOut[23] [6]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _9763_ (
    .CLK(clk_bF$buf90),
    .D(_1433_[7]),
    .Q(\datapath_1.regfile_1.regOut[23] [7]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _9764_ (
    .CLK(clk_bF$buf89),
    .D(_1433_[8]),
    .Q(\datapath_1.regfile_1.regOut[23] [8]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _9765_ (
    .CLK(clk_bF$buf88),
    .D(_1433_[9]),
    .Q(\datapath_1.regfile_1.regOut[23] [9]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _9766_ (
    .CLK(clk_bF$buf87),
    .D(_1433_[10]),
    .Q(\datapath_1.regfile_1.regOut[23] [10]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _9767_ (
    .CLK(clk_bF$buf86),
    .D(_1433_[11]),
    .Q(\datapath_1.regfile_1.regOut[23] [11]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _9768_ (
    .CLK(clk_bF$buf85),
    .D(_1433_[12]),
    .Q(\datapath_1.regfile_1.regOut[23] [12]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _9769_ (
    .CLK(clk_bF$buf84),
    .D(_1433_[13]),
    .Q(\datapath_1.regfile_1.regOut[23] [13]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _9770_ (
    .CLK(clk_bF$buf83),
    .D(_1433_[14]),
    .Q(\datapath_1.regfile_1.regOut[23] [14]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _9771_ (
    .CLK(clk_bF$buf82),
    .D(_1433_[15]),
    .Q(\datapath_1.regfile_1.regOut[23] [15]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _9772_ (
    .CLK(clk_bF$buf81),
    .D(_1433_[16]),
    .Q(\datapath_1.regfile_1.regOut[23] [16]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _9773_ (
    .CLK(clk_bF$buf80),
    .D(_1433_[17]),
    .Q(\datapath_1.regfile_1.regOut[23] [17]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _9774_ (
    .CLK(clk_bF$buf79),
    .D(_1433_[18]),
    .Q(\datapath_1.regfile_1.regOut[23] [18]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _9775_ (
    .CLK(clk_bF$buf78),
    .D(_1433_[19]),
    .Q(\datapath_1.regfile_1.regOut[23] [19]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _9776_ (
    .CLK(clk_bF$buf77),
    .D(_1433_[20]),
    .Q(\datapath_1.regfile_1.regOut[23] [20]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _9777_ (
    .CLK(clk_bF$buf76),
    .D(_1433_[21]),
    .Q(\datapath_1.regfile_1.regOut[23] [21]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _9778_ (
    .CLK(clk_bF$buf75),
    .D(_1433_[22]),
    .Q(\datapath_1.regfile_1.regOut[23] [22]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _9779_ (
    .CLK(clk_bF$buf74),
    .D(_1433_[23]),
    .Q(\datapath_1.regfile_1.regOut[23] [23]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _9780_ (
    .CLK(clk_bF$buf73),
    .D(_1433_[24]),
    .Q(\datapath_1.regfile_1.regOut[23] [24]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _9781_ (
    .CLK(clk_bF$buf72),
    .D(_1433_[25]),
    .Q(\datapath_1.regfile_1.regOut[23] [25]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _9782_ (
    .CLK(clk_bF$buf71),
    .D(_1433_[26]),
    .Q(\datapath_1.regfile_1.regOut[23] [26]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _9783_ (
    .CLK(clk_bF$buf70),
    .D(_1433_[27]),
    .Q(\datapath_1.regfile_1.regOut[23] [27]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _9784_ (
    .CLK(clk_bF$buf69),
    .D(_1433_[28]),
    .Q(\datapath_1.regfile_1.regOut[23] [28]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _9785_ (
    .CLK(clk_bF$buf68),
    .D(_1433_[29]),
    .Q(\datapath_1.regfile_1.regOut[23] [29]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _9786_ (
    .CLK(clk_bF$buf67),
    .D(_1433_[30]),
    .Q(\datapath_1.regfile_1.regOut[23] [30]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _9787_ (
    .CLK(clk_bF$buf66),
    .D(_1433_[31]),
    .Q(\datapath_1.regfile_1.regOut[23] [31]),
    .R(rst_bF$buf66),
    .S(vdd)
);

INVX1 _9788_ (
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_1561_)
);

NAND2X1 _9789_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .Y(_1562_)
);

OAI21X1 _9790_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1561_),
    .C(_1562_),
    .Y(_1498_[0])
);

INVX1 _9791_ (
    .A(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_1499_)
);

NAND2X1 _9792_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1500_)
);

OAI21X1 _9793_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1499_),
    .C(_1500_),
    .Y(_1498_[1])
);

INVX1 _9794_ (
    .A(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_1501_)
);

NAND2X1 _9795_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1502_)
);

OAI21X1 _9796_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1501_),
    .C(_1502_),
    .Y(_1498_[2])
);

INVX1 _9797_ (
    .A(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_1503_)
);

NAND2X1 _9798_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1504_)
);

OAI21X1 _9799_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1503_),
    .C(_1504_),
    .Y(_1498_[3])
);

INVX1 _9800_ (
    .A(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_1505_)
);

NAND2X1 _9801_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1506_)
);

OAI21X1 _9802_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1505_),
    .C(_1506_),
    .Y(_1498_[4])
);

INVX1 _9803_ (
    .A(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_1507_)
);

NAND2X1 _9804_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1508_)
);

OAI21X1 _9805_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1507_),
    .C(_1508_),
    .Y(_1498_[5])
);

INVX1 _9806_ (
    .A(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_1509_)
);

NAND2X1 _9807_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1510_)
);

OAI21X1 _9808_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1509_),
    .C(_1510_),
    .Y(_1498_[6])
);

INVX1 _9809_ (
    .A(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_1511_)
);

NAND2X1 _9810_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1512_)
);

OAI21X1 _9811_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1511_),
    .C(_1512_),
    .Y(_1498_[7])
);

INVX1 _9812_ (
    .A(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_1513_)
);

NAND2X1 _9813_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1514_)
);

OAI21X1 _9814_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1513_),
    .C(_1514_),
    .Y(_1498_[8])
);

INVX1 _9815_ (
    .A(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_1515_)
);

NAND2X1 _9816_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1516_)
);

OAI21X1 _9817_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1515_),
    .C(_1516_),
    .Y(_1498_[9])
);

INVX1 _9818_ (
    .A(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_1517_)
);

NAND2X1 _9819_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1518_)
);

OAI21X1 _9820_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1517_),
    .C(_1518_),
    .Y(_1498_[10])
);

INVX1 _9821_ (
    .A(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_1519_)
);

NAND2X1 _9822_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1520_)
);

OAI21X1 _9823_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1519_),
    .C(_1520_),
    .Y(_1498_[11])
);

INVX1 _9824_ (
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_1521_)
);

NAND2X1 _9825_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1522_)
);

OAI21X1 _9826_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1521_),
    .C(_1522_),
    .Y(_1498_[12])
);

INVX1 _9827_ (
    .A(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_1523_)
);

NAND2X1 _9828_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1524_)
);

OAI21X1 _9829_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1523_),
    .C(_1524_),
    .Y(_1498_[13])
);

INVX1 _9830_ (
    .A(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_1525_)
);

NAND2X1 _9831_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1526_)
);

OAI21X1 _9832_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1525_),
    .C(_1526_),
    .Y(_1498_[14])
);

INVX1 _9833_ (
    .A(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_1527_)
);

NAND2X1 _9834_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1528_)
);

OAI21X1 _9835_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1527_),
    .C(_1528_),
    .Y(_1498_[15])
);

INVX1 _9836_ (
    .A(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_1529_)
);

NAND2X1 _9837_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1530_)
);

OAI21X1 _9838_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1529_),
    .C(_1530_),
    .Y(_1498_[16])
);

INVX1 _9839_ (
    .A(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_1531_)
);

NAND2X1 _9840_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1532_)
);

OAI21X1 _9841_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1531_),
    .C(_1532_),
    .Y(_1498_[17])
);

INVX1 _9842_ (
    .A(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_1533_)
);

NAND2X1 _9843_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1534_)
);

OAI21X1 _9844_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1533_),
    .C(_1534_),
    .Y(_1498_[18])
);

INVX1 _9845_ (
    .A(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_1535_)
);

NAND2X1 _9846_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1536_)
);

OAI21X1 _9847_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1535_),
    .C(_1536_),
    .Y(_1498_[19])
);

INVX1 _9848_ (
    .A(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_1537_)
);

NAND2X1 _9849_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1538_)
);

OAI21X1 _9850_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1537_),
    .C(_1538_),
    .Y(_1498_[20])
);

INVX1 _9851_ (
    .A(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_1539_)
);

NAND2X1 _9852_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1540_)
);

OAI21X1 _9853_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1539_),
    .C(_1540_),
    .Y(_1498_[21])
);

INVX1 _9854_ (
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_1541_)
);

NAND2X1 _9855_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1542_)
);

OAI21X1 _9856_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1541_),
    .C(_1542_),
    .Y(_1498_[22])
);

INVX1 _9857_ (
    .A(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_1543_)
);

NAND2X1 _9858_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1544_)
);

OAI21X1 _9859_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1543_),
    .C(_1544_),
    .Y(_1498_[23])
);

INVX1 _9860_ (
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .Y(_1545_)
);

NAND2X1 _9861_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1546_)
);

OAI21X1 _9862_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1545_),
    .C(_1546_),
    .Y(_1498_[24])
);

INVX1 _9863_ (
    .A(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_1547_)
);

NAND2X1 _9864_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1548_)
);

OAI21X1 _9865_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1547_),
    .C(_1548_),
    .Y(_1498_[25])
);

INVX1 _9866_ (
    .A(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_1549_)
);

NAND2X1 _9867_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1550_)
);

OAI21X1 _9868_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1549_),
    .C(_1550_),
    .Y(_1498_[26])
);

INVX1 _9869_ (
    .A(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_1551_)
);

NAND2X1 _9870_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1552_)
);

OAI21X1 _9871_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1551_),
    .C(_1552_),
    .Y(_1498_[27])
);

INVX1 _9872_ (
    .A(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_1553_)
);

NAND2X1 _9873_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1554_)
);

OAI21X1 _9874_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(_1553_),
    .C(_1554_),
    .Y(_1498_[28])
);

INVX1 _9875_ (
    .A(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_1555_)
);

NAND2X1 _9876_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1556_)
);

OAI21X1 _9877_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(_1555_),
    .C(_1556_),
    .Y(_1498_[29])
);

INVX1 _9878_ (
    .A(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_1557_)
);

NAND2X1 _9879_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1558_)
);

OAI21X1 _9880_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(_1557_),
    .C(_1558_),
    .Y(_1498_[30])
);

INVX1 _9881_ (
    .A(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_1559_)
);

NAND2X1 _9882_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1560_)
);

OAI21X1 _9883_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(_1559_),
    .C(_1560_),
    .Y(_1498_[31])
);

DFFSR _9884_ (
    .CLK(clk_bF$buf65),
    .D(_1498_[0]),
    .Q(\datapath_1.regfile_1.regOut[24] [0]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _9885_ (
    .CLK(clk_bF$buf64),
    .D(_1498_[1]),
    .Q(\datapath_1.regfile_1.regOut[24] [1]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _9886_ (
    .CLK(clk_bF$buf63),
    .D(_1498_[2]),
    .Q(\datapath_1.regfile_1.regOut[24] [2]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _9887_ (
    .CLK(clk_bF$buf62),
    .D(_1498_[3]),
    .Q(\datapath_1.regfile_1.regOut[24] [3]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _9888_ (
    .CLK(clk_bF$buf61),
    .D(_1498_[4]),
    .Q(\datapath_1.regfile_1.regOut[24] [4]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _9889_ (
    .CLK(clk_bF$buf60),
    .D(_1498_[5]),
    .Q(\datapath_1.regfile_1.regOut[24] [5]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _9890_ (
    .CLK(clk_bF$buf59),
    .D(_1498_[6]),
    .Q(\datapath_1.regfile_1.regOut[24] [6]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _9891_ (
    .CLK(clk_bF$buf58),
    .D(_1498_[7]),
    .Q(\datapath_1.regfile_1.regOut[24] [7]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _9892_ (
    .CLK(clk_bF$buf57),
    .D(_1498_[8]),
    .Q(\datapath_1.regfile_1.regOut[24] [8]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _9893_ (
    .CLK(clk_bF$buf56),
    .D(_1498_[9]),
    .Q(\datapath_1.regfile_1.regOut[24] [9]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _9894_ (
    .CLK(clk_bF$buf55),
    .D(_1498_[10]),
    .Q(\datapath_1.regfile_1.regOut[24] [10]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _9895_ (
    .CLK(clk_bF$buf54),
    .D(_1498_[11]),
    .Q(\datapath_1.regfile_1.regOut[24] [11]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _9896_ (
    .CLK(clk_bF$buf53),
    .D(_1498_[12]),
    .Q(\datapath_1.regfile_1.regOut[24] [12]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _9897_ (
    .CLK(clk_bF$buf52),
    .D(_1498_[13]),
    .Q(\datapath_1.regfile_1.regOut[24] [13]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _9898_ (
    .CLK(clk_bF$buf51),
    .D(_1498_[14]),
    .Q(\datapath_1.regfile_1.regOut[24] [14]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _9899_ (
    .CLK(clk_bF$buf50),
    .D(_1498_[15]),
    .Q(\datapath_1.regfile_1.regOut[24] [15]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _9900_ (
    .CLK(clk_bF$buf49),
    .D(_1498_[16]),
    .Q(\datapath_1.regfile_1.regOut[24] [16]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _9901_ (
    .CLK(clk_bF$buf48),
    .D(_1498_[17]),
    .Q(\datapath_1.regfile_1.regOut[24] [17]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _9902_ (
    .CLK(clk_bF$buf47),
    .D(_1498_[18]),
    .Q(\datapath_1.regfile_1.regOut[24] [18]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _9903_ (
    .CLK(clk_bF$buf46),
    .D(_1498_[19]),
    .Q(\datapath_1.regfile_1.regOut[24] [19]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _9904_ (
    .CLK(clk_bF$buf45),
    .D(_1498_[20]),
    .Q(\datapath_1.regfile_1.regOut[24] [20]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _9905_ (
    .CLK(clk_bF$buf44),
    .D(_1498_[21]),
    .Q(\datapath_1.regfile_1.regOut[24] [21]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _9906_ (
    .CLK(clk_bF$buf43),
    .D(_1498_[22]),
    .Q(\datapath_1.regfile_1.regOut[24] [22]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _9907_ (
    .CLK(clk_bF$buf42),
    .D(_1498_[23]),
    .Q(\datapath_1.regfile_1.regOut[24] [23]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _9908_ (
    .CLK(clk_bF$buf41),
    .D(_1498_[24]),
    .Q(\datapath_1.regfile_1.regOut[24] [24]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _9909_ (
    .CLK(clk_bF$buf40),
    .D(_1498_[25]),
    .Q(\datapath_1.regfile_1.regOut[24] [25]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _9910_ (
    .CLK(clk_bF$buf39),
    .D(_1498_[26]),
    .Q(\datapath_1.regfile_1.regOut[24] [26]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _9911_ (
    .CLK(clk_bF$buf38),
    .D(_1498_[27]),
    .Q(\datapath_1.regfile_1.regOut[24] [27]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _9912_ (
    .CLK(clk_bF$buf37),
    .D(_1498_[28]),
    .Q(\datapath_1.regfile_1.regOut[24] [28]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _9913_ (
    .CLK(clk_bF$buf36),
    .D(_1498_[29]),
    .Q(\datapath_1.regfile_1.regOut[24] [29]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _9914_ (
    .CLK(clk_bF$buf35),
    .D(_1498_[30]),
    .Q(\datapath_1.regfile_1.regOut[24] [30]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _9915_ (
    .CLK(clk_bF$buf34),
    .D(_1498_[31]),
    .Q(\datapath_1.regfile_1.regOut[24] [31]),
    .R(rst_bF$buf34),
    .S(vdd)
);

INVX1 _9916_ (
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_1626_)
);

NAND2X1 _9917_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .Y(_1627_)
);

OAI21X1 _9918_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1626_),
    .C(_1627_),
    .Y(_1563_[0])
);

INVX1 _9919_ (
    .A(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_1564_)
);

NAND2X1 _9920_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1565_)
);

OAI21X1 _9921_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1564_),
    .C(_1565_),
    .Y(_1563_[1])
);

INVX1 _9922_ (
    .A(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_1566_)
);

NAND2X1 _9923_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1567_)
);

OAI21X1 _9924_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1566_),
    .C(_1567_),
    .Y(_1563_[2])
);

INVX1 _9925_ (
    .A(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_1568_)
);

NAND2X1 _9926_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1569_)
);

OAI21X1 _9927_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1568_),
    .C(_1569_),
    .Y(_1563_[3])
);

INVX1 _9928_ (
    .A(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_1570_)
);

NAND2X1 _9929_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1571_)
);

OAI21X1 _9930_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1570_),
    .C(_1571_),
    .Y(_1563_[4])
);

INVX1 _9931_ (
    .A(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_1572_)
);

NAND2X1 _9932_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1573_)
);

OAI21X1 _9933_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1572_),
    .C(_1573_),
    .Y(_1563_[5])
);

INVX1 _9934_ (
    .A(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_1574_)
);

NAND2X1 _9935_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1575_)
);

OAI21X1 _9936_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1574_),
    .C(_1575_),
    .Y(_1563_[6])
);

INVX1 _9937_ (
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_1576_)
);

NAND2X1 _9938_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1577_)
);

OAI21X1 _9939_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1576_),
    .C(_1577_),
    .Y(_1563_[7])
);

INVX1 _9940_ (
    .A(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_1578_)
);

NAND2X1 _9941_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1579_)
);

OAI21X1 _9942_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1578_),
    .C(_1579_),
    .Y(_1563_[8])
);

INVX1 _9943_ (
    .A(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_1580_)
);

NAND2X1 _9944_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1581_)
);

OAI21X1 _9945_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1580_),
    .C(_1581_),
    .Y(_1563_[9])
);

INVX1 _9946_ (
    .A(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_1582_)
);

NAND2X1 _9947_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1583_)
);

OAI21X1 _9948_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1582_),
    .C(_1583_),
    .Y(_1563_[10])
);

INVX1 _9949_ (
    .A(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_1584_)
);

NAND2X1 _9950_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1585_)
);

OAI21X1 _9951_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1584_),
    .C(_1585_),
    .Y(_1563_[11])
);

INVX1 _9952_ (
    .A(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_1586_)
);

NAND2X1 _9953_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1587_)
);

OAI21X1 _9954_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1586_),
    .C(_1587_),
    .Y(_1563_[12])
);

INVX1 _9955_ (
    .A(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_1588_)
);

NAND2X1 _9956_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1589_)
);

OAI21X1 _9957_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1588_),
    .C(_1589_),
    .Y(_1563_[13])
);

INVX1 _9958_ (
    .A(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_1590_)
);

NAND2X1 _9959_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1591_)
);

OAI21X1 _9960_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1590_),
    .C(_1591_),
    .Y(_1563_[14])
);

INVX1 _9961_ (
    .A(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_1592_)
);

NAND2X1 _9962_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1593_)
);

OAI21X1 _9963_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1592_),
    .C(_1593_),
    .Y(_1563_[15])
);

INVX1 _9964_ (
    .A(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_1594_)
);

NAND2X1 _9965_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1595_)
);

OAI21X1 _9966_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1594_),
    .C(_1595_),
    .Y(_1563_[16])
);

INVX1 _9967_ (
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_1596_)
);

NAND2X1 _9968_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1597_)
);

OAI21X1 _9969_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1596_),
    .C(_1597_),
    .Y(_1563_[17])
);

INVX1 _9970_ (
    .A(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_1598_)
);

NAND2X1 _9971_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1599_)
);

OAI21X1 _9972_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1598_),
    .C(_1599_),
    .Y(_1563_[18])
);

INVX1 _9973_ (
    .A(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_1600_)
);

NAND2X1 _9974_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1601_)
);

OAI21X1 _9975_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1600_),
    .C(_1601_),
    .Y(_1563_[19])
);

INVX1 _9976_ (
    .A(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_1602_)
);

NAND2X1 _9977_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1603_)
);

OAI21X1 _9978_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1602_),
    .C(_1603_),
    .Y(_1563_[20])
);

INVX1 _9979_ (
    .A(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_1604_)
);

NAND2X1 _9980_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1605_)
);

OAI21X1 _9981_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1604_),
    .C(_1605_),
    .Y(_1563_[21])
);

INVX1 _9982_ (
    .A(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_1606_)
);

NAND2X1 _9983_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1607_)
);

OAI21X1 _9984_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1606_),
    .C(_1607_),
    .Y(_1563_[22])
);

INVX1 _9985_ (
    .A(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_1608_)
);

NAND2X1 _9986_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1609_)
);

OAI21X1 _9987_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1608_),
    .C(_1609_),
    .Y(_1563_[23])
);

INVX1 _9988_ (
    .A(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_1610_)
);

NAND2X1 _9989_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1611_)
);

OAI21X1 _9990_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(_1610_),
    .C(_1611_),
    .Y(_1563_[24])
);

INVX1 _9991_ (
    .A(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_1612_)
);

NAND2X1 _9992_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1613_)
);

OAI21X1 _9993_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(_1612_),
    .C(_1613_),
    .Y(_1563_[25])
);

INVX1 _9994_ (
    .A(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_1614_)
);

NAND2X1 _9995_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1615_)
);

OAI21X1 _9996_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(_1614_),
    .C(_1615_),
    .Y(_1563_[26])
);

INVX1 _9997_ (
    .A(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_1616_)
);

NAND2X1 _9998_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1617_)
);

OAI21X1 _9999_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(_1616_),
    .C(_1617_),
    .Y(_1563_[27])
);

endmodule
