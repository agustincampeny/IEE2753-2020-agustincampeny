/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module mips(
    output MemRead,
    output MemWrite,
    input clk,
    output [31:0] memoryAddress,
    input [31:0] memoryOutData,
    output [31:0] memoryWriteData,
    input rst
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf2  ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire [31:0] _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire IRWrite_bF$buf0 ;
wire _1486_ ;
wire IRWrite_bF$buf1 ;
wire _1066_ ;
wire IRWrite_bF$buf2 ;
wire IRWrite_bF$buf3 ;
wire IRWrite_bF$buf4 ;
wire IRWrite_bF$buf5 ;
wire IRWrite_bF$buf6 ;
wire IRWrite_bF$buf7 ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _2712_ ;
wire _5515__bF$buf0 ;
wire _5515__bF$buf1 ;
wire _5515__bF$buf2 ;
wire _5515__bF$buf3 ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf1  ;
wire \datapath_1.mux_wd3.dout_11_bF$buf4  ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf0  ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf4  ;
wire _57_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf0  ;
wire _6504_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _3884__bF$buf0 ;
wire _3884__bF$buf1 ;
wire _3884__bF$buf2 ;
wire _3884__bF$buf3 ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf4  ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf2  ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6542_ ;
wire _6122_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf3  ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf0  ;
wire _6771_ ;
wire _6351_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf7  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf3  ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf7  ;
wire _6580_ ;
wire _6160_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf5  ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _3947__bF$buf0 ;
wire _3947__bF$buf1 ;
wire _3947__bF$buf2 ;
wire _3947__bF$buf3 ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf3  ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire [31:0] \datapath_1.regfile_1.regOut[13]  ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _5503__bF$buf0 ;
wire _5503__bF$buf1 ;
wire _5503__bF$buf2 ;
wire _5503__bF$buf3 ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire \datapath_1.PCJump_27_bF$buf2  ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _2341__bF$buf0 ;
wire _2341__bF$buf1 ;
wire _2341__bF$buf2 ;
wire _2341__bF$buf3 ;
wire _4643_ ;
wire _4223_ ;
wire [31:0] \datapath_1.regfile_1.regOut[7]  ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf2  ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _5495__bF$buf0 ;
wire _5495__bF$buf1 ;
wire _5495__bF$buf2 ;
wire _5495__bF$buf3 ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf1  ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _3966__bF$buf0 ;
wire _3966__bF$buf1 ;
wire _3966__bF$buf2 ;
wire _3966__bF$buf3 ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf5  ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _5518__bF$buf0 ;
wire _5518__bF$buf1 ;
wire _5518__bF$buf2 ;
wire _5518__bF$buf3 ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf1  ;
wire _54_ ;
wire _6501_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf4  ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf1  ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf0  ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf0  ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire PCWrite ;
wire _4678_ ;
wire _4258_ ;
wire _6824_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf4  ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf2  ;
wire _3282_ ;
wire RegWrite_bF$buf0 ;
wire RegWrite_bF$buf1 ;
wire RegWrite_bF$buf2 ;
wire RegWrite_bF$buf3 ;
wire RegWrite_bF$buf4 ;
wire RegWrite_bF$buf5 ;
wire RegWrite_bF$buf6 ;
wire RegWrite_bF$buf7 ;
wire _4487_ ;
wire _4067_ ;
wire _3891__bF$buf0 ;
wire _3891__bF$buf1 ;
wire _3891__bF$buf2 ;
wire _3891__bF$buf3 ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6442_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf0  ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf3  ;
wire _5713_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _2591_ ;
wire _2171_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf7  ;
wire _3796_ ;
wire _3376_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf3  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire \datapath_1.PCJump_22_bF$buf3  ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf7  ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf3  ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _4411_ ;
wire _3954__bF$buf0 ;
wire _3954__bF$buf1 ;
wire _3954__bF$buf2 ;
wire _3954__bF$buf3 ;
wire _3954__bF$buf4 ;
wire \datapath_1.regfile_1.regEn_8_bF$buf7  ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6574_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf2  ;
wire _5939_ ;
wire _5519_ ;
wire _2344__bF$buf0 ;
wire _2344__bF$buf1 ;
wire _2344__bF$buf2 ;
wire _2344__bF$buf3 ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf2  ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf1  ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf5  ;
wire _1286_ ;
wire _197_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf1  ;
wire _3717_ ;
wire _6189_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf4  ;
wire _3902__bF$buf0 ;
wire _3902__bF$buf1 ;
wire _3902__bF$buf2 ;
wire _3902__bF$buf3 ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _2741_ ;
wire _2321_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf1  ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf4  ;
wire _7_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf0  ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf4  ;
wire _3793_ ;
wire _3373_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf0  ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire Branch ;
wire \datapath_1.PCJump_22_bF$buf0  ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf4  ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6533_ ;
wire _6113_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf3  ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf0  ;
wire _6762_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf4  ;
wire _5613_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf7  ;
wire _6818_ ;
wire [31:0] _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6571_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire rst_bF$buf110 ;
wire rst_bF$buf111 ;
wire rst_bF$buf112 ;
wire rst_bF$buf113 ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire RegDst ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6474_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire clk_bF$buf80 ;
wire clk_bF$buf81 ;
wire clk_bF$buf82 ;
wire clk_bF$buf83 ;
wire clk_bF$buf84 ;
wire clk_bF$buf85 ;
wire [31:0] _3620_ ;
wire clk_bF$buf86 ;
wire _3200_ ;
wire clk_bF$buf87 ;
wire clk_bF$buf88 ;
wire clk_bF$buf89 ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _5783_ ;
wire _5363_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf2  ;
wire _2347__bF$buf0 ;
wire _2347__bF$buf1 ;
wire _2347__bF$buf2 ;
wire _2347__bF$buf3 ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf1  ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf5  ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf1  ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf5  ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _3905__bF$buf0 ;
wire _3905__bF$buf1 ;
wire _3905__bF$buf2 ;
wire _3905__bF$buf3 ;
wire _45_ ;
wire _5532__bF$buf0 ;
wire _5532__bF$buf1 ;
wire _5532__bF$buf2 ;
wire _5532__bF$buf3 ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf1  ;
wire _3790_ ;
wire _3370_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf4  ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf5  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf1  ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire _4193_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf0  ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf1  ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf4  ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6433_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _5704_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire _1853_ ;
wire [31:0] _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6471_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf2  ;
wire [31:0] \datapath_1.regfile_1.regOut[2]  ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6565_ ;
wire _6145_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf2  ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire [31:0] \datapath_1.regfile_1.regOut[25]  ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf2  ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire [31:0] _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _5683_ ;
wire _5263_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf2  ;
wire _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire rst_bF$buf0 ;
wire rst_bF$buf1 ;
wire rst_bF$buf2 ;
wire rst_bF$buf3 ;
wire rst_bF$buf4 ;
wire _5968_ ;
wire rst_bF$buf5 ;
wire _5548_ ;
wire rst_bF$buf6 ;
wire _5128_ ;
wire rst_bF$buf7 ;
wire rst_bF$buf8 ;
wire rst_bF$buf9 ;
wire _42_ ;
wire [31:0] _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf1  ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf2  ;
wire _4628_ ;
wire _4208_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf5  ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _3983__bF$buf0 ;
wire _3983__bF$buf1 ;
wire _3983__bF$buf2 ;
wire _3983__bF$buf3 ;
wire _3983__bF$buf4 ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _5535__bF$buf0 ;
wire _5535__bF$buf1 ;
wire _5535__bF$buf2 ;
wire _5535__bF$buf3 ;
wire _5535__bF$buf4 ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf1  ;
wire _6812_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf4  ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf5  ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf4  ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6430_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire [31:0] _3555_ ;
wire _3135_ ;
wire rst_bF$buf90 ;
wire rst_bF$buf91 ;
wire rst_bF$buf92 ;
wire rst_bF$buf93 ;
wire rst_bF$buf94 ;
wire rst_bF$buf95 ;
wire rst_bF$buf96 ;
wire rst_bF$buf97 ;
wire rst_bF$buf98 ;
wire rst_bF$buf99 ;
wire _5701_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire IorD ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6524_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6562_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf2  ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _3967__bF$buf0 ;
wire _3967__bF$buf1 ;
wire _3967__bF$buf2 ;
wire _3967__bF$buf3 ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf5  ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire [31:0] \datapath_1.regfile_1.regOut[15]  ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf4  ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf2  ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf6  ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire [31:0] \datapath_1.regfile_1.regOut[9]  ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf1  ;
wire _1788_ ;
wire [31:0] _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf2  ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf1  ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf5  ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire rst_bF$buf60 ;
wire rst_bF$buf61 ;
wire rst_bF$buf62 ;
wire rst_bF$buf63 ;
wire rst_bF$buf64 ;
wire rst_bF$buf65 ;
wire rst_bF$buf66 ;
wire rst_bF$buf67 ;
wire rst_bF$buf68 ;
wire rst_bF$buf69 ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf5  ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire RegWrite ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6521_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf3  ;
wire _5601_ ;
wire [31:0] \datapath_1.mux_pcsrc.dout  ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _5459__bF$buf0 ;
wire _5459__bF$buf1 ;
wire _4910_ ;
wire _5459__bF$buf2 ;
wire _5459__bF$buf3 ;
wire [31:0] \datapath_1.regfile_1.regOut[30]  ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _5463__bF$buf0 ;
wire _5463__bF$buf1 ;
wire _5463__bF$buf2 ;
wire [5:0] \control_1.op  ;
wire _5463__bF$buf3 ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _3032__bF$buf0 ;
wire _3032__bF$buf1 ;
wire _3032__bF$buf2 ;
wire _3032__bF$buf3 ;
wire _3032__bF$buf4 ;
wire _755_ ;
wire _335_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf2  ;
wire _2629_ ;
wire _2209_ ;
wire _6462_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf1  ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf5  ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf2  ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf3  ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _5526__bF$buf0 ;
wire _5526__bF$buf1 ;
wire _5526__bF$buf2 ;
wire _5526__bF$buf3 ;
wire _5526__bF$buf4 ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf4  ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _5530__bF$buf0 ;
wire _5530__bF$buf1 ;
wire _5530__bF$buf2 ;
wire _5530__bF$buf3 ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _5674_ ;
wire _5254_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf2  ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_31_bF$buf2  ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire rst_bF$buf30 ;
wire rst_bF$buf31 ;
wire rst_bF$buf32 ;
wire rst_bF$buf33 ;
wire rst_bF$buf34 ;
wire rst_bF$buf35 ;
wire rst_bF$buf36 ;
wire rst_bF$buf37 ;
wire rst_bF$buf38 ;
wire rst_bF$buf39 ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _2462__bF$buf0 ;
wire _2462__bF$buf1 ;
wire _2462__bF$buf2 ;
wire _2462__bF$buf3 ;
wire _6497_ ;
wire _6077_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf2  ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf0  ;
wire _4657_ ;
wire _4237_ ;
wire _6803_ ;
wire _5545__bF$buf0 ;
wire _5545__bF$buf1 ;
wire _5545__bF$buf2 ;
wire _5545__bF$buf3 ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire [31:0] _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6421_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf3  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire [31:0] _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf2  ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire [31:0] _68_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf6  ;
wire [31:0] \datapath_1.Data  ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire [31:0] \datapath_1.regfile_1.regOut[20]  ;
wire _5466__bF$buf0 ;
wire _5466__bF$buf1 ;
wire _5466__bF$buf2 ;
wire _5466__bF$buf3 ;
wire _5466__bF$buf4 ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6553_ ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf2  ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf0  ;
wire _5633_ ;
wire _5213_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf1  ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _5918_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf5  ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6456_ ;
wire _6036_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf2  ;
wire _1591_ ;
wire _1171_ ;
wire _3977__bF$buf0 ;
wire _3977__bF$buf1 ;
wire _3977__bF$buf2 ;
wire _3977__bF$buf3 ;
wire _3977__bF$buf4 ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf5  ;
wire _5727_ ;
wire _5307_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf3  ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire [31:0] _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _2185_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire MemRead ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire \datapath_1.PCJump_17_bF$buf4  ;
wire _4616_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _3200__bF$buf0 ;
wire _3200__bF$buf1 ;
wire _3200__bF$buf2 ;
wire \datapath_1.regfile_1.regEn_7_bF$buf6  ;
wire _3200__bF$buf3 ;
wire _3200__bF$buf4 ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire clk_hier0_bF$buf8 ;
wire clk_hier0_bF$buf9 ;
wire _2088_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf4  ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf0  ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire clk_bF$buf110 ;
wire clk_bF$buf111 ;
wire clk_bF$buf112 ;
wire clk_bF$buf113 ;
wire _5548__bF$buf0 ;
wire _5548__bF$buf1 ;
wire _5548__bF$buf2 ;
wire _5548__bF$buf3 ;
wire _5548__bF$buf4 ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _6703_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _5552__bF$buf0 ;
wire _5552__bF$buf1 ;
wire _5552__bF$buf2 ;
wire _5552__bF$buf3 ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6512_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf3  ;
wire _3637_ ;
wire _3217_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf3  ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6550_ ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf2  ;
wire _5821_ ;
wire _5401_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf6  ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _5469__bF$buf0 ;
wire _5469__bF$buf1 ;
wire _5469__bF$buf2 ;
wire _5469__bF$buf3 ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire [31:0] \datapath_1.regfile_1.regOut[10]  ;
wire \datapath_1.regfile_1.regEn_18_bF$buf2  ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6453_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf2  ;
wire _5724_ ;
wire _5304_ ;
wire _6509_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf0  ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf7  ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4005__bF$buf0 ;
wire _4005__bF$buf1 ;
wire _4005__bF$buf2 ;
wire _4005__bF$buf3 ;
wire \datapath_1.PCJump_17_bF$buf1  ;
wire _4613_ ;
wire [31:0] \datapath_1.regfile_1.regOut[4]  ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf5  ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf3  ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire [31:0] _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _4707_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_0_bF$buf1  ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire [31:0] \datapath_1.regfile_1.regOut[27]  ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf4  ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf0  ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf0  ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _6603_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf3  ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire MemToReg ;
wire _6641_ ;
wire _6221_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf2  ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6450_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf6  ;
wire _59_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf2  ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf6  ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf4  ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire [31:0] \datapath_1.rd1  ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf2  ;
wire _6773_ ;
wire _6353_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf0  ;
wire _2693_ ;
wire _2273_ ;
wire _5480__bF$buf0 ;
wire _5480__bF$buf1 ;
wire _5480__bF$buf2 ;
wire _5480__bF$buf3 ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _4079__bF$buf0 ;
wire _4079__bF$buf1 ;
wire _4079__bF$buf2 ;
wire _4079__bF$buf3 ;
wire _5624_ ;
wire _5204_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire [5:0] \aluControl_1.inst  ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf7  ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf1  ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf5  ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire PCEn_bF$buf0 ;
wire PCEn_bF$buf1 ;
wire PCEn_bF$buf2 ;
wire PCEn_bF$buf3 ;
wire PCEn_bF$buf4 ;
wire PCEn_bF$buf5 ;
wire PCEn_bF$buf6 ;
wire PCEn_bF$buf7 ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _5539__bF$buf0 ;
wire _5539__bF$buf1 ;
wire _5539__bF$buf2 ;
wire _5539__bF$buf3 ;
wire _5539__bF$buf4 ;
wire _6485_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf1  ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire [31:0] \datapath_1.regfile_1.regOut[17]  ;
wire \datapath_1.PCJump_27_bF$buf4  ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf4  ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_11_bF$buf3  ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf7  ;
wire _3198__bF$buf0 ;
wire _3198__bF$buf1 ;
wire _3198__bF$buf2 ;
wire _3198__bF$buf3 ;
wire _3198__bF$buf4 ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _3935__bF$buf0 ;
wire _3935__bF$buf1 ;
wire _3935__bF$buf2 ;
wire _4777_ ;
wire _3935__bF$buf3 ;
wire _4357_ ;
wire _3935__bF$buf4 ;
wire \datapath_1.regfile_1.regEn_16_bF$buf3  ;
wire _56_ ;
wire _6503_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf3  ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf1  ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6541_ ;
wire _6121_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf2  ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire [31:0] \datapath_1.alu_1.ALUInB  ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf6  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf2  ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_5_bF$buf4  ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire [3:0] \control_1.reg_state.dout  ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf2  ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _5483__bF$buf0 ;
wire _5483__bF$buf1 ;
wire _5483__bF$buf2 ;
wire _5483__bF$buf3 ;
wire _5483__bF$buf4 ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire \datapath_1.PCJump_27_bF$buf1  ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire [31:0] _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf1  ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf0  ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf4  ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf4  ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _4774_ ;
wire _4354_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf0  ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6500_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf3  ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _4583_ ;
wire _4163_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf0  ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf7  ;
wire _1288_ ;
wire _199_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf3  ;
wire _3719_ ;
wire _5565__bF$buf0 ;
wire _5565__bF$buf1 ;
wire _5565__bF$buf2 ;
wire _5565__bF$buf3 ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _6823_ ;
wire _6403_ ;
wire _3942__bF$buf0 ;
wire _3942__bF$buf1 ;
wire _3942__bF$buf2 ;
wire _3942__bF$buf3 ;
wire _2743_ ;
wire _2323_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf3  ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf1  ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire [31:0] _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire ALUOp_0_bF$buf0 ;
wire ALUOp_0_bF$buf1 ;
wire ALUOp_0_bF$buf2 ;
wire ALUOp_0_bF$buf3 ;
wire _2608_ ;
wire ALUOp_0_bF$buf4 ;
wire ALUOp_0_bF$buf5 ;
wire _6441_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf2  ;
wire _5712_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _2590_ ;
wire _2170_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf6  ;
wire _3795_ ;
wire _3375_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf2  ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire \datapath_1.PCJump_22_bF$buf2  ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf6  ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf2  ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _3201__bF$buf0 ;
wire _3201__bF$buf1 ;
wire \datapath_1.regfile_1.regEn_8_bF$buf6  ;
wire _3201__bF$buf2 ;
wire _3201__bF$buf3 ;
wire _3201__bF$buf4 ;
wire _5615_ ;
wire [31:0] \datapath_1.regfile_1.regOut[22]  ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6573_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _2470__bF$buf0 ;
wire _2470__bF$buf1 ;
wire _2470__bF$buf2 ;
wire _2470__bF$buf3 ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf1  ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf1  ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5549__bF$buf0 ;
wire _5549__bF$buf1 ;
wire _5747_ ;
wire _5549__bF$buf2 ;
wire _5327_ ;
wire _5549__bF$buf3 ;
wire _5549__bF$buf4 ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf0  ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf4  ;
wire _1285_ ;
wire _196_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _3882__bF$buf0 ;
wire _3882__bF$buf1 ;
wire _3882__bF$buf2 ;
wire _3882__bF$buf3 ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf0  ;
wire _3716_ ;
wire _6188_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf3  ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf0  ;
wire \datapath_1.regfile_1.regEn_17_bF$buf7  ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf3  ;
wire _6_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf7  ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf3  ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf7  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf3  ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6532_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _5803_ ;
wire _1723_ ;
wire [31:0] _1303_ ;
wire _4195_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf2  ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf3  ;
wire _5612_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf6  ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6570_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire rst_bF$buf100 ;
wire rst_bF$buf101 ;
wire rst_bF$buf102 ;
wire rst_bF$buf103 ;
wire rst_bF$buf104 ;
wire rst_bF$buf105 ;
wire rst_bF$buf106 ;
wire rst_bF$buf107 ;
wire rst_bF$buf108 ;
wire rst_bF$buf109 ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _5489__bF$buf0 ;
wire _5489__bF$buf1 ;
wire _5489__bF$buf2 ;
wire _5489__bF$buf3 ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire rst ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire [31:0] \datapath_1.regfile_1.regOut[12]  ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6473_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf4  ;
wire MemWrite ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire clk_bF$buf76 ;
wire clk_bF$buf77 ;
wire clk_bF$buf78 ;
wire clk_bF$buf79 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf1  ;
wire _6567_ ;
wire _6147_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf4  ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire [31:0] \datapath_1.regfile_1.regOut[6]  ;
wire _5838_ ;
wire _5418_ ;
wire [31:0] _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf0  ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf4  ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf0  ;
wire [31:0] _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [31:0] \datapath_1.regfile_1.regOut[29]  ;
wire _1185_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf4  ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _2199_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_24_bF$buf3  ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire [31:0] _3425_ ;
wire _3005_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf4  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf0  ;
wire \datapath_1.regfile_1.regEn_24_bF$buf7  ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf0  ;
wire _4668_ ;
wire _4248_ ;
wire [4:0] \datapath_1.a3  ;
wire \datapath_1.regfile_1.regEn_29_bF$buf3  ;
wire _6814_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf7  ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _5504__bF$buf0 ;
wire _5504__bF$buf1 ;
wire _5504__bF$buf2 ;
wire _5504__bF$buf3 ;
wire _5504__bF$buf4 ;
wire _6432_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _5703_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6470_ ;
wire _6050_ ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf1  ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6564_ ;
wire _6144_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf1  ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _2293_ ;
wire _3971__bF$buf0 ;
wire _3971__bF$buf1 ;
wire _3971__bF$buf2 ;
wire _3971__bF$buf3 ;
wire _3498_ ;
wire _3971__bF$buf4 ;
wire _3078_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf4  ;
wire _5644_ ;
wire _5224_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf1  ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf7  ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf1  ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire [31:0] _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf0  ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf1  ;
wire _4627_ ;
wire _4207_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf4  ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire [31:0] \datapath_1.regfile_1.regOut[19]  ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf0  ;
wire _6811_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf3  ;
wire _2731_ ;
wire _2311_ ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf4  ;
wire [31:0] _913_ ;
wire _5679_ ;
wire _5259_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf7  ;
wire _6620_ ;
wire _6200_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf3  ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4051__bF$buf0 ;
wire _4283_ ;
wire _4051__bF$buf1 ;
wire _4051__bF$buf2 ;
wire _4051__bF$buf3 ;
wire _722_ ;
wire _302_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf7  ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire rst_bF$buf80 ;
wire rst_bF$buf81 ;
wire rst_bF$buf82 ;
wire rst_bF$buf83 ;
wire rst_bF$buf84 ;
wire rst_bF$buf85 ;
wire rst_bF$buf86 ;
wire rst_bF$buf87 ;
wire rst_bF$buf88 ;
wire rst_bF$buf89 ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _6714_ ;
wire _3955__bF$buf0 ;
wire _3955__bF$buf1 ;
wire _3955__bF$buf2 ;
wire _3955__bF$buf3 ;
wire _3955__bF$buf4 ;
wire _760_ ;
wire _340_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf7  ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6523_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6561_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf1  ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _5499__bF$buf0 ;
wire _6655_ ;
wire _5499__bF$buf1 ;
wire _6235_ ;
wire _5499__bF$buf2 ;
wire _5499__bF$buf3 ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf4  ;
wire _6464_ ;
wire _6044_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _2193_ ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf3  ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire _6558_ ;
wire _6138_ ;
wire [31:0] _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf7  ;
wire _4624_ ;
wire _4204_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf1  ;
wire _5829_ ;
wire _5409_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf4  ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf5  ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf0  ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf1  ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf0  ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _4280_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf4  ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire rst_bF$buf50 ;
wire rst_bF$buf51 ;
wire rst_bF$buf52 ;
wire rst_bF$buf53 ;
wire rst_bF$buf54 ;
wire rst_bF$buf55 ;
wire rst_bF$buf56 ;
wire rst_bF$buf57 ;
wire rst_bF$buf58 ;
wire rst_bF$buf59 ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _3780_ ;
wire [31:0] _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf4  ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf2  ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6423_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf1  ;
wire _2628_ ;
wire _2208_ ;
wire _6461_ ;
wire _6041_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf4  ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _2190_ ;
wire [31:0] \datapath_1.regfile_1.regOut[1]  ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf0  ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire [31:0] _848_ ;
wire _428_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf4  ;
wire _4621_ ;
wire _4201_ ;
wire _5826_ ;
wire _5406_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf1  ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6784_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf2  ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire [31:0] \datapath_1.regfile_1.regOut[24]  ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf3  ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _4038__bF$buf0 ;
wire _4038__bF$buf1 ;
wire _4038__bF$buf2 ;
wire _4038__bF$buf3 ;
wire \datapath_1.regfile_1.regEn_18_bF$buf7  ;
wire _5673_ ;
wire _5253_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf1  ;
wire _6458_ ;
wire _6038_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf4  ;
wire _1593_ ;
wire [31:0] _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf7  ;
wire _5729_ ;
wire _5309_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf5  ;
wire _1649_ ;
wire _1229_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf1  ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire rst_bF$buf20 ;
wire rst_bF$buf21 ;
wire rst_bF$buf22 ;
wire rst_bF$buf23 ;
wire rst_bF$buf24 ;
wire rst_bF$buf25 ;
wire rst_bF$buf26 ;
wire rst_bF$buf27 ;
wire rst_bF$buf28 ;
wire rst_bF$buf29 ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire [31:0] \datapath_1.mux_wd3.dout  ;
wire _1687_ ;
wire _1267_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf1  ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf2  ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf1  ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf5  ;
wire _3639_ ;
wire _3219_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _5521__bF$buf0 ;
wire _5521__bF$buf1 ;
wire _5521__bF$buf2 ;
wire _5521__bF$buf3 ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6552_ ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf1  ;
wire _3677_ ;
wire _3257_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf4  ;
wire _5823_ ;
wire _5403_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf0  ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf4  ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire [31:0] _328_ ;
wire _6455_ ;
wire _6035_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf1  ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf4  ;
wire _5726_ ;
wire _5306_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf2  ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire [31:0] \datapath_1.regfile_1.regOut[14]  ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire \datapath_1.PCJump_17_bF$buf3  ;
wire _4615_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf7  ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf5  ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire _4653_ ;
wire [31:0] memoryWriteData ;
wire _4233_ ;
wire [31:0] \datapath_1.regfile_1.regOut[8]  ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf3  ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire clk_bF$buf100 ;
wire clk_bF$buf101 ;
wire clk_bF$buf102 ;
wire clk_bF$buf103 ;
wire clk_bF$buf104 ;
wire clk_bF$buf105 ;
wire clk_bF$buf106 ;
wire clk_bF$buf107 ;
wire clk_bF$buf108 ;
wire clk_bF$buf109 ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6511_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf2  ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf2  ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _3674_ ;
wire _3254_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf1  ;
wire ALUSrcA ;
wire [1:0] ALUSrcB ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf5  ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _3972__bF$buf0 ;
wire _3972__bF$buf1 ;
wire _3972__bF$buf2 ;
wire _3972__bF$buf3 ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _5524__bF$buf0 ;
wire _5524__bF$buf1 ;
wire _5524__bF$buf2 ;
wire _5524__bF$buf3 ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf1  ;
wire _1834_ ;
wire _1414_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf4  ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6452_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf1  ;
wire _5723_ ;
wire _5303_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf4  ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire PCSource_1_bF$buf0 ;
wire \datapath_1.regfile_1.regEn_2_bF$buf6  ;
wire PCSource_1_bF$buf1 ;
wire PCSource_1_bF$buf2 ;
wire PCSource_1_bF$buf3 ;
wire PCSource_1_bF$buf4 ;
wire [31:0] _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire \datapath_1.PCJump_17_bF$buf0  ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf4  ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf2  ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _3893__bF$buf0 ;
wire _3893__bF$buf1 ;
wire _3893__bF$buf2 ;
wire _3893__bF$buf3 ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _4706_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf3  ;
wire \datapath_1.mux_wd3.dout_0_bF$buf0  ;
wire _3098_ ;
wire _5664_ ;
wire _5244_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf7  ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf3  ;
wire _1678_ ;
wire _1258_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire BranchNe ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf2  ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire ALUZero ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf1  ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf5  ;
wire _58_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf1  ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf5  ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf3  ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _5527__bF$buf0 ;
wire _5527__bF$buf1 ;
wire _5527__bF$buf2 ;
wire _5527__bF$buf3 ;
wire _5527__bF$buf4 ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6543_ ;
wire _6123_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf4  ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5531__bF$buf0 ;
wire _5531__bF$buf1 ;
wire _5531__bF$buf2 ;
wire _5531__bF$buf3 ;
wire _5531__bF$buf4 ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire [31:0] \datapath_1.a  ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf1  ;
wire _6772_ ;
wire _6352_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf4  ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf6  ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire [31:0] _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf0  ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf4  ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf0  ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire \datapath_1.PCJump_27_bF$buf3  ;
wire [31:0] _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf3  ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf2  ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf6  ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [31:0] ALUOut ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _3036__bF$buf0 ;
wire _3036__bF$buf1 ;
wire _3036__bF$buf2 ;
wire _3036__bF$buf3 ;
wire _3036__bF$buf4 ;
wire \datapath_1.regfile_1.regEn_16_bF$buf2  ;
wire _55_ ;
wire _6502_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _5471__bF$buf0 ;
wire _5471__bF$buf1 ;
wire _5471__bF$buf2 ;
wire _5471__bF$buf3 ;
wire _5471__bF$buf4 ;
wire _5471__bF$buf5 ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf2  ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf0  ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf1  ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire [31:0] \datapath_1.alu_1.ALUInA  ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf1  ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf5  ;
wire \datapath_1.regfile_1.regEn_5_bF$buf3  ;
wire ALUSrcB_1_bF$buf0 ;
wire ALUSrcB_1_bF$buf1 ;
wire ALUSrcB_1_bF$buf2 ;
wire ALUSrcB_1_bF$buf3 ;
wire ALUSrcB_1_bF$buf4 ;
wire _3283_ ;
wire _3982__bF$buf0 ;
wire _3982__bF$buf1 ;
wire _3982__bF$buf2 ;
wire _3982__bF$buf3 ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _5534__bF$buf0 ;
wire _5534__bF$buf1 ;
wire _5534__bF$buf2 ;
wire _5534__bF$buf3 ;
wire _5534__bF$buf4 ;
wire _736_ ;
wire _316_ ;
wire _6443_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf1  ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf4  ;
wire _5714_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf4  ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire [31:0] \datapath_1.regfile_1.regOut[3]  ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire \datapath_1.PCJump_27_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_1_bF$buf4  ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire [1:1] PCSource ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _3997__bF$buf0 ;
wire _3997__bF$buf1 ;
wire _3997__bF$buf2 ;
wire _3997__bF$buf3 ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf0  ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire [2:0] ALUControl ;
wire _5655_ ;
wire _5235_ ;
wire [31:0] \datapath_1.regfile_1.regOut[26]  ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _3930__bF$buf0 ;
wire _3930__bF$buf1 ;
wire _3930__bF$buf2 ;
wire _3930__bF$buf3 ;
wire _4735_ ;
wire _4315_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf3  ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf3  ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf2  ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf6  ;
wire _1287_ ;
wire [31:0] _198_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf2  ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _2742_ ;
wire _2322_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf2  ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf0  ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6440_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf1  ;
wire _5711_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf5  ;
wire _3794_ ;
wire _3374_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf1  ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire \datapath_1.PCJump_22_bF$buf1  ;
wire MemToReg_bF$buf0 ;
wire MemToReg_bF$buf1 ;
wire MemToReg_bF$buf2 ;
wire MemToReg_bF$buf3 ;
wire MemToReg_bF$buf4 ;
wire MemToReg_bF$buf5 ;
wire MemToReg_bF$buf6 ;
wire MemToReg_bF$buf7 ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf5  ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6534_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf4  ;
wire _636_ ;
wire _216_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf1  ;
wire _6763_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf5  ;
wire _5614_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6572_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _5708_ ;
wire [31:0] _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf0  ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf0  ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _3196__bF$buf0 ;
wire _3196__bF$buf1 ;
wire _3196__bF$buf2 ;
wire _3196__bF$buf3 ;
wire _3196__bF$buf4 ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire [31:0] \datapath_1.regfile_1.regOut[16]  ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire clk_bF$buf90 ;
wire clk_bF$buf91 ;
wire clk_bF$buf92 ;
wire clk_bF$buf93 ;
wire clk_bF$buf94 ;
wire clk_bF$buf95 ;
wire _3621_ ;
wire clk_bF$buf96 ;
wire clk_bF$buf97 ;
wire _3201_ ;
wire clk_bF$buf98 ;
wire clk_bF$buf99 ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _5784_ ;
wire _5364_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf3  ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf2  ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf6  ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf2  ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf6  ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf2  ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf2  ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6531_ ;
wire _6111_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire _4194_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf1  ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf2  ;
wire _5611_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf5  ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6434_ ;
wire _6014_ ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5544__bF$buf0 ;
wire _5544__bF$buf1 ;
wire _5544__bF$buf2 ;
wire _5544__bF$buf3 ;
wire _5705_ ;
wire [31:0] \datapath_1.regfile_1.regOut[31]  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6472_ ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf3  ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire [31:0] _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf0  ;
wire _859_ ;
wire _439_ ;
wire _6566_ ;
wire _6146_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf3  ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire IRWrite ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _3034__bF$buf0 ;
wire _3034__bF$buf1 ;
wire _3034__bF$buf2 ;
wire _3034__bF$buf3 ;
wire _3034__bF$buf4 ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _3936__bF$buf0 ;
wire _3936__bF$buf1 ;
wire _3936__bF$buf2 ;
wire _3936__bF$buf3 ;
wire _3936__bF$buf4 ;
wire _286_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf3  ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire [31:0] _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf3  ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire rst_hier0_bF$buf0 ;
wire rst_hier0_bF$buf1 ;
wire rst_hier0_bF$buf2 ;
wire rst_hier0_bF$buf3 ;
wire rst_hier0_bF$buf4 ;
wire rst_hier0_bF$buf5 ;
wire rst_hier0_bF$buf6 ;
wire rst_hier0_bF$buf7 ;
wire rst_hier0_bF$buf8 ;
wire rst_hier0_bF$buf9 ;
wire _4001__bF$buf0 ;
wire _4001__bF$buf1 ;
wire _4001__bF$buf2 ;
wire _4001__bF$buf3 ;
wire \datapath_1.mux_wd3.dout_24_bF$buf2  ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf3  ;
wire _4629_ ;
wire _4209_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf6  ;
wire ALUSrcB_0_bF$buf0 ;
wire ALUSrcB_0_bF$buf1 ;
wire ALUSrcB_0_bF$buf2 ;
wire ALUSrcB_0_bF$buf3 ;
wire ALUSrcB_0_bF$buf4 ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf2  ;
wire _6813_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf6  ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire [3:0] \control_1.next  ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6431_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire _533_ ;
wire ALUSrcA_bF$buf0 ;
wire _113_ ;
wire ALUSrcA_bF$buf1 ;
wire ALUSrcA_bF$buf2 ;
wire ALUSrcA_bF$buf3 ;
wire ALUSrcA_bF$buf4 ;
wire ALUSrcA_bF$buf5 ;
wire _2827_ ;
wire ALUSrcA_bF$buf6 ;
wire _2407_ ;
wire ALUSrcA_bF$buf7 ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _3995__bF$buf0 ;
wire _3995__bF$buf1 ;
wire _3995__bF$buf2 ;
wire _3995__bF$buf3 ;
wire _3995__bF$buf4 ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf0  ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _3924__bF$buf0 ;
wire _3924__bF$buf1 ;
wire _3924__bF$buf2 ;
wire _3924__bF$buf3 ;
wire _5605_ ;
wire [31:0] \datapath_1.regfile_1.regOut[21]  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6563_ ;
wire _6143_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf0  ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf3  ;
wire _5643_ ;
wire _5223_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire [31:0] _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf0  ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf6  ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf0  ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3037__bF$buf0 ;
wire _3037__bF$buf1 ;
wire _3037__bF$buf2 ;
wire _3037__bF$buf3 ;
wire _3037__bF$buf4 ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _5472__bF$buf0 ;
wire _5472__bF$buf1 ;
wire _5472__bF$buf2 ;
wire _5472__bF$buf3 ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf0  ;
wire _4626_ ;
wire _4206_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf3  ;
wire _5570__bF$buf0 ;
wire _5570__bF$buf1 ;
wire _5570__bF$buf2 ;
wire _5570__bF$buf3 ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf7  ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire [3:0] _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf2  ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf3  ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf6  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf2  ;
wire _1598_ ;
wire _1178_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf6  ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire rst_bF$buf70 ;
wire rst_bF$buf71 ;
wire rst_bF$buf72 ;
wire rst_bF$buf73 ;
wire rst_bF$buf74 ;
wire rst_bF$buf75 ;
wire rst_bF$buf76 ;
wire rst_bF$buf77 ;
wire rst_bF$buf78 ;
wire rst_bF$buf79 ;
wire [31:1] \datapath_1.regfile_1.regEn  ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf6  ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6522_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6751_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf4  ;
wire _5602_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6560_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire [31:0] _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _3998__bF$buf0 ;
wire _3998__bF$buf1 ;
wire _3998__bF$buf2 ;
wire _3998__bF$buf3 ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _3494_ ;
wire _3074_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf0  ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire [31:0] _718_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire [31:0] \datapath_1.regfile_1.regOut[11]  ;
wire _1845_ ;
wire _3931__bF$buf0 ;
wire _1425_ ;
wire _3931__bF$buf1 ;
wire _1005_ ;
wire _3931__bF$buf2 ;
wire _3931__bF$buf3 ;
wire _756_ ;
wire _336_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf3  ;
wire _6463_ ;
wire _6043_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire [31:0] _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf2  ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf6  ;
wire _4623_ ;
wire _4203_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf0  ;
wire [31:0] \datapath_1.regfile_1.regOut[5]  ;
wire _5828_ ;
wire _5408_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf3  ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf4  ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire [31:0] \datapath_1.ALUResult  ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf0  ;
wire _5675_ ;
wire _5255_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf3  ;
wire [31:0] \datapath_1.regfile_1.regOut[28]  ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _3950__bF$buf0 ;
wire _3950__bF$buf1 ;
wire _3950__bF$buf2 ;
wire _3950__bF$buf3 ;
wire \datapath_1.regfile_1.regEn_4_bF$buf7  ;
wire \datapath_1.regfile_1.regEn_31_bF$buf3  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire rst_bF$buf40 ;
wire rst_bF$buf41 ;
wire rst_bF$buf42 ;
wire rst_bF$buf43 ;
wire rst_bF$buf44 ;
wire rst_bF$buf45 ;
wire rst_bF$buf46 ;
wire rst_bF$buf47 ;
wire rst_bF$buf48 ;
wire rst_bF$buf49 ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _1689_ ;
wire _1269_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf3  ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire [31:0] _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [31:0] memoryAddress ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf1  ;
wire _4658_ ;
wire _4238_ ;
wire _6804_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire PCEn ;
wire _906_ ;
wire _6613_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6422_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf4  ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf0  ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6460_ ;
wire _6040_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf3  ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf7  ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire [31:8] \datapath_1.PCJump  ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf3  ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf0  ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf1  ;
wire _5634_ ;
wire _5214_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf2  ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf6  ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf0  ;
wire _6457_ ;
wire _6037_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf3  ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf6  ;
wire _5728_ ;
wire _5308_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf4  ;
wire _1648_ ;
wire _1228_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf0  ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire rst_bF$buf10 ;
wire rst_bF$buf11 ;
wire rst_bF$buf12 ;
wire rst_bF$buf13 ;
wire rst_bF$buf14 ;
wire rst_bF$buf15 ;
wire rst_bF$buf16 ;
wire rst_bF$buf17 ;
wire rst_bF$buf18 ;
wire rst_bF$buf19 ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _5478__bF$buf0 ;
wire _5478__bF$buf1 ;
wire _5478__bF$buf2 ;
wire _5478__bF$buf3 ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf0  ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire [31:0] \datapath_1.regfile_1.regOut[18]  ;
wire _1495_ ;
wire _1075_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf7  ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf1  ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire [27:0] \datapath_1.mux_iord.din0  ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _6704_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf0  ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6513_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf4  ;
wire _3638_ ;
wire _3218_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf4  ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _2481__bF$buf0 ;
wire _2481__bF$buf1 ;
wire _6551_ ;
wire _2481__bF$buf2 ;
wire _6131_ ;
wire _2481__bF$buf3 ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf0  ;
wire _3676_ ;
wire _3256_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf3  ;
wire _5822_ ;
wire _5402_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire [31:0] _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _2280_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf7  ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf3  ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6454_ ;
wire _6034_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf0  ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf3  ;
wire _5725_ ;
wire _5305_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf1  ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire \datapath_1.PCJump_17_bF$buf2  ;
wire _4614_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf6  ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf4  ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf2  ;
wire _5485__bF$buf0 ;
wire _5485__bF$buf1 ;
wire _5485__bF$buf2 ;
wire _5485__bF$buf3 ;
wire _5485__bF$buf4 ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf1  ;
wire _3635_ ;
wire _3215_ ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf1  ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _3673_ ;
wire _3253_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf0  ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _6604_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf4  ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf0  ;
wire _1833_ ;
wire _1413_ ;
wire IorD_bF$buf0 ;
wire IorD_bF$buf1 ;
wire IorD_bF$buf2 ;
wire IorD_bF$buf3 ;
wire IorD_bF$buf4 ;
wire IorD_bF$buf5 ;
wire \datapath_1.mux_wd3.dout_16_bF$buf3  ;
wire IorD_bF$buf6 ;
wire IorD_bF$buf7 ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6451_ ;
wire _6031_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf0  ;
wire _5722_ ;
wire _5302_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf7  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf3  ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire [31:0] _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _2180_ ;
wire [31:0] \datapath_1.regfile_1.regOut[0]  ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf7  ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf5  ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire [31:0] \datapath_1.rd2  ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _3944__bF$buf0 ;
wire _3944__bF$buf1 ;
wire _3944__bF$buf2 ;
wire _3944__bF$buf3 ;
wire _3944__bF$buf4 ;
wire _647_ ;
wire _227_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf3  ;
wire _6774_ ;
wire _6354_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf1  ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire [31:0] \datapath_1.regfile_1.regOut[23]  ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire [31:0] memoryOutData ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire [1:0] ALUOp ;
wire _5500__bF$buf0 ;
wire _685_ ;
wire _5500__bF$buf1 ;
wire _265_ ;
wire _5500__bF$buf2 ;
wire _5500__bF$buf3 ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _4705_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf2  ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf6  ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;

FILL FILL_4__13745_ (
);

FILL FILL_4__13325_ (
);

FILL FILL_3__7095_ (
);

AOI21X1 _11689_ (
    .A(_2779_),
    .B(_2780_),
    .C(_2789_),
    .Y(_2790_)
);

INVX2 _11269_ (
    .A(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2388_)
);

FILL FILL_3__12738_ (
);

FILL FILL_1__13772_ (
);

FILL FILL_3__12318_ (
);

FILL FILL_1__13352_ (
);

FILL SFILL84280x62050 (
);

FILL FILL_0__12765_ (
);

INVX1 _12630_ (
    .A(\datapath_1.Data [21]),
    .Y(_3466_)
);

FILL FILL_0__12345_ (
);

OAI21X1 _12210_ (
    .A(_3192_),
    .B(ALUSrcA_bF$buf5),
    .C(_3193_),
    .Y(\datapath_1.alu_1.ALUInA [31])
);

FILL FILL_5__8382_ (
);

FILL FILL_5__15957_ (
);

FILL FILL_5__15537_ (
);

FILL FILL_5__15117_ (
);

DFFSR _9837_ (
    .Q(\datapath_1.regfile_1.regOut[23] [23]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1433_[23])
);

FILL FILL_3__16151_ (
);

OAI21X1 _9417_ (
    .A(_1291_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .C(_1292_),
    .Y(_1238_[27])
);

FILL FILL_5__10672_ (
);

FILL SFILL23960x58050 (
);

FILL FILL_1__8374_ (
);

FILL FILL_5__10252_ (
);

FILL FILL_2__15984_ (
);

FILL FILL_2__15564_ (
);

FILL FILL_2__15144_ (
);

FILL FILL_1__14977_ (
);

FILL FILL_1__14557_ (
);

FILL FILL_1__14137_ (
);

FILL SFILL84200x60050 (
);

FILL FILL_3__9661_ (
);

INVX1 _13835_ (
    .A(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_4340_)
);

FILL FILL_3__9241_ (
);

NOR2X1 _13415_ (
    .A(_3926_),
    .B(_3921_),
    .Y(_3927_)
);

FILL FILL_5__9167_ (
);

FILL FILL_6__12464_ (
);

FILL FILL_6__12044_ (
);

FILL FILL_0__14911_ (
);

FILL SFILL109480x60050 (
);

FILL FILL_5__11877_ (
);

FILL FILL_1__9999_ (
);

FILL FILL_5__11457_ (
);

FILL FILL_3__12491_ (
);

FILL FILL_5__11037_ (
);

FILL FILL_1__9159_ (
);

FILL FILL_3__12071_ (
);

FILL FILL_2__16349_ (
);

FILL FILL_4__7584_ (
);

FILL SFILL23960x13050 (
);

FILL SFILL79800x8050 (
);

FILL FILL_4__7164_ (
);

FILL FILL_2__11484_ (
);

FILL FILL_2__11064_ (
);

FILL FILL_1__10897_ (
);

FILL FILL_1__10057_ (
);

FILL FILL_4__11811_ (
);

FILL FILL_5__15290_ (
);

FILL FILL_0__7484_ (
);

FILL FILL_0__7064_ (
);

INVX1 _9590_ (
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_1431_)
);

OAI21X1 _9170_ (
    .A(_1167_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1168_),
    .Y(_1108_[30])
);

FILL FILL_6__13669_ (
);

FILL FILL_3__10804_ (
);

FILL FILL_6__13249_ (
);

FILL FILL_4__14283_ (
);

FILL FILL_2__8863_ (
);

FILL FILL_0__10831_ (
);

FILL FILL_2__8443_ (
);

FILL FILL_3__13696_ (
);

FILL FILL_3__13276_ (
);

FILL FILL_0__10411_ (
);

FILL FILL_6__14610_ (
);

FILL FILL_0_BUFX2_insert900 (
);

FILL FILL_4__8789_ (
);

FILL FILL_4__8369_ (
);

FILL FILL_0_BUFX2_insert901 (
);

FILL FILL_0_BUFX2_insert902 (
);

FILL FILL_0_BUFX2_insert903 (
);

FILL FILL_0_BUFX2_insert904 (
);

FILL FILL_2__12269_ (
);

FILL FILL_0_BUFX2_insert905 (
);

FILL FILL_0_BUFX2_insert906 (
);

FILL FILL_5__13603_ (
);

FILL FILL_0_BUFX2_insert907 (
);

FILL FILL_0_BUFX2_insert908 (
);

FILL FILL_0_BUFX2_insert909 (
);

DFFSR _7903_ (
    .Q(\datapath_1.regfile_1.regOut[8] [9]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_458_[9])
);

FILL FILL_1__6860_ (
);

FILL FILL_4__9730_ (
);

FILL FILL_2__13630_ (
);

FILL FILL_2__13210_ (
);

FILL FILL_5__16075_ (
);

FILL FILL_0__8269_ (
);

FILL SFILL13560x42050 (
);

FILL FILL_1__12623_ (
);

FILL FILL_4__15488_ (
);

FILL FILL_1__12203_ (
);

FILL FILL_4__15068_ (
);

FILL FILL_2__9648_ (
);

FILL FILL_0__9630_ (
);

FILL FILL_2__9228_ (
);

OAI21X1 _11901_ (
    .A(_2974_),
    .B(IorD_bF$buf3),
    .C(_2975_),
    .Y(_1_[4])
);

FILL FILL_0__9210_ (
);

FILL FILL_0__11616_ (
);

FILL FILL_1__15095_ (
);

FILL FILL_6_CLKBUF1_insert1078 (
);

FILL FILL_5__7233_ (
);

AOI22X1 _14793_ (
    .A(_4154_),
    .B(\datapath_1.regfile_1.regOut[14] [28]),
    .C(\datapath_1.regfile_1.regOut[31] [28]),
    .D(_3995__bF$buf3),
    .Y(_5277_)
);

OAI22X1 _14373_ (
    .A(_3949_),
    .B(_4864_),
    .C(_3977__bF$buf0),
    .D(_4865_),
    .Y(_4866_)
);

FILL FILL_0__14088_ (
);

FILL FILL_5__14808_ (
);

FILL FILL_3__15842_ (
);

FILL FILL_3__15422_ (
);

FILL FILL_3__15002_ (
);

FILL FILL_1__7225_ (
);

FILL FILL_2__14835_ (
);

FILL FILL_2__14415_ (
);

FILL FILL_1__13828_ (
);

FILL FILL_1__13408_ (
);

FILL FILL_3__8512_ (
);

FILL SFILL104360x48050 (
);

FILL FILL_5__8858_ (
);

FILL FILL_5__8438_ (
);

FILL FILL_5__8018_ (
);

NOR2X1 _15998_ (
    .A(_6453_),
    .B(_6454_),
    .Y(_6455_)
);

OAI22X1 _15578_ (
    .A(_5527__bF$buf2),
    .B(_4609_),
    .C(_6044_),
    .D(_5532__bF$buf2),
    .Y(_6045_)
);

INVX1 _15158_ (
    .A(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_5636_)
);

FILL FILL_3__16207_ (
);

INVX1 _10293_ (
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_1734_)
);

FILL FILL_5__10308_ (
);

FILL FILL_3__11762_ (
);

FILL FILL_3__11342_ (
);

FILL FILL_4__6855_ (
);

FILL FILL_0__16234_ (
);

FILL FILL_2__10755_ (
);

FILL FILL_5__14981_ (
);

FILL FILL_5__14561_ (
);

FILL FILL_5__14141_ (
);

FILL FILL112440x54050 (
);

INVX1 _8861_ (
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_1003_)
);

FILL FILL_6__7302_ (
);

INVX1 _8441_ (
    .A(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_784_)
);

OAI21X1 _8021_ (
    .A(_584_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_585_),
    .Y(_523_[31])
);

FILL FILL_4__13974_ (
);

FILL FILL_4__13554_ (
);

FILL FILL_4__13134_ (
);

INVX2 _11498_ (
    .A(_2442_),
    .Y(_2611_)
);

INVX2 _11078_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .Y(_2197_)
);

FILL FILL_2__7714_ (
);

FILL FILL_3__12967_ (
);

FILL SFILL108600x54050 (
);

FILL FILL_3__12127_ (
);

FILL FILL_1__13581_ (
);

FILL FILL_1__13161_ (
);

FILL FILL_0__12994_ (
);

FILL FILL_3_CLKBUF1_insert180 (
);

FILL FILL_0__12574_ (
);

FILL FILL_3_CLKBUF1_insert181 (
);

FILL FILL_0__12154_ (
);

FILL FILL_3_CLKBUF1_insert182 (
);

FILL FILL_3_CLKBUF1_insert183 (
);

FILL FILL_3_CLKBUF1_insert184 (
);

FILL FILL_5__8191_ (
);

FILL FILL_3_CLKBUF1_insert185 (
);

FILL FILL_3_CLKBUF1_insert186 (
);

FILL FILL_3_CLKBUF1_insert187 (
);

FILL FILL_3_CLKBUF1_insert188 (
);

FILL FILL_5_BUFX2_insert300 (
);

FILL FILL_3_CLKBUF1_insert189 (
);

FILL FILL_5_BUFX2_insert301 (
);

FILL FILL_2__12901_ (
);

FILL FILL_5__15766_ (
);

FILL FILL_5_BUFX2_insert302 (
);

FILL FILL_5__15346_ (
);

FILL FILL_5_BUFX2_insert303 (
);

FILL FILL_3__16380_ (
);

FILL FILL_5_BUFX2_insert304 (
);

OAI21X1 _9646_ (
    .A(_1403_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .C(_1404_),
    .Y(_1368_[18])
);

OAI21X1 _9226_ (
    .A(_1184_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1185_),
    .Y(_1173_[6])
);

FILL FILL_5_BUFX2_insert305 (
);

FILL FILL_5_BUFX2_insert306 (
);

FILL FILL_5__10061_ (
);

FILL FILL_1__8183_ (
);

FILL FILL_5_BUFX2_insert307 (
);

FILL FILL_5_BUFX2_insert308 (
);

FILL FILL_4__14759_ (
);

FILL FILL_2__15793_ (
);

FILL FILL_4__14339_ (
);

FILL FILL_5_BUFX2_insert309 (
);

FILL FILL_2__15373_ (
);

FILL FILL_0__8901_ (
);

FILL FILL_1__14786_ (
);

FILL FILL_1__14366_ (
);

FILL FILL_5__6924_ (
);

FILL FILL_4__15700_ (
);

FILL FILL_3__9890_ (
);

FILL FILL_0__13779_ (
);

FILL FILL_3__9470_ (
);

FILL FILL_0__13359_ (
);

NOR2X1 _13644_ (
    .A(_4151_),
    .B(_4148_),
    .Y(_4152_)
);

NAND2X1 _13224_ (
    .A(\datapath_1.a3 [4]),
    .B(_3754_),
    .Y(_3767_)
);

FILL FILL_5__9396_ (
);

FILL FILL_1__6916_ (
);

FILL FILL_0__14720_ (
);

FILL FILL_0__14300_ (
);

FILL FILL_5__11686_ (
);

FILL FILL_1__9388_ (
);

FILL FILL_5__11266_ (
);

FILL SFILL49240x19050 (
);

FILL FILL_2__16158_ (
);

FILL FILL_4__10679_ (
);

FILL FILL_4__10259_ (
);

FILL FILL_2__11293_ (
);

FILL FILL_5__7709_ (
);

FILL FILL_2_BUFX2_insert430 (
);

FILL FILL_2_BUFX2_insert431 (
);

FILL FILL_1__10286_ (
);

FILL FILL_2_BUFX2_insert432 (
);

FILL FILL_2_BUFX2_insert433 (
);

NOR2X1 _14849_ (
    .A(_5331_),
    .B(_3971__bF$buf1),
    .Y(_5332_)
);

FILL FILL_2_BUFX2_insert434 (
);

OAI22X1 _14429_ (
    .A(_3983__bF$buf1),
    .B(_4919_),
    .C(_3971__bF$buf0),
    .D(_4920_),
    .Y(_4921_)
);

FILL FILL_4__11620_ (
);

INVX1 _14009_ (
    .A(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_4510_)
);

FILL FILL_2_BUFX2_insert435 (
);

FILL FILL_4__11200_ (
);

FILL FILL_2_BUFX2_insert436 (
);

FILL FILL_2_BUFX2_insert437 (
);

FILL FILL_0__7293_ (
);

FILL FILL_2_BUFX2_insert438 (
);

FILL FILL_2_BUFX2_insert439 (
);

FILL FILL_0_CLKBUF1_insert130 (
);

FILL FILL_0_CLKBUF1_insert131 (
);

FILL FILL_4__14092_ (
);

FILL FILL_0__15925_ (
);

FILL FILL_0_CLKBUF1_insert132 (
);

FILL FILL_0_CLKBUF1_insert133 (
);

FILL FILL_0__15505_ (
);

FILL SFILL94280x14050 (
);

FILL FILL_0_CLKBUF1_insert134 (
);

FILL FILL_0_CLKBUF1_insert135 (
);

FILL FILL_0_CLKBUF1_insert136 (
);

FILL FILL_0__10640_ (
);

FILL FILL_2__8252_ (
);

FILL FILL_0_CLKBUF1_insert137 (
);

FILL FILL_3__13085_ (
);

FILL FILL_0_CLKBUF1_insert138 (
);

FILL FILL_0_CLKBUF1_insert139 (
);

FILL FILL_4__8598_ (
);

FILL FILL_2__12498_ (
);

FILL FILL_2__12078_ (
);

FILL FILL_5__13832_ (
);

FILL FILL_5__13412_ (
);

FILL SFILL8680x76050 (
);

INVX1 _7712_ (
    .A(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_420_)
);

FILL FILL_4__12825_ (
);

FILL FILL_4__12405_ (
);

FILL FILL_0__8498_ (
);

FILL FILL_0__8078_ (
);

INVX1 _10769_ (
    .A(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_1970_)
);

DFFSR _10349_ (
    .Q(\datapath_1.regfile_1.regOut[27] [23]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_1693_[23])
);

FILL FILL_3__11818_ (
);

FILL FILL_1__12852_ (
);

FILL FILL_1__12432_ (
);

FILL FILL_4__15297_ (
);

FILL FILL_1__12012_ (
);

FILL SFILL84280x57050 (
);

FILL FILL_2__9877_ (
);

FILL FILL_0__11845_ (
);

FILL FILL_2__9037_ (
);

FILL FILL_0__11425_ (
);

AND2X2 _11710_ (
    .A(_2807_),
    .B(_2808_),
    .Y(_2809_)
);

FILL FILL_0__11005_ (
);

FILL FILL_5__7882_ (
);

FILL FILL_6__15204_ (
);

FILL FILL_5__7462_ (
);

FILL FILL_5__7042_ (
);

NAND3X1 _14182_ (
    .A(_4677_),
    .B(_4678_),
    .C(_4676_),
    .Y(_4679_)
);

FILL FILL_5__14617_ (
);

FILL FILL_3__15651_ (
);

FILL SFILL8600x74050 (
);

FILL FILL_3__15231_ (
);

OAI21X1 _8917_ (
    .A(_1039_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .C(_1040_),
    .Y(_978_[31])
);

FILL FILL_1__7874_ (
);

FILL FILL_1__7454_ (
);

FILL FILL_1__7034_ (
);

FILL SFILL48840x81050 (
);

FILL SFILL8680x31050 (
);

FILL FILL_2__14644_ (
);

FILL FILL_2__14224_ (
);

FILL FILL_1__13637_ (
);

FILL FILL_1__13217_ (
);

FILL SFILL84200x55050 (
);

FILL FILL_1_BUFX2_insert450 (
);

FILL FILL_3__8741_ (
);

FILL FILL_1_BUFX2_insert451 (
);

FILL FILL_3__8321_ (
);

OAI21X1 _12915_ (
    .A(_3614_),
    .B(vdd),
    .C(_3615_),
    .Y(_3555_[30])
);

FILL FILL_1_BUFX2_insert452 (
);

FILL FILL_1_BUFX2_insert453 (
);

FILL FILL_1_BUFX2_insert454 (
);

FILL SFILL84280x12050 (
);

FILL FILL_1_BUFX2_insert455 (
);

FILL FILL_1_BUFX2_insert456 (
);

FILL FILL_5__8247_ (
);

FILL FILL_1_BUFX2_insert457 (
);

FILL FILL_1_BUFX2_insert458 (
);

FILL FILL_1_BUFX2_insert459 (
);

FILL SFILL13640x75050 (
);

NOR2X1 _15387_ (
    .A(_5858_),
    .B(_5856_),
    .Y(_5859_)
);

FILL FILL_6__11124_ (
);

FILL SFILL69000x35050 (
);

FILL SFILL109480x55050 (
);

FILL FILL_3__16016_ (
);

FILL FILL_5__10957_ (
);

FILL FILL_3__11991_ (
);

FILL FILL_1__8659_ (
);

FILL FILL_5__10537_ (
);

FILL FILL_1__8239_ (
);

FILL FILL_3__11571_ (
);

FILL FILL_5__10117_ (
);

FILL FILL_3__11151_ (
);

FILL FILL_2__15849_ (
);

FILL FILL_2__15429_ (
);

FILL FILL_2__15009_ (
);

FILL FILL_0__16043_ (
);

FILL FILL_2__10564_ (
);

FILL FILL_2__10144_ (
);

FILL FILL_1__9600_ (
);

FILL FILL_3__9526_ (
);

FILL FILL_3__9106_ (
);

FILL FILL_5__14790_ (
);

FILL SFILL109880x24050 (
);

FILL FILL_5__14370_ (
);

FILL FILL_0__6984_ (
);

FILL SFILL74280x55050 (
);

DFFSR _8670_ (
    .Q(\datapath_1.regfile_1.regOut[14] [8]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_848_[8])
);

OAI21X1 _8250_ (
    .A(_696_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .C(_697_),
    .Y(_653_[22])
);

FILL FILL_4__13783_ (
);

FILL FILL_4__13363_ (
);

FILL SFILL13640x30050 (
);

FILL FILL_2__7943_ (
);

FILL FILL_3__12776_ (
);

FILL FILL_2__7103_ (
);

FILL FILL_3__12356_ (
);

FILL FILL_1__13390_ (
);

FILL SFILL109480x10050 (
);

FILL FILL_4__7869_ (
);

FILL FILL_4__7449_ (
);

FILL FILL_2__11769_ (
);

FILL FILL_2__11349_ (
);

FILL FILL_0__12383_ (
);

FILL FILL_2_CLKBUF1_insert170 (
);

FILL FILL_2_CLKBUF1_insert171 (
);

FILL FILL_5__15995_ (
);

FILL FILL_2_CLKBUF1_insert172 (
);

FILL FILL_2_CLKBUF1_insert173 (
);

FILL FILL_2__12710_ (
);

FILL FILL_5__15575_ (
);

FILL SFILL74200x53050 (
);

FILL FILL_2_CLKBUF1_insert174 (
);

FILL FILL_5__15155_ (
);

FILL FILL_0__7349_ (
);

OAI21X1 _9875_ (
    .A(_1515_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .C(_1516_),
    .Y(_1498_[9])
);

FILL FILL_2_CLKBUF1_insert175 (
);

FILL FILL_2_CLKBUF1_insert176 (
);

DFFSR _9455_ (
    .Q(\datapath_1.regfile_1.regOut[20] [25]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_1238_[25])
);

NAND2X1 _9035_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1099_)
);

FILL FILL_2_CLKBUF1_insert177 (
);

FILL FILL_2_CLKBUF1_insert178 (
);

FILL FILL_5__10290_ (
);

FILL FILL_2_CLKBUF1_insert179 (
);

FILL FILL_4__14988_ (
);

FILL SFILL74280x10050 (
);

FILL FILL_4__14568_ (
);

FILL FILL_1__11703_ (
);

FILL FILL_4__14148_ (
);

FILL FILL_2__15182_ (
);

FILL FILL_2__8728_ (
);

FILL FILL_0__8710_ (
);

FILL FILL_1__14595_ (
);

FILL FILL_1__14175_ (
);

FILL FILL_6_BUFX2_insert1053 (
);

FILL FILL_0__13588_ (
);

NAND3X1 _13873_ (
    .A(_4368_),
    .B(_4369_),
    .C(_4376_),
    .Y(_4377_)
);

FILL FILL_0__13168_ (
);

INVX1 _13453_ (
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_3965_)
);

NAND2X1 _13033_ (
    .A(vdd),
    .B(\datapath_1.rd2 [27]),
    .Y(_3674_)
);

FILL FILL_6_BUFX2_insert1058 (
);

FILL FILL_3__14922_ (
);

FILL FILL_3__14502_ (
);

FILL FILL_2__13915_ (
);

FILL FILL_5__11495_ (
);

FILL FILL112120x73050 (
);

FILL FILL_5__11075_ (
);

FILL FILL_1__12908_ (
);

FILL FILL_2__16387_ (
);

FILL FILL_4__10488_ (
);

FILL FILL_0__9915_ (
);

FILL FILL_4__10068_ (
);

FILL FILL_5__7938_ (
);

AOI22X1 _14658_ (
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .B(_4005__bF$buf0),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_5145_)
);

INVX1 _14238_ (
    .A(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_4734_)
);

FILL FILL_3__15707_ (
);

FILL FILL_1__16321_ (
);

FILL FILL_3__10422_ (
);

FILL FILL_3__10002_ (
);

FILL FILL_0__15734_ (
);

FILL FILL_0__15314_ (
);

FILL FILL_2__8481_ (
);

FILL FILL_2__8061_ (
);

FILL SFILL64200x51050 (
);

FILL FILL_5__13641_ (
);

FILL FILL112440x49050 (
);

FILL FILL_5__13221_ (
);

INVX1 _7941_ (
    .A(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_532_)
);

DFFSR _7521_ (
    .Q(\datapath_1.regfile_1.regOut[5] [11]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_263_[11])
);

OAI21X1 _7101_ (
    .A(_113_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_114_),
    .Y(_68_[23])
);

FILL FILL_4__12634_ (
);

FILL FILL_4__12214_ (
);

INVX2 _10998_ (
    .A(_2116_),
    .Y(_2117_)
);

OAI21X1 _10578_ (
    .A(_1882_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1883_),
    .Y(_1823_[30])
);

FILL SFILL33720x67050 (
);

OAI21X1 _10158_ (
    .A(_1663_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1664_),
    .Y(_1628_[18])
);

FILL FILL_3__11627_ (
);

FILL FILL_1__12661_ (
);

FILL FILL_3__11207_ (
);

FILL FILL_1__12241_ (
);

FILL FILL_2__9266_ (
);

FILL FILL_0__11654_ (
);

FILL FILL_0__11234_ (
);

FILL FILL_3__14099_ (
);

FILL FILL_6__15853_ (
);

FILL FILL_5__7691_ (
);

FILL FILL_5__14846_ (
);

FILL FILL_5__14426_ (
);

FILL FILL_3__15880_ (
);

FILL FILL_5__14006_ (
);

FILL FILL_3__15460_ (
);

FILL FILL_3__15040_ (
);

OAI21X1 _8726_ (
    .A(_932_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .C(_933_),
    .Y(_913_[10])
);

DFFSR _8306_ (
    .Q(\datapath_1.regfile_1.regOut[11] [28]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_653_[28])
);

FILL FILL_1__7683_ (
);

FILL FILL_4__13839_ (
);

FILL FILL_2__14873_ (
);

FILL FILL_4__13419_ (
);

FILL FILL_2__14453_ (
);

FILL FILL_2__14033_ (
);

FILL FILL_3__7189_ (
);

FILL FILL_1__13866_ (
);

FILL FILL_1__13446_ (
);

FILL FILL_1__13026_ (
);

FILL SFILL33720x22050 (
);

FILL FILL_3__8970_ (
);

FILL FILL_0__12859_ (
);

OAI21X1 _12724_ (
    .A(_3507_),
    .B(IRWrite_bF$buf3),
    .C(_3508_),
    .Y(_3490_[9])
);

FILL FILL_0__12439_ (
);

FILL FILL_3__8130_ (
);

FILL FILL_0__12019_ (
);

NAND3X1 _12304_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf0),
    .Y(_3267_)
);

FILL FILL_5__8896_ (
);

FILL FILL_5__8476_ (
);

FILL SFILL58920x71050 (
);

FILL FILL_5__8056_ (
);

FILL FILL_6__11773_ (
);

NAND2X1 _15196_ (
    .A(_5669_),
    .B(_5672_),
    .Y(_5673_)
);

FILL FILL_0__13800_ (
);

FILL FILL_3__16245_ (
);

FILL FILL_5__10766_ (
);

FILL FILL_1__8888_ (
);

FILL FILL_1__8468_ (
);

FILL FILL_3__11380_ (
);

FILL FILL_2__15658_ (
);

FILL FILL_4__6893_ (
);

FILL FILL_2__15238_ (
);

FILL FILL_0__16272_ (
);

FILL FILL_2__10793_ (
);

FILL FILL_2__10373_ (
);

FILL FILL_3__9755_ (
);

FILL SFILL103960x60050 (
);

FILL FILL_3__9335_ (
);

NOR2X1 _13929_ (
    .A(_4421_),
    .B(_4431_),
    .Y(_4432_)
);

FILL FILL_4__10700_ (
);

INVX1 _13509_ (
    .A(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_4020_)
);

FILL FILL_4__13592_ (
);

FILL FILL_4__13172_ (
);

FILL SFILL109640x81050 (
);

FILL FILL_2__7752_ (
);

FILL FILL_3__12585_ (
);

FILL FILL_2__7332_ (
);

FILL FILL_3__12165_ (
);

FILL FILL_4__7678_ (
);

FILL FILL_2__11998_ (
);

FILL FILL_2__11578_ (
);

FILL FILL_2__11158_ (
);

FILL FILL_0__12192_ (
);

FILL FILL_5__12912_ (
);

FILL FILL_6__16391_ (
);

FILL FILL_4__11905_ (
);

FILL SFILL23720x20050 (
);

FILL FILL_0__7998_ (
);

FILL FILL_5__15384_ (
);

FILL FILL_0__7578_ (
);

FILL FILL_0__7158_ (
);

NAND2X1 _9684_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1430_)
);

NAND2X1 _9264_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1211_)
);

FILL FILL_1_CLKBUF1_insert160 (
);

FILL FILL_1_CLKBUF1_insert161 (
);

FILL FILL_1__11932_ (
);

FILL FILL_4__14797_ (
);

FILL FILL_1_CLKBUF1_insert162 (
);

FILL FILL_4__14377_ (
);

FILL FILL_1_CLKBUF1_insert163 (
);

FILL FILL_1__11512_ (
);

FILL FILL_1_CLKBUF1_insert164 (
);

FILL FILL_1_CLKBUF1_insert165 (
);

FILL FILL_1_CLKBUF1_insert166 (
);

FILL FILL_1_CLKBUF1_insert167 (
);

FILL FILL_1_CLKBUF1_insert168 (
);

FILL FILL_2__8957_ (
);

FILL FILL_0__10925_ (
);

FILL FILL_1_CLKBUF1_insert169 (
);

FILL FILL_2__8117_ (
);

FILL FILL_0__10505_ (
);

FILL FILL_5__6962_ (
);

AOI22X1 _13682_ (
    .A(_3882__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[29] [4]),
    .C(\datapath_1.regfile_1.regOut[25] [4]),
    .D(_4040_),
    .Y(_4190_)
);

FILL FILL_0__13397_ (
);

NAND2X1 _13262_ (
    .A(_3751_),
    .B(_3804_),
    .Y(_3805_)
);

FILL FILL_3__14731_ (
);

FILL FILL_3__14311_ (
);

FILL FILL_1__6954_ (
);

FILL FILL_4__9404_ (
);

FILL SFILL13720x63050 (
);

FILL FILL_2__13724_ (
);

FILL FILL_2__13304_ (
);

FILL FILL_5__16169_ (
);

FILL SFILL109560x43050 (
);

FILL FILL_1__12717_ (
);

FILL FILL_2__16196_ (
);

FILL FILL_4__10297_ (
);

FILL FILL_3__7821_ (
);

FILL FILL_0__9724_ (
);

FILL FILL_1__15189_ (
);

FILL FILL_5__7747_ (
);

FILL FILL_2_BUFX2_insert810 (
);

FILL FILL_5__7327_ (
);

FILL FILL_2_BUFX2_insert811 (
);

FILL FILL_4__16103_ (
);

FILL FILL_2_BUFX2_insert812 (
);

FILL FILL_2_BUFX2_insert813 (
);

OAI22X1 _14887_ (
    .A(_5367_),
    .B(_3967__bF$buf1),
    .C(_3920_),
    .D(_5368_),
    .Y(_5369_)
);

NOR2X1 _14467_ (
    .A(_4957_),
    .B(_4954_),
    .Y(_4958_)
);

FILL FILL_2_BUFX2_insert814 (
);

NAND3X1 _14047_ (
    .A(_4537_),
    .B(_4538_),
    .C(_4546_),
    .Y(_4547_)
);

FILL FILL_2_BUFX2_insert815 (
);

FILL FILL_2_BUFX2_insert816 (
);

FILL FILL_3__15936_ (
);

FILL FILL_3__15516_ (
);

FILL FILL_2_BUFX2_insert817 (
);

FILL FILL_2_BUFX2_insert818 (
);

FILL FILL_1__16130_ (
);

FILL FILL_2_BUFX2_insert819 (
);

FILL FILL_1__7739_ (
);

FILL FILL_1__7319_ (
);

FILL FILL_3__10651_ (
);

FILL SFILL8600x24050 (
);

FILL FILL_3__10231_ (
);

FILL FILL_2__14929_ (
);

FILL FILL_2__14509_ (
);

FILL FILL_0__15963_ (
);

FILL FILL_0__15543_ (
);

FILL FILL_0__15123_ (
);

FILL FILL_5__12089_ (
);

FILL FILL_3__8606_ (
);

FILL FILL_5__13870_ (
);

FILL FILL_5__13450_ (
);

FILL FILL_5__13030_ (
);

OAI21X1 _7750_ (
    .A(_444_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_445_),
    .Y(_393_[26])
);

OAI21X1 _7330_ (
    .A(_225_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_226_),
    .Y(_198_[14])
);

FILL FILL_4__12863_ (
);

FILL FILL_4__12443_ (
);

FILL FILL_4__12023_ (
);

FILL SFILL13640x25050 (
);

OAI21X1 _10387_ (
    .A(_1775_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1776_),
    .Y(_1758_[9])
);

FILL FILL_3__11856_ (
);

FILL FILL_1__12890_ (
);

FILL FILL_3__11436_ (
);

FILL FILL_1__12470_ (
);

FILL FILL_3__11016_ (
);

FILL FILL_1__12050_ (
);

FILL FILL_4__6949_ (
);

FILL FILL_0__16328_ (
);

FILL SFILL38840x74050 (
);

FILL FILL_2__10429_ (
);

FILL FILL_0__11883_ (
);

FILL FILL_2__9495_ (
);

FILL FILL_2__10009_ (
);

FILL FILL_0__11463_ (
);

FILL FILL_0__11043_ (
);

FILL FILL_5__7080_ (
);

FILL SFILL43800x57050 (
);

FILL SFILL74200x48050 (
);

FILL FILL_5__14655_ (
);

FILL FILL_5__14235_ (
);

FILL FILL_0__6849_ (
);

OAI21X1 _8955_ (
    .A(_1044_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1045_),
    .Y(_1043_[1])
);

DFFSR _8535_ (
    .Q(\datapath_1.regfile_1.regOut[13] [1]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_783_[1])
);

NAND2X1 _8115_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_628_)
);

FILL FILL_1__7492_ (
);

FILL FILL_1__7072_ (
);

FILL FILL_4__13648_ (
);

FILL FILL_4__13228_ (
);

FILL FILL_2__14682_ (
);

FILL FILL_2__14262_ (
);

FILL FILL_2__7808_ (
);

FILL FILL112200x61050 (
);

FILL FILL_1__13675_ (
);

FILL SFILL99480x54050 (
);

FILL FILL_1__13255_ (
);

FILL FILL_1_BUFX2_insert830 (
);

FILL FILL_1_BUFX2_insert831 (
);

FILL FILL_1_BUFX2_insert832 (
);

OAI21X1 _12953_ (
    .A(_3683_),
    .B(vdd),
    .C(_3684_),
    .Y(_3620_[0])
);

NAND2X1 _12533_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [31]),
    .Y(_3422_)
);

FILL FILL_0__12248_ (
);

FILL FILL_1_BUFX2_insert833 (
);

AOI22X1 _12113_ (
    .A(\datapath_1.ALUResult [31]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3131_)
);

FILL FILL_1_BUFX2_insert834 (
);

FILL FILL_1_BUFX2_insert835 (
);

FILL FILL_1_BUFX2_insert836 (
);

FILL FILL_6__16027_ (
);

FILL FILL_1_BUFX2_insert837 (
);

FILL FILL_1_BUFX2_insert838 (
);

FILL FILL_1_BUFX2_insert839 (
);

FILL FILL_3__16054_ (
);

FILL FILL_5__10995_ (
);

FILL FILL112120x68050 (
);

FILL FILL_5__10575_ (
);

FILL FILL_1__8697_ (
);

FILL FILL_5__10155_ (
);

FILL FILL_1__8277_ (
);

FILL FILL_2__15887_ (
);

FILL FILL_2__15467_ (
);

FILL FILL_2__15047_ (
);

FILL FILL_0__16081_ (
);

FILL FILL_2__10182_ (
);

FILL FILL_3__9984_ (
);

FILL FILL_3__9144_ (
);

NOR2X1 _13738_ (
    .A(_4244_),
    .B(_4234_),
    .Y(_4245_)
);

NOR2X1 _13318_ (
    .A(_3781_),
    .B(_3849_),
    .Y(\datapath_1.regfile_1.regEn [12])
);

FILL FILL_1__15821_ (
);

FILL SFILL28840x72050 (
);

FILL FILL_1__15401_ (
);

FILL FILL_6__12367_ (
);

FILL FILL_0__14814_ (
);

FILL FILL_2__7981_ (
);

FILL FILL_2__7561_ (
);

BUFX2 BUFX2_insert500 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf107)
);

FILL SFILL64200x46050 (
);

BUFX2 BUFX2_insert501 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf106)
);

FILL FILL_3__12394_ (
);

BUFX2 BUFX2_insert502 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf105)
);

BUFX2 BUFX2_insert503 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf104)
);

BUFX2 BUFX2_insert504 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf103)
);

FILL FILL_4__7487_ (
);

BUFX2 BUFX2_insert505 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf102)
);

BUFX2 BUFX2_insert506 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf101)
);

FILL FILL_4__7067_ (
);

BUFX2 BUFX2_insert507 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf100)
);

BUFX2 BUFX2_insert508 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf99)
);

FILL FILL_2__11387_ (
);

BUFX2 BUFX2_insert509 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf98)
);

FILL FILL_5__12721_ (
);

FILL FILL_5__12301_ (
);

FILL FILL_4__11714_ (
);

FILL FILL_5__15193_ (
);

FILL FILL_6__8774_ (
);

NAND2X1 _9493_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1323_)
);

DFFSR _9073_ (
    .Q(\datapath_1.regfile_1.regOut[17] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1043_[27])
);

FILL FILL_3__10707_ (
);

FILL FILL_1__11741_ (
);

FILL FILL_4__14186_ (
);

FILL FILL_1__11321_ (
);

FILL FILL_2__8766_ (
);

FILL FILL_3__13599_ (
);

FILL FILL_2__8346_ (
);

FILL FILL_0__10314_ (
);

FILL FILL_0_BUFX2_insert20 (
);

FILL FILL_0_BUFX2_insert21 (
);

FILL FILL_6__14933_ (
);

FILL FILL_6__14513_ (
);

FILL FILL_0_BUFX2_insert22 (
);

FILL SFILL33800x10050 (
);

FILL FILL_0_BUFX2_insert23 (
);

FILL FILL_0_BUFX2_insert24 (
);

FILL FILL_0_BUFX2_insert25 (
);

FILL FILL_0_BUFX2_insert26 (
);

FILL FILL_0_BUFX2_insert27 (
);

INVX1 _13491_ (
    .A(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_4002_)
);

FILL FILL_0_BUFX2_insert28 (
);

DFFSR _13071_ (
    .Q(_2_[24]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3620_[24])
);

FILL FILL_5__13926_ (
);

FILL FILL_0_BUFX2_insert29 (
);

FILL FILL_3__14960_ (
);

FILL FILL_5__13506_ (
);

FILL FILL_3__14540_ (
);

FILL FILL_3__14120_ (
);

OAI21X1 _7806_ (
    .A(_461_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_462_),
    .Y(_458_[2])
);

FILL FILL_4_BUFX2_insert340 (
);

FILL FILL_4__9633_ (
);

FILL FILL_4_BUFX2_insert341 (
);

FILL FILL_4_BUFX2_insert342 (
);

FILL FILL_4__9213_ (
);

FILL FILL_2__13953_ (
);

FILL FILL_4_BUFX2_insert343 (
);

FILL FILL_4_BUFX2_insert344 (
);

FILL FILL_2__13533_ (
);

FILL FILL_5__16398_ (
);

FILL FILL_2__13113_ (
);

FILL FILL_4_BUFX2_insert345 (
);

FILL FILL_6__9979_ (
);

FILL FILL_4_BUFX2_insert346 (
);

FILL FILL_4_BUFX2_insert347 (
);

FILL FILL_4_BUFX2_insert348 (
);

FILL FILL_4_BUFX2_insert349 (
);

FILL FILL_1__12526_ (
);

FILL FILL_1__12106_ (
);

FILL FILL_0__9533_ (
);

FILL FILL_3__7630_ (
);

FILL FILL_0__11939_ (
);

FILL FILL_0__9113_ (
);

FILL FILL_3__7210_ (
);

OAI21X1 _11804_ (
    .A(_2560_),
    .B(_2344__bF$buf3),
    .C(_2895_),
    .Y(_2896_)
);

FILL FILL_0__11519_ (
);

FILL FILL_5__7976_ (
);

FILL FILL_5__7556_ (
);

FILL FILL_4__16332_ (
);

FILL SFILL79880x64050 (
);

INVX1 _14696_ (
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_5182_)
);

INVX1 _14276_ (
    .A(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_4771_)
);

FILL FILL_3__15745_ (
);

FILL FILL_3__15325_ (
);

FILL FILL_1__7968_ (
);

FILL SFILL13720x5050 (
);

FILL FILL_3__10880_ (
);

FILL FILL_1__7548_ (
);

FILL FILL_3__10040_ (
);

FILL FILL_2__14738_ (
);

FILL FILL_2__14318_ (
);

FILL FILL_0__15772_ (
);

FILL FILL_0__15352_ (
);

FILL FILL_3__8835_ (
);

FILL FILL_4__12252_ (
);

NAND2X1 _10196_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1690_)
);

FILL FILL_3__11665_ (
);

FILL FILL_3__11245_ (
);

FILL FILL_0__16137_ (
);

DFFSR _16422_ (
    .Q(\datapath_1.regfile_1.regOut[0] [5]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_6769_[5])
);

OAI22X1 _16002_ (
    .A(_5549__bF$buf4),
    .B(_5040_),
    .C(_5466__bF$buf3),
    .D(_6458_),
    .Y(_6459_)
);

FILL FILL_2__10658_ (
);

FILL FILL_2__10238_ (
);

FILL FILL_0__11692_ (
);

FILL FILL_0__11272_ (
);

FILL FILL_3_BUFX2_insert360 (
);

FILL SFILL23720x15050 (
);

FILL FILL_3_BUFX2_insert361 (
);

FILL FILL_5__14884_ (
);

FILL FILL_3_BUFX2_insert362 (
);

FILL FILL_5__14464_ (
);

FILL FILL_3_BUFX2_insert363 (
);

FILL FILL_5__14044_ (
);

FILL FILL_3_BUFX2_insert364 (
);

NAND2X1 _8764_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_959_)
);

FILL FILL_3_BUFX2_insert365 (
);

NAND2X1 _8344_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_740_)
);

FILL FILL_3_BUFX2_insert366 (
);

FILL FILL_3_BUFX2_insert367 (
);

FILL FILL_3_BUFX2_insert368 (
);

FILL FILL_4__13877_ (
);

FILL FILL_3_BUFX2_insert369 (
);

FILL FILL_4__13457_ (
);

FILL FILL_2__14491_ (
);

FILL FILL_4__13037_ (
);

FILL FILL_2__14071_ (
);

FILL FILL_2__7617_ (
);

FILL FILL_1__13484_ (
);

FILL FILL_0__12897_ (
);

NAND2X1 _12762_ (
    .A(IRWrite_bF$buf5),
    .B(memoryOutData[22]),
    .Y(_3534_)
);

FILL FILL_0__12477_ (
);

FILL FILL_0__12057_ (
);

NAND3X1 _12342_ (
    .A(_3293_),
    .B(_3294_),
    .C(_3295_),
    .Y(\datapath_1.alu_1.ALUInB [31])
);

FILL FILL_3__13811_ (
);

FILL FILL_5__8094_ (
);

FILL FILL_4__8904_ (
);

FILL SFILL13720x58050 (
);

FILL SFILL44120x49050 (
);

FILL FILL_5__15669_ (
);

FILL FILL_5__15249_ (
);

FILL FILL_3__16283_ (
);

DFFSR _9969_ (
    .Q(\datapath_1.regfile_1.regOut[24] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1498_[27])
);

INVX1 _9549_ (
    .A(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_1360_)
);

INVX1 _9129_ (
    .A(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_1141_)
);

FILL FILL_5__10384_ (
);

FILL FILL_1__8086_ (
);

FILL FILL_2__15696_ (
);

FILL FILL_2__15276_ (
);

FILL FILL_3__6901_ (
);

FILL FILL_1__14689_ (
);

FILL FILL_1__14269_ (
);

FILL FILL_0_BUFX2_insert490 (
);

FILL FILL_0_BUFX2_insert491 (
);

FILL FILL_4__15603_ (
);

FILL FILL_0_BUFX2_insert492 (
);

FILL FILL_0_BUFX2_insert493 (
);

FILL FILL_3__9793_ (
);

FILL FILL_0_BUFX2_insert494 (
);

INVX1 _13967_ (
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_4469_)
);

FILL FILL_3__9373_ (
);

FILL FILL_0_BUFX2_insert495 (
);

OAI22X1 _13547_ (
    .A(_3982__bF$buf2),
    .B(_4055_),
    .C(_3971__bF$buf3),
    .D(_4056_),
    .Y(_4057_)
);

FILL FILL_0_BUFX2_insert496 (
);

INVX1 _13127_ (
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_3716_)
);

FILL FILL_0_BUFX2_insert497 (
);

FILL FILL_0_BUFX2_insert498 (
);

FILL FILL_1__15630_ (
);

FILL FILL_5__9299_ (
);

FILL FILL_0_BUFX2_insert499 (
);

FILL FILL_1__15210_ (
);

FILL SFILL8600x19050 (
);

FILL FILL_0__14623_ (
);

FILL FILL_0__14203_ (
);

FILL SFILL13720x13050 (
);

FILL FILL_5__11589_ (
);

FILL FILL_2__7370_ (
);

FILL FILL_5__11169_ (
);

FILL FILL_4__7296_ (
);

FILL FILL_2__11196_ (
);

FILL FILL_5__12530_ (
);

FILL FILL_5__12110_ (
);

FILL FILL_1__10189_ (
);

FILL FILL_4__11943_ (
);

FILL FILL_4__11523_ (
);

FILL FILL_4__11103_ (
);

FILL FILL_0__7196_ (
);

FILL FILL_6__8583_ (
);

FILL FILL_1__16415_ (
);

FILL FILL_3__10936_ (
);

FILL FILL_1__11970_ (
);

FILL FILL_3__10516_ (
);

FILL FILL_1__11550_ (
);

FILL FILL_1__11130_ (
);

FILL FILL_0__15828_ (
);

FILL FILL_0__15408_ (
);

FILL FILL_2__8995_ (
);

FILL FILL_2__8575_ (
);

FILL FILL_0__10963_ (
);

FILL FILL_0__10543_ (
);

FILL FILL_0__10123_ (
);

FILL SFILL3560x61050 (
);

FILL FILL_5__13735_ (
);

FILL FILL_5__13315_ (
);

NAND2X1 _7615_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_376_)
);

FILL FILL_1__6992_ (
);

FILL FILL_4__9862_ (
);

FILL FILL_4__12728_ (
);

FILL FILL_4__9022_ (
);

FILL FILL_2__13762_ (
);

FILL FILL_4__12308_ (
);

FILL FILL_2__13342_ (
);

FILL FILL112200x56050 (
);

FILL SFILL99480x49050 (
);

FILL FILL_1__12755_ (
);

FILL FILL_1__12335_ (
);

FILL FILL_0__9762_ (
);

FILL FILL_0__11748_ (
);

FILL FILL_0__9342_ (
);

INVX1 _11613_ (
    .A(_2718_),
    .Y(\datapath_1.ALUResult [18])
);

FILL FILL_0__11328_ (
);

FILL FILL_5__7365_ (
);

FILL FILL_4__16141_ (
);

FILL FILL_6__10662_ (
);

NAND3X1 _14085_ (
    .A(_4575_),
    .B(_4576_),
    .C(_4583_),
    .Y(_4584_)
);

FILL FILL_3__15974_ (
);

FILL FILL_3__15554_ (
);

FILL FILL_3__15134_ (
);

FILL SFILL28920x60050 (
);

FILL FILL_1__7357_ (
);

FILL SFILL59080x50 (
);

FILL FILL_2__14967_ (
);

FILL FILL_2__14547_ (
);

FILL FILL_2__14127_ (
);

FILL FILL_0__15581_ (
);

FILL FILL_0__15161_ (
);

FILL FILL112200x11050 (
);

FILL FILL_3__8644_ (
);

DFFSR _12818_ (
    .Q(\control_1.op [1]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3490_[27])
);

FILL FILL_3__8224_ (
);

FILL SFILL28840x67050 (
);

FILL FILL_1__14901_ (
);

FILL FILL_4__12481_ (
);

FILL FILL_4__12061_ (
);

FILL FILL_3__16339_ (
);

FILL FILL_5__9931_ (
);

FILL FILL_3__11894_ (
);

FILL FILL_5__9511_ (
);

FILL FILL_3__11474_ (
);

FILL FILL_3__11054_ (
);

FILL FILL112120x18050 (
);

FILL FILL_4__6987_ (
);

FILL FILL_0__16366_ (
);

NAND2X1 _16231_ (
    .A(_6677_),
    .B(_6681_),
    .Y(_6682_)
);

FILL FILL_2__10887_ (
);

FILL FILL_2__10047_ (
);

FILL FILL_0__11081_ (
);

FILL FILL_5__11801_ (
);

FILL FILL_1__9923_ (
);

FILL FILL_1__9503_ (
);

FILL FILL_6__15280_ (
);

FILL FILL_3__9849_ (
);

FILL FILL_3__9429_ (
);

FILL FILL_3__9009_ (
);

FILL FILL_5__14693_ (
);

FILL FILL_5__14273_ (
);

FILL FILL_0__6887_ (
);

NAND2X1 _8993_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1071_)
);

FILL FILL_6__7854_ (
);

NAND2X1 _8573_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_852_)
);

DFFSR _8153_ (
    .Q(\datapath_1.regfile_1.regOut[10] [3]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_588_[3])
);

FILL FILL_4__13686_ (
);

FILL FILL_1__10821_ (
);

FILL SFILL79560x83050 (
);

FILL SFILL28840x22050 (
);

FILL FILL_4__13266_ (
);

FILL FILL_1__10401_ (
);

FILL FILL_2__7846_ (
);

FILL FILL_2__7426_ (
);

FILL FILL_3__12259_ (
);

FILL FILL_1__13293_ (
);

NAND2X1 _12991_ (
    .A(vdd),
    .B(\datapath_1.rd2 [13]),
    .Y(_3646_)
);

NAND2X1 _12571_ (
    .A(vdd),
    .B(memoryOutData[1]),
    .Y(_3427_)
);

FILL FILL_0__12286_ (
);

INVX1 _12151_ (
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_3154_)
);

FILL FILL_3__13620_ (
);

FILL FILL_4__8713_ (
);

FILL FILL_5__15898_ (
);

FILL SFILL103640x74050 (
);

FILL FILL_2__12613_ (
);

FILL FILL_5__15478_ (
);

FILL FILL_5__15058_ (
);

FILL FILL_3__16092_ (
);

INVX1 _9778_ (
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_1472_)
);

INVX1 _9358_ (
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_1253_)
);

FILL FILL_5__10193_ (
);

FILL FILL_1__11606_ (
);

FILL SFILL18840x65050 (
);

FILL FILL_2__15085_ (
);

FILL FILL_0__8613_ (
);

FILL FILL_1__14498_ (
);

FILL FILL_1__14078_ (
);

FILL FILL_4__15832_ (
);

FILL FILL_4__15412_ (
);

INVX1 _13776_ (
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_4282_)
);

NOR2X1 _13356_ (
    .A(_3872_),
    .B(_3871_),
    .Y(\datapath_1.regfile_1.regEn [27])
);

FILL FILL_3__14825_ (
);

FILL FILL_3__14405_ (
);

FILL FILL_4__9918_ (
);

FILL FILL_2__13818_ (
);

FILL FILL_0__14852_ (
);

FILL FILL_0__14432_ (
);

FILL FILL_0__14012_ (
);

CLKBUF1 CLKBUF1_insert1074 (
    .A(clk),
    .Y(clk_hier0_bF$buf9)
);

CLKBUF1 CLKBUF1_insert1075 (
    .A(clk),
    .Y(clk_hier0_bF$buf8)
);

FILL FILL_5__11398_ (
);

CLKBUF1 CLKBUF1_insert1076 (
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

CLKBUF1 CLKBUF1_insert1077 (
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1078 (
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1079 (
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

FILL SFILL18840x20050 (
);

FILL FILL_4__11752_ (
);

FILL FILL_4__11332_ (
);

FILL FILL_1__16224_ (
);

FILL FILL_3__10745_ (
);

FILL FILL_3__10325_ (
);

OAI22X1 _15922_ (
    .A(_4969_),
    .B(_5548__bF$buf3),
    .C(_5489__bF$buf2),
    .D(_6380_),
    .Y(_6381_)
);

FILL FILL_0__15637_ (
);

FILL FILL_0__15217_ (
);

INVX4 _15502_ (
    .A(_5504__bF$buf0),
    .Y(_5971_)
);

FILL FILL_2__8384_ (
);

FILL FILL_0__10772_ (
);

FILL FILL_5__13964_ (
);

FILL FILL_5__13544_ (
);

FILL FILL_5__13124_ (
);

NAND2X1 _7844_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_488_)
);

FILL SFILL69080x74050 (
);

NAND2X1 _7424_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_269_)
);

DFFSR _7004_ (
    .Q(\datapath_1.regfile_1.regOut[1] [6]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_3_[6])
);

FILL FILL_4_BUFX2_insert720 (
);

FILL FILL_4__9671_ (
);

FILL FILL_4_BUFX2_insert721 (
);

FILL FILL_4__9251_ (
);

FILL FILL_4__12957_ (
);

FILL FILL_4_BUFX2_insert722 (
);

FILL FILL_2__13991_ (
);

FILL FILL_4_BUFX2_insert723 (
);

FILL FILL_4_BUFX2_insert724 (
);

FILL FILL_4__12117_ (
);

FILL FILL_2__13571_ (
);

FILL SFILL44200x37050 (
);

FILL FILL_2__13151_ (
);

FILL FILL_4_BUFX2_insert725 (
);

FILL FILL_4_BUFX2_insert726 (
);

FILL FILL_6__9597_ (
);

FILL FILL_4_BUFX2_insert727 (
);

FILL FILL_4_BUFX2_insert728 (
);

FILL FILL_4_BUFX2_insert729 (
);

FILL FILL_1__12984_ (
);

FILL FILL_1__12144_ (
);

FILL FILL_0__9991_ (
);

FILL FILL_0__11977_ (
);

FILL FILL_0__9151_ (
);

NOR2X1 _11842_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(_2128_),
    .Y(_2930_)
);

FILL FILL_2__9169_ (
);

FILL FILL_0__11557_ (
);

NAND2X1 _11422_ (
    .A(_2321_),
    .B(_2481__bF$buf1),
    .Y(_2538_)
);

FILL FILL_0__11137_ (
);

NOR2X1 _11002_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(_2120_),
    .Y(_2121_)
);

FILL FILL_6__15756_ (
);

FILL FILL_5__7594_ (
);

FILL FILL_4__16370_ (
);

FILL FILL_5__7174_ (
);

FILL FILL_6__10051_ (
);

FILL FILL_5__14749_ (
);

FILL FILL_3__15783_ (
);

FILL FILL_5__14329_ (
);

FILL FILL_3__15363_ (
);

INVX1 _8629_ (
    .A(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_889_)
);

INVX1 _8209_ (
    .A(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_670_)
);

FILL FILL_1__7586_ (
);

FILL FILL_1__7166_ (
);

FILL FILL_2__14776_ (
);

FILL FILL_2__14356_ (
);

FILL FILL_0__15390_ (
);

FILL SFILL48920x14050 (
);

FILL FILL_1__13769_ (
);

FILL FILL_1__13349_ (
);

FILL FILL_3__8873_ (
);

FILL FILL_3__8453_ (
);

INVX1 _12627_ (
    .A(\datapath_1.Data [20]),
    .Y(_3464_)
);

OAI21X1 _12207_ (
    .A(_3190_),
    .B(ALUSrcA_bF$buf5),
    .C(_3191_),
    .Y(\datapath_1.alu_1.ALUInA [30])
);

FILL FILL_5__8379_ (
);

FILL FILL_1__14710_ (
);

FILL FILL_6__11676_ (
);

FILL FILL_4__12290_ (
);

AOI22X1 _15099_ (
    .A(\datapath_1.regfile_1.regOut[12] [1]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_5578_)
);

FILL FILL_0__13703_ (
);

FILL FILL_3__16148_ (
);

FILL FILL_5__10669_ (
);

FILL FILL_2__6870_ (
);

FILL FILL_5__10249_ (
);

FILL FILL_5__9740_ (
);

FILL FILL_3__11283_ (
);

FILL FILL_0__16175_ (
);

INVX1 _16040_ (
    .A(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_6496_)
);

FILL FILL_2__10696_ (
);

FILL SFILL38920x57050 (
);

FILL FILL_2__10276_ (
);

FILL FILL_1__9732_ (
);

FILL FILL_5__11610_ (
);

FILL FILL_3__9658_ (
);

FILL FILL_3_BUFX2_insert740 (
);

FILL FILL_3_BUFX2_insert741 (
);

FILL FILL_3__9238_ (
);

FILL FILL_3_BUFX2_insert742 (
);

FILL FILL_3_BUFX2_insert743 (
);

FILL FILL_3_BUFX2_insert744 (
);

FILL FILL_5__14082_ (
);

FILL FILL_1__15915_ (
);

FILL FILL_3_BUFX2_insert745 (
);

INVX1 _8382_ (
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_765_)
);

FILL FILL_3_BUFX2_insert746 (
);

FILL FILL_3_BUFX2_insert747 (
);

FILL FILL_3_BUFX2_insert748 (
);

FILL FILL_3_BUFX2_insert749 (
);

FILL FILL_4__13495_ (
);

FILL FILL_1__10630_ (
);

FILL FILL_0__14908_ (
);

FILL FILL_3__12488_ (
);

FILL FILL_2__7235_ (
);

FILL FILL_3__12068_ (
);

FILL SFILL59000x70050 (
);

FILL FILL_6__13822_ (
);

FILL SFILL3560x56050 (
);

NAND2X1 _12380_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [12]),
    .Y(_3319_)
);

FILL FILL_0__12095_ (
);

FILL SFILL22840x65050 (
);

FILL SFILL38920x12050 (
);

FILL SFILL104440x73050 (
);

FILL FILL_4__8522_ (
);

FILL FILL_4__8102_ (
);

FILL FILL_4__11808_ (
);

FILL FILL_2__12842_ (
);

FILL FILL_2__12422_ (
);

FILL FILL_5__15287_ (
);

FILL FILL_2__12002_ (
);

DFFSR _9587_ (
    .Q(\datapath_1.regfile_1.regOut[21] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1303_[29])
);

OAI21X1 _9167_ (
    .A(_1165_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .C(_1166_),
    .Y(_1108_[29])
);

FILL FILL_1__11835_ (
);

FILL FILL_1__11415_ (
);

FILL FILL_0__8842_ (
);

FILL FILL_0__10828_ (
);

FILL FILL_0__10408_ (
);

FILL FILL_0__8002_ (
);

FILL SFILL38840x19050 (
);

FILL FILL_5__6865_ (
);

FILL FILL_0_BUFX2_insert870 (
);

FILL FILL_4__15641_ (
);

FILL FILL_0_BUFX2_insert871 (
);

FILL FILL_4__15221_ (
);

FILL FILL_0_BUFX2_insert872 (
);

FILL FILL_0_BUFX2_insert873 (
);

FILL FILL_0_BUFX2_insert874 (
);

INVX1 _13585_ (
    .A(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_4094_)
);

FILL FILL_0_BUFX2_insert875 (
);

OAI21X1 _13165_ (
    .A(_3740_),
    .B(PCEn_bF$buf7),
    .C(_3741_),
    .Y(_3685_[28])
);

FILL FILL_0_BUFX2_insert876 (
);

FILL FILL_0_BUFX2_insert877 (
);

FILL FILL_2__9801_ (
);

FILL FILL_3__14634_ (
);

FILL FILL_0_BUFX2_insert878 (
);

FILL FILL_3__14214_ (
);

FILL FILL_0_BUFX2_insert879 (
);

FILL SFILL28920x55050 (
);

FILL SFILL3560x11050 (
);

FILL FILL_1__6857_ (
);

FILL FILL_4__9727_ (
);

FILL FILL_2__13627_ (
);

FILL FILL_2__13207_ (
);

FILL FILL_0__14661_ (
);

FILL FILL_0__14241_ (
);

FILL FILL_2__16099_ (
);

FILL FILL_0__9627_ (
);

FILL FILL_3__7724_ (
);

FILL FILL_3__7304_ (
);

FILL FILL_0__9207_ (
);

FILL FILL_4__16006_ (
);

FILL FILL_4__11981_ (
);

FILL FILL_6__10527_ (
);

FILL FILL_4__11561_ (
);

FILL FILL_4__11141_ (
);

FILL FILL_3__15839_ (
);

FILL FILL_3__15419_ (
);

FILL FILL_1__16033_ (
);

FILL FILL_3__10974_ (
);

FILL FILL_3__10554_ (
);

FILL FILL_3__10134_ (
);

FILL SFILL28920x10050 (
);

FILL FILL_0__15866_ (
);

FILL FILL_6_BUFX2_insert254 (
);

NOR3X1 _15731_ (
    .A(_6172_),
    .B(_6184_),
    .C(_6194_),
    .Y(_6195_)
);

FILL FILL_0__15446_ (
);

NOR2X1 _15311_ (
    .A(_5509_),
    .B(_5688_),
    .Y(_5785_)
);

FILL FILL_0__15026_ (
);

FILL FILL_2__8193_ (
);

FILL FILL_0__10581_ (
);

FILL FILL_0__10161_ (
);

BUFX2 BUFX2_insert30 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf3 )
);

BUFX2 BUFX2_insert31 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf2 )
);

FILL FILL_6__14360_ (
);

BUFX2 BUFX2_insert32 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf1 )
);

BUFX2 BUFX2_insert33 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf0 )
);

BUFX2 BUFX2_insert34 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf7 )
);

BUFX2 BUFX2_insert35 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf6 )
);

FILL FILL_3__8509_ (
);

BUFX2 BUFX2_insert36 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf5 )
);

FILL FILL_5__13773_ (
);

BUFX2 BUFX2_insert37 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf4 )
);

FILL FILL_5__13353_ (
);

BUFX2 BUFX2_insert38 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf3 )
);

BUFX2 BUFX2_insert39 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf2 )
);

FILL FILL_6__6934_ (
);

DFFSR _7653_ (
    .Q(\datapath_1.regfile_1.regOut[6] [15]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_328_[15])
);

INVX1 _7233_ (
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_182_)
);

FILL FILL_4__9480_ (
);

FILL FILL_4__12766_ (
);

FILL FILL_4__12346_ (
);

FILL FILL_2__13380_ (
);

FILL SFILL114600x1050 (
);

FILL FILL_2__6926_ (
);

FILL FILL_3__11759_ (
);

FILL FILL_3__11339_ (
);

FILL FILL_1__12373_ (
);

FILL SFILL18920x53050 (
);

FILL FILL_0__9380_ (
);

FILL FILL_2__9398_ (
);

FILL FILL_0__11786_ (
);

FILL FILL_0__11366_ (
);

INVX1 _11651_ (
    .A(_2400_),
    .Y(_2754_)
);

INVX1 _11231_ (
    .A(_2114_),
    .Y(_2350_)
);

FILL FILL_3__12700_ (
);

FILL SFILL94760x53050 (
);

FILL FILL_5__14978_ (
);

FILL FILL_5__14558_ (
);

FILL FILL_5__14138_ (
);

FILL FILL_3__15592_ (
);

INVX1 _8858_ (
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_1001_)
);

FILL FILL_3__15172_ (
);

INVX1 _8438_ (
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_846_)
);

OAI21X1 _8018_ (
    .A(_582_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .C(_583_),
    .Y(_523_[30])
);

FILL FILL_2__14585_ (
);

FILL FILL_2__14165_ (
);

FILL FILL_1__13998_ (
);

FILL FILL_1__13578_ (
);

FILL FILL_1__13158_ (
);

FILL FILL_4__14912_ (
);

INVX1 _12856_ (
    .A(\datapath_1.a [11]),
    .Y(_3576_)
);

FILL FILL_3__8262_ (
);

INVX1 _12436_ (
    .A(ALUOut[31]),
    .Y(_3356_)
);

NAND3X1 _12016_ (
    .A(PCSource_1_bF$buf0),
    .B(\aluControl_1.inst [5]),
    .C(_3034__bF$buf0),
    .Y(_3058_)
);

FILL FILL_3__13905_ (
);

FILL FILL_5__8188_ (
);

FILL FILL_5_BUFX2_insert270 (
);

FILL FILL_5_BUFX2_insert271 (
);

FILL FILL_5_BUFX2_insert272 (
);

FILL FILL_0__13932_ (
);

FILL FILL_5_BUFX2_insert273 (
);

FILL FILL_3__16377_ (
);

FILL FILL_0__13512_ (
);

FILL FILL_5_BUFX2_insert274 (
);

FILL FILL_5__10898_ (
);

FILL FILL_5_BUFX2_insert275 (
);

FILL FILL_5_BUFX2_insert276 (
);

FILL FILL_5__10058_ (
);

FILL FILL_5_BUFX2_insert277 (
);

FILL FILL_5_BUFX2_insert1060 (
);

FILL FILL_5_BUFX2_insert278 (
);

FILL FILL_5_BUFX2_insert1061 (
);

FILL FILL_3__11092_ (
);

FILL FILL_5_BUFX2_insert1062 (
);

FILL FILL_5_BUFX2_insert279 (
);

FILL FILL_5_BUFX2_insert1063 (
);

FILL FILL_5_BUFX2_insert1064 (
);

FILL FILL_5_BUFX2_insert1065 (
);

FILL FILL_5_BUFX2_insert1066 (
);

FILL SFILL18840x15050 (
);

FILL FILL_5_BUFX2_insert1067 (
);

FILL SFILL84360x82050 (
);

FILL FILL_5_BUFX2_insert1068 (
);

FILL FILL_5_BUFX2_insert1069 (
);

FILL FILL_1__9541_ (
);

FILL FILL_1__9121_ (
);

FILL FILL_2__16311_ (
);

FILL FILL_3__9887_ (
);

FILL FILL_3__9467_ (
);

FILL FILL_4__10832_ (
);

FILL FILL_4__10412_ (
);

FILL FILL_1__15724_ (
);

FILL FILL_6__7472_ (
);

INVX1 _8191_ (
    .A(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_658_)
);

FILL FILL_1__15304_ (
);

FILL FILL_0__14717_ (
);

FILL FILL_2__7884_ (
);

FILL FILL_2__7464_ (
);

FILL FILL_2__7044_ (
);

FILL FILL_3__12297_ (
);

FILL FILL_5__12624_ (
);

FILL SFILL99400x4050 (
);

FILL FILL_5__12204_ (
);

NAND2X1 _6924_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_17_)
);

FILL FILL_4__8751_ (
);

FILL SFILL99320x9050 (
);

FILL FILL_4__8331_ (
);

FILL FILL_4__11617_ (
);

FILL FILL_2__12651_ (
);

FILL FILL_2__12231_ (
);

FILL FILL_5__15096_ (
);

OAI21X1 _9396_ (
    .A(_1277_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .C(_1278_),
    .Y(_1238_[20])
);

FILL FILL_6__8257_ (
);

FILL SFILL110280x12050 (
);

FILL FILL_1__11644_ (
);

FILL FILL_1__11224_ (
);

FILL FILL_4__14089_ (
);

FILL FILL_0__8651_ (
);

FILL FILL_0__10637_ (
);

FILL FILL_2__8249_ (
);

AND2X2 _10922_ (
    .A(_2061_),
    .B(_2059_),
    .Y(RegWrite)
);

FILL FILL_0__8231_ (
);

FILL SFILL114520x63050 (
);

NAND2X1 _10502_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1833_)
);

FILL FILL_4__15870_ (
);

FILL FILL_6__14416_ (
);

FILL FILL_4__15450_ (
);

FILL FILL_4__15030_ (
);

OAI22X1 _13394_ (
    .A(_3905__bF$buf1),
    .B(_3896_),
    .C(_3902__bF$buf1),
    .D(_3897_),
    .Y(_3906_)
);

FILL FILL_5__13829_ (
);

FILL FILL_2__9610_ (
);

FILL FILL_3__14863_ (
);

FILL FILL_5__13409_ (
);

FILL FILL_3__14443_ (
);

FILL FILL_3__14023_ (
);

INVX1 _7709_ (
    .A(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_418_)
);

FILL FILL_4__9536_ (
);

FILL FILL_4__9116_ (
);

FILL SFILL69080x24050 (
);

FILL FILL_2__13856_ (
);

FILL FILL_2__13436_ (
);

FILL FILL_0__14890_ (
);

FILL FILL_0__14470_ (
);

FILL FILL_2__13016_ (
);

FILL FILL_0__14050_ (
);

FILL FILL_1__12849_ (
);

FILL FILL_1__12429_ (
);

FILL FILL_1__12009_ (
);

FILL FILL_0__9856_ (
);

FILL FILL_3__7953_ (
);

FILL FILL_0__9016_ (
);

FILL FILL_3__7113_ (
);

OAI21X1 _11707_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .C(_2347__bF$buf3),
    .Y(_2806_)
);

FILL FILL_5__7879_ (
);

FILL FILL_5__7459_ (
);

FILL FILL_5__7039_ (
);

FILL FILL_4__16235_ (
);

INVX1 _14599_ (
    .A(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_5087_)
);

FILL FILL_4__11790_ (
);

NOR3X1 _14179_ (
    .A(_4673_),
    .B(_4671_),
    .C(_4675_),
    .Y(_4676_)
);

FILL FILL_4__11370_ (
);

FILL FILL_3__15648_ (
);

FILL FILL_3__15228_ (
);

FILL FILL_1__16262_ (
);

FILL FILL_3__10783_ (
);

FILL FILL_5__8400_ (
);

FILL FILL_3__10363_ (
);

FILL SFILL59080x67050 (
);

FILL FILL_0__15675_ (
);

INVX1 _15960_ (
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_6418_)
);

FILL FILL_0__15255_ (
);

OAI22X1 _15540_ (
    .A(_5549__bF$buf3),
    .B(_4556_),
    .C(_5466__bF$buf2),
    .D(_4528_),
    .Y(_6008_)
);

NAND3X1 _15120_ (
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .B(_5471__bF$buf4),
    .C(_5531__bF$buf3),
    .Y(_5599_)
);

FILL FILL_0__10390_ (
);

FILL FILL_3__8738_ (
);

FILL FILL_3__8318_ (
);

FILL FILL_5__13582_ (
);

FILL FILL_5__13162_ (
);

INVX1 _7882_ (
    .A(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_513_)
);

INVX1 _7462_ (
    .A(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_294_)
);

INVX1 _7042_ (
    .A(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_75_)
);

FILL SFILL43880x51050 (
);

FILL FILL_4__12995_ (
);

FILL FILL_4__12575_ (
);

FILL FILL_4__12155_ (
);

DFFSR _10099_ (
    .Q(\datapath_1.regfile_1.regOut[25] [29]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_1563_[29])
);

FILL FILL_3__11988_ (
);

FILL FILL_3__11568_ (
);

FILL FILL_5__9605_ (
);

FILL FILL_3__11148_ (
);

FILL SFILL59000x65050 (
);

FILL FILL_1__12182_ (
);

NAND2X1 _16325_ (
    .A(gnd),
    .B(gnd),
    .Y(_6771_)
);

FILL SFILL59080x22050 (
);

OAI21X1 _11880_ (
    .A(_2962_),
    .B(RegDst),
    .C(_2963_),
    .Y(\datapath_1.a3 [2])
);

FILL FILL_0__11595_ (
);

FILL FILL_0__11175_ (
);

OAI21X1 _11460_ (
    .A(_2574_),
    .B(_2308_),
    .C(_2289_),
    .Y(_2575_)
);

AOI21X1 _11040_ (
    .A(_2156_),
    .B(_2154_),
    .C(_2158_),
    .Y(_2159_)
);

FILL SFILL104440x68050 (
);

FILL FILL_4__7602_ (
);

FILL FILL_2__11922_ (
);

FILL FILL_5__14787_ (
);

FILL FILL_5__14367_ (
);

FILL FILL_2__11502_ (
);

FILL FILL_6__7948_ (
);

DFFSR _8667_ (
    .Q(\datapath_1.regfile_1.regOut[14] [5]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_848_[5])
);

OAI21X1 _8247_ (
    .A(_694_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .C(_695_),
    .Y(_653_[21])
);

FILL FILL_1__10915_ (
);

FILL FILL_2__14394_ (
);

FILL FILL_0__7502_ (
);

FILL FILL_1__13387_ (
);

FILL FILL_4__14721_ (
);

FILL FILL_4__14301_ (
);

FILL SFILL59000x20050 (
);

FILL SFILL43960x9050 (
);

FILL FILL_3__8491_ (
);

FILL SFILL49080x65050 (
);

DFFSR _12665_ (
    .Q(\datapath_1.Data [2]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3425_[2])
);

FILL FILL_3__8071_ (
);

AOI22X1 _12245_ (
    .A(_2_[7]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf1),
    .D(\aluControl_1.inst [5]),
    .Y(_3223_)
);

FILL FILL_3__13714_ (
);

FILL SFILL73560x76050 (
);

FILL FILL_2__12707_ (
);

FILL FILL_0__13741_ (
);

FILL FILL_0__13321_ (
);

FILL FILL_3__16186_ (
);

FILL FILL_5__10287_ (
);

FILL FILL_2__15599_ (
);

FILL FILL_2__15179_ (
);

FILL FILL_0__8707_ (
);

FILL FILL_1__9770_ (
);

FILL FILL_1__9350_ (
);

FILL FILL_4__15926_ (
);

FILL FILL_4__15506_ (
);

FILL FILL_2__16120_ (
);

FILL SFILL49000x63050 (
);

FILL FILL_3__9276_ (
);

FILL FILL_4__10641_ (
);

FILL FILL_3__14919_ (
);

FILL FILL_1__15953_ (
);

FILL FILL_1__15533_ (
);

FILL FILL_1__15113_ (
);

FILL SFILL94440x72050 (
);

FILL FILL_0__14946_ (
);

NAND3X1 _14811_ (
    .A(_5286_),
    .B(_5287_),
    .C(_5294_),
    .Y(_5295_)
);

FILL FILL_0__14526_ (
);

FILL FILL_0__14106_ (
);

FILL FILL_2__7693_ (
);

FILL FILL_4__7199_ (
);

FILL FILL_2__11099_ (
);

FILL FILL_5__12853_ (
);

FILL FILL_5__12433_ (
);

FILL FILL_5__12013_ (
);

FILL FILL_4__8980_ (
);

FILL SFILL94360x79050 (
);

FILL FILL_4__8140_ (
);

FILL FILL_4__11846_ (
);

FILL FILL_2__12880_ (
);

FILL FILL_4__11426_ (
);

FILL FILL_2__12460_ (
);

FILL FILL_4__11006_ (
);

FILL FILL_2__12040_ (
);

FILL FILL_0__7099_ (
);

FILL FILL_1__16318_ (
);

FILL FILL_1__11873_ (
);

FILL FILL_3__10419_ (
);

FILL FILL_1__11453_ (
);

FILL FILL_1__11033_ (
);

FILL FILL_0__8880_ (
);

FILL FILL_2__8898_ (
);

FILL FILL_0__8460_ (
);

FILL FILL_2__8478_ (
);

DFFSR _10731_ (
    .Q(\datapath_1.regfile_1.regOut[30] [21]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1888_[21])
);

FILL FILL_0__10446_ (
);

FILL FILL_2__8058_ (
);

INVX1 _10311_ (
    .A(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_1746_)
);

FILL FILL_0__10026_ (
);

FILL FILL_5__13638_ (
);

FILL FILL_5__13218_ (
);

FILL FILL_3__14672_ (
);

FILL FILL_3__14252_ (
);

INVX1 _7938_ (
    .A(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_530_)
);

DFFSR _7518_ (
    .Q(\datapath_1.regfile_1.regOut[5] [8]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_263_[8])
);

FILL FILL_1__6895_ (
);

FILL FILL_4__9765_ (
);

FILL FILL_4__9345_ (
);

FILL FILL_2__13665_ (
);

FILL FILL_2__13245_ (
);

FILL SFILL63960x43050 (
);

FILL SFILL39000x61050 (
);

FILL FILL_1__12658_ (
);

FILL FILL_1__12238_ (
);

FILL FILL_3__7762_ (
);

FILL FILL_0__9665_ (
);

NAND2X1 _11936_ (
    .A(IorD_bF$buf0),
    .B(ALUOut[16]),
    .Y(_2999_)
);

FILL FILL_3__7342_ (
);

FILL FILL_0__9245_ (
);

INVX1 _11516_ (
    .A(_2627_),
    .Y(\datapath_1.ALUResult [24])
);

FILL FILL_5__7688_ (
);

FILL SFILL79160x14050 (
);

FILL FILL_4__16044_ (
);

FILL FILL_6__10145_ (
);

FILL FILL_3__15877_ (
);

FILL FILL_3__15457_ (
);

FILL FILL_3__15037_ (
);

FILL FILL_1__16071_ (
);

FILL FILL_3__10172_ (
);

FILL FILL_6_BUFX2_insert633 (
);

FILL FILL_0__15484_ (
);

FILL FILL_0__15064_ (
);

FILL FILL_6_BUFX2_insert638 (
);

FILL FILL_1__8621_ (
);

FILL FILL_1__8201_ (
);

FILL FILL_2__15811_ (
);

FILL FILL_3__8967_ (
);

FILL SFILL79080x9050 (
);

FILL FILL_3__8127_ (
);

FILL FILL_5__13391_ (
);

INVX1 _7691_ (
    .A(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_406_)
);

FILL FILL_1__14804_ (
);

FILL SFILL53560x72050 (
);

FILL FILL_1_BUFX2_insert90 (
);

DFFSR _7271_ (
    .Q(\datapath_1.regfile_1.regOut[3] [17]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_133_[17])
);

FILL FILL_1_BUFX2_insert91 (
);

FILL FILL_1_BUFX2_insert92 (
);

FILL FILL_1_BUFX2_insert93 (
);

FILL FILL_4__12384_ (
);

FILL FILL_1_BUFX2_insert94 (
);

FILL FILL_1_BUFX2_insert95 (
);

FILL SFILL8760x51050 (
);

FILL SFILL78440x6050 (
);

FILL FILL_1_BUFX2_insert96 (
);

FILL FILL_1_BUFX2_insert97 (
);

FILL FILL_1_BUFX2_insert98 (
);

FILL FILL_1_BUFX2_insert99 (
);

FILL FILL_2__6964_ (
);

FILL FILL_3__11797_ (
);

FILL FILL_5__9414_ (
);

FILL FILL_3__11377_ (
);

FILL FILL_0__16269_ (
);

OAI22X1 _16134_ (
    .A(_5569_),
    .B(_5235_),
    .C(_5483__bF$buf0),
    .D(_5264_),
    .Y(_6587_)
);

FILL SFILL114600x51050 (
);

FILL FILL_5__11704_ (
);

FILL SFILL53960x41050 (
);

FILL FILL_1__9406_ (
);

FILL FILL_6__15183_ (
);

FILL FILL_4__7831_ (
);

FILL FILL_5__14596_ (
);

FILL FILL_2__11731_ (
);

FILL FILL_5__14176_ (
);

FILL FILL_2__11311_ (
);

OAI21X1 _8896_ (
    .A(_1025_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .C(_1026_),
    .Y(_978_[24])
);

OAI21X1 _8476_ (
    .A(_806_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .C(_807_),
    .Y(_783_[12])
);

FILL FILL_6__7337_ (
);

OAI21X1 _8056_ (
    .A(_651_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .C(_652_),
    .Y(_588_[0])
);

FILL FILL_4__13589_ (
);

FILL FILL_1__10304_ (
);

FILL FILL_4__13169_ (
);

FILL FILL_0__7731_ (
);

FILL FILL_2__7749_ (
);

FILL FILL_0__7311_ (
);

FILL FILL_2__7329_ (
);

FILL SFILL53880x48050 (
);

FILL FILL_4__14950_ (
);

FILL FILL_4__14530_ (
);

FILL SFILL3720x77050 (
);

FILL FILL_4__14110_ (
);

OAI21X1 _12894_ (
    .A(_3600_),
    .B(vdd),
    .C(_3601_),
    .Y(_3555_[23])
);

FILL FILL_0__12189_ (
);

OAI21X1 _12474_ (
    .A(_3381_),
    .B(vdd),
    .C(_3382_),
    .Y(_3360_[11])
);

NAND3X1 _12054_ (
    .A(_3084_),
    .B(_3085_),
    .C(_3086_),
    .Y(\datapath_1.mux_pcsrc.dout [16])
);

FILL FILL_5__12909_ (
);

FILL FILL_3__13943_ (
);

FILL FILL_3__13523_ (
);

FILL FILL_3__13103_ (
);

FILL FILL_4__8616_ (
);

FILL SFILL69080x19050 (
);

FILL FILL_5_BUFX2_insert650 (
);

FILL FILL_5_BUFX2_insert651 (
);

FILL FILL_5_BUFX2_insert652 (
);

FILL FILL_2__12516_ (
);

FILL FILL_0__13970_ (
);

FILL FILL_5_BUFX2_insert653 (
);

FILL FILL_0__13550_ (
);

FILL FILL_5_BUFX2_insert654 (
);

FILL FILL_0__13130_ (
);

FILL FILL_5_BUFX2_insert655 (
);

FILL FILL_5_BUFX2_insert656 (
);

FILL FILL_5_BUFX2_insert657 (
);

FILL FILL_5_BUFX2_insert658 (
);

FILL FILL_1__11929_ (
);

FILL FILL_5_BUFX2_insert659 (
);

FILL FILL_1__11509_ (
);

FILL FILL_5__16322_ (
);

FILL FILL_0__8516_ (
);

FILL FILL_5__6959_ (
);

FILL FILL_4__15735_ (
);

FILL SFILL114520x13050 (
);

FILL FILL_4__15315_ (
);

INVX1 _13679_ (
    .A(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_4187_)
);

FILL FILL_4__10870_ (
);

FILL FILL_3__9085_ (
);

OAI21X1 _13259_ (
    .A(_3801_),
    .B(_3797_),
    .C(_3798_),
    .Y(_3802_)
);

FILL FILL_4__10450_ (
);

FILL FILL_4__10030_ (
);

FILL SFILL3720x32050 (
);

FILL FILL_3__14728_ (
);

FILL FILL_3__14308_ (
);

FILL FILL_1__15762_ (
);

FILL FILL_1__15342_ (
);

FILL FILL_0__14755_ (
);

INVX1 _14620_ (
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_5108_)
);

FILL FILL_0__14335_ (
);

OAI22X1 _14200_ (
    .A(_4696_),
    .B(_3941_),
    .C(_3960_),
    .D(_4695_),
    .Y(_4697_)
);

FILL FILL_2__7082_ (
);

FILL FILL_3__7818_ (
);

FILL SFILL3640x39050 (
);

FILL FILL_5__12662_ (
);

FILL FILL_5__12242_ (
);

INVX1 _6962_ (
    .A(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_42_)
);

FILL FILL_2_BUFX2_insert780 (
);

FILL SFILL104520x56050 (
);

FILL FILL_2_BUFX2_insert781 (
);

FILL SFILL48920x1050 (
);

FILL FILL_2_BUFX2_insert782 (
);

FILL FILL_2_BUFX2_insert783 (
);

FILL FILL_2_BUFX2_insert784 (
);

FILL FILL_4__11655_ (
);

FILL FILL_2_BUFX2_insert785 (
);

FILL FILL_4__11235_ (
);

FILL FILL_2_BUFX2_insert786 (
);

FILL SFILL48840x6050 (
);

FILL FILL_2_BUFX2_insert787 (
);

FILL FILL_2_BUFX2_insert788 (
);

FILL FILL_2_BUFX2_insert789 (
);

FILL FILL_1__16127_ (
);

FILL FILL_3__10648_ (
);

FILL FILL_1__11682_ (
);

FILL FILL_1__11262_ (
);

NOR2X1 _15825_ (
    .A(_6285_),
    .B(_6280_),
    .Y(_6286_)
);

NOR2X1 _15405_ (
    .A(_5876_),
    .B(_5873_),
    .Y(_5877_)
);

FILL SFILL43480x32050 (
);

FILL SFILL59080x17050 (
);

FILL FILL112280x50050 (
);

NAND2X1 _10960_ (
    .A(_2064_),
    .B(_2085_),
    .Y(_2092_)
);

FILL FILL_0__10675_ (
);

FILL FILL_0__10255_ (
);

INVX1 _10540_ (
    .A(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_1858_)
);

INVX1 _10120_ (
    .A(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_1639_)
);

FILL FILL_5__13867_ (
);

FILL FILL_5__13447_ (
);

FILL FILL_3__14481_ (
);

FILL FILL_5__13027_ (
);

FILL FILL_3__14061_ (
);

OAI21X1 _7747_ (
    .A(_442_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .C(_443_),
    .Y(_393_[25])
);

OAI21X1 _7327_ (
    .A(_223_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .C(_224_),
    .Y(_198_[13])
);

FILL FILL_4__9994_ (
);

FILL FILL_4__9154_ (
);

FILL FILL_2__13894_ (
);

FILL FILL_2__13474_ (
);

FILL SFILL104520x11050 (
);

FILL FILL_1__12887_ (
);

FILL FILL_1__12467_ (
);

FILL FILL_1__12047_ (
);

FILL FILL_4__13801_ (
);

FILL SFILL28600x24050 (
);

FILL FILL_3__7991_ (
);

FILL FILL_0__9894_ (
);

FILL FILL_0__9474_ (
);

FILL FILL_3__7571_ (
);

NAND2X1 _11745_ (
    .A(_2197_),
    .B(_2388_),
    .Y(_2841_)
);

NOR2X1 _11325_ (
    .A(_2443_),
    .B(_2441_),
    .Y(_2444_)
);

FILL FILL_6__15659_ (
);

FILL FILL_6__15239_ (
);

FILL FILL_5__7497_ (
);

FILL FILL_5__7077_ (
);

FILL FILL_4__16273_ (
);

FILL FILL_3__15686_ (
);

FILL FILL_0__12401_ (
);

FILL FILL_3__15266_ (
);

FILL FILL_1__7489_ (
);

FILL FILL_1__7069_ (
);

FILL FILL_2__14679_ (
);

FILL FILL_2__14259_ (
);

FILL FILL_0__15293_ (
);

FILL SFILL108760x26050 (
);

FILL FILL_1__8850_ (
);

FILL FILL_1__8010_ (
);

FILL FILL_2__15620_ (
);

FILL SFILL49000x58050 (
);

FILL FILL_2__15200_ (
);

FILL FILL_3__8776_ (
);

FILL FILL_3__8356_ (
);

FILL SFILL49080x15050 (
);

FILL FILL_1__14613_ (
);

OAI21X1 _7080_ (
    .A(_99_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_100_),
    .Y(_68_[16])
);

FILL FILL_6__11579_ (
);

FILL FILL_6__11159_ (
);

FILL SFILL94440x67050 (
);

FILL FILL_4__12193_ (
);

FILL FILL_0__13606_ (
);

FILL FILL_5__9643_ (
);

FILL FILL_5__9223_ (
);

FILL FILL_3__11186_ (
);

FILL FILL_6__12520_ (
);

FILL SFILL49400x27050 (
);

INVX1 _16363_ (
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_6796_)
);

FILL FILL_0__16078_ (
);

FILL FILL_2__10179_ (
);

FILL FILL_5__11933_ (
);

FILL FILL_1__9635_ (
);

FILL FILL_5__11513_ (
);

FILL FILL_1__9215_ (
);

FILL FILL_2__16405_ (
);

FILL FILL_4__10926_ (
);

FILL FILL_4__7220_ (
);

FILL FILL_2__11960_ (
);

FILL FILL_4__10506_ (
);

FILL FILL_2__11540_ (
);

FILL FILL_2__11120_ (
);

FILL SFILL49000x13050 (
);

FILL FILL_1__15818_ (
);

DFFSR _8285_ (
    .Q(\datapath_1.regfile_1.regOut[11] [7]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_653_[7])
);

FILL FILL_1__10953_ (
);

FILL FILL_1__10533_ (
);

FILL FILL_4__13398_ (
);

FILL FILL_1__10113_ (
);

FILL FILL_0__7960_ (
);

FILL FILL_2__7978_ (
);

FILL SFILL94440x22050 (
);

BUFX2 BUFX2_insert470 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf1 )
);

FILL FILL_2__7558_ (
);

BUFX2 BUFX2_insert471 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf0 )
);

FILL FILL_0__7120_ (
);

BUFX2 BUFX2_insert472 (
    .A(_5521_),
    .Y(_5521__bF$buf3)
);

BUFX2 BUFX2_insert473 (
    .A(_5521_),
    .Y(_5521__bF$buf2)
);

BUFX2 BUFX2_insert474 (
    .A(_5521_),
    .Y(_5521__bF$buf1)
);

FILL FILL_6__13725_ (
);

FILL SFILL18840x5050 (
);

BUFX2 BUFX2_insert475 (
    .A(_5521_),
    .Y(_5521__bF$buf0)
);

BUFX2 BUFX2_insert476 (
    .A(_5518_),
    .Y(_5518__bF$buf3)
);

BUFX2 BUFX2_insert477 (
    .A(_5518_),
    .Y(_5518__bF$buf2)
);

BUFX2 BUFX2_insert478 (
    .A(_5518_),
    .Y(_5518__bF$buf1)
);

BUFX2 BUFX2_insert479 (
    .A(_5518_),
    .Y(_5518__bF$buf0)
);

NAND3X1 _12283_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3251_)
);

FILL FILL_5__12718_ (
);

FILL SFILL23880x42050 (
);

FILL FILL_3__13752_ (
);

FILL FILL_3__13332_ (
);

FILL FILL_4__8845_ (
);

FILL SFILL4120x62050 (
);

FILL FILL_4__8005_ (
);

FILL FILL_2__12745_ (
);

FILL FILL_2__12325_ (
);

FILL SFILL94360x29050 (
);

FILL FILL_1__11738_ (
);

FILL FILL_1__11318_ (
);

FILL FILL_3__6842_ (
);

FILL FILL_5__16131_ (
);

FILL FILL_0__8745_ (
);

FILL FILL_0__8325_ (
);

FILL FILL_4__15964_ (
);

FILL FILL_4__15544_ (
);

FILL FILL_4__15124_ (
);

AOI22X1 _13488_ (
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .B(_3998__bF$buf0),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_3999_)
);

DFFSR _13068_ (
    .Q(_2_[21]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3620_[21])
);

FILL FILL_3__14957_ (
);

FILL FILL_1__15991_ (
);

FILL FILL_3__14537_ (
);

FILL SFILL44280x76050 (
);

FILL FILL_1__15571_ (
);

FILL FILL_3__14117_ (
);

FILL FILL_1__15151_ (
);

FILL FILL_0__14984_ (
);

FILL FILL_0__14564_ (
);

FILL FILL_0__14144_ (
);

FILL FILL111800x13050 (
);

FILL SFILL39000x11050 (
);

FILL FILL_1__7701_ (
);

FILL FILL_3__7627_ (
);

FILL FILL_3__7207_ (
);

FILL FILL_5__12891_ (
);

FILL FILL_5__12471_ (
);

FILL FILL_5__12051_ (
);

FILL FILL_4__16329_ (
);

FILL FILL_4__11884_ (
);

FILL FILL_4__11464_ (
);

FILL SFILL8760x46050 (
);

FILL FILL_4__11044_ (
);

FILL SFILL13800x83050 (
);

FILL FILL_1__16356_ (
);

FILL FILL_3__10877_ (
);

FILL FILL_5__8914_ (
);

FILL FILL_3__10037_ (
);

FILL FILL_1__11491_ (
);

FILL FILL_1__11071_ (
);

FILL FILL_0__15769_ (
);

FILL FILL_0__15349_ (
);

NOR2X1 _15634_ (
    .A(_6098_),
    .B(_6099_),
    .Y(_6100_)
);

NOR2X1 _15214_ (
    .A(_4161_),
    .B(_5549__bF$buf4),
    .Y(_5690_)
);

FILL FILL_2__8096_ (
);

FILL FILL_0__10064_ (
);

FILL SFILL53960x36050 (
);

FILL FILL_1__8906_ (
);

FILL SFILL84360x27050 (
);

FILL FILL_4__6911_ (
);

FILL FILL_2__10811_ (
);

FILL FILL_5__13676_ (
);

FILL FILL_5__13256_ (
);

OAI21X1 _7976_ (
    .A(_554_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .C(_555_),
    .Y(_523_[16])
);

FILL FILL_6__6837_ (
);

FILL FILL_3__14290_ (
);

OAI21X1 _7556_ (
    .A(_335_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_336_),
    .Y(_328_[4])
);

DFFSR _7136_ (
    .Q(\datapath_1.regfile_1.regOut[2] [10]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_68_[10])
);

FILL FILL_4__9383_ (
);

FILL FILL_4__12249_ (
);

FILL FILL_2__13283_ (
);

FILL FILL_1__12696_ (
);

FILL FILL_1__12276_ (
);

FILL FILL_4__13610_ (
);

DFFSR _16419_ (
    .Q(\datapath_1.regfile_1.regOut[0] [2]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_6769_[2])
);

INVX1 _11974_ (
    .A(\datapath_1.PCJump [29]),
    .Y(_3024_)
);

FILL FILL_3__7380_ (
);

FILL FILL_0__11689_ (
);

FILL FILL_0__9283_ (
);

FILL FILL_0__11269_ (
);

AOI22X1 _11554_ (
    .A(_2478_),
    .B(_2231_),
    .C(_2230_),
    .D(_2341__bF$buf0),
    .Y(_2663_)
);

FILL FILL_5_CLKBUF1_insert220 (
);

NAND2X1 _11134_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2253_)
);

FILL SFILL43960x79050 (
);

FILL FILL_5_CLKBUF1_insert221 (
);

FILL FILL_3__12603_ (
);

FILL FILL_5_CLKBUF1_insert222 (
);

FILL FILL_5_CLKBUF1_insert223 (
);

FILL FILL_5_CLKBUF1_insert224 (
);

FILL FILL_4__16082_ (
);

FILL FILL_0__12630_ (
);

FILL FILL_3__15495_ (
);

FILL FILL_3__15075_ (
);

FILL FILL_0__12210_ (
);

FILL FILL_1__7298_ (
);

FILL FILL112360x83050 (
);

FILL FILL_2__14488_ (
);

FILL FILL_2__14068_ (
);

FILL FILL_5__15822_ (
);

FILL FILL_5__15402_ (
);

DFFSR _9702_ (
    .Q(\datapath_1.regfile_1.regOut[22] [16]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1368_[16])
);

FILL SFILL19400x66050 (
);

FILL FILL_4__14815_ (
);

FILL SFILL28680x1050 (
);

FILL FILL_3__8585_ (
);

NAND2X1 _12759_ (
    .A(IRWrite_bF$buf1),
    .B(memoryOutData[21]),
    .Y(_3532_)
);

NAND3X1 _12339_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3293_)
);

FILL SFILL3720x27050 (
);

FILL FILL_3__13808_ (
);

FILL SFILL64840x75050 (
);

FILL FILL_1__14842_ (
);

FILL FILL_1__14422_ (
);

FILL FILL_1__14002_ (
);

FILL SFILL43960x34050 (
);

FILL FILL_0__13835_ (
);

FILL FILL_0__13415_ (
);

INVX1 _13700_ (
    .A(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_4207_)
);

FILL FILL_5__9872_ (
);

FILL FILL_5__9032_ (
);

FILL SFILL108920x52050 (
);

NAND3X1 _16172_ (
    .A(_6617_),
    .B(_6618_),
    .C(_6623_),
    .Y(_6624_)
);

FILL FILL_1__9864_ (
);

FILL FILL_5__11742_ (
);

FILL FILL_5__11322_ (
);

FILL FILL_1__9024_ (
);

FILL FILL_2__16214_ (
);

FILL FILL_4__10315_ (
);

FILL FILL_1__15627_ (
);

FILL SFILL94280x50 (
);

FILL FILL_1__15207_ (
);

NAND2X1 _8094_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_614_)
);

FILL FILL_1__10762_ (
);

NOR2X1 _14905_ (
    .A(_5386_),
    .B(_5383_),
    .Y(_5387_)
);

FILL FILL_2__7367_ (
);

NAND3X1 _12092_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [26]),
    .C(_3034__bF$buf2),
    .Y(_3115_)
);

FILL FILL_5__12527_ (
);

FILL FILL_3__13981_ (
);

FILL FILL_5__12107_ (
);

FILL FILL_3__13561_ (
);

FILL FILL_3__13141_ (
);

FILL FILL_4__8654_ (
);

FILL FILL_4__8234_ (
);

FILL FILL_2__12974_ (
);

FILL FILL_2__12134_ (
);

INVX1 _9299_ (
    .A(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_1234_)
);

FILL FILL_1__11967_ (
);

FILL FILL_1__11547_ (
);

FILL FILL_1__11127_ (
);

FILL FILL_0__8974_ (
);

FILL FILL_5__16360_ (
);

FILL FILL_0__8134_ (
);

OAI21X1 _10825_ (
    .A(_2006_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_2007_),
    .Y(_1953_[27])
);

OAI21X1 _10405_ (
    .A(_1787_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1788_),
    .Y(_1758_[15])
);

FILL FILL_5__6997_ (
);

FILL FILL_6__14319_ (
);

FILL FILL_4__15773_ (
);

FILL FILL_4__15353_ (
);

NOR3X1 _13297_ (
    .A(_3796_),
    .B(_3833_),
    .C(_3781_),
    .Y(\datapath_1.regfile_1.regEn [7])
);

FILL FILL_2__9933_ (
);

FILL FILL_0__11901_ (
);

FILL FILL_3__14766_ (
);

FILL FILL_2__9513_ (
);

FILL FILL_3__14346_ (
);

FILL FILL_1__15380_ (
);

FILL FILL_1__6989_ (
);

FILL FILL_4__9859_ (
);

FILL FILL_4__9019_ (
);

FILL FILL_2__13759_ (
);

FILL FILL_2__13339_ (
);

FILL FILL_0__14793_ (
);

FILL SFILL33880x39050 (
);

FILL FILL_0__14373_ (
);

FILL FILL_1__7930_ (
);

FILL FILL_2__14700_ (
);

FILL FILL_3__7856_ (
);

FILL FILL_0__9759_ (
);

FILL FILL_3__7436_ (
);

FILL FILL_0__9339_ (
);

FILL FILL_5__12280_ (
);

FILL FILL_4__16138_ (
);

FILL SFILL2840x82050 (
);

FILL FILL_4__11693_ (
);

FILL FILL_4__11273_ (
);

FILL FILL_1__16165_ (
);

FILL FILL_3__10686_ (
);

FILL FILL_5__8723_ (
);

FILL FILL_3__10266_ (
);

FILL FILL_0__15998_ (
);

AOI22X1 _15863_ (
    .A(_5570__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[27] [20]),
    .C(\datapath_1.regfile_1.regOut[26] [20]),
    .D(_5484_),
    .Y(_6323_)
);

FILL FILL_0__15578_ (
);

INVX1 _15443_ (
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_5914_)
);

FILL FILL_0__15158_ (
);

NAND2X1 _15023_ (
    .A(_5462_),
    .B(_5500__bF$buf2),
    .Y(_5503_)
);

FILL FILL_0__10293_ (
);

FILL FILL_1__8715_ (
);

FILL FILL_2__15905_ (
);

FILL FILL_5__13485_ (
);

FILL FILL_2__10620_ (
);

DFFSR _7785_ (
    .Q(\datapath_1.regfile_1.regOut[7] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_393_[19])
);

FILL SFILL28760x50 (
);

NAND2X1 _7365_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_250_)
);

FILL FILL_4__12898_ (
);

FILL FILL_4__12478_ (
);

FILL FILL_4__12058_ (
);

FILL FILL_2__13092_ (
);

FILL SFILL94440x17050 (
);

FILL FILL_5_BUFX2_insert40 (
);

FILL FILL_5_BUFX2_insert41 (
);

FILL FILL_5__9928_ (
);

FILL FILL_5__9508_ (
);

FILL FILL_5_BUFX2_insert42 (
);

FILL FILL_5_BUFX2_insert43 (
);

FILL FILL_1__12085_ (
);

FILL FILL_5_BUFX2_insert44 (
);

FILL FILL_5_BUFX2_insert45 (
);

FILL SFILL23080x54050 (
);

FILL FILL_5_BUFX2_insert46 (
);

OAI22X1 _16228_ (
    .A(_5325_),
    .B(_5544__bF$buf3),
    .C(_5523_),
    .D(_6678_),
    .Y(_6679_)
);

FILL FILL_5_BUFX2_insert47 (
);

FILL FILL_5_BUFX2_insert48 (
);

FILL FILL_5_BUFX2_insert49 (
);

FILL FILL_0__9092_ (
);

OR2X2 _11783_ (
    .A(_2875_),
    .B(_2876_),
    .Y(_2877_)
);

FILL FILL_0__11498_ (
);

NAND2X1 _11363_ (
    .A(_2340_),
    .B(_2336_),
    .Y(_2480_)
);

FILL FILL_0__11078_ (
);

FILL SFILL23880x37050 (
);

FILL SFILL54280x28050 (
);

FILL FILL_3__12832_ (
);

FILL FILL_3__12412_ (
);

FILL FILL_4__7505_ (
);

FILL FILL_4_CLKBUF1_insert210 (
);

FILL FILL_4_CLKBUF1_insert211 (
);

FILL FILL_2__11825_ (
);

FILL FILL_4_CLKBUF1_insert212 (
);

FILL FILL_2__11405_ (
);

FILL FILL_4_CLKBUF1_insert213 (
);

FILL FILL_4_CLKBUF1_insert214 (
);

FILL FILL_4_CLKBUF1_insert215 (
);

FILL FILL_4_CLKBUF1_insert216 (
);

FILL FILL_4_CLKBUF1_insert217 (
);

FILL FILL_4_CLKBUF1_insert218 (
);

FILL FILL_1__10818_ (
);

FILL FILL_4_CLKBUF1_insert219 (
);

FILL FILL_2__14297_ (
);

FILL FILL_5__15631_ (
);

FILL SFILL84920x22050 (
);

FILL FILL_5__15211_ (
);

FILL FILL_0__7825_ (
);

NAND2X1 _9931_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1554_)
);

NAND2X1 _9511_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1335_)
);

FILL FILL_4__14624_ (
);

FILL FILL_4__14204_ (
);

FILL FILL_3__8394_ (
);

NAND2X1 _12988_ (
    .A(vdd),
    .B(\datapath_1.rd2 [12]),
    .Y(_3644_)
);

NAND2X1 _12568_ (
    .A(memoryOutData[0]),
    .B(vdd),
    .Y(_3489_)
);

FILL SFILL23800x35050 (
);

INVX1 _12148_ (
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_3152_)
);

FILL FILL_3__13617_ (
);

FILL FILL_1__14651_ (
);

FILL FILL_1__14231_ (
);

FILL SFILL84040x46050 (
);

FILL FILL_0_BUFX2_insert110 (
);

FILL SFILL8840x34050 (
);

FILL FILL_0__13644_ (
);

FILL FILL_0__13224_ (
);

FILL FILL_3__16089_ (
);

FILL FILL_5__9681_ (
);

FILL FILL_5__9261_ (
);

FILL SFILL74120x82050 (
);

FILL FILL_5__16416_ (
);

FILL FILL_5__11971_ (
);

FILL FILL_1__9673_ (
);

FILL FILL_5__11551_ (
);

FILL FILL_1__9253_ (
);

FILL FILL_5__11131_ (
);

FILL FILL_4__15829_ (
);

FILL FILL_4__15409_ (
);

BUFX2 BUFX2_insert1030 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf4 )
);

BUFX2 BUFX2_insert1031 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf3 )
);

FILL FILL_3__9599_ (
);

FILL FILL_2__16023_ (
);

BUFX2 BUFX2_insert1032 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf2 )
);

BUFX2 BUFX2_insert1033 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf1 )
);

FILL FILL_4__10964_ (
);

BUFX2 BUFX2_insert1034 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf0 )
);

FILL FILL_4__10544_ (
);

BUFX2 BUFX2_insert1035 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf4 )
);

FILL FILL_4__10124_ (
);

BUFX2 BUFX2_insert1036 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf3 )
);

BUFX2 BUFX2_insert1037 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf2 )
);

FILL FILL_1__15856_ (
);

BUFX2 BUFX2_insert1038 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf1 )
);

FILL FILL_1__15436_ (
);

BUFX2 BUFX2_insert1039 (
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf0 )
);

FILL FILL_1__15016_ (
);

FILL FILL_1__10991_ (
);

FILL FILL_1__10571_ (
);

FILL FILL_1__10151_ (
);

FILL FILL_0__14849_ (
);

NAND3X1 _14714_ (
    .A(_5199_),
    .B(_5198_),
    .C(_5195_),
    .Y(_5200_)
);

FILL FILL_0__14429_ (
);

FILL FILL_0__14009_ (
);

BUFX2 BUFX2_insert850 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf5 )
);

FILL FILL_2__7596_ (
);

FILL FILL_2__7176_ (
);

BUFX2 BUFX2_insert851 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf4 )
);

BUFX2 BUFX2_insert852 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf3 )
);

BUFX2 BUFX2_insert853 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf2 )
);

BUFX2 BUFX2_insert854 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf1 )
);

BUFX2 BUFX2_insert855 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf0 )
);

BUFX2 BUFX2_insert856 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf7 )
);

BUFX2 BUFX2_insert857 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf6 )
);

BUFX2 BUFX2_insert858 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf5 )
);

BUFX2 BUFX2_insert859 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf4 )
);

FILL FILL_5__12756_ (
);

FILL FILL_3__13790_ (
);

FILL FILL_5__12336_ (
);

FILL FILL_3__13370_ (
);

FILL FILL_4__8883_ (
);

FILL FILL_4__8463_ (
);

FILL FILL_4__11749_ (
);

FILL FILL_2__12783_ (
);

FILL FILL_4__11329_ (
);

FILL FILL_2__12363_ (
);

FILL SFILL13800x33050 (
);

FILL FILL_1__11776_ (
);

FILL FILL_1__11356_ (
);

INVX1 _15919_ (
    .A(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_6378_)
);

FILL FILL_0__8783_ (
);

FILL FILL_3__6880_ (
);

FILL FILL_0__8363_ (
);

FILL FILL_0__10769_ (
);

OAI21X1 _10634_ (
    .A(_1899_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1900_),
    .Y(_1888_[6])
);

DFFSR _10214_ (
    .Q(\datapath_1.regfile_1.regOut[26] [16]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_1628_[16])
);

FILL FILL_6__14968_ (
);

FILL FILL_4__15582_ (
);

FILL FILL_4__15162_ (
);

FILL FILL_2__9742_ (
);

FILL FILL_3__14995_ (
);

FILL FILL_3__14575_ (
);

FILL FILL_0__11710_ (
);

FILL FILL_3__14155_ (
);

FILL FILL_4_BUFX2_insert690 (
);

FILL FILL_4__9668_ (
);

FILL FILL_4_BUFX2_insert691 (
);

FILL FILL_4__9248_ (
);

FILL FILL_4_BUFX2_insert692 (
);

FILL FILL112360x78050 (
);

FILL FILL_2__13988_ (
);

FILL FILL_4_BUFX2_insert693 (
);

FILL FILL_4_BUFX2_insert694 (
);

FILL FILL_2__13568_ (
);

FILL FILL_4_BUFX2_insert695 (
);

FILL FILL_2__13148_ (
);

FILL FILL_0__14182_ (
);

FILL FILL_4_BUFX2_insert696 (
);

FILL FILL_5__14902_ (
);

FILL FILL_4_BUFX2_insert697 (
);

FILL FILL_4_BUFX2_insert698 (
);

FILL FILL_4_BUFX2_insert699 (
);

FILL FILL_0__9988_ (
);

FILL FILL_0__9148_ (
);

FILL FILL_3__7245_ (
);

NAND2X1 _11839_ (
    .A(_2492_),
    .B(_2927_),
    .Y(_2928_)
);

NAND3X1 _11419_ (
    .A(_2316_),
    .B(_2323_),
    .C(_2304_),
    .Y(_2535_)
);

FILL FILL_1__13922_ (
);

FILL FILL_4__16367_ (
);

FILL FILL_1__13502_ (
);

FILL SFILL43960x29050 (
);

FILL SFILL24360x60050 (
);

FILL FILL_4__11082_ (
);

FILL FILL_0__12915_ (
);

FILL FILL_1__16394_ (
);

FILL FILL_5__8952_ (
);

FILL FILL_3__10495_ (
);

FILL FILL_5__8532_ (
);

FILL FILL_5__8112_ (
);

FILL FILL_0__15387_ (
);

OAI22X1 _15672_ (
    .A(_6135_),
    .B(_5545__bF$buf1),
    .C(_5485__bF$buf4),
    .D(_6136_),
    .Y(_6137_)
);

INVX1 _15252_ (
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_5728_)
);

FILL SFILL104200x25050 (
);

FILL FILL112360x33050 (
);

FILL FILL_3__16301_ (
);

FILL FILL_5__10822_ (
);

FILL FILL_5__10402_ (
);

FILL FILL_1__8524_ (
);

FILL FILL_1__8104_ (
);

FILL FILL_2__15714_ (
);

FILL SFILL64040x42050 (
);

FILL FILL_5__13294_ (
);

FILL FILL_1__14707_ (
);

NAND2X1 _7594_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_362_)
);

FILL FILL_4_BUFX2_insert1070 (
);

FILL FILL_4_BUFX2_insert1071 (
);

NAND2X1 _7174_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_143_)
);

FILL FILL_4_BUFX2_insert1072 (
);

FILL FILL_4_BUFX2_insert1073 (
);

FILL FILL_4__12287_ (
);

FILL FILL_3__9811_ (
);

FILL FILL_2__6867_ (
);

FILL FILL_5__9737_ (
);

FILL FILL_6__12614_ (
);

NAND3X1 _16037_ (
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .B(_5477_),
    .C(_5531__bF$buf4),
    .Y(_6493_)
);

NOR2X1 _11592_ (
    .A(_2698_),
    .B(_2697_),
    .Y(_2699_)
);

INVX2 _11172_ (
    .A(_2290_),
    .Y(_2291_)
);

FILL FILL_1__9729_ (
);

FILL FILL_5__11607_ (
);

FILL FILL_3__12641_ (
);

FILL FILL_6__15086_ (
);

FILL FILL_3__12221_ (
);

FILL FILL_4__7734_ (
);

FILL FILL_4__7314_ (
);

FILL FILL_5__14499_ (
);

FILL FILL_2__11634_ (
);

FILL FILL_2__11214_ (
);

FILL FILL_5__14079_ (
);

DFFSR _8799_ (
    .Q(\datapath_1.regfile_1.regOut[15] [9]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_913_[9])
);

INVX1 _8379_ (
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_763_)
);

FILL FILL_1__10627_ (
);

FILL FILL_5__15860_ (
);

FILL FILL_5__15440_ (
);

FILL FILL_5__15020_ (
);

FILL FILL_0__7634_ (
);

NAND2X1 _9740_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1447_)
);

FILL FILL_0__7214_ (
);

DFFSR _9320_ (
    .Q(\datapath_1.regfile_1.regOut[19] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1173_[18])
);

FILL FILL_1__13099_ (
);

FILL FILL_4__14853_ (
);

FILL FILL_4__14433_ (
);

FILL FILL_4__14013_ (
);

DFFSR _12797_ (
    .Q(\datapath_1.PCJump [8]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[6])
);

NAND2X1 _12377_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [11]),
    .Y(_3317_)
);

FILL FILL_3__13846_ (
);

FILL FILL_1__14880_ (
);

FILL FILL_3__13426_ (
);

FILL FILL_1__14460_ (
);

FILL FILL_3__13006_ (
);

FILL FILL_1__14040_ (
);

FILL FILL_4__8519_ (
);

FILL FILL_2__12839_ (
);

FILL FILL_0__13873_ (
);

FILL FILL_2__12419_ (
);

FILL FILL_0__13453_ (
);

FILL FILL_0__13033_ (
);

FILL FILL_5__9490_ (
);

FILL SFILL54040x40050 (
);

FILL FILL_5__16225_ (
);

FILL FILL_3__6936_ (
);

FILL FILL_0__8839_ (
);

FILL FILL_5__11780_ (
);

FILL FILL_1__9482_ (
);

FILL FILL_5__11360_ (
);

FILL FILL_4__15638_ (
);

FILL FILL_4__15218_ (
);

FILL FILL_2__16252_ (
);

FILL FILL_4__10773_ (
);

FILL FILL_1__15665_ (
);

FILL FILL_1__15245_ (
);

FILL FILL_5__7803_ (
);

FILL FILL_1__10380_ (
);

AOI22X1 _14943_ (
    .A(\datapath_1.regfile_1.regOut[2] [31]),
    .B(_3998__bF$buf3),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_5424_)
);

FILL FILL_0__14658_ (
);

FILL FILL_0__14238_ (
);

INVX1 _14523_ (
    .A(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_5013_)
);

INVX1 _14103_ (
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_4602_)
);

FILL SFILL44040x83050 (
);

FILL FILL_6__13572_ (
);

FILL FILL_5__12985_ (
);

FILL FILL_5__12145_ (
);

BUFX2 _6865_ (
    .A(_1_[27]),
    .Y(memoryAddress[27])
);

FILL FILL_4__11978_ (
);

FILL FILL_4__8272_ (
);

FILL FILL_4__11558_ (
);

FILL FILL_2__12592_ (
);

FILL FILL_4__11138_ (
);

FILL FILL_2__12172_ (
);

FILL FILL_1__11585_ (
);

FILL FILL_1__11165_ (
);

OAI22X1 _15728_ (
    .A(_5463__bF$buf3),
    .B(_6191_),
    .C(_5526__bF$buf2),
    .D(_4725_),
    .Y(_6192_)
);

NOR2X1 _15308_ (
    .A(_5781_),
    .B(_5780_),
    .Y(_5782_)
);

FILL FILL_0__8592_ (
);

FILL FILL_0__10998_ (
);

FILL FILL_0__10578_ (
);

DFFSR _10863_ (
    .Q(\datapath_1.regfile_1.regOut[31] [25]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_1953_[25])
);

NAND2X1 _10443_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1814_)
);

FILL FILL_0__10158_ (
);

NAND2X1 _10023_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1595_)
);

FILL FILL_3__11912_ (
);

FILL FILL_4__15391_ (
);

FILL FILL_2__10905_ (
);

FILL FILL112440x9050 (
);

FILL FILL_2__9551_ (
);

FILL FILL_3__14384_ (
);

FILL FILL_2__9131_ (
);

FILL FILL_4__9897_ (
);

FILL SFILL84120x34050 (
);

FILL FILL_4__9477_ (
);

FILL FILL_2__13797_ (
);

FILL FILL_2__13377_ (
);

FILL FILL112120x3050 (
);

FILL FILL_5__14711_ (
);

FILL FILL111800x6050 (
);

FILL FILL_0__6905_ (
);

FILL SFILL109320x77050 (
);

FILL FILL_4__13704_ (
);

FILL FILL_0__9797_ (
);

FILL FILL_0__9377_ (
);

FILL FILL_3__7474_ (
);

FILL FILL_3__7054_ (
);

AOI21X1 _11648_ (
    .A(_2404_),
    .B(_2750_),
    .C(_2749_),
    .Y(_2751_)
);

NAND3X1 _11228_ (
    .A(_2333_),
    .B(ALUControl[0]),
    .C(_2343_),
    .Y(_2347_)
);

FILL FILL_1__13731_ (
);

FILL FILL_1__13311_ (
);

FILL FILL_4__16176_ (
);

FILL FILL_6__10697_ (
);

FILL FILL_0__12724_ (
);

FILL FILL_3__15589_ (
);

FILL FILL_3__15169_ (
);

FILL FILL_0__12304_ (
);

FILL FILL_5__8761_ (
);

FILL FILL_5__8341_ (
);

FILL FILL_0__15196_ (
);

NAND3X1 _15481_ (
    .A(_5944_),
    .B(_5950_),
    .C(_5947_),
    .Y(_5951_)
);

FILL FILL_5__15916_ (
);

NAND3X1 _15061_ (
    .A(\datapath_1.PCJump [26]),
    .B(_5470_),
    .C(_5468_),
    .Y(_5541_)
);

FILL FILL_3__16110_ (
);

FILL FILL_1__8753_ (
);

FILL FILL_5__10631_ (
);

FILL FILL_1__8333_ (
);

FILL FILL_4__14909_ (
);

FILL FILL_2__15943_ (
);

FILL FILL_2__15523_ (
);

FILL FILL_2__15103_ (
);

FILL FILL_3__8259_ (
);

FILL FILL_1__14936_ (
);

FILL FILL_1__14516_ (
);

FILL FILL_4__12096_ (
);

FILL FILL_3__9620_ (
);

FILL FILL_0__13929_ (
);

FILL FILL_0__13509_ (
);

FILL FILL_5__9546_ (
);

FILL FILL_5__9126_ (
);

FILL FILL_3__11089_ (
);

FILL FILL_6__12423_ (
);

NOR3X1 _16266_ (
    .A(_6713_),
    .B(_6715_),
    .C(_6714_),
    .Y(_6716_)
);

FILL SFILL74120x32050 (
);

FILL FILL_5__11836_ (
);

FILL FILL_3__12870_ (
);

FILL FILL_5__11416_ (
);

FILL FILL_1__9538_ (
);

FILL FILL_3__12450_ (
);

FILL FILL_1__9118_ (
);

FILL FILL_3__12030_ (
);

FILL FILL_4__7963_ (
);

FILL FILL_2__16308_ (
);

FILL SFILL99320x81050 (
);

FILL FILL_4__7543_ (
);

FILL FILL_4__10829_ (
);

FILL FILL_4__7123_ (
);

FILL FILL_4__10409_ (
);

FILL FILL_2__11863_ (
);

FILL FILL_2__11443_ (
);

FILL FILL_2__11023_ (
);

INVX1 _8188_ (
    .A(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_656_)
);

FILL SFILL13800x28050 (
);

FILL FILL_1__10436_ (
);

FILL FILL_1__10016_ (
);

FILL FILL_0__7863_ (
);

FILL FILL_0__7443_ (
);

FILL FILL_6__13628_ (
);

FILL FILL_6__13208_ (
);

FILL FILL_4__14662_ (
);

FILL FILL_4__14242_ (
);

OAI21X1 _12186_ (
    .A(_3176_),
    .B(ALUSrcA_bF$buf6),
    .C(_3177_),
    .Y(\datapath_1.alu_1.ALUInA [23])
);

FILL FILL_2__8822_ (
);

FILL FILL_3__13655_ (
);

FILL FILL_2__8402_ (
);

FILL FILL_3__13235_ (
);

FILL FILL_4__8748_ (
);

FILL FILL_4__8328_ (
);

FILL FILL_2__12648_ (
);

FILL FILL_0__13682_ (
);

FILL FILL_2__12228_ (
);

FILL FILL_0__13262_ (
);

FILL FILL_6_BUFX2_insert91 (
);

FILL FILL_5__16034_ (
);

FILL FILL_0__8648_ (
);

FILL FILL_0__8228_ (
);

NOR2X1 _10919_ (
    .A(_2060_),
    .B(_2053_),
    .Y(RegDst)
);

FILL FILL_6_BUFX2_insert96 (
);

FILL FILL_1__9291_ (
);

FILL FILL_4__15867_ (
);

FILL FILL_4__15447_ (
);

FILL FILL_4__15027_ (
);

FILL FILL_2__16061_ (
);

FILL FILL_4__10162_ (
);

FILL SFILL99240x43050 (
);

FILL FILL_2__9607_ (
);

FILL SFILL64120x30050 (
);

FILL FILL_1__15894_ (
);

FILL FILL_1__15474_ (
);

FILL FILL_1__15054_ (
);

FILL FILL_5__7612_ (
);

FILL FILL_0__14887_ (
);

FILL FILL_0__14467_ (
);

OAI22X1 _14752_ (
    .A(_3967__bF$buf2),
    .B(_5235_),
    .C(_3935__bF$buf0),
    .D(_5236_),
    .Y(_5237_)
);

FILL FILL_0__14047_ (
);

NAND3X1 _14332_ (
    .A(_4817_),
    .B(_4818_),
    .C(_4825_),
    .Y(_4826_)
);

FILL FILL112360x28050 (
);

FILL FILL_3__15801_ (
);

FILL FILL_1__7604_ (
);

FILL SFILL64040x37050 (
);

FILL FILL_5__12374_ (
);

FILL FILL_4__11787_ (
);

FILL FILL_4__8081_ (
);

FILL FILL_4__11367_ (
);

FILL SFILL54120x73050 (
);

FILL FILL_1__16259_ (
);

FILL FILL_1__11394_ (
);

INVX1 _15957_ (
    .A(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_6415_)
);

AOI22X1 _15537_ (
    .A(_5570__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .C(\datapath_1.regfile_1.regOut[9] [12]),
    .D(_5560_),
    .Y(_6005_)
);

INVX1 _15117_ (
    .A(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_5596_)
);

NAND2X1 _10672_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1926_)
);

FILL FILL_0__10387_ (
);

NAND2X1 _10252_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1707_)
);

FILL FILL_3__11721_ (
);

FILL FILL_3__11301_ (
);

FILL FILL_5__13999_ (
);

FILL FILL_2__9780_ (
);

FILL FILL_5__13579_ (
);

FILL FILL_2__9360_ (
);

FILL FILL_5__13159_ (
);

FILL FILL_3__14193_ (
);

INVX1 _7879_ (
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_511_)
);

INVX1 _7459_ (
    .A(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_292_)
);

INVX1 _7039_ (
    .A(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_73_)
);

FILL FILL_4__9286_ (
);

FILL FILL_5__14940_ (
);

FILL FILL_5__14520_ (
);

FILL FILL_5__14100_ (
);

DFFSR _8820_ (
    .Q(\datapath_1.regfile_1.regOut[15] [30]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_913_[30])
);

FILL FILL_1__12599_ (
);

INVX1 _8400_ (
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_777_)
);

FILL FILL_1__12179_ (
);

FILL FILL_4__13933_ (
);

FILL FILL_4__13513_ (
);

OAI21X1 _11877_ (
    .A(_2960_),
    .B(RegDst),
    .C(_2961_),
    .Y(\datapath_1.a3 [1])
);

NAND3X1 _11457_ (
    .A(_2540_),
    .B(_2536_),
    .C(_2572_),
    .Y(\datapath_1.ALUResult [28])
);

NOR2X1 _11037_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(_2155_),
    .Y(_2156_)
);

FILL FILL_3__12506_ (
);

FILL FILL_1__13960_ (
);

FILL SFILL18680x61050 (
);

FILL FILL_1__13540_ (
);

FILL FILL_1__13120_ (
);

FILL FILL_2__11919_ (
);

FILL FILL_0__12953_ (
);

FILL FILL_3__15398_ (
);

FILL FILL_0__12533_ (
);

FILL FILL_0__12113_ (
);

FILL FILL_5__8990_ (
);

FILL SFILL54040x35050 (
);

FILL FILL_5__8570_ (
);

INVX1 _15290_ (
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_5765_)
);

FILL FILL_5__15725_ (
);

FILL FILL_5__15305_ (
);

INVX1 _9605_ (
    .A(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_1377_)
);

FILL FILL_1__8982_ (
);

FILL FILL_5__10440_ (
);

FILL FILL_5__10020_ (
);

FILL FILL_1__8142_ (
);

FILL FILL_4__14718_ (
);

FILL FILL_2__15752_ (
);

FILL FILL_2__15332_ (
);

FILL FILL_3__8488_ (
);

FILL FILL_3__8068_ (
);

FILL FILL_1__14745_ (
);

FILL FILL_1__14325_ (
);

FILL FILL_0__13738_ (
);

FILL FILL_0__13318_ (
);

INVX1 _13603_ (
    .A(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_4112_)
);

FILL FILL_5__9775_ (
);

FILL SFILL44040x78050 (
);

FILL FILL_5__9355_ (
);

NAND3X1 _16075_ (
    .A(_6523_),
    .B(_6529_),
    .C(_6525_),
    .Y(_6530_)
);

FILL FILL_1__9767_ (
);

FILL FILL_5__11645_ (
);

FILL FILL_1__9347_ (
);

FILL FILL_5__11225_ (
);

FILL FILL_2__16117_ (
);

FILL FILL_4__7352_ (
);

FILL FILL_4__10638_ (
);

FILL FILL_2__11672_ (
);

FILL FILL_2__11252_ (
);

FILL FILL_1__10665_ (
);

FILL FILL_1__10245_ (
);

INVX1 _14808_ (
    .A(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_5292_)
);

FILL FILL_0__7672_ (
);

FILL FILL_0__7252_ (
);

FILL FILL_4__14891_ (
);

FILL FILL_4__14471_ (
);

FILL FILL_6__13017_ (
);

FILL FILL_4__14051_ (
);

FILL SFILL54040x6050 (
);

FILL FILL_2__8631_ (
);

FILL FILL_3__13884_ (
);

FILL FILL_3__13464_ (
);

FILL FILL_2__8211_ (
);

FILL SFILL94280x4050 (
);

FILL FILL_3__13044_ (
);

FILL FILL_4__8977_ (
);

FILL FILL_4__8137_ (
);

FILL FILL_2__12877_ (
);

FILL FILL_2__12457_ (
);

FILL FILL_2__12037_ (
);

FILL FILL_0__13491_ (
);

FILL FILL_3__6974_ (
);

FILL FILL_5__16263_ (
);

FILL FILL_0__8877_ (
);

FILL FILL_0__8457_ (
);

DFFSR _10728_ (
    .Q(\datapath_1.regfile_1.regOut[30] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_1888_[18])
);

INVX1 _10308_ (
    .A(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_1744_)
);

FILL SFILL104520x2050 (
);

FILL FILL_4__15676_ (
);

FILL FILL_4__15256_ (
);

FILL FILL_2__16290_ (
);

FILL SFILL104440x7050 (
);

FILL SFILL109400x20050 (
);

FILL FILL_4__10391_ (
);

FILL FILL_2__9416_ (
);

FILL FILL_0__11804_ (
);

FILL FILL_3__14669_ (
);

FILL FILL_3__14249_ (
);

FILL FILL_1__15283_ (
);

FILL FILL_5__7841_ (
);

FILL FILL_5__7421_ (
);

NOR2X1 _14981_ (
    .A(\datapath_1.PCJump [24]),
    .B(_5460_),
    .Y(_5461_)
);

FILL FILL_0__14696_ (
);

AOI22X1 _14561_ (
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .B(_4038__bF$buf3),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_5050_)
);

FILL FILL_0__14276_ (
);

OAI22X1 _14141_ (
    .A(_3902__bF$buf0),
    .B(_4637_),
    .C(_4638_),
    .D(_3935__bF$buf1),
    .Y(_4639_)
);

FILL FILL_3__15610_ (
);

FILL FILL_1__7833_ (
);

FILL FILL_2__14603_ (
);

FILL FILL_3__7759_ (
);

FILL FILL_3__7339_ (
);

FILL FILL_5__12183_ (
);

FILL FILL_4__11596_ (
);

FILL FILL_4__11176_ (
);

FILL FILL_3__8700_ (
);

FILL SFILL34040x31050 (
);

FILL FILL_1__16068_ (
);

FILL FILL_5__8626_ (
);

FILL FILL_5__8206_ (
);

FILL FILL_3__10169_ (
);

OAI22X1 _15766_ (
    .A(_5485__bF$buf2),
    .B(_4790_),
    .C(_5483__bF$buf1),
    .D(_4802_),
    .Y(_6229_)
);

FILL SFILL74120x27050 (
);

OAI22X1 _15346_ (
    .A(_5472__bF$buf1),
    .B(_4328_),
    .C(_4327_),
    .D(_5552__bF$buf0),
    .Y(_5819_)
);

FILL FILL_0__10196_ (
);

DFFSR _10481_ (
    .Q(\datapath_1.regfile_1.regOut[28] [27]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1758_[27])
);

INVX1 _10061_ (
    .A(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_1620_)
);

FILL FILL_5__10916_ (
);

FILL FILL_3__11950_ (
);

FILL FILL_1__8618_ (
);

FILL FILL_6__14395_ (
);

FILL FILL_3__11530_ (
);

FILL FILL_3__11110_ (
);

FILL FILL_2__15808_ (
);

FILL SFILL104680x83050 (
);

FILL FILL_0__16002_ (
);

FILL FILL_2__10943_ (
);

FILL FILL_5__13388_ (
);

FILL FILL_2__10523_ (
);

FILL FILL_2__10103_ (
);

INVX1 _7688_ (
    .A(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_404_)
);

DFFSR _7268_ (
    .Q(\datapath_1.regfile_1.regOut[3] [14]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_133_[14])
);

FILL FILL_4__9095_ (
);

FILL FILL_3__9905_ (
);

FILL FILL_0__6943_ (
);

FILL FILL_4__13742_ (
);

FILL FILL_4__13322_ (
);

FILL FILL_3__7092_ (
);

NOR2X1 _11686_ (
    .A(_2786_),
    .B(_2785_),
    .Y(_2787_)
);

NOR2X1 _11266_ (
    .A(_2384_),
    .B(_2195_),
    .Y(_2385_)
);

FILL FILL_3__12735_ (
);

FILL FILL_3__12315_ (
);

FILL FILL_4__7828_ (
);

FILL SFILL24440x43050 (
);

FILL FILL_2__11728_ (
);

FILL FILL_0__12762_ (
);

FILL FILL_2__11308_ (
);

FILL SFILL99320x31050 (
);

FILL FILL_0__12342_ (
);

FILL SFILL23800x3050 (
);

FILL SFILL23720x8050 (
);

FILL FILL_5__15954_ (
);

FILL SFILL63960x6050 (
);

FILL FILL_5__15534_ (
);

FILL FILL_0__7728_ (
);

FILL FILL_5__15114_ (
);

FILL SFILL28760x51050 (
);

FILL SFILL8680x50 (
);

FILL FILL_0__7308_ (
);

DFFSR _9834_ (
    .Q(\datapath_1.regfile_1.regOut[23] [20]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1433_[20])
);

FILL SFILL59160x42050 (
);

OAI21X1 _9414_ (
    .A(_1289_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1290_),
    .Y(_1238_[26])
);

FILL FILL_1__8371_ (
);

FILL FILL_4__14947_ (
);

FILL FILL_2__15981_ (
);

FILL FILL_4__14527_ (
);

FILL FILL_2__15561_ (
);

FILL FILL_4__14107_ (
);

FILL FILL_2__15141_ (
);

FILL SFILL64120x25050 (
);

FILL SFILL3640x4050 (
);

FILL FILL_1__14974_ (
);

FILL FILL_1__14554_ (
);

FILL FILL_1__14134_ (
);

FILL FILL_0__13967_ (
);

INVX1 _13832_ (
    .A(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_4337_)
);

FILL FILL_0__13547_ (
);

NAND2X1 _13412_ (
    .A(_3888_),
    .B(_3917_),
    .Y(_3924_)
);

FILL FILL_0__13127_ (
);

FILL FILL_5__9164_ (
);

FILL FILL_5__16319_ (
);

FILL FILL_1__9996_ (
);

FILL FILL_5__11874_ (
);

FILL FILL_5__11454_ (
);

FILL FILL_1__9156_ (
);

FILL FILL_5__11034_ (
);

FILL FILL_2__16346_ (
);

FILL FILL_4__7581_ (
);

FILL FILL_4__7161_ (
);

FILL SFILL114280x3050 (
);

FILL FILL_4__10447_ (
);

FILL FILL_4__10027_ (
);

FILL FILL_2__11481_ (
);

FILL SFILL54120x68050 (
);

FILL FILL_2__11061_ (
);

FILL FILL_1__15759_ (
);

FILL FILL_1__15339_ (
);

FILL FILL_1__10894_ (
);

FILL FILL_1__10054_ (
);

NAND3X1 _14617_ (
    .A(_5096_),
    .B(_5097_),
    .C(_5104_),
    .Y(_5105_)
);

FILL FILL_2__7499_ (
);

FILL FILL_0__7481_ (
);

FILL FILL_2__7079_ (
);

FILL FILL_0__7061_ (
);

FILL FILL_3__10801_ (
);

FILL FILL_4__14280_ (
);

FILL FILL_5__12659_ (
);

FILL FILL_2__8860_ (
);

FILL FILL_2__8440_ (
);

FILL FILL_5__12239_ (
);

FILL FILL_3__13693_ (
);

FILL FILL_3__13273_ (
);

INVX1 _6959_ (
    .A(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_40_)
);

FILL FILL_2__8020_ (
);

FILL FILL_4__8786_ (
);

FILL FILL_4__8366_ (
);

FILL FILL_2__12266_ (
);

FILL FILL_5__13600_ (
);

DFFSR _7900_ (
    .Q(\datapath_1.regfile_1.regOut[8] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_458_[6])
);

FILL SFILL54120x23050 (
);

FILL FILL_1__11679_ (
);

FILL FILL_1__11259_ (
);

FILL FILL_5__16072_ (
);

NAND2X1 _10957_ (
    .A(\control_1.op [3]),
    .B(_2071_),
    .Y(_2089_)
);

FILL FILL_0__8266_ (
);

FILL FILL_6__9653_ (
);

INVX1 _10537_ (
    .A(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_1856_)
);

INVX1 _10117_ (
    .A(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_1637_)
);

FILL SFILL79320x72050 (
);

FILL SFILL18680x56050 (
);

FILL FILL_1__12620_ (
);

FILL FILL_4__15485_ (
);

FILL FILL_4__15065_ (
);

FILL FILL_1__12200_ (
);

FILL FILL_2__9645_ (
);

FILL FILL_3__14898_ (
);

FILL FILL_3__14478_ (
);

FILL FILL_2__9225_ (
);

FILL FILL_0__11613_ (
);

FILL FILL_3__14058_ (
);

FILL FILL_1__15092_ (
);

FILL FILL_6__15812_ (
);

FILL FILL_5__7230_ (
);

NOR2X1 _14790_ (
    .A(_5274_),
    .B(_5260_),
    .Y(_5275_)
);

OAI22X1 _14370_ (
    .A(_4862_),
    .B(_3941_),
    .C(_3978_),
    .D(_4861_),
    .Y(_4863_)
);

FILL FILL_0__14085_ (
);

FILL FILL_5__14805_ (
);

FILL FILL_1__7222_ (
);

FILL FILL_2__14832_ (
);

FILL FILL_2__14412_ (
);

FILL FILL_3__7988_ (
);

FILL FILL_3__7568_ (
);

FILL FILL_1__13825_ (
);

FILL FILL_1__13405_ (
);

FILL SFILL18680x11050 (
);

FILL FILL_1__16297_ (
);

FILL FILL_5__8855_ (
);

FILL FILL_3__10398_ (
);

FILL FILL_5__8015_ (
);

NAND3X1 _15995_ (
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .B(_5477_),
    .C(_5531__bF$buf2),
    .Y(_6452_)
);

FILL FILL_6__11732_ (
);

AOI22X1 _15575_ (
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .B(_5567_),
    .C(_5565__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_6042_)
);

NOR2X1 _15155_ (
    .A(_5630_),
    .B(_5632_),
    .Y(_5633_)
);

FILL FILL_3__16204_ (
);

INVX1 _10290_ (
    .A(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_1732_)
);

FILL FILL_1__8847_ (
);

FILL FILL_5__10305_ (
);

FILL FILL_1__8007_ (
);

FILL SFILL79240x34050 (
);

FILL FILL_2__15617_ (
);

FILL FILL_4__6852_ (
);

FILL FILL_0__16231_ (
);

FILL FILL_2__10752_ (
);

OAI21X1 _7497_ (
    .A(_316_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_317_),
    .Y(_263_[27])
);

OAI21X1 _7077_ (
    .A(_97_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .C(_98_),
    .Y(_68_[15])
);

FILL SFILL109320x4050 (
);

FILL FILL_4__13971_ (
);

FILL SFILL44040x28050 (
);

FILL FILL_4__13551_ (
);

FILL FILL_4__13131_ (
);

AOI22X1 _11495_ (
    .A(_2294_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf0),
    .D(_2295_),
    .Y(_2608_)
);

XNOR2X1 _11075_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2194_)
);

FILL FILL_3__12964_ (
);

FILL FILL_2__7711_ (
);

FILL FILL_3__12124_ (
);

FILL FILL_4__7637_ (
);

FILL FILL_4__7217_ (
);

FILL FILL_2__11957_ (
);

FILL FILL_0__12991_ (
);

FILL FILL_2__11537_ (
);

FILL FILL_0__12571_ (
);

FILL FILL_3_CLKBUF1_insert150 (
);

FILL FILL_2__11117_ (
);

FILL FILL_0__12151_ (
);

FILL FILL_3_CLKBUF1_insert151 (
);

FILL FILL_3_CLKBUF1_insert152 (
);

FILL FILL_3_CLKBUF1_insert153 (
);

FILL FILL_6__16350_ (
);

FILL FILL_3_CLKBUF1_insert154 (
);

FILL FILL_3_CLKBUF1_insert155 (
);

FILL FILL_3_CLKBUF1_insert156 (
);

FILL FILL_3_CLKBUF1_insert157 (
);

FILL FILL_3_CLKBUF1_insert158 (
);

FILL FILL_3_CLKBUF1_insert159 (
);

FILL FILL_5__15763_ (
);

FILL FILL_5__15343_ (
);

FILL FILL_0__7957_ (
);

FILL FILL_0__7117_ (
);

OAI21X1 _9643_ (
    .A(_1401_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .C(_1402_),
    .Y(_1368_[17])
);

OAI21X1 _9223_ (
    .A(_1182_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .C(_1183_),
    .Y(_1173_[5])
);

FILL FILL_4__14756_ (
);

FILL FILL_2__15790_ (
);

FILL FILL_4__14336_ (
);

FILL FILL_2__15370_ (
);

FILL SFILL109400x15050 (
);

FILL FILL_2__8916_ (
);

FILL FILL_3__13749_ (
);

FILL FILL_3__13329_ (
);

FILL FILL_1__14783_ (
);

FILL FILL_1__14363_ (
);

FILL FILL_5__6921_ (
);

FILL FILL_0__13776_ (
);

FILL SFILL69240x32050 (
);

FILL FILL_0__13356_ (
);

INVX1 _13641_ (
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_4149_)
);

NOR2X1 _13221_ (
    .A(\datapath_1.a3 [0]),
    .B(_3763_),
    .Y(_3764_)
);

FILL FILL_5__9393_ (
);

FILL FILL_1__6913_ (
);

FILL FILL_6__12270_ (
);

FILL FILL_3__6839_ (
);

FILL FILL_5__16128_ (
);

FILL FILL_5__11683_ (
);

FILL FILL_1__9385_ (
);

FILL FILL_5__11263_ (
);

FILL FILL_2__16155_ (
);

FILL SFILL99400x64050 (
);

FILL SFILL38760x48050 (
);

FILL FILL_4__10676_ (
);

FILL SFILL69160x39050 (
);

FILL FILL_4__10256_ (
);

FILL FILL_2__11290_ (
);

FILL FILL_1__15988_ (
);

FILL FILL_1__15568_ (
);

FILL FILL_1__15148_ (
);

FILL FILL_5__7706_ (
);

FILL FILL_2_BUFX2_insert400 (
);

FILL FILL_2_BUFX2_insert401 (
);

FILL FILL_1__10283_ (
);

FILL FILL_2_BUFX2_insert402 (
);

NAND3X1 _14846_ (
    .A(_5318_),
    .B(_5321_),
    .C(_5328_),
    .Y(_5329_)
);

FILL FILL_2_BUFX2_insert403 (
);

FILL FILL_2_BUFX2_insert404 (
);

OAI22X1 _14426_ (
    .A(_4916_),
    .B(_3955__bF$buf4),
    .C(_3924__bF$buf2),
    .D(_4917_),
    .Y(_4918_)
);

INVX1 _14006_ (
    .A(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_4507_)
);

FILL FILL_2_BUFX2_insert405 (
);

FILL FILL_2_BUFX2_insert406 (
);

FILL FILL_2_BUFX2_insert407 (
);

FILL FILL_0__7290_ (
);

FILL FILL_2_BUFX2_insert408 (
);

FILL FILL_2_BUFX2_insert409 (
);

FILL FILL_0__15922_ (
);

FILL FILL_0__15502_ (
);

FILL FILL_5__12888_ (
);

FILL FILL_5__12468_ (
);

FILL FILL_5__12048_ (
);

FILL FILL_3__13082_ (
);

FILL SFILL69080x5050 (
);

FILL FILL_4__8595_ (
);

FILL FILL_2__12495_ (
);

FILL FILL_2__12075_ (
);

FILL SFILL8520x1050 (
);

FILL FILL_1__11488_ (
);

FILL FILL_1__11068_ (
);

FILL FILL_4__12402_ (
);

FILL FILL_0__8495_ (
);

INVX1 _10766_ (
    .A(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_1968_)
);

FILL FILL_0__8075_ (
);

FILL FILL_6__9462_ (
);

DFFSR _10346_ (
    .Q(\datapath_1.regfile_1.regOut[27] [20]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1693_[20])
);

FILL FILL_3__11815_ (
);

FILL FILL_4__15294_ (
);

FILL FILL_4__6908_ (
);

FILL FILL_2__10808_ (
);

FILL FILL_2__9874_ (
);

FILL SFILL99320x26050 (
);

FILL FILL_0__11842_ (
);

FILL FILL_2__9034_ (
);

FILL FILL_3__14287_ (
);

FILL FILL_0__11422_ (
);

FILL FILL_0__11002_ (
);

FILL SFILL89400x62050 (
);

FILL FILL_5__14614_ (
);

FILL SFILL28760x46050 (
);

FILL SFILL59160x37050 (
);

OAI21X1 _8914_ (
    .A(_1037_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1038_),
    .Y(_978_[30])
);

FILL FILL_1__7871_ (
);

FILL FILL_1__7451_ (
);

FILL FILL_1__7031_ (
);

FILL FILL_4__13607_ (
);

FILL FILL_2__14641_ (
);

FILL FILL_2__14221_ (
);

FILL FILL_3__7377_ (
);

FILL FILL_5_CLKBUF1_insert190 (
);

FILL FILL_5_CLKBUF1_insert191 (
);

FILL FILL_5_CLKBUF1_insert192 (
);

FILL FILL_5_CLKBUF1_insert193 (
);

FILL FILL_1__13634_ (
);

FILL FILL_1__13214_ (
);

FILL FILL_5_CLKBUF1_insert194 (
);

FILL FILL_4__16079_ (
);

FILL FILL_5_CLKBUF1_insert195 (
);

FILL FILL_5_CLKBUF1_insert196 (
);

FILL FILL_5_CLKBUF1_insert197 (
);

FILL FILL_5_CLKBUF1_insert198 (
);

FILL FILL_1_BUFX2_insert420 (
);

FILL FILL_5_CLKBUF1_insert199 (
);

FILL FILL_1_BUFX2_insert421 (
);

FILL SFILL89320x69050 (
);

FILL FILL_0__12627_ (
);

OAI21X1 _12912_ (
    .A(_3612_),
    .B(vdd),
    .C(_3613_),
    .Y(_3555_[29])
);

FILL FILL_1_BUFX2_insert422 (
);

FILL FILL_0__12207_ (
);

FILL FILL_1_BUFX2_insert423 (
);

FILL FILL_1_BUFX2_insert424 (
);

FILL FILL_1_BUFX2_insert425 (
);

FILL FILL_6__16406_ (
);

FILL FILL_1_BUFX2_insert426 (
);

FILL FILL_1_BUFX2_insert427 (
);

FILL FILL_6_BUFX2_insert981 (
);

FILL FILL_5__8244_ (
);

FILL FILL_1_BUFX2_insert428 (
);

FILL FILL_1_BUFX2_insert429 (
);

OAI22X1 _15384_ (
    .A(_5526__bF$buf3),
    .B(_4385_),
    .C(_4360_),
    .D(_5527__bF$buf4),
    .Y(_5856_)
);

FILL FILL_0__15099_ (
);

FILL FILL_6_BUFX2_insert986 (
);

FILL FILL_5__15819_ (
);

FILL FILL_3__16013_ (
);

FILL FILL_5__10954_ (
);

FILL FILL_5__10534_ (
);

FILL FILL_1__8656_ (
);

FILL FILL_5__10114_ (
);

FILL FILL_1__8236_ (
);

FILL FILL_2__15846_ (
);

FILL FILL_2__15426_ (
);

FILL FILL_2__15006_ (
);

FILL FILL_0__16040_ (
);

FILL FILL_2__10981_ (
);

FILL FILL_2__10561_ (
);

FILL FILL_2__10141_ (
);

FILL FILL_1__14839_ (
);

FILL FILL_1__14419_ (
);

FILL FILL_3__9523_ (
);

FILL FILL_3__9103_ (
);

FILL SFILL33960x64050 (
);

FILL FILL_0__6981_ (
);

FILL FILL_5__9869_ (
);

FILL FILL_5__9029_ (
);

FILL FILL_4__13780_ (
);

FILL FILL_6__12326_ (
);

FILL FILL_4__13360_ (
);

INVX1 _16169_ (
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_6621_)
);

FILL FILL_2__7940_ (
);

FILL FILL_5__11739_ (
);

FILL FILL_3__12773_ (
);

FILL FILL_5__11319_ (
);

FILL FILL_2__7100_ (
);

FILL FILL_3__12353_ (
);

FILL SFILL18760x44050 (
);

FILL FILL_4__7866_ (
);

FILL FILL_4__7446_ (
);

FILL FILL_2__11766_ (
);

FILL FILL_2__11346_ (
);

FILL FILL_0__12380_ (
);

FILL SFILL54120x18050 (
);

FILL FILL_1__10759_ (
);

FILL FILL_2_CLKBUF1_insert140 (
);

FILL FILL_2_CLKBUF1_insert141 (
);

FILL FILL_2_CLKBUF1_insert142 (
);

FILL FILL_5__15992_ (
);

FILL FILL_2_CLKBUF1_insert143 (
);

FILL FILL_5__15572_ (
);

FILL FILL_2_CLKBUF1_insert144 (
);

FILL FILL_5__15152_ (
);

OAI21X1 _9872_ (
    .A(_1513_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1514_),
    .Y(_1498_[8])
);

FILL FILL_2_CLKBUF1_insert145 (
);

FILL FILL_0__7346_ (
);

FILL FILL_6__8733_ (
);

FILL FILL_2_CLKBUF1_insert146 (
);

DFFSR _9452_ (
    .Q(\datapath_1.regfile_1.regOut[20] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1238_[22])
);

FILL SFILL79320x67050 (
);

NAND2X1 _9032_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1097_)
);

FILL FILL_2_CLKBUF1_insert147 (
);

FILL FILL_2_CLKBUF1_insert148 (
);

FILL FILL_2_CLKBUF1_insert149 (
);

FILL FILL_4__14985_ (
);

FILL FILL_4__14565_ (
);

FILL FILL_1__11700_ (
);

FILL FILL_4__14145_ (
);

AOI22X1 _12089_ (
    .A(\datapath_1.ALUResult [25]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3113_)
);

FILL FILL_3__13978_ (
);

FILL FILL_2__8725_ (
);

FILL FILL_3__13558_ (
);

FILL FILL_1__14592_ (
);

FILL FILL_3__13138_ (
);

FILL FILL_1__14172_ (
);

FILL SFILL39160x78050 (
);

FILL FILL_6_BUFX2_insert1022 (
);

FILL FILL_0__13585_ (
);

INVX1 _13870_ (
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_4374_)
);

FILL FILL_0__13165_ (
);

NOR2X1 _13450_ (
    .A(_3961_),
    .B(_3956_),
    .Y(_3962_)
);

NAND2X1 _13030_ (
    .A(vdd),
    .B(\datapath_1.rd2 [26]),
    .Y(_3672_)
);

FILL FILL_6_BUFX2_insert1027 (
);

FILL FILL_2__13912_ (
);

FILL FILL_5__16357_ (
);

FILL FILL_5__11492_ (
);

FILL FILL_5__11072_ (
);

FILL FILL_1__12905_ (
);

FILL FILL_2__16384_ (
);

FILL SFILL79320x22050 (
);

FILL FILL_0__9912_ (
);

FILL FILL_4__10065_ (
);

FILL FILL_1__15797_ (
);

FILL FILL_1__15377_ (
);

FILL FILL_5__7935_ (
);

AOI22X1 _14655_ (
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_5142_)
);

INVX1 _14235_ (
    .A(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_4731_)
);

FILL FILL_3__15704_ (
);

FILL FILL_1__7927_ (
);

FILL FILL_1__7507_ (
);

FILL SFILL79240x29050 (
);

FILL FILL_0__15731_ (
);

FILL FILL_0__15311_ (
);

FILL FILL_5__12697_ (
);

FILL FILL_5__12277_ (
);

OAI21X1 _6997_ (
    .A(_64_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_65_),
    .Y(_3_[31])
);

FILL FILL_1__11297_ (
);

FILL FILL_4__12631_ (
);

FILL FILL_4__12211_ (
);

NOR2X1 _10995_ (
    .A(_2112_),
    .B(_2113_),
    .Y(_2114_)
);

OAI21X1 _10575_ (
    .A(_1880_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .C(_1881_),
    .Y(_1823_[29])
);

OAI21X1 _10155_ (
    .A(_1661_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1662_),
    .Y(_1628_[17])
);

FILL FILL_3__11624_ (
);

FILL FILL_3__11204_ (
);

FILL FILL_3_BUFX2_insert1084 (
);

FILL FILL_3_BUFX2_insert1085 (
);

FILL FILL_3_BUFX2_insert1086 (
);

FILL FILL_3_BUFX2_insert1087 (
);

FILL FILL_3_BUFX2_insert1088 (
);

FILL FILL_3_BUFX2_insert1089 (
);

FILL FILL_2__9683_ (
);

FILL FILL_2__10617_ (
);

FILL FILL_2__9263_ (
);

FILL FILL_0__11651_ (
);

FILL FILL_0__11231_ (
);

FILL FILL_3__14096_ (
);

FILL FILL_2__13089_ (
);

FILL FILL_5__14843_ (
);

FILL FILL_5__14423_ (
);

FILL FILL_5__14003_ (
);

OAI21X1 _8723_ (
    .A(_930_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_931_),
    .Y(_913_[9])
);

DFFSR _8303_ (
    .Q(\datapath_1.regfile_1.regOut[11] [25]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_653_[25])
);

FILL FILL_1__7680_ (
);

FILL FILL_4__13836_ (
);

FILL FILL_2__14870_ (
);

FILL FILL_4__13416_ (
);

FILL FILL_2__14450_ (
);

FILL FILL_2__14030_ (
);

FILL FILL_0__9089_ (
);

FILL FILL_3__7186_ (
);

FILL FILL_3__12829_ (
);

FILL FILL_1__13863_ (
);

FILL FILL_3__12409_ (
);

FILL FILL_1__13443_ (
);

FILL FILL_1__13023_ (
);

FILL FILL_4_CLKBUF1_insert180 (
);

FILL FILL_4_CLKBUF1_insert181 (
);

FILL SFILL69240x27050 (
);

FILL FILL_0__12856_ (
);

FILL FILL_4_CLKBUF1_insert182 (
);

OAI21X1 _12721_ (
    .A(_3505_),
    .B(IRWrite_bF$buf1),
    .C(_3506_),
    .Y(_3490_[8])
);

FILL FILL_0__12436_ (
);

FILL FILL_4_CLKBUF1_insert183 (
);

FILL FILL_0__12016_ (
);

FILL FILL_4_CLKBUF1_insert184 (
);

AOI22X1 _12301_ (
    .A(_2_[21]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3265_)
);

FILL FILL_4_CLKBUF1_insert185 (
);

FILL FILL_4_CLKBUF1_insert186 (
);

FILL FILL_5__8893_ (
);

FILL FILL_4_CLKBUF1_insert187 (
);

FILL FILL_5__8473_ (
);

FILL FILL_4_CLKBUF1_insert188 (
);

FILL FILL_4_CLKBUF1_insert189 (
);

OAI22X1 _15193_ (
    .A(_4106_),
    .B(_5539__bF$buf4),
    .C(_5527__bF$buf4),
    .D(_4112_),
    .Y(_5670_)
);

FILL FILL_5__15628_ (
);

FILL FILL_5__15208_ (
);

FILL FILL_3__16242_ (
);

NAND2X1 _9928_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1552_)
);

NAND2X1 _9508_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1333_)
);

FILL FILL_5__10763_ (
);

FILL FILL_1__8885_ (
);

FILL FILL_1__8465_ (
);

FILL FILL_2__15655_ (
);

FILL SFILL99400x59050 (
);

FILL FILL_2__15235_ (
);

FILL FILL_4__6890_ (
);

FILL FILL_2__10790_ (
);

FILL FILL_2__10370_ (
);

FILL FILL_1__14648_ (
);

FILL FILL_1__14228_ (
);

FILL FILL_3__9752_ (
);

AOI22X1 _13926_ (
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .B(_4154_),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_4429_)
);

INVX1 _13506_ (
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_4017_)
);

FILL SFILL99000x45050 (
);

FILL FILL_5__9678_ (
);

FILL SFILL104360x52050 (
);

FILL FILL_5__9258_ (
);

OAI21X1 _16398_ (
    .A(_6818_),
    .B(gnd),
    .C(_6819_),
    .Y(_6769_[25])
);

FILL FILL_5__11968_ (
);

FILL FILL_5__11548_ (
);

FILL SFILL3800x47050 (
);

FILL FILL_3__12582_ (
);

FILL FILL_5__11128_ (
);

FILL FILL_3__12162_ (
);

FILL FILL_4__7675_ (
);

FILL FILL_2__11995_ (
);

FILL FILL_2__11575_ (
);

FILL FILL_2__11155_ (
);

FILL SFILL99400x14050 (
);

FILL FILL_1__10988_ (
);

FILL FILL_1__10568_ (
);

FILL FILL_1__10148_ (
);

FILL FILL_4__11902_ (
);

FILL FILL_5__15381_ (
);

FILL FILL_0__7995_ (
);

FILL FILL_0__7575_ (
);

NAND2X1 _9681_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1428_)
);

NAND2X1 _9261_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1209_)
);

FILL FILL_1_CLKBUF1_insert130 (
);

FILL FILL_1_CLKBUF1_insert131 (
);

FILL FILL_4__14794_ (
);

FILL FILL_1_CLKBUF1_insert132 (
);

FILL FILL_1_CLKBUF1_insert133 (
);

FILL FILL_4__14374_ (
);

FILL FILL_1_CLKBUF1_insert134 (
);

FILL FILL_1_CLKBUF1_insert135 (
);

FILL FILL_1_CLKBUF1_insert136 (
);

FILL FILL_1_CLKBUF1_insert137 (
);

FILL FILL_1_CLKBUF1_insert138 (
);

FILL FILL_2__8954_ (
);

FILL FILL_0__10922_ (
);

FILL FILL_3__13787_ (
);

FILL FILL_1_CLKBUF1_insert139 (
);

FILL FILL_3__13367_ (
);

FILL FILL_2__8114_ (
);

FILL FILL_0__10502_ (
);

FILL FILL_0__13394_ (
);

FILL SFILL89400x57050 (
);

FILL FILL_1__6951_ (
);

FILL FILL_4__9401_ (
);

FILL FILL_2__13721_ (
);

FILL FILL_2__13301_ (
);

FILL FILL_3__6877_ (
);

FILL FILL_5__16166_ (
);

FILL FILL_4__15999_ (
);

FILL FILL_1__12714_ (
);

FILL FILL_4__15579_ (
);

FILL FILL_4__15159_ (
);

FILL FILL_2__16193_ (
);

FILL FILL_4__10294_ (
);

FILL FILL_2__9739_ (
);

FILL FILL_0__9721_ (
);

FILL FILL_0__9301_ (
);

FILL FILL_0__11707_ (
);

FILL FILL_1__15186_ (
);

FILL FILL_5__7744_ (
);

FILL FILL_5__7324_ (
);

FILL FILL_4__16100_ (
);

FILL FILL_0__14599_ (
);

OAI22X1 _14884_ (
    .A(_3884__bF$buf2),
    .B(_5364_),
    .C(_5365_),
    .D(_3925_),
    .Y(_5366_)
);

FILL FILL_6__10621_ (
);

INVX1 _14464_ (
    .A(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_4955_)
);

FILL FILL_0__14179_ (
);

INVX1 _14044_ (
    .A(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_4544_)
);

FILL FILL_3__15933_ (
);

FILL FILL_3__15513_ (
);

FILL SFILL89400x12050 (
);

FILL FILL_1__7736_ (
);

FILL FILL_1__7316_ (
);

FILL SFILL94280x63050 (
);

FILL FILL_2__14926_ (
);

FILL FILL_0__15960_ (
);

FILL FILL_2__14506_ (
);

FILL FILL_0__15540_ (
);

FILL FILL_0__15120_ (
);

FILL FILL_5__12086_ (
);

FILL FILL_1__13919_ (
);

FILL FILL_4__11499_ (
);

FILL FILL_4__11079_ (
);

FILL FILL_3__8603_ (
);

FILL SFILL33960x59050 (
);

FILL SFILL89320x19050 (
);

FILL FILL_5__8529_ (
);

FILL FILL_5__8109_ (
);

NAND2X1 _15669_ (
    .A(\datapath_1.regfile_1.regOut[23] [15]),
    .B(_5649_),
    .Y(_6134_)
);

FILL FILL_4__12860_ (
);

OAI22X1 _15249_ (
    .A(_4183_),
    .B(_5548__bF$buf3),
    .C(_5489__bF$buf2),
    .D(_5724_),
    .Y(_5725_)
);

FILL FILL_4__12440_ (
);

FILL FILL_4__12020_ (
);

OAI21X1 _10384_ (
    .A(_1773_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1774_),
    .Y(_1758_[8])
);

FILL FILL_6__9080_ (
);

FILL FILL_5__10819_ (
);

FILL FILL_3__11853_ (
);

FILL SFILL94200x61050 (
);

FILL SFILL18760x39050 (
);

FILL FILL_6__14298_ (
);

FILL FILL_3__11433_ (
);

FILL FILL_3__11013_ (
);

FILL FILL_4__6946_ (
);

FILL FILL_0__16325_ (
);

FILL FILL_0__11880_ (
);

FILL FILL_2__10426_ (
);

FILL FILL_2__9492_ (
);

FILL FILL_0__11460_ (
);

FILL FILL_2__10006_ (
);

FILL FILL_0__11040_ (
);

FILL FILL_3__9808_ (
);

FILL FILL_5__14652_ (
);

FILL FILL_5__14232_ (
);

FILL FILL_0__6846_ (
);

OAI21X1 _8952_ (
    .A(_1106_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .C(_1107_),
    .Y(_1043_[0])
);

FILL FILL_6__7813_ (
);

NAND2X1 _8532_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_845_)
);

FILL SFILL8680x80050 (
);

NAND2X1 _8112_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_626_)
);

FILL FILL_4__13645_ (
);

FILL FILL_4__13225_ (
);

NAND3X1 _11589_ (
    .A(_2462__bF$buf1),
    .B(_2695_),
    .C(_2690_),
    .Y(_2696_)
);

NOR2X1 _11169_ (
    .A(_2285_),
    .B(_2287_),
    .Y(_2288_)
);

FILL FILL_2__7805_ (
);

FILL FILL_3__12638_ (
);

FILL FILL_1__13672_ (
);

FILL FILL_3__12218_ (
);

FILL FILL_1__13252_ (
);

FILL FILL_1_BUFX2_insert800 (
);

FILL FILL_1_BUFX2_insert801 (
);

DFFSR _12950_ (
    .Q(\datapath_1.a [31]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_3555_[31])
);

FILL FILL_1_BUFX2_insert802 (
);

NAND2X1 _12530_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [30]),
    .Y(_3420_)
);

FILL FILL_0__12245_ (
);

FILL FILL_1_BUFX2_insert803 (
);

NAND3X1 _12110_ (
    .A(_3126_),
    .B(_3127_),
    .C(_3128_),
    .Y(\datapath_1.mux_pcsrc.dout [30])
);

FILL FILL_1_BUFX2_insert804 (
);

FILL FILL_1_BUFX2_insert805 (
);

FILL FILL_1_BUFX2_insert806 (
);

FILL FILL_1_BUFX2_insert807 (
);

FILL FILL_1_BUFX2_insert808 (
);

FILL FILL_1_BUFX2_insert809 (
);

FILL FILL_5__15857_ (
);

FILL FILL_5__15437_ (
);

FILL FILL_5__15017_ (
);

NAND2X1 _9737_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1445_)
);

FILL FILL_3__16051_ (
);

DFFSR _9317_ (
    .Q(\datapath_1.regfile_1.regOut[19] [15]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_1173_[15])
);

FILL FILL_5__10992_ (
);

FILL FILL_5__10572_ (
);

FILL FILL_1__8694_ (
);

FILL FILL_5__10152_ (
);

FILL FILL_1__8274_ (
);

FILL FILL_2__15884_ (
);

FILL FILL_2__15464_ (
);

FILL FILL_2__15044_ (
);

FILL FILL_1__14877_ (
);

FILL FILL_1__14457_ (
);

FILL FILL_1__14037_ (
);

FILL FILL_3__9981_ (
);

FILL FILL_3__9141_ (
);

AOI22X1 _13735_ (
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .B(_3891__bF$buf2),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_4242_)
);

NAND2X1 _13315_ (
    .A(_3834_),
    .B(_3785_),
    .Y(_3847_)
);

FILL FILL_5__9487_ (
);

FILL FILL_6__12784_ (
);

FILL SFILL114840x56050 (
);

FILL FILL_0__14811_ (
);

FILL FILL_1__9899_ (
);

FILL FILL_5__11777_ (
);

FILL FILL_5__11357_ (
);

FILL FILL_1__9479_ (
);

FILL FILL_3__12391_ (
);

FILL FILL_2__16249_ (
);

FILL FILL_4__7484_ (
);

FILL FILL_4__7064_ (
);

FILL FILL_2__11384_ (
);

FILL SFILL114440x42050 (
);

FILL FILL_1__10797_ (
);

FILL FILL_1__10377_ (
);

FILL FILL_4__11711_ (
);

FILL FILL_5__15190_ (
);

NAND2X1 _9490_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1321_)
);

FILL FILL_6__8351_ (
);

DFFSR _9070_ (
    .Q(\datapath_1.regfile_1.regOut[17] [24]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_1043_[24])
);

FILL FILL_3__10704_ (
);

FILL FILL_4__14183_ (
);

FILL FILL_2__8763_ (
);

FILL FILL_3__13596_ (
);

FILL FILL_2__8343_ (
);

FILL FILL_0__10311_ (
);

FILL SFILL74600x71050 (
);

FILL FILL_4__8269_ (
);

FILL FILL_2__12589_ (
);

FILL FILL_2__12169_ (
);

FILL FILL_5__13923_ (
);

FILL FILL_5__13503_ (
);

OAI21X1 _7803_ (
    .A(_459_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_460_),
    .Y(_458_[1])
);

FILL FILL_4_BUFX2_insert310 (
);

FILL FILL_4_BUFX2_insert311 (
);

FILL FILL_4__9630_ (
);

FILL FILL_4__12916_ (
);

FILL FILL_4__9210_ (
);

FILL FILL_4_BUFX2_insert312 (
);

FILL FILL_4_BUFX2_insert313 (
);

FILL FILL_2__13950_ (
);

FILL FILL_5__16395_ (
);

FILL FILL_4_BUFX2_insert314 (
);

FILL FILL_2__13530_ (
);

FILL FILL_0__8589_ (
);

FILL FILL_2__13110_ (
);

FILL FILL_4_BUFX2_insert315 (
);

FILL FILL_4_BUFX2_insert316 (
);

FILL FILL_4_BUFX2_insert317 (
);

FILL FILL_6__9136_ (
);

FILL FILL_4_BUFX2_insert318 (
);

FILL FILL_3__11909_ (
);

FILL FILL_4_BUFX2_insert319 (
);

FILL FILL_4__15388_ (
);

FILL FILL_1__12523_ (
);

FILL FILL_1__12103_ (
);

FILL FILL_2__9548_ (
);

FILL FILL_0__11936_ (
);

FILL FILL_0__9530_ (
);

FILL FILL_0__11516_ (
);

FILL FILL_2__9128_ (
);

NAND2X1 _11801_ (
    .A(_2368_),
    .B(_2850_),
    .Y(_2893_)
);

FILL FILL_0__9110_ (
);

FILL FILL_5__7973_ (
);

FILL FILL_6__15715_ (
);

FILL FILL_5__7553_ (
);

AOI22X1 _14693_ (
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .B(_4154_),
    .C(_4051__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_5179_)
);

AOI22X1 _14273_ (
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .B(_3891__bF$buf2),
    .C(_4051__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_4768_)
);

FILL FILL_5__14708_ (
);

FILL FILL_3__15742_ (
);

FILL FILL_3__15322_ (
);

FILL FILL_1__7965_ (
);

FILL FILL_1__7545_ (
);

FILL FILL_1__7125_ (
);

FILL FILL_2__14735_ (
);

FILL FILL_2__14315_ (
);

FILL FILL_1__13728_ (
);

FILL FILL_1__13308_ (
);

FILL FILL_3__8832_ (
);

FILL SFILL104360x47050 (
);

FILL FILL_5__8758_ (
);

FILL FILL_5__8338_ (
);

INVX1 _15898_ (
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_6357_)
);

FILL FILL_6__11635_ (
);

INVX1 _15478_ (
    .A(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_5948_)
);

NAND2X1 _15058_ (
    .A(_5537_),
    .B(_5529_),
    .Y(_5538_)
);

FILL FILL_3__16107_ (
);

NAND2X1 _10193_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1688_)
);

FILL FILL_5__10628_ (
);

FILL FILL_3__11662_ (
);

FILL FILL_3__11242_ (
);

FILL FILL_0__16134_ (
);

FILL FILL_2__10655_ (
);

FILL FILL_2__10235_ (
);

FILL SFILL3400x28050 (
);

FILL FILL_3_BUFX2_insert330 (
);

FILL FILL_3__9617_ (
);

FILL FILL_3_BUFX2_insert331 (
);

FILL FILL_5__14881_ (
);

FILL FILL_3_BUFX2_insert332 (
);

FILL FILL_5__14461_ (
);

FILL FILL_3_BUFX2_insert333 (
);

FILL FILL_5__14041_ (
);

FILL FILL_3_BUFX2_insert334 (
);

FILL FILL112440x53050 (
);

NAND2X1 _8761_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_957_)
);

FILL FILL_3_BUFX2_insert335 (
);

FILL FILL_3_BUFX2_insert336 (
);

NAND2X1 _8341_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_738_)
);

FILL FILL_3_BUFX2_insert337 (
);

FILL FILL_3_BUFX2_insert338 (
);

FILL FILL_4__13874_ (
);

FILL FILL_3_BUFX2_insert339 (
);

FILL FILL_4__13454_ (
);

FILL FILL_4__13034_ (
);

FILL SFILL89960x9050 (
);

OAI21X1 _11398_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(_2206_),
    .C(_2514_),
    .Y(_2515_)
);

FILL FILL_2__7614_ (
);

FILL FILL_3__12867_ (
);

FILL FILL_3__12447_ (
);

FILL FILL_3__12027_ (
);

FILL FILL_1__13481_ (
);

FILL FILL_0__12894_ (
);

FILL FILL_0__12474_ (
);

FILL FILL_0__12054_ (
);

FILL FILL_5__8091_ (
);

FILL FILL_4__8901_ (
);

FILL FILL_5__15666_ (
);

FILL FILL_5__15246_ (
);

DFFSR _9966_ (
    .Q(\datapath_1.regfile_1.regOut[24] [24]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1498_[24])
);

FILL FILL_3__16280_ (
);

INVX1 _9546_ (
    .A(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_1358_)
);

INVX1 _9126_ (
    .A(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_1139_)
);

FILL FILL_5__10381_ (
);

FILL FILL_1__8083_ (
);

FILL FILL_4__14659_ (
);

FILL FILL_4__14239_ (
);

FILL FILL_2__15693_ (
);

FILL FILL_2__15273_ (
);

FILL FILL_1__14686_ (
);

FILL FILL_1__14266_ (
);

FILL FILL_0_BUFX2_insert460 (
);

FILL FILL_0_BUFX2_insert461 (
);

FILL FILL_4__15600_ (
);

FILL FILL_0_BUFX2_insert462 (
);

FILL FILL_3__9790_ (
);

FILL FILL_0_BUFX2_insert463 (
);

FILL FILL_0__13679_ (
);

FILL FILL_3__9370_ (
);

FILL FILL_0_BUFX2_insert464 (
);

INVX1 _13964_ (
    .A(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_4466_)
);

FILL FILL_0__13259_ (
);

NAND3X1 _13544_ (
    .A(_4052_),
    .B(_4053_),
    .C(_4050_),
    .Y(_4054_)
);

FILL FILL_0_BUFX2_insert465 (
);

FILL FILL_0_BUFX2_insert466 (
);

INVX1 _13124_ (
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_3714_)
);

FILL FILL_0_BUFX2_insert467 (
);

FILL FILL_0_BUFX2_insert468 (
);

FILL FILL_0_BUFX2_insert469 (
);

FILL FILL_5__9296_ (
);

FILL SFILL94280x58050 (
);

FILL FILL_6__12593_ (
);

FILL FILL_0__14620_ (
);

FILL FILL_0__14200_ (
);

FILL FILL_5__11586_ (
);

FILL FILL_1__9288_ (
);

FILL FILL_5__11166_ (
);

FILL FILL_2__16058_ (
);

FILL FILL_4__10999_ (
);

FILL FILL_4__7293_ (
);

FILL FILL_4__10579_ (
);

FILL FILL_4__10159_ (
);

FILL FILL_2__11193_ (
);

FILL FILL_5__7609_ (
);

FILL FILL_1__10186_ (
);

FILL FILL_4__11940_ (
);

OAI22X1 _14749_ (
    .A(_5233_),
    .B(_3936__bF$buf4),
    .C(_3905__bF$buf0),
    .D(_5232_),
    .Y(_5234_)
);

INVX1 _14329_ (
    .A(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_4823_)
);

FILL FILL_4__11520_ (
);

FILL FILL_4__11100_ (
);

FILL FILL_0__7193_ (
);

FILL FILL_1__16412_ (
);

FILL FILL_3__10933_ (
);

FILL FILL_3__10513_ (
);

FILL FILL_0__15825_ (
);

FILL FILL_0__15405_ (
);

FILL SFILL94280x13050 (
);

FILL FILL_2__8992_ (
);

FILL FILL_0__10960_ (
);

FILL FILL_2__8572_ (
);

FILL FILL_0__10540_ (
);

FILL FILL_0__10120_ (
);

FILL FILL_4__8498_ (
);

FILL FILL_4__8078_ (
);

FILL FILL_2__12398_ (
);

FILL FILL_5__13732_ (
);

FILL FILL_5__13312_ (
);

FILL SFILL8680x75050 (
);

NAND2X1 _7612_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_374_)
);

FILL FILL_4__12725_ (
);

FILL FILL_4__12305_ (
);

FILL FILL_0__8398_ (
);

NAND2X1 _10669_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1924_)
);

NAND2X1 _10249_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1705_)
);

FILL FILL_3__11718_ (
);

FILL FILL_1__12752_ (
);

FILL FILL_4__15197_ (
);

FILL FILL_1__12332_ (
);

FILL SFILL84280x56050 (
);

FILL FILL_2__9777_ (
);

FILL FILL_2__9357_ (
);

FILL FILL_0__11745_ (
);

FILL FILL_0__11325_ (
);

NAND2X1 _11610_ (
    .A(_2715_),
    .B(_2701_),
    .Y(_2716_)
);

FILL FILL_5__7362_ (
);

FILL FILL_5__14937_ (
);

INVX1 _14082_ (
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_4581_)
);

FILL FILL_3__15971_ (
);

FILL FILL_5__14517_ (
);

FILL FILL_3__15551_ (
);

FILL SFILL8600x73050 (
);

DFFSR _8817_ (
    .Q(\datapath_1.regfile_1.regOut[15] [27]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_913_[27])
);

FILL FILL_3__15131_ (
);

FILL FILL_1__7354_ (
);

FILL FILL_2__14964_ (
);

FILL SFILL8680x30050 (
);

FILL FILL_2__14544_ (
);

FILL FILL_2__14124_ (
);

FILL FILL_1__13957_ (
);

FILL FILL_1__13537_ (
);

FILL FILL_1__13117_ (
);

FILL SFILL23560x38050 (
);

FILL FILL_3__8641_ (
);

DFFSR _12815_ (
    .Q(\datapath_1.PCJump [26]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3490_[24])
);

FILL FILL_3__8221_ (
);

FILL SFILL84280x11050 (
);

FILL FILL_5__8987_ (
);

FILL FILL_5__8567_ (
);

FILL FILL_6__16309_ (
);

FILL FILL_5__8147_ (
);

FILL SFILL13640x74050 (
);

INVX1 _15287_ (
    .A(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_5762_)
);

FILL FILL_3__16336_ (
);

FILL FILL_1__8979_ (
);

FILL FILL_5__10437_ (
);

FILL FILL_3__11891_ (
);

FILL FILL_5__10017_ (
);

FILL FILL_1__8139_ (
);

FILL FILL_3__11471_ (
);

FILL FILL_3__11051_ (
);

FILL FILL_2__15749_ (
);

FILL FILL_2__15329_ (
);

FILL FILL_4__6984_ (
);

FILL FILL_0__16363_ (
);

FILL FILL_2__10884_ (
);

FILL SFILL114440x37050 (
);

FILL FILL_2__10044_ (
);

FILL FILL_1__9920_ (
);

FILL FILL_1__9500_ (
);

FILL FILL_3__9846_ (
);

FILL FILL_3__9426_ (
);

FILL SFILL109560x7050 (
);

FILL FILL_3__9006_ (
);

FILL FILL_5__14690_ (
);

FILL FILL_0__6884_ (
);

FILL FILL_5__14270_ (
);

FILL SFILL74280x54050 (
);

NAND2X1 _8990_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1069_)
);

NAND2X1 _8570_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_850_)
);

FILL FILL_6__7431_ (
);

DFFSR _8150_ (
    .Q(\datapath_1.regfile_1.regOut[10] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_588_[0])
);

FILL FILL_6__12649_ (
);

FILL FILL_4__13683_ (
);

FILL FILL_6__12229_ (
);

FILL FILL_4__13263_ (
);

FILL FILL_2__7843_ (
);

FILL FILL_2__7423_ (
);

FILL FILL_3__12256_ (
);

FILL FILL_1__13290_ (
);

FILL FILL_4__7349_ (
);

FILL FILL_2__11669_ (
);

FILL FILL_2__11249_ (
);

FILL FILL_0__12283_ (
);

FILL FILL_4__8710_ (
);

FILL FILL_5__15895_ (
);

FILL FILL_2__12610_ (
);

FILL FILL_5__15475_ (
);

FILL FILL_5__15055_ (
);

FILL SFILL13560x36050 (
);

INVX1 _9775_ (
    .A(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_1470_)
);

FILL FILL_0__7249_ (
);

INVX1 _9355_ (
    .A(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_1251_)
);

FILL FILL_6__8216_ (
);

FILL FILL_5__10190_ (
);

FILL FILL_4__14888_ (
);

FILL FILL_4__14468_ (
);

FILL FILL_1__11603_ (
);

FILL FILL_4__14048_ (
);

FILL FILL_2__15082_ (
);

FILL FILL_0__8610_ (
);

FILL FILL_2__8628_ (
);

FILL FILL_2__8208_ (
);

FILL SFILL78520x60050 (
);

FILL FILL_1__14495_ (
);

FILL FILL_1__14075_ (
);

INVX1 _13773_ (
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_4279_)
);

FILL FILL_0__13488_ (
);

NAND3X1 _13353_ (
    .A(\datapath_1.a3 [3]),
    .B(_3856_),
    .C(_3767_),
    .Y(_3870_)
);

FILL FILL_3__14822_ (
);

FILL FILL_3__14402_ (
);

FILL FILL_4__9915_ (
);

FILL FILL_2__13815_ (
);

FILL FILL_5__11395_ (
);

FILL FILL_1__9097_ (
);

FILL FILL_2__16287_ (
);

FILL FILL_4__10388_ (
);

FILL FILL_5__7838_ (
);

FILL FILL_5__7418_ (
);

AOI21X1 _14978_ (
    .A(_5458_),
    .B(_5433_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [31])
);

AOI22X1 _14558_ (
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_5047_)
);

OAI22X1 _14138_ (
    .A(_4634_),
    .B(_3931__bF$buf2),
    .C(_3959_),
    .D(_4635_),
    .Y(_4636_)
);

FILL FILL_3__15607_ (
);

FILL FILL_1__16221_ (
);

FILL FILL_3__10742_ (
);

FILL FILL_3__10322_ (
);

FILL FILL_0__15634_ (
);

FILL FILL_0__15214_ (
);

FILL FILL_2__8381_ (
);

FILL SFILL64200x50050 (
);

FILL FILL_5__13961_ (
);

FILL FILL_5__13541_ (
);

FILL FILL112440x48050 (
);

FILL FILL_5__13121_ (
);

NAND2X1 _7841_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_486_)
);

NAND2X1 _7421_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_267_)
);

DFFSR _7001_ (
    .Q(\datapath_1.regfile_1.regOut[1] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_3_[3])
);

FILL FILL_4__12954_ (
);

FILL FILL_4__12534_ (
);

FILL FILL_4__12114_ (
);

NAND2X1 _10898_ (
    .A(\control_1.reg_state.dout [3]),
    .B(_2046_),
    .Y(_2047_)
);

DFFSR _10478_ (
    .Q(\datapath_1.regfile_1.regOut[28] [24]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_1758_[24])
);

INVX1 _10058_ (
    .A(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_1618_)
);

FILL FILL_3__11947_ (
);

FILL FILL_1__12981_ (
);

FILL FILL_3__11527_ (
);

FILL FILL_3__11107_ (
);

FILL FILL_1__12141_ (
);

FILL FILL112040x34050 (
);

FILL FILL_0__11974_ (
);

FILL FILL_2__9166_ (
);

FILL FILL_0__11554_ (
);

FILL FILL_0__11134_ (
);

FILL FILL_5__7591_ (
);

FILL FILL_5__7171_ (
);

FILL FILL_5__14746_ (
);

FILL FILL_3__15780_ (
);

FILL FILL_5__14326_ (
);

FILL FILL_3__15360_ (
);

INVX1 _8626_ (
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_887_)
);

INVX1 _8206_ (
    .A(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_668_)
);

FILL FILL_1__7583_ (
);

FILL FILL_1__7163_ (
);

FILL FILL_4__13739_ (
);

FILL FILL_4__13319_ (
);

FILL FILL_2__14773_ (
);

FILL FILL_2__14353_ (
);

FILL FILL_3__7089_ (
);

FILL FILL_1__13766_ (
);

FILL FILL_1__13346_ (
);

FILL FILL_3__8870_ (
);

FILL FILL_0__12759_ (
);

FILL FILL_3__8450_ (
);

INVX1 _12624_ (
    .A(\datapath_1.Data [19]),
    .Y(_3462_)
);

FILL FILL_0__12339_ (
);

OAI21X1 _12204_ (
    .A(_3188_),
    .B(ALUSrcA_bF$buf6),
    .C(_3189_),
    .Y(\datapath_1.alu_1.ALUInA [29])
);

FILL FILL_5__8376_ (
);

AOI21X1 _15096_ (
    .A(\datapath_1.regfile_1.regOut[3] [1]),
    .B(_5494_),
    .C(_5574_),
    .Y(_5575_)
);

FILL FILL_0__13700_ (
);

FILL FILL_3__16145_ (
);

FILL FILL_5__10666_ (
);

FILL FILL_1__8788_ (
);

FILL FILL_1__8368_ (
);

FILL FILL_5__10246_ (
);

FILL FILL_3__11280_ (
);

FILL FILL_2__15978_ (
);

FILL FILL_2__15558_ (
);

FILL FILL_2__15138_ (
);

FILL FILL_0__16172_ (
);

FILL FILL_2__10693_ (
);

FILL FILL_2__10273_ (
);

FILL SFILL23720x64050 (
);

FILL FILL_3__9655_ (
);

FILL FILL_3_BUFX2_insert710 (
);

NOR2X1 _13829_ (
    .A(_4333_),
    .B(_3971__bF$buf1),
    .Y(_4334_)
);

FILL FILL_3_BUFX2_insert711 (
);

FILL FILL_3__9235_ (
);

FILL SFILL33240x14050 (
);

OAI22X1 _13409_ (
    .A(_3915_),
    .B(_3916_),
    .C(_3920_),
    .D(_3914_),
    .Y(_3921_)
);

FILL FILL_3_BUFX2_insert712 (
);

FILL FILL_3_BUFX2_insert713 (
);

FILL FILL_3_BUFX2_insert714 (
);

FILL FILL_1__15912_ (
);

FILL FILL_3_BUFX2_insert715 (
);

FILL FILL_3_BUFX2_insert716 (
);

FILL FILL_3_BUFX2_insert717 (
);

FILL FILL_3_BUFX2_insert718 (
);

FILL FILL_3_BUFX2_insert719 (
);

FILL FILL_4__13492_ (
);

FILL FILL_0__14905_ (
);

FILL SFILL23320x50050 (
);

FILL FILL_2__7232_ (
);

FILL FILL_3__12485_ (
);

FILL FILL_3__12065_ (
);

FILL SFILL105240x79050 (
);

FILL FILL_4__7998_ (
);

FILL FILL_4__7578_ (
);

FILL FILL_4__7158_ (
);

FILL FILL_2__11898_ (
);

FILL FILL_2__11478_ (
);

FILL FILL_2__11058_ (
);

FILL FILL_0__12092_ (
);

FILL FILL_4__11805_ (
);

FILL FILL_5__15284_ (
);

FILL FILL_0__7478_ (
);

DFFSR _9584_ (
    .Q(\datapath_1.regfile_1.regOut[21] [26]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_1303_[26])
);

FILL FILL_0__7058_ (
);

FILL SFILL74040x3050 (
);

OAI21X1 _9164_ (
    .A(_1163_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1164_),
    .Y(_1108_[28])
);

FILL FILL_4__14697_ (
);

FILL FILL_1__11832_ (
);

FILL FILL_4__14277_ (
);

FILL FILL_1__11412_ (
);

FILL FILL_2__8857_ (
);

FILL FILL_0__10825_ (
);

FILL FILL_0__10405_ (
);

FILL FILL_2__8017_ (
);

FILL FILL_5__6862_ (
);

FILL FILL_0_BUFX2_insert840 (
);

FILL FILL_0_BUFX2_insert841 (
);

FILL FILL_0_BUFX2_insert842 (
);

FILL FILL_0_BUFX2_insert843 (
);

FILL FILL_0_BUFX2_insert844 (
);

FILL FILL_0__13297_ (
);

NAND3X1 _13582_ (
    .A(_4089_),
    .B(_4091_),
    .C(_4088_),
    .Y(_4092_)
);

FILL FILL_0_BUFX2_insert845 (
);

OAI21X1 _13162_ (
    .A(_3738_),
    .B(PCEn_bF$buf0),
    .C(_3739_),
    .Y(_3685_[27])
);

FILL FILL_0_BUFX2_insert846 (
);

FILL FILL_0_BUFX2_insert847 (
);

FILL SFILL8600x68050 (
);

FILL FILL_3__14631_ (
);

FILL FILL_0_BUFX2_insert848 (
);

FILL FILL_3__14211_ (
);

FILL FILL_0_BUFX2_insert849 (
);

FILL FILL_1__6854_ (
);

FILL FILL_4__9724_ (
);

FILL SFILL8680x25050 (
);

FILL SFILL13720x62050 (
);

FILL FILL_2__13624_ (
);

FILL FILL_5__16069_ (
);

FILL SFILL109560x42050 (
);

FILL FILL_1__12617_ (
);

FILL FILL_2__16096_ (
);

FILL FILL_4__10197_ (
);

FILL FILL_0__9624_ (
);

FILL FILL_3__7721_ (
);

FILL FILL_3__7301_ (
);

FILL FILL_1__15089_ (
);

FILL FILL_5__7227_ (
);

FILL FILL_4__16003_ (
);

FILL SFILL13640x69050 (
);

NOR2X1 _14787_ (
    .A(_5271_),
    .B(_3954__bF$buf4),
    .Y(_5272_)
);

FILL FILL_6__10104_ (
);

NAND3X1 _14367_ (
    .A(_4851_),
    .B(_4852_),
    .C(_4859_),
    .Y(_4860_)
);

FILL SFILL69000x29050 (
);

FILL FILL_3__15836_ (
);

FILL SFILL109480x49050 (
);

FILL FILL_3__15416_ (
);

FILL FILL_1__16450_ (
);

FILL FILL_1__16030_ (
);

FILL FILL_3__10971_ (
);

FILL FILL_3__10551_ (
);

FILL FILL_1__7219_ (
);

FILL SFILL8600x23050 (
);

FILL FILL_3__10131_ (
);

FILL FILL_2__14829_ (
);

FILL FILL_2__14409_ (
);

FILL FILL_0__15863_ (
);

FILL FILL_0__15443_ (
);

FILL FILL_0__15023_ (
);

FILL FILL_2__8190_ (
);

FILL FILL_6_BUFX2_insert229 (
);

FILL SFILL109080x35050 (
);

FILL FILL_3__8506_ (
);

FILL FILL_5__13770_ (
);

FILL SFILL74280x49050 (
);

FILL FILL_5__13350_ (
);

DFFSR _7650_ (
    .Q(\datapath_1.regfile_1.regOut[6] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_328_[12])
);

INVX1 _7230_ (
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_180_)
);

FILL FILL_4__12763_ (
);

FILL FILL_4__12343_ (
);

INVX1 _10287_ (
    .A(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_1730_)
);

FILL FILL_2__6923_ (
);

FILL FILL_3__11756_ (
);

FILL FILL_1__12790_ (
);

FILL FILL_3__11336_ (
);

FILL FILL_1__12370_ (
);

FILL FILL_4__6849_ (
);

FILL FILL_0__16228_ (
);

FILL FILL_2__10749_ (
);

FILL SFILL38840x73050 (
);

FILL FILL_2__9395_ (
);

FILL FILL_0__11783_ (
);

FILL FILL_0__11363_ (
);

FILL FILL_6__15562_ (
);

FILL FILL_6__15142_ (
);

FILL FILL_5__14975_ (
);

FILL SFILL74200x47050 (
);

FILL FILL_5__14555_ (
);

FILL FILL_5__14135_ (
);

INVX1 _8855_ (
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_999_)
);

DFFSR _8435_ (
    .Q(\datapath_1.regfile_1.regOut[12] [29]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_718_[29])
);

OAI21X1 _8015_ (
    .A(_580_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .C(_581_),
    .Y(_523_[29])
);

FILL FILL_4__13968_ (
);

FILL FILL_4__13548_ (
);

FILL FILL_2__14582_ (
);

FILL FILL_4__13128_ (
);

FILL FILL_2__14162_ (
);

FILL SFILL34520x20050 (
);

FILL FILL_2__7708_ (
);

FILL FILL_1__13995_ (
);

FILL FILL112200x60050 (
);

FILL FILL_1__13575_ (
);

FILL SFILL99480x53050 (
);

FILL FILL_1__13155_ (
);

FILL SFILL44040x2050 (
);

FILL FILL_0__12988_ (
);

FILL FILL_0__12568_ (
);

INVX1 _12853_ (
    .A(\datapath_1.a [10]),
    .Y(_3574_)
);

FILL SFILL3480x72050 (
);

FILL FILL_0__12148_ (
);

INVX1 _12433_ (
    .A(ALUOut[30]),
    .Y(_3354_)
);

AOI22X1 _12013_ (
    .A(\datapath_1.ALUResult [6]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3056_)
);

FILL FILL_3__13902_ (
);

FILL FILL_5__8185_ (
);

FILL FILL_6__11482_ (
);

FILL FILL_5_BUFX2_insert240 (
);

FILL FILL_6__11062_ (
);

FILL FILL_5_BUFX2_insert241 (
);

FILL FILL_5_BUFX2_insert242 (
);

FILL FILL_5_BUFX2_insert243 (
);

FILL FILL_3__16374_ (
);

FILL FILL_5_BUFX2_insert244 (
);

FILL FILL_5_BUFX2_insert245 (
);

FILL FILL_5__10895_ (
);

FILL FILL112120x67050 (
);

FILL FILL_5_BUFX2_insert246 (
);

FILL FILL_1__8597_ (
);

FILL FILL_5_BUFX2_insert247 (
);

FILL FILL_5__10055_ (
);

FILL FILL_5_BUFX2_insert1030 (
);

FILL FILL_5_BUFX2_insert248 (
);

FILL FILL_5_BUFX2_insert1031 (
);

FILL FILL_5_BUFX2_insert1032 (
);

FILL FILL_2__15787_ (
);

FILL FILL_5_BUFX2_insert249 (
);

FILL FILL_5_BUFX2_insert1033 (
);

FILL FILL_2__15367_ (
);

FILL FILL_5_BUFX2_insert1034 (
);

FILL FILL_5_BUFX2_insert1035 (
);

FILL FILL_5_BUFX2_insert1036 (
);

FILL FILL_5_BUFX2_insert1037 (
);

FILL FILL_5_BUFX2_insert1038 (
);

FILL FILL_5_BUFX2_insert1039 (
);

FILL FILL_5__6918_ (
);

FILL FILL_3__9884_ (
);

FILL FILL_3__9464_ (
);

FILL SFILL64600x59050 (
);

INVX1 _13638_ (
    .A(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_4146_)
);

FILL FILL_3__9044_ (
);

NAND2X1 _13218_ (
    .A(_3760_),
    .B(_3758_),
    .Y(_3761_)
);

FILL FILL_1__15721_ (
);

FILL SFILL28840x71050 (
);

FILL FILL_1__15301_ (
);

FILL FILL_0__14714_ (
);

FILL FILL_2__7881_ (
);

FILL SFILL33800x54050 (
);

FILL FILL_2__7461_ (
);

FILL SFILL64200x45050 (
);

FILL FILL_2__7041_ (
);

FILL FILL_3__12294_ (
);

FILL FILL112120x22050 (
);

FILL FILL_2__11287_ (
);

FILL FILL_5__12621_ (
);

FILL FILL_5__12201_ (
);

NAND2X1 _6921_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_15_)
);

FILL FILL_2_BUFX2_insert370 (
);

FILL FILL_2_BUFX2_insert371 (
);

FILL FILL_2_BUFX2_insert372 (
);

FILL FILL_2_BUFX2_insert373 (
);

FILL FILL_2_BUFX2_insert374 (
);

FILL FILL_4__11614_ (
);

FILL FILL_2_BUFX2_insert375 (
);

FILL FILL_2_BUFX2_insert376 (
);

FILL FILL_5__15093_ (
);

FILL FILL_0__7287_ (
);

FILL FILL_2_BUFX2_insert377 (
);

OAI21X1 _9393_ (
    .A(_1275_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .C(_1276_),
    .Y(_1238_[19])
);

FILL FILL_2_BUFX2_insert378 (
);

FILL FILL_2_BUFX2_insert379 (
);

FILL FILL_1__11641_ (
);

FILL FILL_1__11221_ (
);

FILL FILL_4__14086_ (
);

FILL FILL_0__15919_ (
);

FILL FILL_2__8246_ (
);

FILL FILL_0__10634_ (
);

FILL FILL_3__13499_ (
);

FILL FILL_3__13079_ (
);

AND2X2 _13391_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3903_)
);

FILL FILL_5__13826_ (
);

FILL FILL_3__14860_ (
);

FILL FILL_5__13406_ (
);

FILL FILL_2_BUFX2_insert1090 (
);

FILL FILL_2_BUFX2_insert1091 (
);

FILL FILL_3__14440_ (
);

FILL FILL_3__14020_ (
);

INVX1 _7706_ (
    .A(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_416_)
);

FILL FILL_2_BUFX2_insert1092 (
);

FILL FILL_2_BUFX2_insert1093 (
);

FILL FILL_4__9533_ (
);

FILL FILL_4__9113_ (
);

FILL FILL_2__13853_ (
);

FILL FILL_2__13433_ (
);

FILL FILL_5__16298_ (
);

FILL FILL_2__13013_ (
);

FILL SFILL54600x57050 (
);

FILL FILL_1__12846_ (
);

FILL FILL_1__12426_ (
);

FILL FILL_1__12006_ (
);

FILL FILL_3__7950_ (
);

FILL FILL_0__9853_ (
);

FILL FILL_0__11839_ (
);

FILL SFILL79080x80050 (
);

FILL FILL_0__9013_ (
);

FILL FILL_3__7110_ (
);

FILL FILL_0__11419_ (
);

OAI21X1 _11704_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2190_),
    .C(_2802_),
    .Y(_2803_)
);

FILL FILL_6__15618_ (
);

FILL FILL_5__7876_ (
);

FILL FILL_5__7456_ (
);

FILL FILL_4__16232_ (
);

FILL FILL_5__7036_ (
);

NOR2X1 _14596_ (
    .A(_5084_),
    .B(_5069_),
    .Y(_5085_)
);

NOR2X1 _14176_ (
    .A(_4672_),
    .B(_3949_),
    .Y(_4673_)
);

FILL FILL_3__15645_ (
);

FILL FILL_3__15225_ (
);

FILL SFILL39000x8050 (
);

FILL FILL_1__7868_ (
);

FILL SFILL13720x4050 (
);

FILL FILL_3__10780_ (
);

FILL FILL_1__7448_ (
);

FILL FILL_3__10360_ (
);

FILL FILL_2__14638_ (
);

FILL FILL_2__14218_ (
);

FILL FILL_0__15672_ (
);

FILL SFILL13640x9050 (
);

FILL FILL_0__15252_ (
);

FILL FILL_1_BUFX2_insert390 (
);

FILL FILL_1_BUFX2_insert391 (
);

FILL FILL_3__8735_ (
);

FILL FILL_1_BUFX2_insert392 (
);

OAI21X1 _12909_ (
    .A(_3610_),
    .B(vdd),
    .C(_3611_),
    .Y(_3555_[28])
);

FILL FILL_3__8315_ (
);

FILL FILL_1_BUFX2_insert393 (
);

FILL FILL_1_BUFX2_insert394 (
);

FILL FILL_1_BUFX2_insert395 (
);

FILL FILL_1_BUFX2_insert396 (
);

FILL FILL_1_BUFX2_insert397 (
);

FILL FILL_1_BUFX2_insert398 (
);

FILL FILL_1_BUFX2_insert399 (
);

FILL FILL_4__12992_ (
);

FILL FILL_6__11538_ (
);

FILL FILL_4__12572_ (
);

FILL FILL_6__11118_ (
);

FILL FILL_4__12152_ (
);

DFFSR _10096_ (
    .Q(\datapath_1.regfile_1.regOut[25] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_1563_[26])
);

FILL FILL_3__11985_ (
);

FILL FILL_5__9602_ (
);

FILL FILL_3__11565_ (
);

FILL FILL_3__11145_ (
);

FILL FILL_0__16037_ (
);

NAND2X1 _16322_ (
    .A(gnd),
    .B(gnd),
    .Y(_6833_)
);

FILL FILL_2__10978_ (
);

FILL FILL_2__10558_ (
);

FILL FILL_2__10138_ (
);

FILL FILL_0__11592_ (
);

FILL FILL_0__11172_ (
);

FILL SFILL23720x14050 (
);

FILL FILL_5__14784_ (
);

FILL FILL_5__14364_ (
);

FILL FILL_0__6978_ (
);

DFFSR _8664_ (
    .Q(\datapath_1.regfile_1.regOut[14] [2]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_848_[2])
);

OAI21X1 _8244_ (
    .A(_692_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_693_),
    .Y(_653_[20])
);

FILL FILL_6__7105_ (
);

FILL FILL_1__10912_ (
);

FILL FILL_4__13777_ (
);

FILL FILL_4__13357_ (
);

FILL SFILL48920x63050 (
);

FILL FILL_2__14391_ (
);

FILL FILL_2__7937_ (
);

FILL FILL_1__13384_ (
);

OAI21X1 _12662_ (
    .A(_3486_),
    .B(vdd),
    .C(_3487_),
    .Y(_3425_[31])
);

FILL FILL_0__12377_ (
);

NAND3X1 _12242_ (
    .A(_3218_),
    .B(_3219_),
    .C(_3220_),
    .Y(\datapath_1.alu_1.ALUInB [6])
);

FILL FILL_3__13711_ (
);

FILL SFILL13720x57050 (
);

FILL FILL_5__15989_ (
);

FILL SFILL44120x48050 (
);

FILL FILL_2__12704_ (
);

FILL FILL_5__15569_ (
);

FILL FILL_5__15149_ (
);

OAI21X1 _9869_ (
    .A(_1511_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1512_),
    .Y(_1498_[7])
);

FILL FILL_3__16183_ (
);

FILL SFILL109560x37050 (
);

DFFSR _9449_ (
    .Q(\datapath_1.regfile_1.regOut[20] [19]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1238_[19])
);

NAND2X1 _9029_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1095_)
);

FILL FILL_5__10284_ (
);

FILL FILL_2__15596_ (
);

FILL FILL_2__15176_ (
);

FILL FILL_0__8704_ (
);

FILL FILL_1__14589_ (
);

FILL FILL_1__14169_ (
);

FILL FILL_4__15923_ (
);

FILL FILL_4__15503_ (
);

INVX1 _13867_ (
    .A(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_4371_)
);

FILL FILL_3__9273_ (
);

NAND3X1 _13447_ (
    .A(_3898_),
    .B(_3904_),
    .C(_3879_),
    .Y(_3959_)
);

NAND2X1 _13027_ (
    .A(vdd),
    .B(\datapath_1.rd2 [25]),
    .Y(_3670_)
);

FILL FILL_3__14916_ (
);

FILL FILL_1__15950_ (
);

FILL FILL_1__15530_ (
);

FILL FILL_1__15110_ (
);

FILL SFILL8600x18050 (
);

FILL FILL_2__13909_ (
);

FILL FILL_0__14943_ (
);

FILL FILL_0__14523_ (
);

FILL FILL_0__14103_ (
);

FILL SFILL13720x12050 (
);

FILL FILL_2__7690_ (
);

FILL FILL_5__11489_ (
);

FILL FILL_5__11069_ (
);

FILL FILL_4__7196_ (
);

FILL FILL_0__9909_ (
);

FILL FILL_2__11096_ (
);

FILL SFILL38920x61050 (
);

FILL FILL_5__12850_ (
);

FILL FILL_5__12430_ (
);

FILL FILL_5__12010_ (
);

FILL FILL_4__11843_ (
);

FILL FILL_4__11423_ (
);

FILL FILL_4__11003_ (
);

FILL SFILL13640x19050 (
);

FILL FILL_0__7096_ (
);

FILL FILL_1__16315_ (
);

FILL FILL_3__10836_ (
);

FILL FILL_1__11870_ (
);

FILL FILL_3__10416_ (
);

FILL FILL_1__11450_ (
);

FILL FILL_1__11030_ (
);

FILL FILL_0__15728_ (
);

FILL FILL_0__15308_ (
);

FILL SFILL38840x68050 (
);

FILL FILL_2__8895_ (
);

FILL FILL_2__8475_ (
);

FILL FILL_0__10443_ (
);

FILL FILL_2__8055_ (
);

FILL FILL_0__10023_ (
);

FILL SFILL3560x60050 (
);

FILL FILL_5__13635_ (
);

FILL FILL_5__13215_ (
);

INVX1 _7935_ (
    .A(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_528_)
);

DFFSR _7515_ (
    .Q(\datapath_1.regfile_1.regOut[5] [5]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_263_[5])
);

FILL FILL_1__6892_ (
);

FILL FILL_4__9762_ (
);

FILL FILL_4__9342_ (
);

FILL FILL_4__12628_ (
);

FILL FILL_2__13662_ (
);

FILL FILL_4__12208_ (
);

FILL FILL_2__13242_ (
);

FILL FILL112200x55050 (
);

FILL SFILL99480x48050 (
);

FILL FILL_1__12655_ (
);

FILL FILL_1__12235_ (
);

FILL FILL_0__9662_ (
);

FILL SFILL3480x67050 (
);

NAND2X1 _11933_ (
    .A(IorD_bF$buf0),
    .B(ALUOut[15]),
    .Y(_2997_)
);

FILL FILL_0__9242_ (
);

FILL FILL_0__11648_ (
);

FILL FILL_0__11228_ (
);

OAI21X1 _11513_ (
    .A(_2437_),
    .B(_2611_),
    .C(_2470__bF$buf2),
    .Y(_2625_)
);

FILL FILL_5__7685_ (
);

FILL FILL_4__16041_ (
);

FILL FILL_3__15874_ (
);

FILL FILL_3__15454_ (
);

FILL FILL_3__15034_ (
);

FILL FILL_1__7677_ (
);

FILL FILL_2__14867_ (
);

FILL FILL_6_BUFX2_insert602 (
);

FILL FILL_2__14447_ (
);

FILL FILL_2__14027_ (
);

FILL FILL_0__15481_ (
);

FILL FILL_0__15061_ (
);

FILL FILL_6_BUFX2_insert607 (
);

FILL FILL112200x10050 (
);

FILL FILL_3__8964_ (
);

FILL FILL_3__8124_ (
);

OAI21X1 _12718_ (
    .A(_3503_),
    .B(IRWrite_bF$buf0),
    .C(_3504_),
    .Y(_3490_[7])
);

FILL SFILL28840x66050 (
);

FILL FILL_1__14801_ (
);

FILL FILL_1_BUFX2_insert60 (
);

FILL FILL_1_BUFX2_insert61 (
);

FILL FILL_1_BUFX2_insert62 (
);

FILL FILL_1_BUFX2_insert63 (
);

FILL FILL_4__12381_ (
);

FILL FILL_1_BUFX2_insert64 (
);

FILL FILL_1_BUFX2_insert65 (
);

FILL FILL_1_BUFX2_insert66 (
);

FILL FILL_3__16239_ (
);

FILL FILL_1_BUFX2_insert67 (
);

FILL FILL_1_BUFX2_insert68 (
);

FILL SFILL33800x49050 (
);

FILL FILL_1_BUFX2_insert69 (
);

FILL FILL_2__6961_ (
);

FILL FILL_3__11794_ (
);

FILL FILL_3__11374_ (
);

FILL FILL_5__9411_ (
);

FILL FILL_4__6887_ (
);

FILL FILL_0__16266_ (
);

NAND3X1 _16131_ (
    .A(_6582_),
    .B(_6583_),
    .C(_6581_),
    .Y(_6584_)
);

FILL FILL_2__10787_ (
);

FILL FILL_2__10367_ (
);

FILL FILL_5__11701_ (
);

FILL FILL_1__9403_ (
);

FILL FILL_3__9749_ (
);

FILL FILL_5__14593_ (
);

FILL FILL_5__14173_ (
);

OAI21X1 _8893_ (
    .A(_1023_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .C(_1024_),
    .Y(_978_[23])
);

OAI21X1 _8473_ (
    .A(_804_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_805_),
    .Y(_783_[11])
);

DFFSR _8053_ (
    .Q(\datapath_1.regfile_1.regOut[9] [31]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_523_[31])
);

FILL FILL_4__13586_ (
);

FILL SFILL28840x21050 (
);

FILL FILL_1__10301_ (
);

FILL FILL_4__13166_ (
);

FILL FILL_3__12999_ (
);

FILL FILL_2__7746_ (
);

FILL FILL_3__12579_ (
);

FILL FILL_2__7326_ (
);

FILL FILL_3__12159_ (
);

OAI21X1 _12891_ (
    .A(_3598_),
    .B(vdd),
    .C(_3599_),
    .Y(_3555_[22])
);

FILL FILL_0__12186_ (
);

OAI21X1 _12471_ (
    .A(_3379_),
    .B(vdd),
    .C(_3380_),
    .Y(_3360_[10])
);

NAND3X1 _12051_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[16]),
    .C(_3032__bF$buf3),
    .Y(_3084_)
);

FILL FILL_5__12906_ (
);

FILL FILL_3__13940_ (
);

FILL FILL_6__16385_ (
);

FILL FILL_3__13520_ (
);

FILL FILL_3__13100_ (
);

FILL FILL_4__8613_ (
);

FILL FILL_5_BUFX2_insert620 (
);

FILL FILL_5__15798_ (
);

FILL FILL_5_BUFX2_insert621 (
);

FILL FILL_5_BUFX2_insert622 (
);

FILL FILL_5__15378_ (
);

FILL FILL_2__12513_ (
);

FILL FILL_5_BUFX2_insert623 (
);

NAND2X1 _9678_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1426_)
);

FILL FILL_5_BUFX2_insert624 (
);

FILL FILL_5_BUFX2_insert625 (
);

NAND2X1 _9258_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1207_)
);

FILL FILL_5_BUFX2_insert626 (
);

FILL FILL_5_BUFX2_insert627 (
);

FILL FILL_5_BUFX2_insert628 (
);

FILL FILL_1__11926_ (
);

FILL FILL_5_BUFX2_insert629 (
);

FILL FILL_1__11506_ (
);

FILL SFILL18840x64050 (
);

FILL FILL_0__10919_ (
);

FILL FILL_0__8513_ (
);

FILL FILL_1__14398_ (
);

FILL FILL_5__6956_ (
);

FILL FILL_4__15732_ (
);

FILL FILL_4__15312_ (
);

INVX1 _13676_ (
    .A(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_4184_)
);

FILL FILL_3__9082_ (
);

INVX2 _13256_ (
    .A(_3777_),
    .Y(_3799_)
);

FILL FILL_3__14725_ (
);

FILL FILL_3__14305_ (
);

FILL FILL_1__6948_ (
);

FILL FILL_2__13718_ (
);

FILL FILL_0__14752_ (
);

FILL FILL_0__14332_ (
);

FILL FILL_5__11298_ (
);

FILL FILL_0__9718_ (
);

FILL FILL_3__7815_ (
);

FILL FILL_2_BUFX2_insert750 (
);

FILL FILL_2_BUFX2_insert751 (
);

FILL FILL_2_BUFX2_insert752 (
);

FILL FILL_2_BUFX2_insert753 (
);

FILL FILL_2_BUFX2_insert754 (
);

FILL FILL_4__11652_ (
);

FILL FILL_2_BUFX2_insert755 (
);

FILL FILL_4__11232_ (
);

FILL FILL_2_BUFX2_insert756 (
);

FILL FILL_2_BUFX2_insert757 (
);

FILL FILL_2_BUFX2_insert758 (
);

FILL FILL_1__16124_ (
);

FILL FILL_2_BUFX2_insert759 (
);

FILL FILL_3__10645_ (
);

FILL FILL_0__15957_ (
);

FILL FILL_0__15537_ (
);

AOI22X1 _15822_ (
    .A(_5567_),
    .B(\datapath_1.regfile_1.regOut[28] [19]),
    .C(\datapath_1.regfile_1.regOut[31] [19]),
    .D(_5571_),
    .Y(_6283_)
);

INVX1 _15402_ (
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_5874_)
);

FILL FILL_0__15117_ (
);

FILL FILL_0__10672_ (
);

FILL FILL_0__10252_ (
);

FILL FILL_6__14871_ (
);

FILL FILL_5__13864_ (
);

FILL FILL_5__13444_ (
);

FILL FILL_5__13024_ (
);

OAI21X1 _7744_ (
    .A(_440_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .C(_441_),
    .Y(_393_[24])
);

OAI21X1 _7324_ (
    .A(_221_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_222_),
    .Y(_198_[12])
);

FILL FILL_4__9991_ (
);

FILL FILL_4__9151_ (
);

FILL FILL_4__12857_ (
);

FILL SFILL48920x58050 (
);

FILL FILL_4__12437_ (
);

FILL FILL_2__13891_ (
);

FILL FILL_4__12017_ (
);

FILL FILL_2__13471_ (
);

FILL FILL_1__12884_ (
);

FILL FILL_1__12464_ (
);

FILL FILL_1__12044_ (
);

FILL FILL_6_CLKBUF1_insert203 (
);

FILL FILL_0__9891_ (
);

FILL FILL_0__9471_ (
);

FILL FILL_0__11877_ (
);

FILL FILL_2__9489_ (
);

FILL FILL_0__11457_ (
);

NOR2X1 _11742_ (
    .A(_2160_),
    .B(_2147_),
    .Y(_2838_)
);

FILL FILL_0__11037_ (
);

INVX1 _11322_ (
    .A(_2440_),
    .Y(_2441_)
);

FILL FILL_6_CLKBUF1_insert208 (
);

FILL FILL_5__7494_ (
);

FILL FILL_5__7074_ (
);

FILL FILL_4__16270_ (
);

FILL FILL_6__10791_ (
);

FILL FILL_5__14649_ (
);

FILL FILL_5__14229_ (
);

FILL FILL_3__15683_ (
);

DFFSR _8949_ (
    .Q(\datapath_1.regfile_1.regOut[16] [31]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_978_[31])
);

FILL FILL_3__15263_ (
);

NAND2X1 _8529_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_843_)
);

NAND2X1 _8109_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_624_)
);

FILL FILL_1__7486_ (
);

FILL FILL_1__7066_ (
);

FILL FILL_2__14676_ (
);

FILL FILL_2__14256_ (
);

FILL FILL_0__15290_ (
);

FILL SFILL48920x13050 (
);

FILL FILL_1__13669_ (
);

FILL FILL_1__13249_ (
);

FILL FILL_1_BUFX2_insert770 (
);

FILL FILL_1_BUFX2_insert771 (
);

FILL FILL_3__8773_ (
);

FILL FILL_3__8353_ (
);

DFFSR _12947_ (
    .Q(\datapath_1.a [28]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3555_[28])
);

FILL FILL_1_BUFX2_insert772 (
);

FILL FILL_1_BUFX2_insert773 (
);

NAND2X1 _12527_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [29]),
    .Y(_3418_)
);

FILL FILL_1_BUFX2_insert774 (
);

NAND3X1 _12107_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[30]),
    .C(_3032__bF$buf1),
    .Y(_3126_)
);

FILL FILL_1_BUFX2_insert775 (
);

FILL FILL_1_BUFX2_insert776 (
);

FILL FILL_5__8699_ (
);

FILL FILL_1__14610_ (
);

FILL FILL_1_BUFX2_insert777 (
);

FILL FILL_1_BUFX2_insert778 (
);

FILL FILL_1_BUFX2_insert779 (
);

FILL FILL_4__12190_ (
);

FILL FILL_0__13603_ (
);

FILL FILL_3__16048_ (
);

FILL FILL_5__10989_ (
);

FILL FILL_5__10569_ (
);

FILL FILL_5__9640_ (
);

FILL FILL_5__10149_ (
);

FILL FILL_5__9220_ (
);

FILL FILL_3__11183_ (
);

FILL SFILL59080x71050 (
);

FILL FILL_0__16075_ (
);

INVX1 _16360_ (
    .A(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_6794_)
);

FILL SFILL38920x56050 (
);

FILL FILL_2__10176_ (
);

FILL FILL_5__11930_ (
);

FILL FILL_1__9632_ (
);

FILL FILL_5__11510_ (
);

FILL FILL_1__9212_ (
);

FILL FILL_3__9978_ (
);

FILL FILL_2__16402_ (
);

FILL FILL_4__10923_ (
);

FILL FILL_3__9138_ (
);

FILL FILL_4__10503_ (
);

FILL FILL_6__7983_ (
);

FILL FILL_1__15815_ (
);

DFFSR _8282_ (
    .Q(\datapath_1.regfile_1.regOut[11] [4]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_653_[4])
);

FILL FILL_1__10950_ (
);

FILL FILL_1__10530_ (
);

FILL FILL_4__13395_ (
);

FILL FILL_1__10110_ (
);

FILL FILL_0__14808_ (
);

FILL FILL_2__7975_ (
);

FILL FILL_2__7555_ (
);

BUFX2 BUFX2_insert440 (
    .A(_5565_),
    .Y(_5565__bF$buf1)
);

FILL FILL_3__12388_ (
);

BUFX2 BUFX2_insert441 (
    .A(_5565_),
    .Y(_5565__bF$buf0)
);

BUFX2 BUFX2_insert442 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf4 )
);

FILL SFILL99560x36050 (
);

BUFX2 BUFX2_insert443 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf3 )
);

BUFX2 BUFX2_insert444 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf2 )
);

BUFX2 BUFX2_insert445 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf1 )
);

BUFX2 BUFX2_insert446 (
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf0 )
);

BUFX2 BUFX2_insert447 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf7 )
);

BUFX2 BUFX2_insert448 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf6 )
);

BUFX2 BUFX2_insert449 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf5 )
);

FILL SFILL3560x55050 (
);

NAND3X1 _12280_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3198__bF$buf2),
    .Y(_3249_)
);

FILL FILL_5__12715_ (
);

FILL SFILL38920x11050 (
);

FILL SFILL104440x72050 (
);

FILL FILL_4__8842_ (
);

FILL FILL_4__8002_ (
);

FILL FILL_4__11708_ (
);

FILL FILL_2__12742_ (
);

FILL FILL_5__15187_ (
);

FILL FILL_2__12322_ (
);

NAND2X1 _9487_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1319_)
);

DFFSR _9067_ (
    .Q(\datapath_1.regfile_1.regOut[17] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_1043_[21])
);

FILL FILL_1__11735_ (
);

FILL FILL_1__11315_ (
);

FILL FILL_0__8742_ (
);

FILL FILL_0__8322_ (
);

FILL FILL_0__10308_ (
);

FILL SFILL89560x79050 (
);

FILL SFILL38840x18050 (
);

FILL FILL_6__14927_ (
);

FILL FILL_4__15961_ (
);

FILL FILL_4__15541_ (
);

FILL FILL_4__15121_ (
);

AOI22X1 _13485_ (
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .B(_3995__bF$buf0),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_3996_)
);

DFFSR _13065_ (
    .Q(_2_[18]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_3620_[18])
);

FILL FILL_3__14954_ (
);

FILL FILL_3__14534_ (
);

FILL FILL_3__14114_ (
);

FILL SFILL28920x54050 (
);

FILL SFILL3560x10050 (
);

FILL FILL_4_BUFX2_insert280 (
);

FILL FILL_4_BUFX2_insert281 (
);

FILL FILL_4__9627_ (
);

FILL FILL_4_BUFX2_insert282 (
);

FILL FILL_4__9207_ (
);

FILL FILL_4_BUFX2_insert283 (
);

FILL FILL_2__13947_ (
);

FILL SFILL89160x65050 (
);

FILL FILL_2__13527_ (
);

FILL FILL_0__14981_ (
);

FILL FILL_4_BUFX2_insert284 (
);

FILL FILL_0__14561_ (
);

FILL FILL_2__13107_ (
);

FILL FILL_4_BUFX2_insert285 (
);

FILL FILL_4_BUFX2_insert286 (
);

FILL FILL_0__14141_ (
);

FILL FILL_4_BUFX2_insert287 (
);

FILL FILL_4_BUFX2_insert288 (
);

FILL FILL_4_BUFX2_insert289 (
);

FILL FILL_0__9527_ (
);

FILL FILL_3__7624_ (
);

FILL FILL_3__7204_ (
);

FILL FILL_0__9107_ (
);

FILL FILL_4__16326_ (
);

FILL FILL_4__11881_ (
);

FILL FILL_4__11461_ (
);

FILL FILL_4__11041_ (
);

FILL FILL_3__15739_ (
);

FILL FILL_3__15319_ (
);

FILL FILL_1__16353_ (
);

FILL FILL_5__8911_ (
);

FILL FILL_3__10874_ (
);

FILL FILL_3__10034_ (
);

FILL FILL_0__15766_ (
);

FILL FILL_0__15346_ (
);

NAND3X1 _15631_ (
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf3),
    .Y(_6097_)
);

NOR2X1 _15211_ (
    .A(_4164_),
    .B(_5534__bF$buf0),
    .Y(_5687_)
);

FILL FILL_2__8093_ (
);

FILL FILL_0__10061_ (
);

FILL FILL_1__8903_ (
);

FILL FILL_3__8829_ (
);

FILL FILL_5__13673_ (
);

FILL FILL_5__13253_ (
);

OAI21X1 _7973_ (
    .A(_552_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .C(_553_),
    .Y(_523_[15])
);

OAI21X1 _7553_ (
    .A(_333_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .C(_334_),
    .Y(_328_[3])
);

DFFSR _7133_ (
    .Q(\datapath_1.regfile_1.regOut[2] [7]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_68_[7])
);

FILL SFILL58600x79050 (
);

FILL FILL_4__9380_ (
);

FILL SFILL94360x83050 (
);

FILL FILL_4__12246_ (
);

FILL FILL_2__13280_ (
);

FILL FILL_3__11659_ (
);

FILL FILL_3__11239_ (
);

FILL FILL_1__12273_ (
);

OAI21X1 _16416_ (
    .A(_6830_),
    .B(gnd),
    .C(_6831_),
    .Y(_6769_[31])
);

FILL FILL_0__9280_ (
);

INVX1 _11971_ (
    .A(\datapath_1.PCJump [28]),
    .Y(_3022_)
);

FILL FILL_0__11686_ (
);

FILL FILL_2__9298_ (
);

FILL SFILL79160x63050 (
);

OAI21X1 _11551_ (
    .A(_2659_),
    .B(_2235_),
    .C(_2430_),
    .Y(_2660_)
);

FILL FILL_0__11266_ (
);

NAND2X1 _11131_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2250_)
);

FILL FILL_3__12600_ (
);

FILL FILL_6__15465_ (
);

FILL FILL_6__15045_ (
);

FILL SFILL90040x30050 (
);

FILL FILL_5__14878_ (
);

FILL FILL_5__14458_ (
);

FILL FILL_5__14038_ (
);

FILL FILL_3__15492_ (
);

NAND2X1 _8758_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_955_)
);

FILL FILL_3__15072_ (
);

NAND2X1 _8338_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_736_)
);

FILL FILL_1__7295_ (
);

FILL SFILL18840x59050 (
);

FILL FILL_2__14485_ (
);

FILL FILL_2__14065_ (
);

FILL FILL_1__13898_ (
);

FILL FILL_1__13478_ (
);

FILL FILL_4__14812_ (
);

FILL FILL_3__8582_ (
);

NAND2X1 _12756_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[20]),
    .Y(_3530_)
);

NAND3X1 _12336_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3198__bF$buf1),
    .Y(_3291_)
);

FILL FILL_3__13805_ (
);

FILL FILL_5__8088_ (
);

FILL FILL_0__13832_ (
);

FILL FILL_0__13412_ (
);

FILL FILL_3__16277_ (
);

FILL FILL_5__10798_ (
);

FILL FILL_5__10378_ (
);

FILL SFILL84360x81050 (
);

FILL FILL_1__9861_ (
);

FILL FILL_1__9021_ (
);

FILL FILL_3__9787_ (
);

FILL FILL_2__16211_ (
);

FILL FILL_3__9367_ (
);

FILL FILL_4__10312_ (
);

FILL FILL_1__15624_ (
);

FILL FILL_1__15204_ (
);

NAND2X1 _8091_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_612_)
);

FILL FILL_0__14617_ (
);

INVX1 _14902_ (
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_5384_)
);

FILL FILL_2__7364_ (
);

FILL FILL_3__12197_ (
);

FILL FILL_6__13531_ (
);

FILL FILL_5__12524_ (
);

FILL SFILL99400x3050 (
);

FILL FILL_5__12104_ (
);

FILL FILL_4__8651_ (
);

FILL FILL_4__8231_ (
);

FILL FILL_4__11937_ (
);

FILL FILL_2__12971_ (
);

FILL FILL_4__11517_ (
);

FILL FILL_6__8997_ (
);

FILL FILL_2__12131_ (
);

FILL FILL_1__16409_ (
);

INVX1 _9296_ (
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_1232_)
);

FILL FILL_1__11964_ (
);

FILL FILL_1__11544_ (
);

FILL FILL_1__11124_ (
);

FILL FILL_0__8971_ (
);

FILL FILL_2__8989_ (
);

FILL FILL_0__10957_ (
);

FILL FILL_2__8569_ (
);

FILL FILL_2__8149_ (
);

OAI21X1 _10822_ (
    .A(_2004_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_2005_),
    .Y(_1953_[26])
);

FILL FILL_0__10537_ (
);

FILL FILL_0__8131_ (
);

FILL SFILL114520x62050 (
);

OAI21X1 _10402_ (
    .A(_1785_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .C(_1786_),
    .Y(_1758_[14])
);

FILL FILL_0__10117_ (
);

FILL FILL_5__6994_ (
);

FILL FILL_4__15770_ (
);

FILL FILL_4__15350_ (
);

FILL SFILL3720x81050 (
);

INVX1 _13294_ (
    .A(_3774_),
    .Y(_3831_)
);

FILL FILL_2__9930_ (
);

FILL FILL_5__13729_ (
);

FILL FILL_5__13309_ (
);

FILL FILL_2__9510_ (
);

FILL FILL_3__14763_ (
);

FILL FILL_3__14343_ (
);

NAND2X1 _7609_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_372_)
);

FILL FILL_1__6986_ (
);

FILL FILL_4__9856_ (
);

FILL FILL_4__9016_ (
);

FILL FILL_2__13756_ (
);

FILL FILL_2__13336_ (
);

FILL FILL_0__14790_ (
);

FILL FILL_0__14370_ (
);

FILL FILL_1__12749_ (
);

FILL FILL_1__12329_ (
);

FILL FILL_0__9756_ (
);

FILL FILL_3__7853_ (
);

FILL FILL_3__7433_ (
);

FILL FILL_0__9336_ (
);

OAI22X1 _11607_ (
    .A(_2240_),
    .B(_2346_),
    .C(_2347__bF$buf1),
    .D(_2239_),
    .Y(_2713_)
);

FILL FILL_5__7359_ (
);

FILL FILL_4__16135_ (
);

NOR2X1 _14499_ (
    .A(_4989_),
    .B(_4974_),
    .Y(_4990_)
);

FILL FILL_4__11690_ (
);

FILL FILL_4__11270_ (
);

INVX1 _14079_ (
    .A(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_4578_)
);

FILL FILL_3__15968_ (
);

FILL FILL_3__15548_ (
);

FILL FILL_3__15128_ (
);

FILL FILL_1__16162_ (
);

FILL FILL_3__10683_ (
);

FILL FILL_5__8720_ (
);

FILL FILL_3__10263_ (
);

FILL SFILL59080x66050 (
);

FILL FILL_0__15995_ (
);

NAND3X1 _15860_ (
    .A(_6318_),
    .B(_6319_),
    .C(_6317_),
    .Y(_6320_)
);

FILL FILL_0__15575_ (
);

FILL FILL_0__15155_ (
);

NAND3X1 _15440_ (
    .A(_5906_),
    .B(_5910_),
    .C(_5908_),
    .Y(_5911_)
);

NOR3X1 _15020_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(\datapath_1.PCJump [24]),
    .C(\datapath_1.PCJump [23]),
    .Y(_5500_)
);

FILL FILL_0__10290_ (
);

FILL FILL_1__8712_ (
);

FILL SFILL83560x77050 (
);

FILL FILL_2__15902_ (
);

FILL FILL_3__8638_ (
);

FILL FILL_3__8218_ (
);

FILL SFILL3640x43050 (
);

FILL FILL_5__13482_ (
);

DFFSR _7782_ (
    .Q(\datapath_1.regfile_1.regOut[7] [16]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_393_[16])
);

NAND2X1 _7362_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_248_)
);

FILL FILL_4__12895_ (
);

FILL FILL_4__12475_ (
);

FILL FILL_4__12055_ (
);

FILL FILL_5_BUFX2_insert10 (
);

FILL FILL_5_BUFX2_insert11 (
);

FILL FILL_3__11888_ (
);

FILL FILL_5__9925_ (
);

FILL FILL_5__9505_ (
);

FILL FILL_5_BUFX2_insert12 (
);

FILL FILL_3__11468_ (
);

FILL SFILL83960x46050 (
);

FILL FILL_5_BUFX2_insert13 (
);

FILL FILL_3__11048_ (
);

FILL SFILL59000x64050 (
);

FILL FILL_1__12082_ (
);

FILL FILL_5_BUFX2_insert14 (
);

FILL FILL_5_BUFX2_insert15 (
);

FILL FILL_5_BUFX2_insert16 (
);

OAI22X1 _16225_ (
    .A(_6675_),
    .B(_5545__bF$buf0),
    .C(_5569_),
    .D(_5356_),
    .Y(_6676_)
);

FILL FILL_5_BUFX2_insert17 (
);

FILL SFILL38120x23050 (
);

FILL FILL_5_BUFX2_insert18 (
);

FILL FILL_5_BUFX2_insert19 (
);

FILL SFILL59080x21050 (
);

NOR2X1 _11780_ (
    .A(_2873_),
    .B(_2872_),
    .Y(_2874_)
);

FILL FILL_0__11495_ (
);

OAI21X1 _11360_ (
    .A(_2475_),
    .B(_2452_),
    .C(_2470__bF$buf3),
    .Y(_2477_)
);

FILL FILL_0__11075_ (
);

FILL FILL_1__9917_ (
);

FILL SFILL104440x67050 (
);

FILL FILL_4__7502_ (
);

FILL FILL_2__11822_ (
);

FILL FILL_5__14687_ (
);

FILL FILL_5__14267_ (
);

FILL FILL_2__11402_ (
);

NAND2X1 _8987_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1067_)
);

NAND2X1 _8567_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .Y(_912_)
);

INVX1 _8147_ (
    .A(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_649_)
);

FILL FILL_1__10815_ (
);

FILL FILL_2__14294_ (
);

FILL FILL_0__7822_ (
);

FILL FILL_1__13287_ (
);

FILL FILL_4__14621_ (
);

FILL FILL_4__14201_ (
);

FILL SFILL43960x8050 (
);

NAND2X1 _12985_ (
    .A(vdd),
    .B(\datapath_1.rd2 [11]),
    .Y(_3642_)
);

FILL FILL_3__8391_ (
);

DFFSR _12565_ (
    .Q(ALUOut[30]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3360_[30])
);

INVX1 _12145_ (
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_3150_)
);

FILL FILL_3__13614_ (
);

FILL FILL_4__8707_ (
);

FILL SFILL104440x22050 (
);

FILL FILL_2__12607_ (
);

FILL FILL_0__13641_ (
);

FILL FILL_0__13221_ (
);

FILL FILL_3__16086_ (
);

FILL FILL_5__10187_ (
);

FILL FILL_2__15499_ (
);

FILL FILL_2__15079_ (
);

FILL FILL_5__16413_ (
);

FILL FILL_0__8607_ (
);

FILL SFILL108760x30050 (
);

FILL FILL_1__9670_ (
);

FILL FILL_1__9250_ (
);

FILL FILL_4__15826_ (
);

FILL FILL_4__15406_ (
);

BUFX2 BUFX2_insert1000 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf4 )
);

BUFX2 BUFX2_insert1001 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf3 )
);

FILL SFILL89560x29050 (
);

FILL FILL_2__16020_ (
);

BUFX2 BUFX2_insert1002 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf2 )
);

FILL FILL_3__9596_ (
);

FILL SFILL49000x62050 (
);

BUFX2 BUFX2_insert1003 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf1 )
);

FILL FILL_4__10961_ (
);

BUFX2 BUFX2_insert1004 (
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf0 )
);

FILL FILL_4__10541_ (
);

FILL FILL_4__10121_ (
);

BUFX2 BUFX2_insert1005 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf4)
);

FILL FILL_3__14819_ (
);

BUFX2 BUFX2_insert1006 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf3)
);

BUFX2 BUFX2_insert1007 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf2)
);

FILL FILL_1__15853_ (
);

BUFX2 BUFX2_insert1008 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf1)
);

FILL FILL_1__15433_ (
);

FILL FILL_1__15013_ (
);

BUFX2 BUFX2_insert1009 (
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf0)
);

FILL SFILL94440x71050 (
);

FILL FILL_0__14846_ (
);

NOR2X1 _14711_ (
    .A(_5196_),
    .B(_3977__bF$buf0),
    .Y(_5197_)
);

FILL FILL_0__14426_ (
);

FILL FILL_0__14006_ (
);

FILL FILL_2__7593_ (
);

BUFX2 BUFX2_insert820 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf1 )
);

FILL FILL_2__7173_ (
);

BUFX2 BUFX2_insert821 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf0 )
);

BUFX2 BUFX2_insert822 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf7 )
);

BUFX2 BUFX2_insert823 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf6 )
);

BUFX2 BUFX2_insert824 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf5 )
);

BUFX2 BUFX2_insert825 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf4 )
);

FILL FILL_4__7099_ (
);

BUFX2 BUFX2_insert826 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf3 )
);

BUFX2 BUFX2_insert827 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf2 )
);

BUFX2 BUFX2_insert828 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf1 )
);

BUFX2 BUFX2_insert829 (
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf0 )
);

FILL FILL_5__12753_ (
);

FILL FILL_5__12333_ (
);

FILL FILL_4__8880_ (
);

FILL FILL_4__8460_ (
);

FILL FILL_4__11746_ (
);

FILL FILL_2__12780_ (
);

FILL FILL_4__11326_ (
);

FILL FILL_2__12360_ (
);

FILL FILL_6__8386_ (
);

FILL FILL_1__16218_ (
);

FILL FILL_3__10319_ (
);

FILL FILL_1__11773_ (
);

FILL FILL_1__11353_ (
);

AOI21X1 _15916_ (
    .A(\datapath_1.regfile_1.regOut[30] [21]),
    .B(_5481_),
    .C(_6374_),
    .Y(_6375_)
);

FILL FILL_0__8780_ (
);

FILL SFILL79160x58050 (
);

FILL FILL_0__8360_ (
);

FILL FILL_0__10766_ (
);

FILL FILL_2__8378_ (
);

OAI21X1 _10631_ (
    .A(_1897_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1898_),
    .Y(_1888_[5])
);

DFFSR _10211_ (
    .Q(\datapath_1.regfile_1.regOut[26] [13]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_1628_[13])
);

FILL FILL_5__13958_ (
);

FILL FILL_3__14992_ (
);

FILL FILL_5__13538_ (
);

FILL FILL_3__14572_ (
);

FILL FILL_5__13118_ (
);

FILL FILL_3__14152_ (
);

NAND2X1 _7838_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_484_)
);

NAND2X1 _7418_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_265_)
);

FILL FILL_4_BUFX2_insert660 (
);

FILL FILL_4_BUFX2_insert661 (
);

FILL FILL_4__9665_ (
);

FILL FILL_4_BUFX2_insert662 (
);

FILL FILL_4__9245_ (
);

FILL FILL_2__13985_ (
);

FILL FILL_4_BUFX2_insert663 (
);

FILL FILL_4_BUFX2_insert664 (
);

FILL FILL_2__13565_ (
);

FILL FILL111800x62050 (
);

FILL FILL_2__13145_ (
);

FILL FILL_4_BUFX2_insert665 (
);

FILL FILL_4_BUFX2_insert666 (
);

FILL FILL_4_BUFX2_insert667 (
);

FILL SFILL39000x60050 (
);

FILL SFILL94360x33050 (
);

FILL FILL_4_BUFX2_insert668 (
);

FILL FILL_4_BUFX2_insert669 (
);

FILL FILL_1__12978_ (
);

FILL FILL_1__12138_ (
);

FILL FILL_0__9985_ (
);

FILL FILL_3__7242_ (
);

FILL FILL_0__9145_ (
);

OAI21X1 _11836_ (
    .A(_2920_),
    .B(_2542_),
    .C(_2924_),
    .Y(_2925_)
);

NOR2X1 _11416_ (
    .A(_2532_),
    .B(_2326_),
    .Y(_2533_)
);

FILL FILL_5__7588_ (
);

FILL SFILL79160x13050 (
);

FILL FILL_5__7168_ (
);

FILL FILL_4__16364_ (
);

FILL FILL111720x69050 (
);

FILL FILL_0__12912_ (
);

FILL FILL_3__15777_ (
);

FILL FILL_3__15357_ (
);

FILL FILL_1__16391_ (
);

FILL FILL_3__10492_ (
);

FILL FILL_0__15384_ (
);

FILL SFILL84360x76050 (
);

FILL FILL_1__8521_ (
);

FILL FILL_1__8101_ (
);

FILL FILL_2__15711_ (
);

FILL FILL_3__8867_ (
);

FILL FILL_3__8447_ (
);

FILL FILL_5__13291_ (
);

NAND2X1 _7591_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_360_)
);

FILL FILL_1__14704_ (
);

FILL FILL_4_BUFX2_insert1040 (
);

NAND2X1 _7171_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_141_)
);

FILL FILL_4_BUFX2_insert1041 (
);

FILL FILL_4_BUFX2_insert1042 (
);

FILL FILL_4_BUFX2_insert1043 (
);

FILL FILL_4_BUFX2_insert1044 (
);

FILL FILL_4__12284_ (
);

FILL FILL_4_BUFX2_insert1045 (
);

FILL FILL_4_BUFX2_insert1046 (
);

FILL FILL_4_BUFX2_insert1047 (
);

FILL FILL_4_BUFX2_insert1048 (
);

FILL FILL_4_BUFX2_insert1049 (
);

FILL FILL_2__6864_ (
);

FILL FILL_5__9734_ (
);

FILL FILL_3__11697_ (
);

FILL FILL_3__11277_ (
);

FILL FILL_0__16169_ (
);

INVX1 _16034_ (
    .A(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_6490_)
);

FILL SFILL114600x50050 (
);

FILL FILL_1__9726_ (
);

FILL FILL_5__11604_ (
);

FILL SFILL53960x40050 (
);

FILL SFILL84360x31050 (
);

FILL FILL_3_BUFX2_insert680 (
);

FILL FILL_4__7731_ (
);

FILL FILL_4__7311_ (
);

FILL FILL_3_BUFX2_insert681 (
);

FILL FILL_3_BUFX2_insert682 (
);

FILL FILL_5__14496_ (
);

FILL FILL_3_BUFX2_insert683 (
);

FILL FILL_2__11631_ (
);

FILL FILL_3_BUFX2_insert684 (
);

FILL FILL_2__11211_ (
);

FILL FILL_5__14076_ (
);

FILL FILL_1__15909_ (
);

DFFSR _8796_ (
    .Q(\datapath_1.regfile_1.regOut[15] [6]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_913_[6])
);

FILL FILL_3_BUFX2_insert685 (
);

INVX1 _8376_ (
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_761_)
);

FILL FILL_3_BUFX2_insert686 (
);

FILL FILL_3_BUFX2_insert687 (
);

FILL FILL_3_BUFX2_insert688 (
);

FILL FILL_3_BUFX2_insert689 (
);

FILL FILL_1__10624_ (
);

FILL FILL_4__13489_ (
);

FILL FILL_0__7631_ (
);

FILL SFILL114520x57050 (
);

FILL FILL_2__7229_ (
);

FILL FILL_0__7211_ (
);

FILL SFILL53880x47050 (
);

FILL FILL_1__13096_ (
);

FILL FILL_4__14850_ (
);

FILL FILL_4__14430_ (
);

FILL SFILL3720x76050 (
);

FILL FILL_4__14010_ (
);

DFFSR _12794_ (
    .Q(\aluControl_1.inst [3]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3490_[3])
);

NAND2X1 _12374_ (
    .A(MemToReg_bF$buf0),
    .B(\datapath_1.Data [10]),
    .Y(_3315_)
);

FILL FILL_0__12089_ (
);

FILL FILL_3__13843_ (
);

FILL SFILL43960x83050 (
);

FILL FILL_3__13423_ (
);

FILL FILL_6__16288_ (
);

FILL FILL_3__13003_ (
);

FILL FILL_4__8516_ (
);

FILL SFILL69080x18050 (
);

FILL FILL_2__12836_ (
);

FILL FILL_2__12416_ (
);

FILL FILL_0__13870_ (
);

FILL FILL_0__13450_ (
);

FILL FILL_0__13030_ (
);

FILL FILL_1__11829_ (
);

FILL FILL_1__11409_ (
);

FILL FILL_5__16222_ (
);

FILL FILL_0__8836_ (
);

FILL FILL_3__6933_ (
);

FILL FILL_5__6859_ (
);

FILL FILL_4__15635_ (
);

FILL SFILL114520x12050 (
);

FILL FILL_4__15215_ (
);

INVX1 _13999_ (
    .A(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_4500_)
);

AOI22X1 _13579_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [2]),
    .C(\datapath_1.regfile_1.regOut[2] [2]),
    .D(_3998__bF$buf0),
    .Y(_4089_)
);

FILL FILL_4__10770_ (
);

OAI21X1 _13159_ (
    .A(_3736_),
    .B(PCEn_bF$buf7),
    .C(_3737_),
    .Y(_3685_[26])
);

FILL SFILL3720x31050 (
);

FILL FILL_3__14628_ (
);

FILL FILL_1__15662_ (
);

FILL FILL_3__14208_ (
);

FILL FILL_1__15242_ (
);

FILL FILL_5__7800_ (
);

INVX1 _14940_ (
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_5421_)
);

FILL FILL_0__14655_ (
);

FILL FILL_0__14235_ (
);

INVX1 _14520_ (
    .A(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_5010_)
);

INVX1 _14100_ (
    .A(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_4599_)
);

FILL FILL_3__7718_ (
);

FILL SFILL49480x8050 (
);

FILL SFILL3640x38050 (
);

FILL FILL_5__12982_ (
);

FILL FILL_5__12142_ (
);

BUFX2 _6862_ (
    .A(_1_[24]),
    .Y(memoryAddress[24])
);

FILL SFILL104520x55050 (
);

FILL FILL_4__11975_ (
);

FILL FILL_4__11555_ (
);

FILL FILL_4__11135_ (
);

FILL FILL_1__16027_ (
);

FILL FILL_3__10968_ (
);

FILL SFILL49080x7050 (
);

FILL FILL_3__10548_ (
);

FILL SFILL59000x59050 (
);

FILL FILL_3__10128_ (
);

FILL FILL_1__11582_ (
);

FILL FILL_1__11162_ (
);

NOR2X1 _15725_ (
    .A(_6188_),
    .B(_6185_),
    .Y(_6189_)
);

AOI22X1 _15305_ (
    .A(_5565__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [6]),
    .C(\datapath_1.regfile_1.regOut[5] [6]),
    .D(_5700_),
    .Y(_5779_)
);

FILL SFILL59080x16050 (
);

FILL FILL_0__10995_ (
);

FILL FILL_0__10575_ (
);

DFFSR _10860_ (
    .Q(\datapath_1.regfile_1.regOut[31] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_1953_[22])
);

FILL FILL_2__8187_ (
);

FILL FILL_0__10155_ (
);

NAND2X1 _10440_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1812_)
);

NAND2X1 _10020_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1593_)
);

FILL FILL_6__14774_ (
);

FILL FILL_6__14354_ (
);

FILL FILL_2__10902_ (
);

FILL FILL_5__13767_ (
);

FILL FILL_5__13347_ (
);

FILL FILL_3__14381_ (
);

DFFSR _7647_ (
    .Q(\datapath_1.regfile_1.regOut[6] [9]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_328_[9])
);

INVX1 _7227_ (
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_178_)
);

FILL FILL_4__9894_ (
);

FILL FILL_4__9474_ (
);

FILL FILL_2__13794_ (
);

FILL FILL_2__13374_ (
);

FILL SFILL104520x10050 (
);

FILL FILL_0__6902_ (
);

FILL FILL_1__12787_ (
);

FILL FILL_1__12367_ (
);

FILL FILL_4__13701_ (
);

FILL SFILL59000x14050 (
);

FILL FILL_3__7891_ (
);

FILL FILL_0__9794_ (
);

FILL FILL_3__7471_ (
);

FILL FILL_0__9374_ (
);

FILL FILL_3__7051_ (
);

NAND2X1 _11645_ (
    .A(_2402_),
    .B(_2481__bF$buf3),
    .Y(_2748_)
);

NAND3X1 _11225_ (
    .A(ALUControl[1]),
    .B(ALUControl[0]),
    .C(_2343_),
    .Y(_2344_)
);

FILL FILL_4__16173_ (
);

FILL FILL_6__10274_ (
);

FILL FILL_0__12721_ (
);

FILL FILL_3__15586_ (
);

FILL FILL_0__12301_ (
);

FILL FILL_3__15166_ (
);

FILL FILL_2__14999_ (
);

FILL FILL_2__14579_ (
);

FILL FILL_2__14159_ (
);

FILL FILL_0__15193_ (
);

FILL SFILL33880x43050 (
);

FILL FILL_5__15913_ (
);

FILL FILL_1__8750_ (
);

FILL FILL_1__8330_ (
);

FILL FILL_4__14906_ (
);

FILL FILL_2__15940_ (
);

FILL FILL_2__15520_ (
);

FILL SFILL49000x57050 (
);

FILL FILL_2__15100_ (
);

FILL FILL_3__8256_ (
);

FILL FILL_1__14933_ (
);

FILL SFILL49080x14050 (
);

FILL FILL_1__14513_ (
);

FILL SFILL94440x66050 (
);

FILL FILL_4__12093_ (
);

FILL FILL_0__13926_ (
);

FILL FILL_0__13506_ (
);

FILL FILL_5__9543_ (
);

FILL FILL_5__9123_ (
);

FILL FILL_3__11086_ (
);

FILL FILL_0__16398_ (
);

NOR3X1 _16263_ (
    .A(_5403_),
    .B(_5459__bF$buf2),
    .C(_5519_),
    .Y(_6713_)
);

FILL FILL_2__10499_ (
);

FILL FILL_5__11833_ (
);

FILL FILL_1__9535_ (
);

FILL FILL_5__11413_ (
);

FILL FILL_1__9115_ (
);

FILL FILL_4__7960_ (
);

FILL FILL_2__16305_ (
);

FILL FILL_4__10826_ (
);

FILL FILL_4__7120_ (
);

FILL FILL_4__10406_ (
);

FILL FILL_2__11860_ (
);

FILL FILL_2__11440_ (
);

FILL FILL_2__11020_ (
);

FILL SFILL49000x12050 (
);

FILL FILL_1__15718_ (
);

FILL SFILL39080x57050 (
);

INVX1 _8185_ (
    .A(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_654_)
);

FILL FILL_4__13298_ (
);

FILL FILL_1__10433_ (
);

FILL FILL_1__10013_ (
);

FILL FILL_2__7878_ (
);

FILL FILL_0__7860_ (
);

FILL FILL_0__7440_ (
);

FILL FILL_2__7458_ (
);

FILL FILL_2__7038_ (
);

FILL SFILL18840x4050 (
);

FILL SFILL18760x9050 (
);

OAI21X1 _12183_ (
    .A(_3174_),
    .B(ALUSrcA_bF$buf5),
    .C(_3175_),
    .Y(\datapath_1.alu_1.ALUInA [22])
);

FILL FILL_5__12618_ (
);

FILL SFILL23880x41050 (
);

FILL FILL_3__13652_ (
);

FILL FILL_3__13232_ (
);

NAND2X1 _6918_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_13_)
);

FILL FILL_4__8745_ (
);

FILL FILL_4__8325_ (
);

FILL FILL_2__12645_ (
);

FILL FILL_2__12225_ (
);

FILL SFILL39000x55050 (
);

FILL SFILL94360x28050 (
);

FILL FILL_1__11638_ (
);

FILL FILL_1__11218_ (
);

FILL FILL_6_BUFX2_insert60 (
);

FILL FILL_5__16451_ (
);

FILL FILL_5__16031_ (
);

FILL FILL_0__8645_ (
);

FILL FILL_6__9612_ (
);

NAND2X1 _10916_ (
    .A(_2047_),
    .B(_2053_),
    .Y(_2059_)
);

FILL FILL_0__8225_ (
);

FILL FILL_6_BUFX2_insert65 (
);

FILL FILL_4__15864_ (
);

FILL FILL_4__15444_ (
);

FILL FILL_4__15024_ (
);

NAND2X1 _13388_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3900_)
);

FILL SFILL39400x24050 (
);

FILL FILL_3__14857_ (
);

FILL FILL_2__9604_ (
);

FILL FILL_3__14437_ (
);

FILL FILL_1__15891_ (
);

FILL FILL_3__14017_ (
);

FILL FILL_1__15471_ (
);

FILL FILL_1__15051_ (
);

FILL FILL_0__14884_ (
);

FILL FILL_0__14464_ (
);

FILL FILL_0__14044_ (
);

FILL FILL111800x12050 (
);

FILL FILL_1__7601_ (
);

FILL FILL_3__7947_ (
);

FILL FILL_3__7107_ (
);

FILL FILL_5__12371_ (
);

FILL FILL_4__16229_ (
);

FILL FILL_4__11784_ (
);

FILL FILL_4__11364_ (
);

FILL SFILL13800x82050 (
);

FILL FILL_1__16256_ (
);

FILL FILL_3__10777_ (
);

FILL FILL_1__11391_ (
);

FILL FILL_0__15669_ (
);

NOR2X1 _15954_ (
    .A(_6409_),
    .B(_6411_),
    .Y(_6412_)
);

FILL FILL_0__15249_ (
);

NAND2X1 _15534_ (
    .A(_6002_),
    .B(_5997_),
    .Y(_6003_)
);

NAND3X1 _15114_ (
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf1),
    .Y(_5593_)
);

FILL FILL_0__10384_ (
);

FILL SFILL114600x45050 (
);

FILL SFILL53960x35050 (
);

FILL SFILL84360x26050 (
);

FILL FILL_5__13996_ (
);

FILL FILL_5__13576_ (
);

FILL FILL_5__13156_ (
);

FILL FILL_3__14190_ (
);

INVX1 _7876_ (
    .A(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_509_)
);

INVX1 _7456_ (
    .A(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_290_)
);

FILL SFILL74440x62050 (
);

INVX1 _7036_ (
    .A(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_71_)
);

FILL FILL_4__12989_ (
);

FILL FILL_4__9283_ (
);

FILL FILL_4__12569_ (
);

FILL FILL_4__12149_ (
);

FILL FILL_1__12596_ (
);

FILL FILL_1__12176_ (
);

FILL FILL_4__13930_ (
);

NOR3X1 _16319_ (
    .A(_6757_),
    .B(_6746_),
    .C(_6767_),
    .Y(_6768_)
);

FILL FILL_4__13510_ (
);

OAI21X1 _11874_ (
    .A(_2958_),
    .B(RegDst),
    .C(_2959_),
    .Y(\datapath_1.a3 [0])
);

FILL FILL_0__11589_ (
);

FILL FILL_0__11169_ (
);

OAI21X1 _11454_ (
    .A(_2569_),
    .B(_2436_),
    .C(_2444_),
    .Y(_2570_)
);

AOI21X1 _11034_ (
    .A(_2152_),
    .B(_2148_),
    .C(_2150_),
    .Y(_2153_)
);

FILL SFILL43960x78050 (
);

FILL FILL_3__12503_ (
);

FILL FILL_2__11916_ (
);

FILL FILL_3__15395_ (
);

FILL FILL_0__12530_ (
);

FILL FILL_0__12110_ (
);

FILL FILL_1__7198_ (
);

FILL FILL_1__10909_ (
);

FILL FILL_2__14388_ (
);

FILL FILL_5__15722_ (
);

FILL FILL_5__15302_ (
);

INVX1 _9602_ (
    .A(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_1375_)
);

FILL FILL_4__14715_ (
);

FILL FILL_3__8485_ (
);

OAI21X1 _12659_ (
    .A(_3484_),
    .B(vdd),
    .C(_3485_),
    .Y(_3425_[30])
);

FILL FILL_3__8065_ (
);

NAND3X1 _12239_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3218_)
);

FILL FILL_3__13708_ (
);

FILL FILL_1__14742_ (
);

FILL FILL_1__14322_ (
);

FILL FILL_0__13735_ (
);

FILL FILL_0__13315_ (
);

INVX1 _13600_ (
    .A(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_4109_)
);

FILL FILL_5__9772_ (
);

FILL FILL_5__9352_ (
);

INVX1 _16072_ (
    .A(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_6527_)
);

FILL FILL_1__9764_ (
);

FILL FILL_5__11642_ (
);

FILL FILL_1__9344_ (
);

FILL FILL_5__11222_ (
);

FILL FILL_2__16114_ (
);

FILL SFILL24280x71050 (
);

FILL FILL_4__10635_ (
);

FILL FILL_1__15947_ (
);

FILL FILL_1__15527_ (
);

FILL FILL_1__15107_ (
);

FILL FILL_1__10662_ (
);

FILL FILL_1__10242_ (
);

INVX1 _14805_ (
    .A(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_5289_)
);

FILL FILL112280x44050 (
);

FILL FILL_2__7687_ (
);

FILL FILL_6__13434_ (
);

FILL FILL_5__12847_ (
);

FILL FILL_3__13881_ (
);

FILL FILL_5__12427_ (
);

FILL FILL_3__13461_ (
);

FILL FILL_5__12007_ (
);

FILL FILL_3__13041_ (
);

FILL FILL_4__8974_ (
);

FILL FILL_4__8134_ (
);

FILL FILL_2__12874_ (
);

FILL FILL_2__12454_ (
);

FILL FILL_2__12034_ (
);

DFFSR _9199_ (
    .Q(\datapath_1.regfile_1.regOut[18] [25]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_1108_[25])
);

FILL FILL_1__11867_ (
);

FILL FILL_1__11447_ (
);

FILL FILL_1__11027_ (
);

FILL FILL_3__6971_ (
);

FILL FILL_5__16260_ (
);

FILL FILL_0__8874_ (
);

FILL FILL_0__8454_ (
);

DFFSR _10725_ (
    .Q(\datapath_1.regfile_1.regOut[30] [15]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_1888_[15])
);

INVX1 _10305_ (
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_1742_)
);

FILL FILL_5__6897_ (
);

FILL FILL_4__15673_ (
);

FILL FILL_4__15253_ (
);

DFFSR _13197_ (
    .Q(\datapath_1.mux_iord.din0 [22]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3685_[22])
);

FILL FILL_2__9413_ (
);

FILL FILL_0__11801_ (
);

FILL FILL_3__14666_ (
);

FILL FILL_3__14246_ (
);

FILL FILL_1__15280_ (
);

FILL FILL_1__6889_ (
);

FILL FILL_4__9759_ (
);

FILL FILL_4__9339_ (
);

FILL FILL_2__13659_ (
);

FILL FILL_2__13239_ (
);

FILL FILL_0__14693_ (
);

FILL SFILL33880x38050 (
);

FILL FILL_0__14273_ (
);

FILL FILL_1__7830_ (
);

FILL FILL_2__14600_ (
);

FILL FILL_0__9659_ (
);

FILL FILL_3__7756_ (
);

FILL FILL_3__7336_ (
);

FILL FILL_0__9239_ (
);

FILL SFILL94120x40050 (
);

FILL FILL_5__12180_ (
);

FILL FILL_4__16038_ (
);

FILL FILL_4__11593_ (
);

FILL FILL_4__11173_ (
);

FILL FILL_1__16065_ (
);

FILL FILL_5__8623_ (
);

FILL FILL_3__10166_ (
);

FILL FILL_5__8203_ (
);

FILL FILL_6_BUFX2_insert572 (
);

FILL FILL_0__15898_ (
);

INVX1 _15763_ (
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_6226_)
);

FILL FILL_0__15478_ (
);

NOR3X1 _15343_ (
    .A(_5813_),
    .B(_5815_),
    .C(_5814_),
    .Y(_5816_)
);

FILL FILL_0__15058_ (
);

FILL FILL_6_BUFX2_insert577 (
);

FILL FILL_0__10193_ (
);

FILL FILL_5__10913_ (
);

FILL FILL_1__8615_ (
);

FILL FILL_2__15805_ (
);

FILL FILL_2__10940_ (
);

FILL SFILL18600x16050 (
);

FILL FILL_5__13385_ (
);

FILL FILL_2__10520_ (
);

INVX1 _7685_ (
    .A(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_402_)
);

DFFSR _7265_ (
    .Q(\datapath_1.regfile_1.regOut[3] [11]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_133_[11])
);

FILL FILL_4__9092_ (
);

FILL FILL_4__12378_ (
);

FILL FILL_3__9902_ (
);

FILL SFILL94440x16050 (
);

FILL FILL_0__6940_ (
);

FILL FILL_2__6958_ (
);

FILL FILL_5__9408_ (
);

FILL SFILL23800x79050 (
);

NOR2X1 _16128_ (
    .A(_6579_),
    .B(_6580_),
    .Y(_6581_)
);

NOR2X1 _11683_ (
    .A(_2781_),
    .B(_2783_),
    .Y(_2784_)
);

FILL FILL_0__11398_ (
);

FILL SFILL84520x52050 (
);

NOR2X1 _11263_ (
    .A(_2380_),
    .B(_2381_),
    .Y(_2382_)
);

FILL SFILL23880x36050 (
);

FILL FILL_3__12732_ (
);

FILL FILL_3__12312_ (
);

FILL FILL_4__7825_ (
);

FILL FILL_2__11725_ (
);

FILL FILL_2__11305_ (
);

FILL FILL_2__14197_ (
);

FILL FILL_5__15951_ (
);

FILL FILL_5__15531_ (
);

FILL FILL_0__7725_ (
);

FILL FILL_5__15111_ (
);

FILL FILL_0__7305_ (
);

DFFSR _9831_ (
    .Q(\datapath_1.regfile_1.regOut[23] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_1433_[17])
);

OAI21X1 _9411_ (
    .A(_1287_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .C(_1288_),
    .Y(_1238_[25])
);

FILL FILL_4__14944_ (
);

FILL FILL_4__14524_ (
);

FILL FILL_4__14104_ (
);

OAI21X1 _12888_ (
    .A(_3596_),
    .B(vdd),
    .C(_3597_),
    .Y(_3555_[21])
);

OAI21X1 _12468_ (
    .A(_3377_),
    .B(vdd),
    .C(_3378_),
    .Y(_3360_[9])
);

NAND3X1 _12048_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [15]),
    .C(_3034__bF$buf0),
    .Y(_3082_)
);

FILL FILL_3__13937_ (
);

FILL FILL_1__14971_ (
);

FILL FILL_3__13517_ (
);

FILL FILL_1__14551_ (
);

FILL FILL_1__14131_ (
);

FILL FILL_5_BUFX2_insert590 (
);

FILL FILL_5_BUFX2_insert591 (
);

FILL FILL_5_BUFX2_insert592 (
);

FILL FILL_0__13964_ (
);

FILL FILL_5_BUFX2_insert593 (
);

FILL FILL_0__13544_ (
);

FILL FILL_5_BUFX2_insert594 (
);

FILL FILL_0__13124_ (
);

FILL FILL_5_BUFX2_insert595 (
);

FILL FILL_5_BUFX2_insert596 (
);

FILL FILL_5_BUFX2_insert597 (
);

FILL FILL_5_BUFX2_insert598 (
);

FILL FILL_5__9161_ (
);

FILL SFILL74120x81050 (
);

FILL FILL_5_BUFX2_insert599 (
);

FILL FILL_5__16316_ (
);

FILL FILL_1__9993_ (
);

FILL FILL_5__11871_ (
);

FILL FILL_5__11451_ (
);

FILL FILL_5__11031_ (
);

FILL FILL_1__9153_ (
);

FILL FILL_4__15729_ (
);

FILL FILL_4__15309_ (
);

FILL FILL_2__16343_ (
);

FILL FILL_3__9499_ (
);

FILL FILL_3__9079_ (
);

FILL FILL_4__10444_ (
);

FILL SFILL13800x77050 (
);

FILL FILL_4__10024_ (
);

FILL FILL_1__15756_ (
);

FILL FILL_1__15336_ (
);

FILL FILL_6__7084_ (
);

FILL FILL_1__10891_ (
);

FILL FILL_1__10051_ (
);

FILL FILL_0__14749_ (
);

INVX1 _14614_ (
    .A(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_5102_)
);

FILL FILL_0__14329_ (
);

FILL FILL_2__7496_ (
);

FILL FILL_2__7076_ (
);

FILL SFILL29000x48050 (
);

FILL FILL_5__12656_ (
);

FILL FILL_5__12236_ (
);

FILL FILL_3__13690_ (
);

FILL FILL_3__13270_ (
);

INVX1 _6956_ (
    .A(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_38_)
);

FILL FILL_4__8783_ (
);

FILL FILL_4__8363_ (
);

FILL FILL_4__11649_ (
);

FILL FILL_4__11229_ (
);

FILL FILL_2__12263_ (
);

FILL SFILL13800x32050 (
);

FILL FILL_1__11676_ (
);

FILL FILL_1__11256_ (
);

NAND3X1 _15819_ (
    .A(_6278_),
    .B(_6279_),
    .C(_6277_),
    .Y(_6280_)
);

FILL SFILL74040x43050 (
);

NOR2X1 _10954_ (
    .A(_2075_),
    .B(_2086_),
    .Y(_2087_)
);

FILL FILL_0__10669_ (
);

FILL FILL_0__8263_ (
);

INVX1 _10534_ (
    .A(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_1854_)
);

FILL FILL_0__10249_ (
);

INVX1 _10114_ (
    .A(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_1635_)
);

FILL FILL_4__15482_ (
);

FILL FILL_4__15062_ (
);

FILL FILL_2__9642_ (
);

FILL FILL_3__14895_ (
);

FILL FILL_3__14475_ (
);

FILL FILL_2__9222_ (
);

FILL FILL_0__11610_ (
);

FILL FILL_3__14055_ (
);

FILL FILL_4__9988_ (
);

FILL FILL_4__9148_ (
);

FILL FILL112360x77050 (
);

FILL FILL_2__13888_ (
);

FILL FILL_2__13468_ (
);

FILL FILL_0__14082_ (
);

FILL FILL_5__14802_ (
);

FILL FILL_6_CLKBUF1_insert173 (
);

FILL FILL_0__9888_ (
);

FILL FILL_3__7985_ (
);

FILL FILL_3__7565_ (
);

FILL FILL_0__9468_ (
);

NOR2X1 _11739_ (
    .A(_2835_),
    .B(_2801_),
    .Y(_2836_)
);

NOR2X1 _11319_ (
    .A(_2292_),
    .B(_2291_),
    .Y(_2438_)
);

FILL FILL_6_CLKBUF1_insert178 (
);

FILL FILL_1__13822_ (
);

FILL FILL_1__13402_ (
);

FILL FILL_4__16267_ (
);

FILL SFILL43960x28050 (
);

FILL FILL_1__16294_ (
);

FILL FILL_5__8852_ (
);

FILL FILL_3__10395_ (
);

FILL FILL_5__8012_ (
);

OAI22X1 _15992_ (
    .A(_5472__bF$buf1),
    .B(_5063_),
    .C(_5071_),
    .D(_5483__bF$buf4),
    .Y(_6449_)
);

NOR3X1 _15572_ (
    .A(_6018_),
    .B(_6039_),
    .C(_6028_),
    .Y(_6040_)
);

FILL FILL_0__15287_ (
);

OAI21X1 _15152_ (
    .A(_4074_),
    .B(_5535__bF$buf1),
    .C(_5629_),
    .Y(_5630_)
);

FILL FILL112360x32050 (
);

FILL FILL_3__16201_ (
);

FILL FILL_1__8844_ (
);

FILL FILL_5__10302_ (
);

FILL FILL_1__8004_ (
);

FILL FILL_2__15614_ (
);

FILL FILL_4_CLKBUF1_insert1074 (
);

FILL FILL_4_CLKBUF1_insert1075 (
);

FILL FILL_4_CLKBUF1_insert1076 (
);

FILL SFILL64040x41050 (
);

FILL FILL_4_CLKBUF1_insert1077 (
);

FILL FILL_4_CLKBUF1_insert1078 (
);

FILL FILL_1__14607_ (
);

OAI21X1 _7494_ (
    .A(_314_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_315_),
    .Y(_263_[26])
);

FILL FILL_4_CLKBUF1_insert1079 (
);

OAI21X1 _7074_ (
    .A(_95_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .C(_96_),
    .Y(_68_[14])
);

FILL FILL_4__12187_ (
);

FILL FILL_5__9637_ (
);

FILL FILL_5__9217_ (
);

INVX1 _16357_ (
    .A(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_6792_)
);

AND2X2 _11492_ (
    .A(_2604_),
    .B(_2297_),
    .Y(_2605_)
);

FILL FILL_5__11927_ (
);

NOR2X1 _11072_ (
    .A(_2189_),
    .B(_2190_),
    .Y(_2191_)
);

FILL FILL_3__12961_ (
);

FILL FILL_5__11507_ (
);

FILL FILL_1__9629_ (
);

FILL FILL_1__9209_ (
);

FILL FILL_3__12121_ (
);

FILL FILL_4__7634_ (
);

FILL FILL_4__7214_ (
);

FILL FILL_2__11954_ (
);

FILL FILL_5__14399_ (
);

FILL FILL_2__11534_ (
);

FILL FILL_3_CLKBUF1_insert120 (
);

FILL FILL_2__11114_ (
);

FILL FILL_3_CLKBUF1_insert121 (
);

OAI21X1 _8699_ (
    .A(_914_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .C(_915_),
    .Y(_913_[1])
);

FILL FILL_3_CLKBUF1_insert122 (
);

DFFSR _8279_ (
    .Q(\datapath_1.regfile_1.regOut[11] [1]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_653_[1])
);

FILL FILL_3_CLKBUF1_insert123 (
);

FILL FILL_3_CLKBUF1_insert124 (
);

FILL FILL_1__10947_ (
);

FILL FILL_3_CLKBUF1_insert125 (
);

FILL FILL_3_CLKBUF1_insert126 (
);

FILL FILL_1__10527_ (
);

FILL FILL_3_CLKBUF1_insert127 (
);

FILL FILL_1__10107_ (
);

FILL FILL_3_CLKBUF1_insert128 (
);

FILL FILL_3_CLKBUF1_insert129 (
);

FILL FILL_5__15760_ (
);

FILL FILL_5__15340_ (
);

FILL FILL_0__7954_ (
);

OAI21X1 _9640_ (
    .A(_1399_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1400_),
    .Y(_1368_[16])
);

FILL FILL_0__7114_ (
);

OAI21X1 _9220_ (
    .A(_1180_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .C(_1181_),
    .Y(_1173_[4])
);

FILL FILL_4__14753_ (
);

FILL FILL_4__14333_ (
);

OAI21X1 _12697_ (
    .A(_3553_),
    .B(IRWrite_bF$buf2),
    .C(_3554_),
    .Y(_3490_[0])
);

AOI22X1 _12277_ (
    .A(_2_[15]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump [15]),
    .Y(_3247_)
);

FILL FILL_2__8913_ (
);

FILL FILL_3__13746_ (
);

FILL FILL_3__13326_ (
);

FILL FILL_1__14780_ (
);

FILL FILL_1__14360_ (
);

FILL FILL_4__8839_ (
);

FILL FILL_2__12739_ (
);

FILL FILL_0__13773_ (
);

FILL FILL_2__12319_ (
);

FILL FILL_0__13353_ (
);

FILL FILL_5__9390_ (
);

FILL FILL_1__6910_ (
);

FILL FILL_3__6836_ (
);

FILL FILL_0__8739_ (
);

FILL FILL_5__16125_ (
);

FILL FILL_0__8319_ (
);

FILL FILL_5__11680_ (
);

FILL FILL_1__9382_ (
);

FILL FILL_5__11260_ (
);

FILL FILL_4__15958_ (
);

FILL FILL_4__15538_ (
);

FILL FILL_4__15118_ (
);

FILL FILL_2__16152_ (
);

FILL FILL_4__10673_ (
);

FILL FILL_4__10253_ (
);

FILL FILL_1__15985_ (
);

FILL FILL_1__15565_ (
);

FILL FILL_1__15145_ (
);

FILL FILL_5__7703_ (
);

FILL FILL_1__10280_ (
);

FILL FILL_0__14978_ (
);

INVX1 _14843_ (
    .A(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_5326_)
);

FILL FILL_0__14558_ (
);

FILL FILL_0__14138_ (
);

NOR2X1 _14423_ (
    .A(_4904_),
    .B(_4914_),
    .Y(_4915_)
);

NOR2X1 _14003_ (
    .A(_4503_),
    .B(_3983__bF$buf4),
    .Y(_4504_)
);

FILL SFILL44040x82050 (
);

FILL FILL_5__12885_ (
);

FILL FILL_5__12465_ (
);

FILL FILL_5__12045_ (
);

FILL FILL_4__8592_ (
);

FILL FILL_4__11878_ (
);

FILL FILL_4__11458_ (
);

FILL FILL_2__12492_ (
);

FILL FILL_4__11038_ (
);

FILL FILL_2__12072_ (
);

FILL FILL_5__8908_ (
);

FILL FILL_1__11485_ (
);

FILL FILL_1__11065_ (
);

NAND3X1 _15628_ (
    .A(_6085_),
    .B(_6086_),
    .C(_6093_),
    .Y(_6094_)
);

AOI21X1 _15208_ (
    .A(_5662_),
    .B(_5684_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [3])
);

FILL FILL_0__10898_ (
);

FILL FILL_0__8492_ (
);

INVX1 _10763_ (
    .A(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_1966_)
);

FILL FILL_0__8072_ (
);

FILL FILL_0__10058_ (
);

DFFSR _10343_ (
    .Q(\datapath_1.regfile_1.regOut[27] [17]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_1693_[17])
);

FILL FILL_3__11812_ (
);

FILL FILL_6__14677_ (
);

FILL FILL_6__14257_ (
);

FILL FILL_4__15291_ (
);

FILL FILL_4__6905_ (
);

FILL FILL_2__9871_ (
);

FILL FILL_2__10805_ (
);

FILL FILL112440x8050 (
);

FILL FILL_3__14284_ (
);

FILL FILL_2__9031_ (
);

FILL FILL_4__9797_ (
);

FILL SFILL84120x33050 (
);

FILL FILL_4__9377_ (
);

FILL FILL_2__13697_ (
);

FILL FILL_2__13277_ (
);

FILL FILL_5__14611_ (
);

OAI21X1 _8911_ (
    .A(_1035_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .C(_1036_),
    .Y(_978_[29])
);

FILL FILL_4__13604_ (
);

FILL SFILL88440x41050 (
);

FILL FILL_3__7374_ (
);

FILL FILL_0__9277_ (
);

INVX1 _11968_ (
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3020_)
);

NAND3X1 _11548_ (
    .A(_2470__bF$buf0),
    .B(_2645_),
    .C(_2657_),
    .Y(_2658_)
);

FILL FILL_5_CLKBUF1_insert160 (
);

INVX1 _11128_ (
    .A(_2246_),
    .Y(_2247_)
);

FILL FILL_5_CLKBUF1_insert161 (
);

FILL FILL_5_CLKBUF1_insert162 (
);

FILL FILL_1__13631_ (
);

FILL FILL_5_CLKBUF1_insert163 (
);

FILL FILL_1__13211_ (
);

FILL FILL_5_CLKBUF1_insert164 (
);

FILL FILL_4__16076_ (
);

FILL FILL_5_CLKBUF1_insert165 (
);

FILL FILL_5_CLKBUF1_insert166 (
);

FILL FILL_5_CLKBUF1_insert167 (
);

FILL FILL_5_CLKBUF1_insert168 (
);

FILL FILL_5_CLKBUF1_insert169 (
);

FILL FILL_0__12624_ (
);

FILL FILL_3__15489_ (
);

FILL FILL_0__12204_ (
);

FILL FILL_3__15069_ (
);

FILL FILL_6_BUFX2_insert950 (
);

FILL FILL_5__8661_ (
);

FILL FILL_5__8241_ (
);

FILL FILL_6_BUFX2_insert955 (
);

NAND3X1 _15381_ (
    .A(_5846_),
    .B(_5852_),
    .C(_5851_),
    .Y(_5853_)
);

FILL FILL_0__15096_ (
);

FILL FILL_5__15816_ (
);

FILL FILL_3__16010_ (
);

FILL FILL_5__10951_ (
);

FILL SFILL8440x14050 (
);

FILL FILL_1__8653_ (
);

FILL FILL_5__10531_ (
);

FILL FILL_5__10111_ (
);

FILL FILL_1__8233_ (
);

FILL FILL_4__14809_ (
);

FILL FILL_2__15843_ (
);

FILL FILL_3__8999_ (
);

FILL FILL_2__15423_ (
);

FILL SFILL109320x31050 (
);

FILL FILL_3__8579_ (
);

FILL FILL_2__15003_ (
);

FILL FILL_1__14836_ (
);

FILL FILL_1__14416_ (
);

FILL FILL_3__9940_ (
);

FILL FILL_0__13829_ (
);

FILL FILL_3__9520_ (
);

FILL FILL_3__9100_ (
);

FILL FILL_0__13409_ (
);

FILL FILL_2__6996_ (
);

FILL FILL_5__9866_ (
);

FILL FILL_5__9026_ (
);

FILL FILL_6__12743_ (
);

AOI22X1 _16166_ (
    .A(_5570__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .C(\datapath_1.regfile_1.regOut[6] [28]),
    .D(_5565__bF$buf3),
    .Y(_6618_)
);

FILL FILL_1__9858_ (
);

FILL FILL_5__11736_ (
);

FILL FILL_3__12770_ (
);

FILL FILL_5__11316_ (
);

FILL FILL_3__12350_ (
);

FILL FILL_1__9018_ (
);

FILL FILL_4__7863_ (
);

FILL FILL_2__16208_ (
);

FILL FILL_4__7443_ (
);

FILL FILL_4__10309_ (
);

FILL FILL_2__11763_ (
);

FILL FILL_2__11343_ (
);

NAND2X1 _8088_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_610_)
);

FILL FILL_1__10756_ (
);

FILL FILL_2_CLKBUF1_insert111 (
);

FILL FILL_2_CLKBUF1_insert112 (
);

FILL FILL_2_CLKBUF1_insert113 (
);

FILL FILL_2_CLKBUF1_insert114 (
);

FILL FILL_0__7763_ (
);

FILL FILL_0__7343_ (
);

FILL FILL_2_CLKBUF1_insert115 (
);

FILL FILL_6__8310_ (
);

FILL FILL_2_CLKBUF1_insert116 (
);

FILL FILL_2_CLKBUF1_insert117 (
);

FILL FILL_2_CLKBUF1_insert118 (
);

FILL FILL_2_CLKBUF1_insert119 (
);

FILL FILL_4__14982_ (
);

FILL FILL_4__14562_ (
);

FILL FILL_4__14142_ (
);

FILL SFILL64120x74050 (
);

NAND3X1 _12086_ (
    .A(_3108_),
    .B(_3109_),
    .C(_3110_),
    .Y(\datapath_1.mux_pcsrc.dout [24])
);

FILL FILL_3__13975_ (
);

FILL FILL_2__8722_ (
);

FILL FILL_3__13555_ (
);

FILL FILL_3__13135_ (
);

FILL FILL_4__8648_ (
);

FILL FILL_4__8228_ (
);

FILL FILL_5_BUFX2_insert970 (
);

FILL FILL_5_BUFX2_insert971 (
);

FILL FILL_2__12968_ (
);

FILL FILL_5_BUFX2_insert972 (
);

FILL FILL_2__12128_ (
);

FILL FILL_5_BUFX2_insert973 (
);

FILL FILL_0__13582_ (
);

FILL FILL_5_BUFX2_insert974 (
);

FILL FILL_0__13162_ (
);

FILL FILL_5_BUFX2_insert975 (
);

FILL FILL_5_BUFX2_insert976 (
);

FILL FILL_5_BUFX2_insert977 (
);

FILL FILL_5_BUFX2_insert978 (
);

FILL FILL_5_BUFX2_insert979 (
);

FILL FILL_0__8968_ (
);

FILL FILL_5__16354_ (
);

FILL FILL_0__8128_ (
);

OAI21X1 _10819_ (
    .A(_2002_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .C(_2003_),
    .Y(_1953_[25])
);

FILL FILL_1__12902_ (
);

FILL FILL_4__15767_ (
);

FILL FILL_4__15347_ (
);

FILL FILL_2__16381_ (
);

FILL FILL_4__10062_ (
);

FILL FILL_2__9927_ (
);

FILL FILL_2__9507_ (
);

FILL FILL_1__15794_ (
);

FILL FILL_1__15374_ (
);

FILL FILL_5__7932_ (
);

FILL FILL_0__14787_ (
);

FILL FILL_0__14367_ (
);

INVX1 _14652_ (
    .A(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_5139_)
);

FILL SFILL104200x19050 (
);

INVX1 _14232_ (
    .A(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_4728_)
);

FILL FILL112360x27050 (
);

FILL FILL_3__15701_ (
);

FILL FILL_1__7504_ (
);

FILL SFILL64040x36050 (
);

FILL FILL_5__12274_ (
);

OAI21X1 _6994_ (
    .A(_62_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_63_),
    .Y(_3_[30])
);

FILL SFILL113880x40050 (
);

FILL FILL_4__11687_ (
);

FILL FILL_4__11267_ (
);

FILL SFILL84120x1050 (
);

FILL FILL_1__16159_ (
);

FILL FILL_5__8717_ (
);

FILL FILL_1__11294_ (
);

AOI22X1 _15857_ (
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [20]),
    .C(\datapath_1.regfile_1.regOut[11] [20]),
    .D(_5496_),
    .Y(_6317_)
);

AOI21X1 _15437_ (
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .B(_5567_),
    .C(_5907_),
    .Y(_5908_)
);

AOI22X1 _15017_ (
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_5497_)
);

INVX2 _10992_ (
    .A(_2110_),
    .Y(_2111_)
);

OAI21X1 _10572_ (
    .A(_1878_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1879_),
    .Y(_1823_[28])
);

FILL FILL_0__10287_ (
);

OAI21X1 _10152_ (
    .A(_1659_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .C(_1660_),
    .Y(_1628_[16])
);

FILL FILL_3_BUFX2_insert1050 (
);

FILL FILL_3_BUFX2_insert1051 (
);

FILL FILL_1__8709_ (
);

FILL FILL_3_BUFX2_insert1052 (
);

FILL FILL_3__11621_ (
);

FILL FILL_3_BUFX2_insert1053 (
);

FILL FILL_3__11201_ (
);

FILL FILL_3_BUFX2_insert1054 (
);

FILL FILL_3_BUFX2_insert1055 (
);

FILL FILL_3_BUFX2_insert1056 (
);

FILL FILL_3_BUFX2_insert1057 (
);

FILL FILL_3_BUFX2_insert1058 (
);

FILL FILL_5__13899_ (
);

FILL FILL_3_BUFX2_insert1059 (
);

FILL FILL_2__10614_ (
);

FILL FILL_5__13479_ (
);

FILL FILL_2__9680_ (
);

FILL FILL_2__9260_ (
);

FILL FILL_3__14093_ (
);

DFFSR _7779_ (
    .Q(\datapath_1.regfile_1.regOut[7] [13]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_393_[13])
);

NAND2X1 _7359_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_246_)
);

FILL FILL_2__13086_ (
);

FILL FILL_5__14840_ (
);

FILL FILL_5__14420_ (
);

FILL FILL_5__14000_ (
);

OAI21X1 _8720_ (
    .A(_928_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_929_),
    .Y(_913_[8])
);

FILL SFILL89240x40050 (
);

DFFSR _8300_ (
    .Q(\datapath_1.regfile_1.regOut[11] [22]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_653_[22])
);

FILL FILL_1__12499_ (
);

FILL FILL_1__12079_ (
);

FILL FILL_4__13833_ (
);

FILL FILL_4__13413_ (
);

FILL FILL_3__7183_ (
);

NAND2X1 _11777_ (
    .A(_2139_),
    .B(_2341__bF$buf3),
    .Y(_2871_)
);

FILL FILL_0__9086_ (
);

INVX1 _11357_ (
    .A(_2322_),
    .Y(_2474_)
);

FILL FILL_3__12826_ (
);

FILL FILL_3__12406_ (
);

FILL FILL_1__13860_ (
);

FILL FILL_1__13440_ (
);

FILL FILL_1__13020_ (
);

FILL FILL_4_CLKBUF1_insert150 (
);

FILL FILL_4_CLKBUF1_insert151 (
);

FILL FILL_2__11819_ (
);

FILL FILL_4_CLKBUF1_insert152 (
);

FILL FILL_0__12853_ (
);

FILL FILL_3__15298_ (
);

FILL FILL_4_CLKBUF1_insert153 (
);

FILL FILL_0__12433_ (
);

FILL FILL_0__12013_ (
);

FILL FILL_4_CLKBUF1_insert154 (
);

FILL FILL_4_CLKBUF1_insert155 (
);

FILL FILL_4_CLKBUF1_insert156 (
);

FILL FILL_5__8890_ (
);

FILL FILL_4_CLKBUF1_insert157 (
);

FILL FILL_6__16212_ (
);

FILL FILL_5__8470_ (
);

FILL FILL_4_CLKBUF1_insert158 (
);

FILL FILL_4_CLKBUF1_insert159 (
);

INVX1 _15190_ (
    .A(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_5667_)
);

FILL FILL_5__15625_ (
);

FILL FILL_0__7819_ (
);

FILL FILL_5__15205_ (
);

NAND2X1 _9925_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1550_)
);

NAND2X1 _9505_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1331_)
);

FILL FILL_5__10760_ (
);

FILL FILL_1__8882_ (
);

FILL FILL_1__8462_ (
);

FILL FILL_4__14618_ (
);

FILL FILL_2__15652_ (
);

FILL FILL_2__15232_ (
);

FILL FILL_3__8388_ (
);

FILL FILL_1__14645_ (
);

FILL FILL_1__14225_ (
);

FILL FILL_0__13638_ (
);

INVX1 _13923_ (
    .A(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_4426_)
);

FILL FILL_0__13218_ (
);

NAND3X1 _13503_ (
    .A(_4004_),
    .B(_4006_),
    .C(_4013_),
    .Y(_4014_)
);

FILL FILL_5__9675_ (
);

FILL SFILL44040x77050 (
);

FILL FILL_5__9255_ (
);

OAI21X1 _16395_ (
    .A(_6816_),
    .B(gnd),
    .C(_6817_),
    .Y(_6769_[24])
);

FILL FILL_5__11965_ (
);

FILL FILL_5__11545_ (
);

FILL FILL_1__9667_ (
);

FILL FILL_1__9247_ (
);

FILL FILL_5__11125_ (
);

FILL FILL_2__16017_ (
);

FILL FILL_4__7672_ (
);

FILL FILL_4__10958_ (
);

FILL FILL_4__7252_ (
);

FILL FILL_2__11992_ (
);

FILL FILL_4__10538_ (
);

FILL FILL_2__11572_ (
);

FILL FILL_4__10118_ (
);

FILL FILL_2__11152_ (
);

FILL FILL_6__7178_ (
);

FILL FILL111880x51050 (
);

FILL FILL_1__10565_ (
);

FILL FILL_1__10145_ (
);

OAI22X1 _14708_ (
    .A(_5193_),
    .B(_3910_),
    .C(_3884__bF$buf0),
    .D(_5192_),
    .Y(_5194_)
);

FILL FILL_0__7992_ (
);

BUFX2 BUFX2_insert790 (
    .A(_5532_),
    .Y(_5532__bF$buf2)
);

FILL FILL_0__7572_ (
);

BUFX2 BUFX2_insert791 (
    .A(_5532_),
    .Y(_5532__bF$buf1)
);

BUFX2 BUFX2_insert792 (
    .A(_5532_),
    .Y(_5532__bF$buf0)
);

BUFX2 BUFX2_insert793 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf7 )
);

FILL SFILL109400x64050 (
);

BUFX2 BUFX2_insert794 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf6 )
);

BUFX2 BUFX2_insert795 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf5 )
);

FILL FILL_4__14791_ (
);

FILL FILL_4__14371_ (
);

BUFX2 BUFX2_insert796 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf4 )
);

BUFX2 BUFX2_insert797 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf3 )
);

FILL SFILL53800x3050 (
);

BUFX2 BUFX2_insert798 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf2 )
);

BUFX2 BUFX2_insert799 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf1 )
);

FILL FILL_2__8951_ (
);

FILL FILL_3__13784_ (
);

FILL FILL_2__8531_ (
);

FILL FILL_3__13364_ (
);

FILL FILL_2__8111_ (
);

FILL SFILL94280x3050 (
);

FILL FILL_4__8877_ (
);

FILL FILL_4__8457_ (
);

FILL FILL_2__12777_ (
);

FILL FILL_2__12357_ (
);

FILL FILL_0__13391_ (
);

FILL FILL_3__6874_ (
);

FILL FILL_5__16163_ (
);

FILL FILL_0__8777_ (
);

FILL FILL_0__8357_ (
);

OAI21X1 _10628_ (
    .A(_1895_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .C(_1896_),
    .Y(_1888_[4])
);

DFFSR _10208_ (
    .Q(\datapath_1.regfile_1.regOut[26] [10]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_1628_[10])
);

FILL FILL_4__15996_ (
);

FILL FILL_1__12711_ (
);

FILL FILL_4__15576_ (
);

FILL FILL_4__15156_ (
);

FILL FILL_2__16190_ (
);

FILL FILL_4__10291_ (
);

FILL FILL_2__9736_ (
);

FILL FILL_3__14989_ (
);

FILL FILL_3__14569_ (
);

FILL FILL_0__11704_ (
);

FILL FILL_3__14149_ (
);

FILL FILL_1__15183_ (
);

FILL FILL_5__7741_ (
);

FILL FILL_5__7321_ (
);

FILL FILL_0__14596_ (
);

AOI21X1 _14881_ (
    .A(_5342_),
    .B(_5363_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [29])
);

INVX1 _14461_ (
    .A(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_4952_)
);

FILL FILL_0__14176_ (
);

INVX1 _14041_ (
    .A(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_4541_)
);

FILL FILL_3__15930_ (
);

FILL FILL_3__15510_ (
);

FILL FILL_1__7733_ (
);

FILL FILL_1__7313_ (
);

FILL FILL_6__13090_ (
);

FILL FILL_2__14923_ (
);

FILL FILL_2__14503_ (
);

FILL FILL_3__7239_ (
);

FILL FILL_5__12083_ (
);

FILL FILL_1__13916_ (
);

FILL FILL_4__11496_ (
);

FILL FILL_4__11076_ (
);

FILL SFILL69160x43050 (
);

FILL FILL_3__8600_ (
);

FILL FILL_0__12909_ (
);

FILL FILL_1__16388_ (
);

FILL FILL_5__8526_ (
);

FILL FILL_3__10489_ (
);

FILL FILL_3__10069_ (
);

FILL FILL_5__8106_ (
);

NOR2X1 _15666_ (
    .A(_6130_),
    .B(_6128_),
    .Y(_6131_)
);

FILL SFILL74120x26050 (
);

NAND3X1 _15246_ (
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5722_)
);

OAI21X1 _10381_ (
    .A(_1771_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .C(_1772_),
    .Y(_1758_[7])
);

FILL FILL_5__10816_ (
);

FILL FILL_1__8518_ (
);

FILL FILL_3__11850_ (
);

FILL FILL_3__11430_ (
);

FILL FILL_3__11010_ (
);

FILL FILL_2__15708_ (
);

FILL SFILL99320x75050 (
);

FILL FILL_4__6943_ (
);

FILL FILL_0__16322_ (
);

FILL FILL_2__10423_ (
);

FILL FILL_5__13288_ (
);

FILL FILL_2__10003_ (
);

NAND2X1 _7588_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_358_)
);

NAND2X1 _7168_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_139_)
);

FILL FILL_3__9805_ (
);

FILL FILL_0__6843_ (
);

FILL FILL_4__13642_ (
);

FILL SFILL64120x69050 (
);

FILL FILL_4__13222_ (
);

AOI21X1 _11586_ (
    .A(_2216_),
    .B(_2176_),
    .C(_2258_),
    .Y(_2693_)
);

NOR2X1 _11166_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2285_)
);

FILL FILL_2__7802_ (
);

FILL FILL_3__12635_ (
);

FILL FILL_3__12215_ (
);

FILL FILL_4__7728_ (
);

FILL FILL_4__7308_ (
);

FILL FILL_2__11628_ (
);

FILL FILL_0__12662_ (
);

FILL FILL_2__11208_ (
);

FILL SFILL99320x30050 (
);

FILL FILL_0__12242_ (
);

FILL SFILL38680x14050 (
);

FILL SFILL23800x2050 (
);

FILL SFILL23720x7050 (
);

FILL FILL_5__15854_ (
);

FILL FILL_5__15434_ (
);

FILL FILL_0__7628_ (
);

FILL FILL_5__15014_ (
);

FILL FILL_0__7208_ (
);

NAND2X1 _9734_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1443_)
);

FILL SFILL59160x41050 (
);

DFFSR _9314_ (
    .Q(\datapath_1.regfile_1.regOut[19] [12]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_1173_[12])
);

FILL FILL_1__8271_ (
);

FILL FILL_4__14847_ (
);

FILL FILL_2__15881_ (
);

FILL FILL_4__14427_ (
);

FILL FILL_4__14007_ (
);

FILL FILL_2__15461_ (
);

FILL FILL_2__15041_ (
);

FILL FILL_3__8197_ (
);

FILL SFILL64120x24050 (
);

FILL SFILL3640x3050 (
);

FILL FILL_1__14874_ (
);

FILL FILL_1__14454_ (
);

FILL FILL_1__14034_ (
);

FILL FILL_0__13867_ (
);

FILL FILL_0__13447_ (
);

INVX1 _13732_ (
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_4239_)
);

FILL SFILL89320x73050 (
);

OAI21X1 _13312_ (
    .A(_3843_),
    .B(_3844_),
    .C(_3750_),
    .Y(_3845_)
);

FILL FILL_0__13027_ (
);

FILL FILL_5__9484_ (
);

FILL FILL_5__16219_ (
);

FILL FILL_1__9896_ (
);

FILL FILL_5__11774_ (
);

FILL FILL_1__9476_ (
);

FILL FILL_5__11354_ (
);

FILL FILL_2__16246_ (
);

FILL FILL_4__7481_ (
);

FILL FILL_4__10767_ (
);

FILL FILL_4__7061_ (
);

FILL FILL_2__11381_ (
);

FILL SFILL54120x67050 (
);

FILL FILL_1__15659_ (
);

FILL FILL_1__15239_ (
);

FILL FILL_1__10794_ (
);

FILL FILL_1__10374_ (
);

OAI22X1 _14937_ (
    .A(_5417_),
    .B(_3890_),
    .C(_3954__bF$buf4),
    .D(_5416_),
    .Y(_5418_)
);

INVX1 _14517_ (
    .A(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_5007_)
);

FILL FILL_0__7381_ (
);

FILL FILL_6__13986_ (
);

FILL FILL_3__10701_ (
);

FILL FILL_6__13146_ (
);

FILL FILL_4__14180_ (
);

FILL FILL_5__12979_ (
);

FILL FILL_2__8760_ (
);

FILL FILL_3__13593_ (
);

FILL FILL_5__12139_ (
);

FILL FILL_2__8340_ (
);

BUFX2 _6859_ (
    .A(_1_[21]),
    .Y(memoryAddress[21])
);

FILL FILL_3__13173_ (
);

FILL FILL_4__8266_ (
);

FILL FILL_2__12586_ (
);

FILL FILL_2__12166_ (
);

FILL FILL_5__13920_ (
);

FILL FILL_5__13500_ (
);

FILL SFILL89240x35050 (
);

FILL FILL_1__11999_ (
);

OAI21X1 _7800_ (
    .A(_521_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .C(_522_),
    .Y(_458_[0])
);

FILL SFILL54120x22050 (
);

FILL FILL_1__11579_ (
);

FILL FILL_1__11159_ (
);

FILL FILL_4__12913_ (
);

FILL FILL_5__16392_ (
);

FILL FILL_0__8586_ (
);

DFFSR _10857_ (
    .Q(\datapath_1.regfile_1.regOut[31] [19]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_1953_[19])
);

NAND2X1 _10437_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1810_)
);

NAND2X1 _10017_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1591_)
);

FILL SFILL79320x71050 (
);

FILL FILL_3__11906_ (
);

FILL SFILL18680x55050 (
);

FILL FILL_4__15385_ (
);

FILL FILL_1__12520_ (
);

FILL FILL_1__12100_ (
);

FILL FILL_0__11933_ (
);

FILL FILL_3__14798_ (
);

FILL FILL_2__9545_ (
);

FILL FILL_2__9125_ (
);

FILL FILL_3__14378_ (
);

FILL FILL_0__11513_ (
);

FILL SFILL54040x29050 (
);

FILL FILL_5__7970_ (
);

FILL FILL_5__7550_ (
);

NAND3X1 _14690_ (
    .A(_5175_),
    .B(_5176_),
    .C(_5174_),
    .Y(_5177_)
);

INVX1 _14270_ (
    .A(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_4765_)
);

FILL FILL_5__14705_ (
);

FILL SFILL79240x78050 (
);

FILL FILL_1__7962_ (
);

FILL FILL_1__7542_ (
);

FILL FILL_1__7122_ (
);

FILL FILL_2__14732_ (
);

FILL FILL_2__14312_ (
);

FILL FILL_3__7888_ (
);

FILL FILL_3__7468_ (
);

FILL FILL_3__7048_ (
);

FILL FILL_1__13725_ (
);

FILL FILL_1__13305_ (
);

FILL SFILL18680x10050 (
);

FILL SFILL33880x9050 (
);

FILL FILL_0__12718_ (
);

FILL FILL_1__16197_ (
);

FILL FILL_5__8755_ (
);

FILL FILL_5__8335_ (
);

FILL FILL_3__10298_ (
);

NOR3X1 _15895_ (
    .A(_4978_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6354_)
);

INVX1 _15475_ (
    .A(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_5945_)
);

NAND3X1 _15055_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5477_),
    .C(_5468_),
    .Y(_5535_)
);

FILL FILL_3__16104_ (
);

NAND2X1 _10190_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1686_)
);

FILL FILL_5__10625_ (
);

FILL FILL_1__8747_ (
);

FILL FILL_1__8327_ (
);

FILL FILL_2__15937_ (
);

FILL FILL_2__15517_ (
);

FILL FILL_0__16131_ (
);

FILL FILL_2__10652_ (
);

FILL FILL_5__13097_ (
);

FILL FILL_2__10232_ (
);

DFFSR _7397_ (
    .Q(\datapath_1.regfile_1.regOut[4] [15]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_198_[15])
);

FILL FILL111880x46050 (
);

FILL FILL_3_BUFX2_insert300 (
);

FILL FILL_3__9614_ (
);

FILL SFILL109320x3050 (
);

FILL FILL_3_BUFX2_insert301 (
);

FILL FILL_3_BUFX2_insert302 (
);

FILL FILL_3_BUFX2_insert303 (
);

FILL FILL_3_BUFX2_insert304 (
);

FILL FILL_3_BUFX2_insert305 (
);

FILL FILL_3_BUFX2_insert306 (
);

FILL FILL_3_BUFX2_insert307 (
);

FILL SFILL48760x49050 (
);

FILL FILL_3_BUFX2_insert308 (
);

FILL FILL_4__13871_ (
);

FILL FILL_3_BUFX2_insert309 (
);

FILL FILL_4__13451_ (
);

FILL FILL_4__13031_ (
);

OAI21X1 _11395_ (
    .A(_2510_),
    .B(_2171_),
    .C(_2511_),
    .Y(_2512_)
);

FILL FILL_2__7611_ (
);

FILL FILL_3__12864_ (
);

FILL FILL_3__12444_ (
);

FILL FILL_3__12024_ (
);

FILL FILL_4__7957_ (
);

FILL FILL_4__7117_ (
);

FILL FILL_2__11857_ (
);

FILL FILL_0__12891_ (
);

FILL FILL_2__11437_ (
);

FILL FILL_0__12471_ (
);

FILL FILL_2__11017_ (
);

FILL FILL_0__12051_ (
);

FILL SFILL109800x28050 (
);

FILL FILL_5__15663_ (
);

FILL FILL_5__15243_ (
);

FILL FILL_0__7857_ (
);

FILL FILL_0__7437_ (
);

DFFSR _9963_ (
    .Q(\datapath_1.regfile_1.regOut[24] [21]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1498_[21])
);

INVX1 _9543_ (
    .A(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_1356_)
);

INVX1 _9123_ (
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_1137_)
);

FILL FILL_1__8080_ (
);

FILL FILL_4__14656_ (
);

FILL FILL_2__15690_ (
);

FILL FILL_4__14236_ (
);

FILL FILL_2__15270_ (
);

FILL SFILL109400x14050 (
);

FILL FILL_3__13649_ (
);

FILL FILL_3__13229_ (
);

FILL FILL_1__14683_ (
);

FILL FILL_1__14263_ (
);

FILL FILL_0_BUFX2_insert430 (
);

FILL FILL_0_BUFX2_insert431 (
);

FILL FILL_0_BUFX2_insert432 (
);

FILL FILL_0_BUFX2_insert433 (
);

FILL FILL_0_BUFX2_insert434 (
);

FILL FILL_0__13676_ (
);

AOI22X1 _13961_ (
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .B(_3891__bF$buf1),
    .C(_3998__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_4463_)
);

FILL SFILL69240x31050 (
);

FILL FILL_0__13256_ (
);

INVX8 _13541_ (
    .A(_3978_),
    .Y(_4051_)
);

FILL FILL_0_BUFX2_insert435 (
);

INVX1 _13121_ (
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_3712_)
);

FILL FILL_0_BUFX2_insert436 (
);

FILL FILL_0_BUFX2_insert437 (
);

FILL FILL_0_BUFX2_insert438 (
);

FILL FILL_5__9293_ (
);

FILL FILL_0_BUFX2_insert439 (
);

FILL FILL_5__16028_ (
);

FILL FILL_5__11583_ (
);

FILL FILL_1__9285_ (
);

FILL FILL_5__11163_ (
);

FILL FILL_2__16055_ (
);

FILL SFILL99400x63050 (
);

FILL FILL_4__10996_ (
);

FILL FILL_4__7290_ (
);

FILL FILL_4__10576_ (
);

FILL SFILL69160x38050 (
);

FILL FILL_4__10156_ (
);

FILL FILL_2__11190_ (
);

FILL FILL_1__15888_ (
);

FILL FILL_1__15468_ (
);

FILL FILL_1__15048_ (
);

FILL FILL_5__7606_ (
);

FILL FILL_1__10183_ (
);

AOI22X1 _14746_ (
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .B(_3894_),
    .C(_4051__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_5231_)
);

INVX1 _14326_ (
    .A(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_4820_)
);

FILL FILL_0__7190_ (
);

FILL FILL_3__10930_ (
);

FILL FILL_3__10510_ (
);

FILL FILL_0__15822_ (
);

FILL SFILL104680x77050 (
);

FILL FILL_0__15402_ (
);

FILL FILL_5__12788_ (
);

FILL FILL_5__12368_ (
);

FILL FILL_4__8495_ (
);

FILL FILL_4__8075_ (
);

FILL FILL_2__12395_ (
);

FILL FILL_1__11388_ (
);

FILL FILL_4__12722_ (
);

FILL FILL_4__12302_ (
);

FILL FILL_6__9782_ (
);

FILL FILL_0__8395_ (
);

NAND2X1 _10666_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1922_)
);

NAND2X1 _10246_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1703_)
);

FILL FILL_3__11715_ (
);

FILL FILL_4__15194_ (
);

FILL FILL_2__10708_ (
);

FILL FILL_2__9774_ (
);

FILL FILL_2__9354_ (
);

FILL FILL_0__11742_ (
);

FILL FILL_3__14187_ (
);

FILL FILL_0__11322_ (
);

FILL FILL_6__15521_ (
);

FILL FILL_6__15101_ (
);

FILL FILL_5__14934_ (
);

FILL SFILL89400x61050 (
);

FILL FILL_5__14514_ (
);

FILL SFILL59160x36050 (
);

DFFSR _8814_ (
    .Q(\datapath_1.regfile_1.regOut[15] [24]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_913_[24])
);

FILL FILL_1__7351_ (
);

FILL FILL_4__13927_ (
);

FILL FILL_2__14961_ (
);

FILL FILL_4__13507_ (
);

FILL FILL_2__14541_ (
);

FILL FILL_3__7697_ (
);

FILL FILL_2__14121_ (
);

FILL SFILL64120x19050 (
);

FILL FILL_1__13954_ (
);

FILL FILL_4__16399_ (
);

FILL FILL_1__13534_ (
);

FILL FILL_1__13114_ (
);

FILL SFILL89320x68050 (
);

DFFSR _12812_ (
    .Q(\datapath_1.PCJump [23]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[21])
);

FILL FILL_0__12527_ (
);

FILL FILL_0__12107_ (
);

FILL FILL_5__8984_ (
);

FILL FILL_5__8144_ (
);

FILL FILL_6__11441_ (
);

FILL FILL_6__11021_ (
);

NOR2X1 _15284_ (
    .A(_5757_),
    .B(_5758_),
    .Y(_5759_)
);

FILL FILL_5__15719_ (
);

FILL FILL_3__16333_ (
);

FILL FILL_1__8976_ (
);

FILL FILL_5__10434_ (
);

FILL FILL_1__8136_ (
);

FILL FILL_5__10014_ (
);

FILL FILL_2__15746_ (
);

FILL FILL_2__15326_ (
);

FILL FILL_4__6981_ (
);

FILL FILL_0__16360_ (
);

FILL FILL_2__10881_ (
);

FILL FILL_2__10041_ (
);

FILL FILL_1__14739_ (
);

FILL FILL_1__14319_ (
);

FILL FILL_3__9423_ (
);

FILL FILL_3__9003_ (
);

FILL FILL_0__6881_ (
);

FILL FILL_2__6899_ (
);

FILL FILL_5__9769_ (
);

FILL FILL_5__9349_ (
);

FILL FILL_4__13680_ (
);

FILL FILL_4__13260_ (
);

OAI22X1 _16069_ (
    .A(_5466__bF$buf4),
    .B(_5147_),
    .C(_5139_),
    .D(_5483__bF$buf2),
    .Y(_6524_)
);

FILL FILL_2__7840_ (
);

FILL FILL_5__11639_ (
);

FILL FILL_5__11219_ (
);

FILL FILL_2__7420_ (
);

FILL FILL_3__12253_ (
);

FILL SFILL18760x43050 (
);

FILL FILL_4__7346_ (
);

FILL FILL_2__11666_ (
);

FILL FILL_2__11246_ (
);

FILL FILL_0__12280_ (
);

FILL FILL_1__10659_ (
);

FILL FILL_1__10239_ (
);

FILL FILL_5__15892_ (
);

FILL FILL_5__15472_ (
);

FILL FILL_5__15052_ (
);

INVX1 _9772_ (
    .A(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_1468_)
);

FILL FILL_0__7246_ (
);

INVX1 _9352_ (
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_1249_)
);

FILL SFILL79320x66050 (
);

FILL FILL_4__14885_ (
);

FILL FILL_4__14465_ (
);

FILL FILL_1__11600_ (
);

FILL FILL_4__14045_ (
);

FILL FILL_3__13878_ (
);

FILL FILL_2__8625_ (
);

FILL FILL_2__8205_ (
);

FILL FILL_3__13458_ (
);

FILL FILL_1__14492_ (
);

FILL FILL_3__13038_ (
);

FILL FILL_1__14072_ (
);

AOI22X1 _13770_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [6]),
    .C(\datapath_1.regfile_1.regOut[6] [6]),
    .D(_4001__bF$buf2),
    .Y(_4276_)
);

FILL FILL_0__13485_ (
);

OAI21X1 _13350_ (
    .A(_3752_),
    .B(_3767_),
    .C(_3868_),
    .Y(_3869_)
);

FILL FILL_4__9912_ (
);

FILL FILL_2__13812_ (
);

FILL FILL_3__6968_ (
);

FILL FILL_5__16257_ (
);

FILL FILL_5__11392_ (
);

FILL FILL_1__9094_ (
);

FILL FILL_2__16284_ (
);

FILL FILL_4__10385_ (
);

FILL FILL_0__9812_ (
);

FILL FILL_1__15697_ (
);

FILL FILL_1__15277_ (
);

FILL FILL_5__7835_ (
);

FILL FILL_5__7415_ (
);

FILL FILL111960x34050 (
);

NOR2X1 _14975_ (
    .A(_5455_),
    .B(_5452_),
    .Y(_5456_)
);

OAI22X1 _14555_ (
    .A(_5042_),
    .B(_3884__bF$buf0),
    .C(_3959_),
    .D(_5043_),
    .Y(_5044_)
);

AOI22X1 _14135_ (
    .A(_4038__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [14]),
    .C(\datapath_1.regfile_1.regOut[27] [14]),
    .D(_4129_),
    .Y(_4633_)
);

FILL FILL_3__15604_ (
);

FILL FILL_1__7827_ (
);

FILL SFILL79240x28050 (
);

FILL FILL_0__15631_ (
);

FILL FILL_0__15211_ (
);

FILL FILL_5__12597_ (
);

FILL FILL_5__12177_ (
);

BUFX2 _6897_ (
    .A(_2_[27]),
    .Y(memoryWriteData[27])
);

FILL FILL_1__11197_ (
);

FILL FILL_6__11917_ (
);

FILL FILL_4__12951_ (
);

FILL FILL_4__12531_ (
);

FILL FILL_4__12111_ (
);

FILL FILL_6__9591_ (
);

OAI21X1 _10895_ (
    .A(_2038_),
    .B(_2040_),
    .C(_2037_),
    .Y(_2041_)
);

DFFSR _10475_ (
    .Q(\datapath_1.regfile_1.regOut[28] [21]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_1758_[21])
);

INVX1 _10055_ (
    .A(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_1616_)
);

FILL FILL_3__11944_ (
);

FILL FILL_3__11524_ (
);

FILL FILL_3__11104_ (
);

FILL FILL_0__16416_ (
);

FILL FILL_2__10937_ (
);

FILL SFILL114360x53050 (
);

FILL FILL_0__11971_ (
);

FILL FILL_2__10517_ (
);

FILL FILL_2__9163_ (
);

FILL FILL_0__11551_ (
);

FILL FILL_0__11131_ (
);

FILL FILL_4__9089_ (
);

FILL FILL_5__14743_ (
);

FILL FILL_0__6937_ (
);

FILL FILL_5__14323_ (
);

INVX1 _8623_ (
    .A(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_885_)
);

INVX1 _8203_ (
    .A(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_666_)
);

FILL FILL_1__7580_ (
);

FILL FILL_1__7160_ (
);

FILL FILL_4__13736_ (
);

FILL FILL_4__13316_ (
);

FILL FILL_2__14770_ (
);

FILL FILL_2__14350_ (
);

FILL FILL_3__7086_ (
);

FILL FILL_3__12729_ (
);

FILL FILL_1__13763_ (
);

FILL FILL_3__12309_ (
);

FILL FILL_1__13343_ (
);

FILL SFILL69240x26050 (
);

FILL FILL_0__12756_ (
);

INVX1 _12621_ (
    .A(\datapath_1.Data [18]),
    .Y(_3460_)
);

FILL FILL_0__12336_ (
);

OAI21X1 _12201_ (
    .A(_3186_),
    .B(ALUSrcA_bF$buf5),
    .C(_3187_),
    .Y(\datapath_1.alu_1.ALUInA [28])
);

FILL FILL_5__8373_ (
);

FILL FILL_5__15948_ (
);

AOI22X1 _15093_ (
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .B(_5571_),
    .C(_5570__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_5572_)
);

FILL FILL_5__15528_ (
);

FILL FILL_5__15108_ (
);

DFFSR _9828_ (
    .Q(\datapath_1.regfile_1.regOut[23] [14]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_1433_[14])
);

FILL FILL_3__16142_ (
);

OAI21X1 _9408_ (
    .A(_1285_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1286_),
    .Y(_1238_[24])
);

FILL FILL_5__10663_ (
);

FILL FILL_1__8785_ (
);

FILL FILL_5__10243_ (
);

FILL FILL_1__8365_ (
);

FILL FILL_2__15975_ (
);

FILL FILL_2__15555_ (
);

FILL SFILL99400x58050 (
);

FILL FILL_2__15135_ (
);

FILL FILL_2__10690_ (
);

FILL FILL_2__10270_ (
);

FILL FILL_1__14968_ (
);

FILL FILL_1__14548_ (
);

FILL FILL_1__14128_ (
);

FILL FILL_3__9652_ (
);

FILL FILL_3__9232_ (
);

NAND3X1 _13826_ (
    .A(_4322_),
    .B(_4323_),
    .C(_4330_),
    .Y(_4331_)
);

INVX1 _13406_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_3918_)
);

FILL FILL_5__9998_ (
);

FILL SFILL104360x51050 (
);

FILL FILL_5__9158_ (
);

NAND3X1 _16298_ (
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf4),
    .Y(_6747_)
);

FILL FILL_0__14902_ (
);

FILL FILL_5__11868_ (
);

FILL FILL_5__11448_ (
);

FILL FILL_3__12482_ (
);

FILL FILL_5__11028_ (
);

FILL FILL_3__12062_ (
);

FILL FILL_4__7995_ (
);

FILL FILL_4__7575_ (
);

FILL FILL_2__11895_ (
);

FILL FILL_2__11475_ (
);

FILL FILL_2__11055_ (
);

FILL SFILL99400x13050 (
);

FILL FILL_1__10888_ (
);

FILL FILL_1__10048_ (
);

FILL SFILL49720x74050 (
);

FILL FILL_4__11802_ (
);

FILL FILL_5__15281_ (
);

FILL FILL_0__7475_ (
);

FILL FILL_6__8862_ (
);

FILL FILL_0__7055_ (
);

DFFSR _9581_ (
    .Q(\datapath_1.regfile_1.regOut[21] [23]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1303_[23])
);

OAI21X1 _9161_ (
    .A(_1161_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .C(_1162_),
    .Y(_1108_[27])
);

FILL FILL_4__14694_ (
);

FILL FILL_4__14274_ (
);

FILL FILL_2__8854_ (
);

FILL FILL_0__10822_ (
);

FILL FILL_3__13687_ (
);

FILL FILL_2__8014_ (
);

FILL FILL_3__13267_ (
);

FILL FILL_0__10402_ (
);

FILL FILL_0_BUFX2_insert810 (
);

FILL FILL_0_BUFX2_insert811 (
);

FILL FILL_0_BUFX2_insert812 (
);

FILL FILL_0_BUFX2_insert813 (
);

FILL FILL_0_BUFX2_insert814 (
);

FILL FILL_0__13294_ (
);

FILL FILL_0_BUFX2_insert815 (
);

FILL SFILL89400x56050 (
);

FILL FILL_0_BUFX2_insert816 (
);

FILL FILL_0_BUFX2_insert817 (
);

FILL FILL_0_BUFX2_insert818 (
);

FILL FILL_0_BUFX2_insert819 (
);

FILL FILL_1__6851_ (
);

FILL FILL_4__9721_ (
);

FILL FILL_4__9301_ (
);

FILL FILL_2__13621_ (
);

FILL FILL_5__16066_ (
);

FILL FILL_4__15899_ (
);

FILL FILL_1__12614_ (
);

FILL FILL_4__15479_ (
);

FILL FILL_4__15059_ (
);

FILL FILL_2__16093_ (
);

FILL FILL_4__10194_ (
);

FILL SFILL73720x78050 (
);

FILL FILL_2__9639_ (
);

FILL FILL_0__9621_ (
);

FILL FILL_2__9219_ (
);

FILL FILL_0__11607_ (
);

FILL FILL_1__15086_ (
);

FILL FILL_5__7224_ (
);

FILL FILL_4__16000_ (
);

FILL FILL_6__10941_ (
);

FILL FILL_0__14499_ (
);

INVX1 _14784_ (
    .A(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_5269_)
);

INVX1 _14364_ (
    .A(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_4857_)
);

FILL FILL_0__14079_ (
);

FILL FILL_3__15833_ (
);

FILL FILL_3__15413_ (
);

FILL FILL_1__7636_ (
);

FILL FILL_1__7216_ (
);

FILL SFILL94280x62050 (
);

FILL FILL_2__14826_ (
);

FILL FILL_0__15860_ (
);

FILL FILL_2__14406_ (
);

FILL FILL_0__15440_ (
);

FILL FILL_0__15020_ (
);

FILL FILL_1__13819_ (
);

FILL FILL_4__11399_ (
);

FILL FILL_3__8503_ (
);

FILL SFILL33960x58050 (
);

FILL FILL_5__8849_ (
);

FILL SFILL89320x18050 (
);

FILL FILL_5__8009_ (
);

FILL SFILL94680x31050 (
);

INVX1 _15989_ (
    .A(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_6446_)
);

FILL FILL_4__12760_ (
);

OAI22X1 _15569_ (
    .A(_5518__bF$buf1),
    .B(_4544_),
    .C(_5469__bF$buf2),
    .D(_4567_),
    .Y(_6037_)
);

FILL FILL_4__12340_ (
);

OAI22X1 _15149_ (
    .A(_4071_),
    .B(_5544__bF$buf0),
    .C(_5499__bF$buf0),
    .D(_5626_),
    .Y(_5627_)
);

INVX1 _10284_ (
    .A(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_1728_)
);

FILL FILL_2__6920_ (
);

FILL FILL_3__11753_ (
);

FILL SFILL18760x38050 (
);

FILL FILL_3__11333_ (
);

FILL SFILL33560x44050 (
);

FILL FILL_4__6846_ (
);

FILL FILL_0__16225_ (
);

FILL FILL_2__10746_ (
);

FILL FILL_2__9392_ (
);

FILL FILL_0__11780_ (
);

FILL FILL_0__11360_ (
);

FILL SFILL23640x80050 (
);

FILL FILL_5__14972_ (
);

FILL FILL_5__14552_ (
);

FILL FILL_5__14132_ (
);

INVX1 _8852_ (
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_997_)
);

DFFSR _8432_ (
    .Q(\datapath_1.regfile_1.regOut[12] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_718_[26])
);

OAI21X1 _8012_ (
    .A(_578_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_579_),
    .Y(_523_[28])
);

FILL FILL_4__13965_ (
);

FILL FILL_4__13545_ (
);

FILL FILL_4__13125_ (
);

INVX1 _11489_ (
    .A(_2301_),
    .Y(_2602_)
);

XNOR2X1 _11069_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2188_)
);

FILL FILL_2__7705_ (
);

FILL FILL_3__12958_ (
);

FILL FILL_1__13992_ (
);

FILL FILL_3__12118_ (
);

FILL FILL_1__13572_ (
);

FILL FILL_1__13152_ (
);

FILL SFILL84280x60050 (
);

FILL FILL_0__12985_ (
);

INVX1 _12850_ (
    .A(\datapath_1.a [9]),
    .Y(_3572_)
);

INVX1 _12430_ (
    .A(ALUOut[29]),
    .Y(_3352_)
);

FILL FILL_0__12145_ (
);

NAND3X1 _12010_ (
    .A(_3051_),
    .B(_3052_),
    .C(_3053_),
    .Y(\datapath_1.mux_pcsrc.dout [5])
);

FILL FILL_5__8182_ (
);

FILL FILL_5__15757_ (
);

FILL FILL_5__15337_ (
);

FILL FILL_3__16371_ (
);

OAI21X1 _9637_ (
    .A(_1397_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .C(_1398_),
    .Y(_1368_[15])
);

OAI21X1 _9217_ (
    .A(_1178_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .C(_1179_),
    .Y(_1173_[3])
);

FILL FILL_5__10892_ (
);

FILL FILL_1__8594_ (
);

FILL FILL_5__10052_ (
);

FILL FILL_5_BUFX2_insert1000 (
);

FILL FILL_5_BUFX2_insert1001 (
);

FILL FILL_2__15784_ (
);

FILL FILL_5_BUFX2_insert1002 (
);

FILL FILL_5_BUFX2_insert1003 (
);

FILL FILL_2__15364_ (
);

FILL FILL_5_BUFX2_insert1004 (
);

FILL FILL_5_BUFX2_insert1005 (
);

FILL FILL_5_BUFX2_insert1006 (
);

FILL FILL_5_BUFX2_insert1007 (
);

FILL FILL_5_BUFX2_insert1008 (
);

FILL FILL_5_BUFX2_insert1009 (
);

FILL FILL_1__14777_ (
);

FILL FILL_1__14357_ (
);

FILL FILL_5__6915_ (
);

FILL FILL_3__9881_ (
);

NAND3X1 _13635_ (
    .A(_4134_),
    .B(_4136_),
    .C(_4143_),
    .Y(_4144_)
);

FILL FILL_3__9041_ (
);

NOR2X1 _13215_ (
    .A(\datapath_1.a3 [2]),
    .B(_3757_),
    .Y(_3758_)
);

FILL FILL_5__9387_ (
);

FILL FILL_1__6907_ (
);

FILL FILL_6__12264_ (
);

FILL FILL_0__14711_ (
);

FILL FILL_1__9799_ (
);

FILL FILL_5__11677_ (
);

FILL FILL_1__9379_ (
);

FILL FILL_5__11257_ (
);

FILL FILL_3__12291_ (
);

FILL SFILL69320x59050 (
);

FILL FILL_2__16149_ (
);

FILL FILL_2__11284_ (
);

FILL SFILL114440x41050 (
);

FILL FILL_2_BUFX2_insert340 (
);

FILL FILL_1__10697_ (
);

FILL FILL_1__10277_ (
);

FILL FILL_2_BUFX2_insert341 (
);

FILL FILL_2_BUFX2_insert342 (
);

FILL FILL_2_BUFX2_insert343 (
);

FILL FILL_2_BUFX2_insert344 (
);

FILL FILL_4__11611_ (
);

FILL FILL_2_BUFX2_insert345 (
);

FILL FILL_5__15090_ (
);

FILL FILL_2_BUFX2_insert346 (
);

FILL FILL_2_BUFX2_insert347 (
);

OAI21X1 _9390_ (
    .A(_1273_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1274_),
    .Y(_1238_[18])
);

FILL FILL_2_BUFX2_insert348 (
);

FILL FILL_2_BUFX2_insert349 (
);

FILL FILL_6__13889_ (
);

FILL FILL_6__13469_ (
);

FILL FILL_4__14083_ (
);

FILL FILL_0__15916_ (
);

FILL FILL_2__8243_ (
);

FILL FILL_3__13496_ (
);

FILL FILL_0__10631_ (
);

FILL FILL_6__14830_ (
);

FILL FILL_4__8589_ (
);

FILL FILL_2__12489_ (
);

FILL FILL_2__12069_ (
);

FILL FILL_5__13823_ (
);

FILL FILL_5__13403_ (
);

FILL FILL_2_BUFX2_insert1060 (
);

FILL FILL_2_BUFX2_insert1061 (
);

INVX1 _7703_ (
    .A(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_414_)
);

FILL FILL_2_BUFX2_insert1062 (
);

FILL FILL_2_BUFX2_insert1063 (
);

FILL FILL_2_BUFX2_insert1064 (
);

FILL FILL_4__9530_ (
);

FILL FILL_2_BUFX2_insert1065 (
);

FILL FILL_2_BUFX2_insert1066 (
);

FILL FILL_4__9110_ (
);

FILL FILL_2__13850_ (
);

FILL FILL_2_BUFX2_insert1067 (
);

FILL FILL_2__13430_ (
);

FILL FILL_2_BUFX2_insert1068 (
);

FILL FILL_5__16295_ (
);

FILL FILL_2__13010_ (
);

FILL FILL_0__8489_ (
);

FILL FILL_2_BUFX2_insert1069 (
);

FILL FILL_0__8069_ (
);

FILL FILL_3__11809_ (
);

FILL FILL_1__12843_ (
);

FILL FILL_1__12423_ (
);

FILL FILL_4__15288_ (
);

FILL FILL_1__12003_ (
);

FILL SFILL104840x53050 (
);

FILL FILL_2__9868_ (
);

FILL FILL_0__9850_ (
);

FILL FILL_0__11836_ (
);

FILL FILL_2__9028_ (
);

FILL FILL_0__11416_ (
);

FILL FILL_0__9010_ (
);

INVX1 _11701_ (
    .A(_2172_),
    .Y(_2800_)
);

FILL FILL_5__7873_ (
);

FILL FILL_5__7453_ (
);

FILL FILL_5__7033_ (
);

FILL FILL_6__10750_ (
);

OAI22X1 _14593_ (
    .A(_5081_),
    .B(_3982__bF$buf3),
    .C(_3983__bF$buf0),
    .D(_5080_),
    .Y(_5082_)
);

INVX1 _14173_ (
    .A(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_4670_)
);

FILL FILL_5__14608_ (
);

FILL FILL_3__15642_ (
);

OAI21X1 _8908_ (
    .A(_1033_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .C(_1034_),
    .Y(_978_[28])
);

FILL FILL_3__15222_ (
);

FILL FILL_1__7865_ (
);

FILL FILL_1__7445_ (
);

FILL FILL_2__14635_ (
);

FILL FILL_2__14215_ (
);

FILL SFILL19160x68050 (
);

FILL FILL_1__13628_ (
);

FILL FILL_1__13208_ (
);

FILL FILL_1_BUFX2_insert360 (
);

FILL FILL_3__8732_ (
);

FILL FILL_1_BUFX2_insert361 (
);

FILL FILL_3__8312_ (
);

OAI21X1 _12906_ (
    .A(_3608_),
    .B(vdd),
    .C(_3609_),
    .Y(_3555_[27])
);

FILL FILL_1_BUFX2_insert362 (
);

FILL FILL_1_BUFX2_insert363 (
);

FILL SFILL83400x54050 (
);

FILL FILL_1_BUFX2_insert364 (
);

FILL FILL_1_BUFX2_insert365 (
);

FILL FILL_1_BUFX2_insert366 (
);

FILL FILL_5__8658_ (
);

FILL FILL_5__8238_ (
);

FILL FILL_1_BUFX2_insert367 (
);

FILL FILL_1_BUFX2_insert368 (
);

FILL FILL_1_BUFX2_insert369 (
);

OAI22X1 _15798_ (
    .A(_6258_),
    .B(_5545__bF$buf1),
    .C(_5466__bF$buf2),
    .D(_6259_),
    .Y(_6260_)
);

NOR2X1 _15378_ (
    .A(_5849_),
    .B(_5535__bF$buf2),
    .Y(_5850_)
);

FILL FILL_3__16007_ (
);

FILL FILL_5__10948_ (
);

DFFSR _10093_ (
    .Q(\datapath_1.regfile_1.regOut[25] [23]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_1563_[23])
);

FILL FILL_5__10528_ (
);

FILL FILL_3__11982_ (
);

FILL FILL_3__11562_ (
);

FILL FILL_5__10108_ (
);

FILL FILL_3__11142_ (
);

FILL SFILL108680x54050 (
);

FILL FILL_0__16034_ (
);

FILL FILL_2__10975_ (
);

FILL FILL_2__10555_ (
);

FILL FILL_2__10135_ (
);

FILL FILL_3__9937_ (
);

FILL FILL_3__9517_ (
);

FILL FILL_5__14781_ (
);

FILL FILL_0__6975_ (
);

FILL FILL_5__14361_ (
);

FILL FILL_6__7942_ (
);

FILL FILL112440x52050 (
);

OAI21X1 _8661_ (
    .A(_909_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_910_),
    .Y(_848_[31])
);

OAI21X1 _8241_ (
    .A(_690_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .C(_691_),
    .Y(_653_[19])
);

FILL FILL_4__13774_ (
);

FILL FILL_4__13354_ (
);

INVX1 _11298_ (
    .A(_2416_),
    .Y(_2417_)
);

FILL FILL_2__7934_ (
);

FILL FILL_3__12767_ (
);

FILL FILL_3__12347_ (
);

FILL FILL_1__13381_ (
);

FILL FILL_0__12374_ (
);

FILL FILL_5__15986_ (
);

FILL FILL_2__12701_ (
);

FILL FILL_5__15566_ (
);

FILL FILL_5__15146_ (
);

OAI21X1 _9866_ (
    .A(_1509_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .C(_1510_),
    .Y(_1498_[6])
);

FILL FILL_3__16180_ (
);

DFFSR _9446_ (
    .Q(\datapath_1.regfile_1.regOut[20] [16]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_1238_[16])
);

NAND2X1 _9026_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1093_)
);

FILL FILL_5__10281_ (
);

FILL FILL_4__14979_ (
);

FILL FILL_4__14559_ (
);

FILL FILL_4__14139_ (
);

FILL FILL_2__15593_ (
);

FILL FILL_2__15173_ (
);

FILL FILL_2__8719_ (
);

FILL FILL_0__8701_ (
);

FILL FILL_1__14586_ (
);

FILL FILL_1__14166_ (
);

FILL FILL_4__15920_ (
);

FILL FILL_4__15500_ (
);

FILL FILL_0__13999_ (
);

AOI22X1 _13864_ (
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .B(_4154_),
    .C(_4051__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_4368_)
);

FILL FILL_3__9270_ (
);

FILL FILL_0__13579_ (
);

FILL FILL_0__13159_ (
);

OAI22X1 _13444_ (
    .A(_3952_),
    .B(_3955__bF$buf1),
    .C(_3954__bF$buf4),
    .D(_3953_),
    .Y(_3956_)
);

NAND2X1 _13024_ (
    .A(vdd),
    .B(\datapath_1.rd2 [24]),
    .Y(_3668_)
);

FILL FILL_3__14913_ (
);

FILL FILL_2__13906_ (
);

FILL FILL_0__14940_ (
);

FILL FILL_0__14520_ (
);

FILL FILL_0__14100_ (
);

FILL FILL_5__11486_ (
);

FILL FILL_5__11066_ (
);

FILL FILL_2__16378_ (
);

FILL FILL_4__10899_ (
);

FILL FILL_4__7193_ (
);

FILL FILL_4__10059_ (
);

FILL FILL_0__9906_ (
);

FILL FILL_2__11093_ (
);

FILL FILL_5__7929_ (
);

FILL FILL_5__7509_ (
);

FILL FILL_6__10806_ (
);

FILL FILL_4__11840_ (
);

INVX1 _14649_ (
    .A(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_5136_)
);

INVX1 _14229_ (
    .A(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_4725_)
);

FILL FILL_4__11420_ (
);

FILL FILL_4__11000_ (
);

FILL FILL_0__7093_ (
);

FILL FILL_6__8480_ (
);

FILL SFILL98920x77050 (
);

FILL FILL_1__16312_ (
);

FILL FILL_3__10833_ (
);

FILL FILL_3__10413_ (
);

FILL FILL_0__15725_ (
);

FILL FILL_0__15305_ (
);

FILL FILL_2__8892_ (
);

FILL FILL_2__8472_ (
);

FILL FILL_0__10440_ (
);

FILL FILL_0__10020_ (
);

FILL SFILL23640x75050 (
);

FILL FILL_4__8398_ (
);

FILL FILL_2__12298_ (
);

FILL FILL_5__13632_ (
);

FILL FILL_5__13212_ (
);

INVX1 _7932_ (
    .A(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_526_)
);

FILL SFILL8680x74050 (
);

DFFSR _7512_ (
    .Q(\datapath_1.regfile_1.regOut[5] [2]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_263_[2])
);

FILL FILL_4__12625_ (
);

FILL FILL_4__12205_ (
);

NAND2X1 _10989_ (
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2108_)
);

FILL FILL_6__9265_ (
);

OAI21X1 _10569_ (
    .A(_1876_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .C(_1877_),
    .Y(_1823_[27])
);

OAI21X1 _10149_ (
    .A(_1657_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1658_),
    .Y(_1628_[15])
);

FILL FILL_3__11618_ (
);

FILL FILL_1__12652_ (
);

FILL FILL_4__15097_ (
);

FILL FILL_1__12232_ (
);

FILL SFILL84280x55050 (
);

FILL FILL_2__9677_ (
);

NAND2X1 _11930_ (
    .A(IorD_bF$buf4),
    .B(ALUOut[14]),
    .Y(_2995_)
);

FILL FILL_2__9257_ (
);

FILL FILL_0__11645_ (
);

FILL FILL_0__11225_ (
);

OAI21X1 _11510_ (
    .A(_2611_),
    .B(_2344__bF$buf2),
    .C(_2621_),
    .Y(_2622_)
);

FILL FILL_5__7682_ (
);

FILL FILL_6__15424_ (
);

FILL FILL_6__15004_ (
);

FILL SFILL23640x30050 (
);

FILL FILL_5__14837_ (
);

FILL FILL_5__14417_ (
);

FILL FILL_3__15871_ (
);

FILL FILL_3__15451_ (
);

OAI21X1 _8717_ (
    .A(_926_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_927_),
    .Y(_913_[7])
);

FILL FILL_3__15031_ (
);

FILL FILL_1__7674_ (
);

FILL FILL_2__14864_ (
);

FILL FILL_2__14444_ (
);

FILL FILL_2__14024_ (
);

FILL SFILL94360x50 (
);

FILL FILL_1__13857_ (
);

FILL FILL_1__13437_ (
);

FILL FILL_1__13017_ (
);

FILL SFILL88920x75050 (
);

FILL SFILL84200x53050 (
);

FILL FILL_3__8961_ (
);

OAI21X1 _12715_ (
    .A(_3501_),
    .B(IRWrite_bF$buf6),
    .C(_3502_),
    .Y(_3490_[6])
);

FILL FILL_3__8121_ (
);

FILL FILL_5__8887_ (
);

FILL FILL_5__8467_ (
);

FILL FILL_1_BUFX2_insert30 (
);

FILL FILL_1_BUFX2_insert31 (
);

FILL FILL_1_BUFX2_insert32 (
);

FILL FILL_1_BUFX2_insert33 (
);

FILL FILL_6__11344_ (
);

FILL SFILL13640x73050 (
);

FILL FILL_1_BUFX2_insert34 (
);

NOR3X1 _15187_ (
    .A(_5515__bF$buf1),
    .B(_5663_),
    .C(_5521__bF$buf0),
    .Y(_5664_)
);

FILL FILL_1_BUFX2_insert35 (
);

FILL FILL_1_BUFX2_insert36 (
);

FILL SFILL69000x33050 (
);

FILL FILL_3__16236_ (
);

FILL FILL_1_BUFX2_insert37 (
);

FILL FILL_1_BUFX2_insert38 (
);

FILL FILL_1__8879_ (
);

FILL FILL_1_BUFX2_insert39 (
);

FILL FILL_5__10757_ (
);

FILL FILL_1__8459_ (
);

FILL FILL_3__11791_ (
);

FILL FILL_3__11371_ (
);

FILL FILL_2__15649_ (
);

FILL FILL_2__15229_ (
);

FILL FILL_4__6884_ (
);

FILL FILL_0__16263_ (
);

FILL FILL_2__10784_ (
);

FILL SFILL114440x36050 (
);

FILL FILL_2__10364_ (
);

FILL FILL_1__9400_ (
);

FILL SFILL109640x1050 (
);

FILL FILL_3__9746_ (
);

FILL FILL_5__14590_ (
);

FILL FILL_5__14170_ (
);

FILL SFILL74280x53050 (
);

OAI21X1 _8890_ (
    .A(_1021_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .C(_1022_),
    .Y(_978_[22])
);

FILL FILL_6__7751_ (
);

OAI21X1 _8470_ (
    .A(_802_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_803_),
    .Y(_783_[10])
);

DFFSR _8050_ (
    .Q(\datapath_1.regfile_1.regOut[9] [28]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_523_[28])
);

FILL FILL_4__13583_ (
);

FILL FILL_4__13163_ (
);

FILL FILL_2__7743_ (
);

FILL FILL_3__12996_ (
);

FILL FILL_3__12576_ (
);

FILL FILL_2__7323_ (
);

FILL FILL_3__12156_ (
);

FILL FILL_4__7249_ (
);

FILL FILL_2__11989_ (
);

FILL FILL_2__11569_ (
);

FILL FILL_2__11149_ (
);

FILL FILL_0__12183_ (
);

FILL FILL_5__12903_ (
);

FILL FILL_4__8610_ (
);

FILL FILL_5__15795_ (
);

FILL FILL_0__7989_ (
);

FILL FILL_5__15375_ (
);

FILL FILL_2__12510_ (
);

FILL SFILL74200x51050 (
);

FILL FILL_0__7569_ (
);

FILL FILL_6__8956_ (
);

NAND2X1 _9675_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1424_)
);

NAND2X1 _9255_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1205_)
);

FILL FILL_1__11923_ (
);

FILL FILL_4__14788_ (
);

FILL FILL_4__14368_ (
);

FILL FILL_1__11503_ (
);

FILL FILL_0__10916_ (
);

FILL FILL_0__8510_ (
);

FILL FILL_2__8528_ (
);

FILL FILL_2__8108_ (
);

FILL FILL_1__14395_ (
);

FILL FILL_5__6953_ (
);

FILL SFILL54040x50 (
);

NOR2X1 _13673_ (
    .A(_4177_),
    .B(_4180_),
    .Y(_4181_)
);

FILL FILL_0__13388_ (
);

NAND2X1 _13253_ (
    .A(_3788_),
    .B(_3795_),
    .Y(_3796_)
);

FILL FILL_3__14722_ (
);

FILL FILL_3__14302_ (
);

FILL FILL_1__6945_ (
);

FILL FILL_2__13715_ (
);

FILL FILL_5__11295_ (
);

FILL FILL112120x71050 (
);

FILL FILL_1__12708_ (
);

FILL FILL_2__16187_ (
);

FILL FILL_4__10288_ (
);

FILL FILL_3__7812_ (
);

FILL FILL_5__7738_ (
);

FILL FILL_5__7318_ (
);

FILL FILL_2_BUFX2_insert720 (
);

FILL FILL_2_BUFX2_insert721 (
);

FILL FILL_2_BUFX2_insert722 (
);

AOI22X1 _14878_ (
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .B(_4001__bF$buf0),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_5361_)
);

FILL FILL_2_BUFX2_insert723 (
);

AOI22X1 _14458_ (
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .B(_4102_),
    .C(_3942__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_4949_)
);

FILL FILL_2_BUFX2_insert724 (
);

AOI22X1 _14038_ (
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .B(_3885_),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_4538_)
);

FILL FILL_2_BUFX2_insert725 (
);

FILL FILL_2_BUFX2_insert726 (
);

FILL FILL_3__15927_ (
);

FILL FILL_2_BUFX2_insert727 (
);

FILL FILL_3__15507_ (
);

FILL FILL_2_BUFX2_insert728 (
);

FILL FILL112040x78050 (
);

FILL FILL_1__16121_ (
);

FILL FILL_2_BUFX2_insert729 (
);

FILL FILL_3__10642_ (
);

FILL FILL_0__15954_ (
);

FILL FILL_0__15534_ (
);

FILL FILL_0__15114_ (
);

FILL FILL_5__13861_ (
);

FILL FILL_5__13441_ (
);

FILL FILL112440x47050 (
);

FILL FILL_5__13021_ (
);

OAI21X1 _7741_ (
    .A(_438_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_439_),
    .Y(_393_[23])
);

OAI21X1 _7321_ (
    .A(_219_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_220_),
    .Y(_198_[11])
);

FILL FILL_4__12854_ (
);

FILL FILL_4__12434_ (
);

FILL FILL_4__12014_ (
);

OAI21X1 _10798_ (
    .A(_1988_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1989_),
    .Y(_1953_[18])
);

OAI21X1 _10378_ (
    .A(_1769_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1770_),
    .Y(_1758_[6])
);

FILL SFILL33720x65050 (
);

FILL FILL_3__11847_ (
);

FILL FILL_1__12881_ (
);

FILL FILL_3__11427_ (
);

FILL FILL_1__12461_ (
);

FILL FILL_3__11007_ (
);

FILL FILL_1__12041_ (
);

FILL FILL112040x33050 (
);

FILL FILL_0__16319_ (
);

FILL FILL_2__9486_ (
);

FILL FILL_0__11874_ (
);

FILL FILL_0__11454_ (
);

FILL FILL_0__11034_ (
);

FILL FILL_5__7491_ (
);

FILL FILL_5__7071_ (
);

FILL FILL_5__14646_ (
);

FILL FILL_3__15680_ (
);

FILL FILL_5__14226_ (
);

DFFSR _8946_ (
    .Q(\datapath_1.regfile_1.regOut[16] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_978_[28])
);

FILL FILL_3__15260_ (
);

NAND2X1 _8526_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_841_)
);

NAND2X1 _8106_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_622_)
);

FILL FILL_1__7483_ (
);

FILL FILL_1__7063_ (
);

FILL FILL_4__13639_ (
);

FILL FILL_4__13219_ (
);

FILL FILL_2__14673_ (
);

FILL FILL_2__14253_ (
);

FILL FILL_1__13666_ (
);

FILL FILL_1__13246_ (
);

FILL FILL_1_BUFX2_insert740 (
);

FILL FILL_1_BUFX2_insert741 (
);

FILL FILL_3__8770_ (
);

FILL FILL_0__12659_ (
);

FILL FILL_1_BUFX2_insert742 (
);

DFFSR _12944_ (
    .Q(\datapath_1.a [25]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_3555_[25])
);

FILL FILL_3__8350_ (
);

NAND2X1 _12524_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [28]),
    .Y(_3416_)
);

FILL FILL_1_BUFX2_insert743 (
);

FILL FILL_0__12239_ (
);

NAND3X1 _12104_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [29]),
    .C(_3034__bF$buf0),
    .Y(_3124_)
);

FILL FILL_1_BUFX2_insert744 (
);

FILL FILL_1_BUFX2_insert745 (
);

FILL FILL_1_BUFX2_insert746 (
);

FILL FILL_5__8696_ (
);

FILL FILL_5__8276_ (
);

FILL FILL_1_BUFX2_insert747 (
);

FILL FILL_1_BUFX2_insert748 (
);

FILL FILL_1_BUFX2_insert749 (
);

FILL FILL_6__11993_ (
);

FILL FILL_0__13600_ (
);

FILL FILL_3__16045_ (
);

FILL FILL_5__10566_ (
);

FILL FILL_1__8268_ (
);

FILL FILL_5__10146_ (
);

FILL FILL_3__11180_ (
);

FILL FILL_2__15878_ (
);

FILL FILL_2__15458_ (
);

FILL FILL_2__15038_ (
);

FILL FILL_0__16072_ (
);

FILL FILL_2__10173_ (
);

FILL SFILL58840x76050 (
);

FILL FILL_3__9975_ (
);

FILL FILL_3__9555_ (
);

FILL FILL_4__10920_ (
);

FILL FILL_3__9135_ (
);

INVX1 _13729_ (
    .A(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_4236_)
);

NOR2X1 _13309_ (
    .A(_3781_),
    .B(_3842_),
    .Y(\datapath_1.regfile_1.regEn [10])
);

FILL FILL_4__10500_ (
);

FILL FILL_6__7560_ (
);

FILL FILL_1__15812_ (
);

FILL FILL_4__13392_ (
);

FILL FILL_0__14805_ (
);

FILL FILL_2__7972_ (
);

FILL FILL_2__7552_ (
);

BUFX2 BUFX2_insert410 (
    .A(_3995_),
    .Y(_3995__bF$buf4)
);

FILL FILL_3__12385_ (
);

BUFX2 BUFX2_insert411 (
    .A(_3995_),
    .Y(_3995__bF$buf3)
);

BUFX2 BUFX2_insert412 (
    .A(_3995_),
    .Y(_3995__bF$buf2)
);

BUFX2 BUFX2_insert413 (
    .A(_3995_),
    .Y(_3995__bF$buf1)
);

BUFX2 BUFX2_insert414 (
    .A(_3995_),
    .Y(_3995__bF$buf0)
);

FILL FILL_4__7478_ (
);

BUFX2 BUFX2_insert415 (
    .A(_5530_),
    .Y(_5530__bF$buf3)
);

BUFX2 BUFX2_insert416 (
    .A(_5530_),
    .Y(_5530__bF$buf2)
);

FILL FILL_4__7058_ (
);

BUFX2 BUFX2_insert417 (
    .A(_5530_),
    .Y(_5530__bF$buf1)
);

FILL FILL_2__11798_ (
);

BUFX2 BUFX2_insert418 (
    .A(_5530_),
    .Y(_5530__bF$buf0)
);

FILL FILL_2__11378_ (
);

BUFX2 BUFX2_insert419 (
    .A(_5471_),
    .Y(_5471__bF$buf5)
);

FILL FILL_5__12712_ (
);

FILL SFILL8680x69050 (
);

FILL FILL_6__16191_ (
);

FILL FILL_4__11705_ (
);

FILL FILL_5__15184_ (
);

FILL FILL_0__7798_ (
);

FILL FILL_0__7378_ (
);

NAND2X1 _9484_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1317_)
);

FILL FILL_6__8345_ (
);

DFFSR _9064_ (
    .Q(\datapath_1.regfile_1.regOut[17] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_1043_[18])
);

FILL FILL_4__14597_ (
);

FILL FILL_1__11732_ (
);

FILL FILL_4__14177_ (
);

FILL FILL_1__11312_ (
);

FILL FILL_2__8757_ (
);

FILL FILL_2__8337_ (
);

FILL FILL_0__10305_ (
);

OAI22X1 _13482_ (
    .A(_3991_),
    .B(_3936__bF$buf4),
    .C(_3935__bF$buf2),
    .D(_3992_),
    .Y(_3993_)
);

DFFSR _13062_ (
    .Q(_2_[15]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3620_[15])
);

FILL FILL_5__13917_ (
);

FILL FILL_3__14951_ (
);

FILL SFILL8600x67050 (
);

FILL FILL_3__14531_ (
);

FILL FILL_3__14111_ (
);

FILL FILL_4_BUFX2_insert250 (
);

FILL FILL_4__9624_ (
);

FILL FILL_4_BUFX2_insert251 (
);

FILL FILL_4_BUFX2_insert252 (
);

FILL SFILL8680x24050 (
);

FILL FILL_4_BUFX2_insert253 (
);

FILL FILL_2__13944_ (
);

FILL SFILL13720x61050 (
);

FILL FILL_4_BUFX2_insert254 (
);

FILL FILL_5__16389_ (
);

FILL FILL_2__13524_ (
);

FILL FILL_2__13104_ (
);

FILL FILL_4_BUFX2_insert255 (
);

FILL FILL_4_BUFX2_insert256 (
);

FILL FILL_4_BUFX2_insert257 (
);

FILL FILL_4_BUFX2_insert258 (
);

FILL FILL_4_BUFX2_insert259 (
);

FILL FILL_1__12517_ (
);

FILL SFILL84200x48050 (
);

FILL FILL_3__7621_ (
);

FILL FILL_0__9524_ (
);

FILL FILL_0__9104_ (
);

FILL FILL_3__7201_ (
);

FILL FILL_5__7967_ (
);

FILL FILL_5__7547_ (
);

FILL FILL_4__16323_ (
);

FILL FILL_6__10424_ (
);

NOR2X1 _14687_ (
    .A(_5170_),
    .B(_5173_),
    .Y(_5174_)
);

INVX1 _14267_ (
    .A(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_4762_)
);

FILL FILL_3__15736_ (
);

FILL SFILL109480x48050 (
);

FILL FILL_3__15316_ (
);

FILL FILL_1__16350_ (
);

FILL FILL_1__7959_ (
);

FILL FILL_3__10871_ (
);

FILL FILL_1__7119_ (
);

FILL FILL_3__10451_ (
);

FILL SFILL8600x22050 (
);

FILL FILL_3__10031_ (
);

FILL FILL_2__14729_ (
);

FILL FILL_0__15763_ (
);

FILL FILL_2__14309_ (
);

FILL FILL_0__15343_ (
);

FILL FILL_2__8090_ (
);

FILL FILL_1__8900_ (
);

FILL FILL_3__8826_ (
);

FILL FILL_5__13670_ (
);

FILL FILL_5__13250_ (
);

OAI21X1 _7970_ (
    .A(_550_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_551_),
    .Y(_523_[14])
);

OAI21X1 _7550_ (
    .A(_331_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .C(_332_),
    .Y(_328_[2])
);

DFFSR _7130_ (
    .Q(\datapath_1.regfile_1.regOut[2] [4]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_68_[4])
);

FILL FILL_4__12243_ (
);

FILL SFILL13640x23050 (
);

NAND2X1 _10187_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1684_)
);

FILL FILL_3__11656_ (
);

FILL FILL_3__11236_ (
);

FILL FILL_1__12270_ (
);

FILL FILL_0__16128_ (
);

OAI21X1 _16413_ (
    .A(_6828_),
    .B(gnd),
    .C(_6829_),
    .Y(_6769_[30])
);

FILL FILL_2__10649_ (
);

FILL SFILL38840x72050 (
);

FILL FILL_2__9295_ (
);

FILL FILL_0__11683_ (
);

FILL FILL_0__11263_ (
);

FILL FILL_3_BUFX2_insert270 (
);

FILL FILL_3_BUFX2_insert271 (
);

FILL FILL_5__14875_ (
);

FILL FILL_3_BUFX2_insert272 (
);

FILL SFILL74200x46050 (
);

FILL FILL_3_BUFX2_insert273 (
);

FILL FILL_5__14455_ (
);

FILL FILL_3_BUFX2_insert274 (
);

FILL FILL_5__14035_ (
);

FILL FILL_6__7616_ (
);

FILL FILL_3_BUFX2_insert275 (
);

NAND2X1 _8755_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_953_)
);

NAND2X1 _8335_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_734_)
);

FILL FILL_3_BUFX2_insert276 (
);

FILL FILL_3_BUFX2_insert277 (
);

FILL FILL_3_BUFX2_insert278 (
);

FILL FILL_1__7292_ (
);

FILL FILL_4__13868_ (
);

FILL FILL_3_BUFX2_insert279 (
);

FILL FILL_4__13448_ (
);

FILL FILL_2__14482_ (
);

FILL FILL_4__13028_ (
);

FILL FILL_2__14062_ (
);

FILL FILL_2__7608_ (
);

FILL FILL_1__13895_ (
);

FILL FILL_1__13475_ (
);

FILL SFILL44040x1050 (
);

FILL SFILL43720x4050 (
);

FILL FILL_0__12888_ (
);

NAND2X1 _12753_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[19]),
    .Y(_3528_)
);

FILL FILL_0__12468_ (
);

FILL SFILL3480x71050 (
);

FILL FILL_0__12048_ (
);

AOI22X1 _12333_ (
    .A(_2_[29]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3289_)
);

FILL FILL_3__13802_ (
);

FILL FILL_6__16247_ (
);

FILL FILL_5__8085_ (
);

FILL FILL_3__16274_ (
);

FILL FILL_5__10795_ (
);

FILL FILL112120x66050 (
);

FILL FILL_1__8497_ (
);

FILL FILL_5__10375_ (
);

FILL FILL_1__8077_ (
);

FILL FILL_2__15687_ (
);

FILL FILL_2__15267_ (
);

FILL FILL_3__9784_ (
);

FILL FILL_3__9364_ (
);

INVX1 _13958_ (
    .A(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_4460_)
);

INVX1 _13538_ (
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_4048_)
);

INVX1 _13118_ (
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_3710_)
);

FILL FILL_1__15621_ (
);

FILL SFILL28840x70050 (
);

FILL FILL_1__15201_ (
);

FILL FILL_6__12167_ (
);

FILL FILL_0__14614_ (
);

FILL FILL_2__7361_ (
);

FILL SFILL64200x44050 (
);

FILL FILL_3__12194_ (
);

FILL SFILL85160x42050 (
);

FILL FILL112120x21050 (
);

FILL FILL_4__7287_ (
);

FILL FILL_2__11187_ (
);

FILL FILL_5__12521_ (
);

FILL FILL_5__12101_ (
);

FILL FILL_4__11934_ (
);

FILL FILL_4__11514_ (
);

FILL FILL_2_BUFX2_insert80 (
);

FILL FILL_0__7187_ (
);

INVX1 _9293_ (
    .A(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_1230_)
);

FILL FILL_1__16406_ (
);

FILL FILL_2_BUFX2_insert81 (
);

FILL FILL_2_BUFX2_insert82 (
);

FILL FILL_3__10927_ (
);

FILL FILL_2_BUFX2_insert83 (
);

FILL FILL_3__10507_ (
);

FILL FILL_1__11961_ (
);

FILL FILL_2_BUFX2_insert84 (
);

FILL FILL_2_BUFX2_insert85 (
);

FILL FILL_1__11541_ (
);

FILL FILL112040x28050 (
);

FILL FILL_2_BUFX2_insert86 (
);

FILL FILL_1__11121_ (
);

FILL FILL_2_BUFX2_insert87 (
);

FILL FILL_0__15819_ (
);

FILL FILL_2_BUFX2_insert88 (
);

FILL FILL_2_BUFX2_insert89 (
);

FILL FILL_2__8986_ (
);

FILL FILL_0__10954_ (
);

FILL FILL_2__8566_ (
);

FILL FILL_0__10534_ (
);

FILL FILL_3__13399_ (
);

FILL FILL_2__8146_ (
);

FILL FILL_0__10114_ (
);

FILL FILL_5__6991_ (
);

FILL FILL_6__14733_ (
);

NAND2X1 _13291_ (
    .A(_3821_),
    .B(_3828_),
    .Y(_3829_)
);

FILL FILL_5__13726_ (
);

FILL FILL_5__13306_ (
);

FILL FILL_3__14760_ (
);

FILL FILL_3__14340_ (
);

NAND2X1 _7606_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_370_)
);

FILL FILL_1__6983_ (
);

FILL FILL_4__9853_ (
);

FILL FILL_4__12719_ (
);

FILL FILL_4__9013_ (
);

FILL FILL_2__13753_ (
);

FILL FILL_2__13333_ (
);

FILL FILL_5__16198_ (
);

FILL FILL_6__9359_ (
);

FILL FILL_1__12746_ (
);

FILL FILL_1__12326_ (
);

FILL SFILL33720x15050 (
);

FILL FILL_0__9753_ (
);

FILL FILL_3__7850_ (
);

FILL FILL_3__7430_ (
);

FILL FILL_0__11739_ (
);

FILL FILL_0__11319_ (
);

AOI21X1 _11604_ (
    .A(_2263_),
    .B(_2708_),
    .C(_2709_),
    .Y(_2710_)
);

FILL FILL_5__7356_ (
);

FILL FILL_4__16132_ (
);

FILL SFILL54200x42050 (
);

OAI22X1 _14496_ (
    .A(_3967__bF$buf0),
    .B(_4985_),
    .C(_4986_),
    .D(_3972__bF$buf1),
    .Y(_4987_)
);

FILL FILL_6__10233_ (
);

AOI22X1 _14076_ (
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .B(_4005__bF$buf0),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_4575_)
);

FILL FILL_3__15965_ (
);

FILL FILL_3__15545_ (
);

FILL FILL_3__15125_ (
);

FILL SFILL39000x7050 (
);

FILL SFILL13720x3050 (
);

FILL FILL_3__10680_ (
);

FILL FILL_1__7348_ (
);

FILL FILL_3__10260_ (
);

FILL FILL_2__14958_ (
);

FILL FILL_0__15992_ (
);

FILL FILL_2__14538_ (
);

FILL FILL_0__15572_ (
);

FILL FILL_2__14118_ (
);

FILL SFILL13640x8050 (
);

FILL FILL_0__15152_ (
);

FILL FILL_3__8635_ (
);

DFFSR _12809_ (
    .Q(\datapath_1.PCJump [20]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3490_[18])
);

FILL FILL_3__8215_ (
);

FILL FILL_4__12892_ (
);

FILL FILL_4__12472_ (
);

FILL FILL_4__12052_ (
);

FILL FILL_3__11885_ (
);

FILL FILL_5__9922_ (
);

FILL FILL_3__11465_ (
);

FILL FILL_5__9502_ (
);

FILL FILL_3__11045_ (
);

FILL FILL_4__6978_ (
);

FILL FILL_0__16357_ (
);

INVX1 _16222_ (
    .A(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_6673_)
);

FILL FILL_2__10878_ (
);

FILL FILL_2__10038_ (
);

FILL FILL_0__11492_ (
);

FILL FILL_0__11072_ (
);

FILL FILL_1__9914_ (
);

FILL FILL_5__14684_ (
);

FILL FILL_5__14264_ (
);

FILL FILL_0__6878_ (
);

NAND2X1 _8984_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1065_)
);

DFFSR _8564_ (
    .Q(\datapath_1.regfile_1.regOut[13] [30]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_783_[30])
);

INVX1 _8144_ (
    .A(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_647_)
);

FILL FILL_1__10812_ (
);

FILL FILL_4__13677_ (
);

FILL FILL_4__13257_ (
);

FILL SFILL48920x62050 (
);

FILL FILL_2__14291_ (
);

FILL FILL_2__7837_ (
);

FILL FILL_2__7417_ (
);

FILL FILL_1__13284_ (
);

FILL FILL_0__12697_ (
);

NAND2X1 _12982_ (
    .A(vdd),
    .B(\datapath_1.rd2 [10]),
    .Y(_3640_)
);

DFFSR _12562_ (
    .Q(ALUOut[27]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3360_[27])
);

FILL FILL_0__12277_ (
);

INVX1 _12142_ (
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_3148_)
);

FILL FILL_3__13611_ (
);

FILL FILL_4__8704_ (
);

FILL SFILL8680x19050 (
);

FILL SFILL13720x56050 (
);

FILL FILL_5__15889_ (
);

FILL FILL_2__12604_ (
);

FILL FILL_5__15469_ (
);

FILL FILL_5__15049_ (
);

INVX1 _9769_ (
    .A(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_1466_)
);

FILL FILL_3__16083_ (
);

INVX1 _9349_ (
    .A(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_1247_)
);

FILL FILL_5__10184_ (
);

FILL FILL_2__15496_ (
);

FILL FILL_2__15076_ (
);

FILL FILL_5__16410_ (
);

FILL FILL_0__8604_ (
);

FILL FILL_1__14489_ (
);

FILL FILL_1__14069_ (
);

FILL FILL_4__15823_ (
);

FILL FILL_4__15403_ (
);

FILL FILL_3__9593_ (
);

INVX1 _13767_ (
    .A(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_4273_)
);

FILL FILL_3__9173_ (
);

AOI21X1 _13347_ (
    .A(\datapath_1.a3 [3]),
    .B(_3865_),
    .C(_3750_),
    .Y(_3866_)
);

FILL FILL_3__14816_ (
);

FILL FILL_1__15850_ (
);

FILL FILL_5__9099_ (
);

FILL FILL_1__15430_ (
);

FILL FILL_1__15010_ (
);

FILL FILL_4__9909_ (
);

FILL SFILL8600x17050 (
);

FILL FILL_2__13809_ (
);

FILL FILL_0__14843_ (
);

FILL FILL_0__14423_ (
);

FILL FILL_0__14003_ (
);

FILL SFILL48840x24050 (
);

FILL SFILL13720x11050 (
);

FILL FILL_2__7590_ (
);

FILL FILL_5__11389_ (
);

FILL FILL_2__7170_ (
);

FILL FILL_4__7096_ (
);

FILL FILL_0__9809_ (
);

FILL SFILL38920x60050 (
);

FILL FILL_5__12750_ (
);

FILL FILL_5__12330_ (
);

FILL FILL_4__11743_ (
);

FILL FILL_4__11323_ (
);

FILL SFILL13640x18050 (
);

FILL FILL_1__16215_ (
);

FILL FILL_3__10316_ (
);

FILL FILL_1__11770_ (
);

FILL FILL_1__11350_ (
);

AOI21X1 _15913_ (
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .B(_5567_),
    .C(_6371_),
    .Y(_6372_)
);

FILL FILL_0__15628_ (
);

FILL FILL_0__15208_ (
);

FILL FILL_2__8375_ (
);

FILL FILL_0__10763_ (
);

FILL FILL_5__13955_ (
);

FILL FILL_5__13535_ (
);

FILL FILL_5__13115_ (
);

NAND2X1 _7835_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_482_)
);

NAND2X1 _7415_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .Y(_327_)
);

FILL FILL_4_BUFX2_insert630 (
);

FILL FILL_4__9662_ (
);

FILL FILL_4_BUFX2_insert631 (
);

FILL FILL_4_BUFX2_insert632 (
);

FILL FILL_4__9242_ (
);

FILL FILL_4_BUFX2_insert633 (
);

FILL FILL_4__12528_ (
);

FILL FILL_2__13982_ (
);

FILL FILL_4_BUFX2_insert634 (
);

FILL FILL_4__12108_ (
);

FILL FILL_2__13562_ (
);

FILL FILL_4_BUFX2_insert635 (
);

FILL FILL_2__13142_ (
);

FILL FILL_4_BUFX2_insert636 (
);

FILL FILL_4_BUFX2_insert637 (
);

FILL FILL_4_BUFX2_insert638 (
);

FILL FILL_4_BUFX2_insert639 (
);

FILL FILL112200x54050 (
);

FILL FILL_1__12975_ (
);

FILL FILL_1__12135_ (
);

FILL FILL_0__9982_ (
);

FILL FILL_0__11968_ (
);

FILL FILL_0__9142_ (
);

AOI22X1 _11833_ (
    .A(_2491_),
    .B(_2481__bF$buf1),
    .C(_2620_),
    .D(_2130_),
    .Y(_2922_)
);

FILL FILL_0__11548_ (
);

OAI21X1 _11413_ (
    .A(_2528_),
    .B(_2529_),
    .C(_2324_),
    .Y(_2530_)
);

FILL FILL_0__11128_ (
);

FILL SFILL38840x22050 (
);

FILL FILL_5__7585_ (
);

FILL FILL_4__16361_ (
);

FILL FILL_5__7165_ (
);

FILL FILL_3__15774_ (
);

FILL FILL_3__15354_ (
);

FILL FILL_1__7997_ (
);

FILL FILL_1__7577_ (
);

FILL FILL_2__14767_ (
);

FILL FILL_2__14347_ (
);

FILL FILL_0__15381_ (
);

FILL SFILL89960x52050 (
);

FILL FILL_3__8864_ (
);

FILL FILL_3__8444_ (
);

INVX1 _12618_ (
    .A(\datapath_1.Data [17]),
    .Y(_3458_)
);

FILL FILL_4_BUFX2_insert1010 (
);

FILL FILL_1__14701_ (
);

FILL FILL_4_BUFX2_insert1011 (
);

FILL FILL_4_BUFX2_insert1012 (
);

FILL FILL_4_BUFX2_insert1013 (
);

FILL FILL_4_BUFX2_insert1014 (
);

FILL FILL_4__12281_ (
);

FILL FILL_4_BUFX2_insert1015 (
);

FILL FILL_4_BUFX2_insert1016 (
);

FILL FILL_4_BUFX2_insert1017 (
);

FILL FILL_4_BUFX2_insert1018 (
);

FILL FILL_3__16139_ (
);

FILL FILL_4_BUFX2_insert1019 (
);

FILL SFILL33800x48050 (
);

FILL FILL_2__6861_ (
);

FILL SFILL64200x39050 (
);

FILL FILL_5__9731_ (
);

FILL FILL_3__11694_ (
);

FILL FILL_3__11274_ (
);

OAI21X1 _16451_ (
    .A(_6834_),
    .B(ALUZero),
    .C(_6835_),
    .Y(PCEn)
);

FILL FILL_0__16166_ (
);

OAI22X1 _16031_ (
    .A(_5485__bF$buf4),
    .B(_5087_),
    .C(_5483__bF$buf3),
    .D(_5122_),
    .Y(_6487_)
);

FILL FILL_2__10687_ (
);

FILL FILL_2__10267_ (
);

FILL FILL_1__9723_ (
);

FILL FILL_5__11601_ (
);

FILL FILL_3_BUFX2_insert650 (
);

FILL FILL_3__9649_ (
);

FILL FILL_3__9229_ (
);

FILL FILL_3_BUFX2_insert651 (
);

FILL FILL_3_BUFX2_insert652 (
);

FILL FILL_5__14493_ (
);

FILL FILL_3_BUFX2_insert653 (
);

FILL FILL_3_BUFX2_insert654 (
);

FILL FILL_5__14073_ (
);

DFFSR _8793_ (
    .Q(\datapath_1.regfile_1.regOut[15] [3]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_913_[3])
);

FILL FILL_1__15906_ (
);

FILL FILL_3_BUFX2_insert655 (
);

INVX1 _8373_ (
    .A(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_759_)
);

FILL FILL_3_BUFX2_insert656 (
);

FILL FILL_6__7234_ (
);

FILL FILL_3_BUFX2_insert657 (
);

FILL FILL_3_BUFX2_insert658 (
);

FILL FILL_3_BUFX2_insert659 (
);

FILL FILL_4__13486_ (
);

FILL FILL_1__10621_ (
);

FILL FILL_3__12899_ (
);

FILL FILL_2__7226_ (
);

FILL FILL_3__12479_ (
);

FILL FILL_3__12059_ (
);

FILL FILL_1__13093_ (
);

DFFSR _12791_ (
    .Q(\aluControl_1.inst [0]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3490_[0])
);

FILL FILL_0__12086_ (
);

NAND2X1 _12371_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [9]),
    .Y(_3313_)
);

FILL FILL_3__13840_ (
);

FILL FILL_3__13420_ (
);

FILL FILL_3__13000_ (
);

FILL SFILL79960x50050 (
);

FILL FILL_4__8513_ (
);

FILL FILL_5__15698_ (
);

FILL FILL_2__12833_ (
);

FILL FILL_2__12413_ (
);

FILL FILL_5__15278_ (
);

INVX1 _9998_ (
    .A(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_1578_)
);

FILL FILL_6__8439_ (
);

DFFSR _9578_ (
    .Q(\datapath_1.regfile_1.regOut[21] [20]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1303_[20])
);

OAI21X1 _9158_ (
    .A(_1159_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1160_),
    .Y(_1108_[26])
);

FILL FILL_6__8019_ (
);

FILL FILL_1__11826_ (
);

FILL FILL_1__11406_ (
);

FILL SFILL18840x63050 (
);

FILL FILL_0__8833_ (
);

FILL FILL_3__6930_ (
);

FILL FILL_0__10819_ (
);

FILL FILL_1__14298_ (
);

FILL FILL_5__6856_ (
);

FILL FILL_0_BUFX2_insert780 (
);

FILL FILL_4__15632_ (
);

FILL FILL_0_BUFX2_insert781 (
);

FILL FILL_4__15212_ (
);

FILL FILL_0_BUFX2_insert782 (
);

FILL FILL_0_BUFX2_insert783 (
);

NOR2X1 _13996_ (
    .A(_4496_),
    .B(_4493_),
    .Y(_4497_)
);

FILL FILL_0_BUFX2_insert784 (
);

FILL FILL_0_BUFX2_insert785 (
);

INVX1 _13576_ (
    .A(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_4086_)
);

OAI21X1 _13156_ (
    .A(_3734_),
    .B(PCEn_bF$buf3),
    .C(_3735_),
    .Y(_3685_[25])
);

FILL FILL_0_BUFX2_insert786 (
);

FILL FILL_0_BUFX2_insert787 (
);

FILL FILL_3__14625_ (
);

FILL FILL_0_BUFX2_insert788 (
);

FILL FILL_3__14205_ (
);

FILL FILL_0_BUFX2_insert789 (
);

FILL FILL_1__6848_ (
);

FILL FILL_4__9718_ (
);

FILL FILL_2__13618_ (
);

FILL FILL_0__14652_ (
);

FILL FILL_0__14232_ (
);

FILL FILL_5__11198_ (
);

FILL FILL_3__7715_ (
);

FILL FILL_0__9618_ (
);

FILL FILL_4__11972_ (
);

FILL FILL_4__11552_ (
);

FILL FILL_4__11132_ (
);

FILL FILL_1__16024_ (
);

FILL FILL_3__10965_ (
);

FILL FILL_3__10545_ (
);

FILL FILL_3__10125_ (
);

FILL FILL_0__15857_ (
);

INVX1 _15722_ (
    .A(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_6186_)
);

FILL FILL_0__15437_ (
);

NOR2X1 _15302_ (
    .A(_5775_),
    .B(_5773_),
    .Y(_5776_)
);

FILL FILL_0__15017_ (
);

FILL FILL_0__10992_ (
);

FILL FILL_0__10572_ (
);

FILL FILL_2__8184_ (
);

FILL FILL_0__10152_ (
);

FILL SFILL8760x50 (
);

FILL FILL_5__13764_ (
);

FILL FILL_5__13344_ (
);

DFFSR _7644_ (
    .Q(\datapath_1.regfile_1.regOut[6] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_328_[6])
);

INVX1 _7224_ (
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_176_)
);

FILL FILL_4__9891_ (
);

FILL FILL_4__9471_ (
);

FILL FILL_4__12757_ (
);

FILL SFILL48920x57050 (
);

FILL FILL_2__13791_ (
);

FILL FILL_4__12337_ (
);

FILL FILL_2__13371_ (
);

FILL FILL_2__6917_ (
);

FILL FILL_1__12784_ (
);

FILL FILL_1__12364_ (
);

FILL FILL_0__9791_ (
);

FILL FILL_0__9371_ (
);

FILL FILL_2__9389_ (
);

FILL FILL_0__11777_ (
);

FILL FILL_0__11357_ (
);

NOR2X1 _11642_ (
    .A(_2211_),
    .B(_2744_),
    .Y(_2745_)
);

AND2X2 _11222_ (
    .A(_2336_),
    .B(_2340_),
    .Y(_2341_)
);

FILL FILL_6__15976_ (
);

FILL FILL_4__16170_ (
);

FILL FILL_5__14969_ (
);

FILL FILL_5__14549_ (
);

FILL FILL_5__14129_ (
);

FILL FILL_3__15583_ (
);

FILL FILL_3__15163_ (
);

INVX1 _8849_ (
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_995_)
);

DFFSR _8429_ (
    .Q(\datapath_1.regfile_1.regOut[12] [23]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_718_[23])
);

OAI21X1 _8009_ (
    .A(_576_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_577_),
    .Y(_523_[27])
);

FILL FILL_2__14996_ (
);

FILL FILL_2__14576_ (
);

FILL FILL_2__14156_ (
);

FILL FILL_0__15190_ (
);

FILL FILL_5__15910_ (
);

FILL SFILL48920x12050 (
);

FILL FILL_1__13989_ (
);

FILL FILL_1__13569_ (
);

FILL FILL_1__13149_ (
);

FILL FILL_4__14903_ (
);

FILL FILL_3__8253_ (
);

INVX1 _12847_ (
    .A(\datapath_1.a [8]),
    .Y(_3570_)
);

INVX1 _12427_ (
    .A(ALUOut[28]),
    .Y(_3350_)
);

NAND3X1 _12007_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[5]),
    .C(_3032__bF$buf1),
    .Y(_3051_)
);

FILL FILL_5__8599_ (
);

FILL FILL_1__14930_ (
);

FILL FILL_1__14510_ (
);

FILL FILL_6__11896_ (
);

FILL FILL_4__12090_ (
);

FILL FILL_0__13923_ (
);

FILL FILL_3__16368_ (
);

FILL FILL_0__13503_ (
);

FILL FILL_5__10889_ (
);

FILL FILL_5__9540_ (
);

FILL FILL_5__10049_ (
);

FILL FILL_5__9120_ (
);

FILL FILL_3__11083_ (
);

FILL SFILL59080x70050 (
);

FILL FILL_0__16395_ (
);

AOI22X1 _16260_ (
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .B(_5693_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_6710_)
);

FILL FILL_2__10496_ (
);

FILL SFILL38920x55050 (
);

FILL FILL_5__11830_ (
);

FILL FILL_1__9532_ (
);

FILL FILL_5__11410_ (
);

FILL FILL_1__9112_ (
);

FILL FILL_2__16302_ (
);

FILL FILL_3__9878_ (
);

FILL FILL_3__9038_ (
);

FILL FILL_4__10823_ (
);

FILL FILL_4__10403_ (
);

FILL FILL_1__15715_ (
);

FILL FILL_6__7043_ (
);

INVX1 _8182_ (
    .A(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_716_)
);

FILL FILL_4__13295_ (
);

FILL FILL_1__10430_ (
);

FILL FILL_1__10010_ (
);

FILL FILL_0__14708_ (
);

FILL FILL_2_CLKBUF1_insert1080 (
);

FILL FILL_2_CLKBUF1_insert1081 (
);

FILL FILL_2_CLKBUF1_insert1082 (
);

FILL FILL_2_CLKBUF1_insert1083 (
);

FILL FILL_2__7875_ (
);

FILL FILL_2__7455_ (
);

FILL FILL_3__12288_ (
);

FILL FILL_2__7035_ (
);

FILL SFILL3560x54050 (
);

OAI21X1 _12180_ (
    .A(_3172_),
    .B(ALUSrcA_bF$buf6),
    .C(_3173_),
    .Y(\datapath_1.alu_1.ALUInA [21])
);

FILL FILL_5__12615_ (
);

NAND2X1 _6915_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_11_)
);

FILL FILL_6__16094_ (
);

FILL SFILL104440x71050 (
);

FILL FILL_4__8742_ (
);

FILL FILL_4__8322_ (
);

FILL FILL_4__11608_ (
);

FILL FILL_2__12642_ (
);

FILL FILL_2__12222_ (
);

FILL FILL_5__15087_ (
);

OAI21X1 _9387_ (
    .A(_1271_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1272_),
    .Y(_1238_[17])
);

FILL FILL112200x49050 (
);

FILL FILL_1__11635_ (
);

FILL FILL_1__11215_ (
);

FILL FILL_0__8642_ (
);

NOR2X1 _10913_ (
    .A(_2051_),
    .B(_2057_),
    .Y(IRWrite)
);

FILL FILL_0__10628_ (
);

FILL FILL_0__8222_ (
);

FILL FILL_6_BUFX2_insert35 (
);

FILL FILL_4__15861_ (
);

FILL FILL_4__15441_ (
);

FILL FILL_4__15021_ (
);

INVX1 _13385_ (
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_3897_)
);

FILL FILL_2__9601_ (
);

FILL FILL_3__14854_ (
);

FILL FILL_3__14434_ (
);

FILL FILL_3__14014_ (
);

FILL SFILL28920x53050 (
);

FILL SFILL24200x31050 (
);

FILL FILL_4__9527_ (
);

FILL FILL_4__9107_ (
);

FILL FILL_2__13847_ (
);

FILL FILL_0__14881_ (
);

FILL FILL_2__13427_ (
);

FILL FILL_0__14461_ (
);

FILL FILL_2__13007_ (
);

FILL FILL_0__14041_ (
);

FILL FILL_3__7944_ (
);

FILL FILL_0__9847_ (
);

FILL FILL_0__9427_ (
);

FILL FILL_3__7104_ (
);

FILL FILL_0__9007_ (
);

FILL FILL_4__16226_ (
);

FILL SFILL89560x33050 (
);

FILL FILL_4__11781_ (
);

FILL FILL_4__11361_ (
);

FILL FILL_3__15639_ (
);

FILL FILL_3__15219_ (
);

FILL FILL_1__16253_ (
);

FILL FILL_3__10774_ (
);

FILL FILL_0__15666_ (
);

OAI21X1 _15951_ (
    .A(_5006_),
    .B(_5535__bF$buf4),
    .C(_6408_),
    .Y(_6409_)
);

FILL FILL_0__15246_ (
);

INVX1 _15531_ (
    .A(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_6000_)
);

OAI22X1 _15111_ (
    .A(_5489__bF$buf3),
    .B(_4035_),
    .C(_4031_),
    .D(_5504__bF$buf0),
    .Y(_5590_)
);

FILL FILL_0__10381_ (
);

FILL FILL_6__14580_ (
);

FILL FILL_6__14160_ (
);

FILL FILL_3__8729_ (
);

FILL FILL_5__13993_ (
);

FILL FILL_5__13573_ (
);

FILL FILL_5__13153_ (
);

INVX1 _7873_ (
    .A(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_507_)
);

INVX1 _7453_ (
    .A(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_288_)
);

INVX1 _7033_ (
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_69_)
);

FILL SFILL115160x7050 (
);

FILL FILL_4__9280_ (
);

FILL FILL_4__12986_ (
);

FILL SFILL28840x15050 (
);

FILL SFILL94360x82050 (
);

FILL FILL_4__12146_ (
);

FILL FILL_3__11979_ (
);

FILL FILL_3__11559_ (
);

FILL FILL_1__12593_ (
);

FILL FILL_3__11139_ (
);

FILL FILL_1__12173_ (
);

OAI22X1 _16316_ (
    .A(_6764_),
    .B(_5544__bF$buf0),
    .C(_5523_),
    .D(_5438_),
    .Y(_6765_)
);

NOR3X1 _11871_ (
    .A(\datapath_1.ALUResult [31]),
    .B(_2952_),
    .C(_2957_),
    .Y(ALUZero)
);

FILL FILL_0__11586_ (
);

FILL SFILL79160x62050 (
);

FILL FILL_0__11166_ (
);

NOR2X1 _11451_ (
    .A(_2416_),
    .B(_2566_),
    .Y(_2567_)
);

NOR2X1 _11031_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(_2149_),
    .Y(_2150_)
);

FILL FILL_3__12500_ (
);

FILL FILL_2__11913_ (
);

FILL FILL_5__14778_ (
);

FILL FILL_5__14358_ (
);

FILL FILL_3__15392_ (
);

OAI21X1 _8658_ (
    .A(_907_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .C(_908_),
    .Y(_848_[30])
);

OAI21X1 _8238_ (
    .A(_688_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_689_),
    .Y(_653_[18])
);

FILL FILL_1__7195_ (
);

FILL FILL_1__10906_ (
);

FILL SFILL18840x58050 (
);

FILL FILL_2__14385_ (
);

FILL FILL_1__13798_ (
);

FILL FILL_1__13378_ (
);

FILL FILL_4__14712_ (
);

FILL FILL_3__8482_ (
);

OAI21X1 _12656_ (
    .A(_3482_),
    .B(vdd),
    .C(_3483_),
    .Y(_3425_[29])
);

FILL FILL_3__8062_ (
);

NAND3X1 _12236_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\aluControl_1.inst [5]),
    .C(_3198__bF$buf3),
    .Y(_3216_)
);

FILL FILL_3__13705_ (
);

FILL FILL111720x73050 (
);

FILL FILL_0__13732_ (
);

FILL FILL_0__13312_ (
);

FILL FILL_3__16177_ (
);

FILL FILL_5__10698_ (
);

FILL FILL_5__10278_ (
);

FILL SFILL18840x13050 (
);

FILL SFILL84360x80050 (
);

FILL FILL_1__9761_ (
);

FILL FILL_1__9341_ (
);

FILL FILL_4__15917_ (
);

FILL FILL_2__16111_ (
);

FILL FILL_3__9267_ (
);

FILL FILL_4__10632_ (
);

FILL FILL_1__15944_ (
);

FILL SFILL103560x29050 (
);

FILL FILL_1__15524_ (
);

FILL FILL_1__15104_ (
);

FILL FILL_0__14937_ (
);

AOI22X1 _14802_ (
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .B(_4038__bF$buf1),
    .C(_4079__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_5286_)
);

FILL FILL_0__14517_ (
);

FILL FILL_2__7684_ (
);

FILL FILL_3__12097_ (
);

FILL FILL_6__13011_ (
);

FILL FILL_5__12844_ (
);

FILL FILL_5__12424_ (
);

FILL FILL_5__12004_ (
);

FILL FILL_4__8971_ (
);

FILL FILL_4__11837_ (
);

FILL FILL_4__8131_ (
);

FILL FILL_2__12871_ (
);

FILL FILL_4__11417_ (
);

FILL FILL_2__12451_ (
);

FILL FILL_2__12031_ (
);

FILL SFILL93560x78050 (
);

DFFSR _9196_ (
    .Q(\datapath_1.regfile_1.regOut[18] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1108_[22])
);

FILL FILL_1__16309_ (
);

FILL FILL_1__11864_ (
);

FILL FILL_1__11444_ (
);

FILL FILL_1__11024_ (
);

FILL FILL_0__8871_ (
);

FILL FILL_2__8889_ (
);

FILL FILL_0__8451_ (
);

FILL FILL_2__8469_ (
);

FILL SFILL70040x70050 (
);

FILL FILL_0__10437_ (
);

DFFSR _10722_ (
    .Q(\datapath_1.regfile_1.regOut[30] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_1888_[12])
);

FILL SFILL114520x61050 (
);

INVX1 _10302_ (
    .A(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_1740_)
);

FILL FILL_0__10017_ (
);

FILL FILL_6__14636_ (
);

FILL FILL_5__6894_ (
);

FILL FILL_4__15670_ (
);

FILL FILL_6__14216_ (
);

FILL FILL_4__15250_ (
);

DFFSR _13194_ (
    .Q(\datapath_1.mux_iord.din0 [19]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3685_[19])
);

FILL FILL_5__13629_ (
);

FILL FILL_5__13209_ (
);

FILL FILL_3__14663_ (
);

FILL FILL_2__9410_ (
);

FILL FILL_3__14243_ (
);

INVX1 _7929_ (
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_524_)
);

OAI21X1 _7509_ (
    .A(_324_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_325_),
    .Y(_263_[31])
);

FILL FILL_1__6886_ (
);

FILL FILL_4__9756_ (
);

FILL FILL_4__9336_ (
);

FILL FILL_2__13656_ (
);

FILL FILL_2__13236_ (
);

FILL FILL_0__14690_ (
);

FILL FILL_0__14270_ (
);

FILL FILL_1__12649_ (
);

FILL FILL_1__12229_ (
);

FILL FILL_0__9656_ (
);

FILL FILL_3__7753_ (
);

FILL FILL_3__7333_ (
);

NAND2X1 _11927_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[13]),
    .Y(_2993_)
);

FILL FILL_0__9236_ (
);

AOI21X1 _11507_ (
    .A(_2617_),
    .B(_2442_),
    .C(_2618_),
    .Y(_2619_)
);

FILL FILL_5__7679_ (
);

FILL FILL_4__16035_ (
);

FILL FILL_6__10976_ (
);

AOI22X1 _14399_ (
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .B(_4005__bF$buf2),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_4892_)
);

FILL FILL_4__11590_ (
);

FILL FILL_4__11170_ (
);

FILL FILL_3__15868_ (
);

FILL FILL_3__15448_ (
);

FILL FILL_3__15028_ (
);

FILL FILL_1__16062_ (
);

FILL FILL_5__8620_ (
);

FILL FILL_5__8200_ (
);

FILL FILL_3__10163_ (
);

FILL FILL_6_BUFX2_insert541 (
);

FILL SFILL59080x65050 (
);

FILL FILL_0__15895_ (
);

OAI21X1 _15760_ (
    .A(_5524__bF$buf2),
    .B(_4798_),
    .C(_6222_),
    .Y(_6223_)
);

FILL FILL_0__15475_ (
);

NOR2X1 _15340_ (
    .A(_4299_),
    .B(_5549__bF$buf4),
    .Y(_5813_)
);

FILL FILL_0__15055_ (
);

FILL FILL_6_BUFX2_insert546 (
);

FILL FILL_0__10190_ (
);

FILL FILL_5__10910_ (
);

FILL FILL_1__8612_ (
);

FILL FILL_2__15802_ (
);

FILL FILL_3__8958_ (
);

FILL FILL_3__8118_ (
);

FILL SFILL3640x42050 (
);

FILL FILL_5__13382_ (
);

INVX1 _7682_ (
    .A(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_400_)
);

DFFSR _7262_ (
    .Q(\datapath_1.regfile_1.regOut[3] [8]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_133_[8])
);

FILL FILL_4__12375_ (
);

FILL FILL_2__6955_ (
);

FILL FILL_3__11788_ (
);

FILL FILL_5__9405_ (
);

FILL FILL_3__11368_ (
);

FILL SFILL59000x63050 (
);

FILL FILL_6__12702_ (
);

INVX1 _16125_ (
    .A(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_6578_)
);

FILL SFILL3560x49050 (
);

FILL SFILL59080x20050 (
);

OAI22X1 _11680_ (
    .A(_2181_),
    .B(_2344__bF$buf1),
    .C(_2480_),
    .D(_2399_),
    .Y(_2781_)
);

FILL FILL_0__11395_ (
);

NOR2X1 _11260_ (
    .A(_2377_),
    .B(_2378_),
    .Y(_2379_)
);

FILL SFILL104440x66050 (
);

FILL FILL_4__7822_ (
);

FILL FILL_5__14587_ (
);

FILL FILL_2__11722_ (
);

FILL FILL_5__14167_ (
);

FILL FILL_2__11302_ (
);

OAI21X1 _8887_ (
    .A(_1019_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1020_),
    .Y(_978_[21])
);

OAI21X1 _8467_ (
    .A(_800_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_801_),
    .Y(_783_[9])
);

DFFSR _8047_ (
    .Q(\datapath_1.regfile_1.regOut[9] [25]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_523_[25])
);

FILL SFILL49480x77050 (
);

FILL FILL_2__14194_ (
);

FILL FILL_0__7722_ (
);

FILL FILL_0__7302_ (
);

FILL FILL_4__14941_ (
);

FILL FILL_4__14521_ (
);

FILL FILL_4__14101_ (
);

FILL SFILL43960x7050 (
);

OAI21X1 _12885_ (
    .A(_3594_),
    .B(vdd),
    .C(_3595_),
    .Y(_3555_[20])
);

FILL SFILL49080x63050 (
);

OAI21X1 _12465_ (
    .A(_3375_),
    .B(vdd),
    .C(_3376_),
    .Y(_3360_[8])
);

AOI22X1 _12045_ (
    .A(\datapath_1.ALUResult [14]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3080_)
);

FILL FILL_3__13934_ (
);

FILL FILL_3__13514_ (
);

FILL SFILL28920x48050 (
);

FILL FILL_4__8607_ (
);

FILL FILL_5_BUFX2_insert560 (
);

FILL SFILL73560x74050 (
);

FILL FILL_5_BUFX2_insert561 (
);

FILL SFILL104440x21050 (
);

FILL FILL_5_BUFX2_insert562 (
);

FILL FILL_2__12507_ (
);

FILL FILL_0__13961_ (
);

FILL FILL_5_BUFX2_insert563 (
);

FILL FILL_0__13541_ (
);

FILL FILL_0__13121_ (
);

FILL FILL_5_BUFX2_insert564 (
);

FILL FILL_5_BUFX2_insert565 (
);

FILL FILL_5_BUFX2_insert566 (
);

FILL FILL_5_BUFX2_insert567 (
);

FILL FILL_5_BUFX2_insert568 (
);

FILL FILL_1_BUFX2_insert0 (
);

FILL FILL_5_BUFX2_insert569 (
);

FILL FILL_1_BUFX2_insert1 (
);

FILL FILL_2__15399_ (
);

FILL FILL_1_BUFX2_insert2 (
);

FILL FILL_1_BUFX2_insert3 (
);

FILL FILL_1_BUFX2_insert4 (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_5__16313_ (
);

FILL FILL_0__8507_ (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

FILL FILL_1__9990_ (
);

FILL FILL_1__9150_ (
);

FILL FILL_4__15726_ (
);

FILL FILL_1_BUFX2_insert1090 (
);

FILL FILL_4__15306_ (
);

FILL FILL_1_BUFX2_insert1091 (
);

FILL FILL_2__16340_ (
);

FILL FILL_1_BUFX2_insert1092 (
);

FILL SFILL73960x43050 (
);

FILL FILL_3__9496_ (
);

FILL FILL_1_BUFX2_insert1093 (
);

FILL SFILL49000x61050 (
);

FILL FILL_4__10441_ (
);

FILL FILL_4__10021_ (
);

FILL FILL_3__14719_ (
);

FILL FILL_1__15753_ (
);

FILL FILL_1__15333_ (
);

FILL SFILL94440x70050 (
);

FILL FILL_0__14746_ (
);

INVX1 _14611_ (
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_5099_)
);

FILL FILL_0__14326_ (
);

FILL FILL_2__7493_ (
);

FILL FILL_2__7073_ (
);

FILL FILL_3__7809_ (
);

FILL FILL_5__12653_ (
);

FILL FILL_5__12233_ (
);

INVX1 _6953_ (
    .A(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_36_)
);

FILL FILL_2_BUFX2_insert690 (
);

FILL FILL_2_BUFX2_insert691 (
);

FILL FILL_4__8780_ (
);

FILL FILL_2_BUFX2_insert692 (
);

FILL FILL_4__8360_ (
);

FILL FILL_2_BUFX2_insert693 (
);

FILL SFILL94360x77050 (
);

FILL FILL_2_BUFX2_insert694 (
);

FILL FILL_4__11646_ (
);

FILL FILL_2_BUFX2_insert695 (
);

FILL FILL_4__11226_ (
);

FILL FILL_2_BUFX2_insert696 (
);

FILL FILL_2__12260_ (
);

FILL FILL_2_BUFX2_insert697 (
);

FILL FILL_2_BUFX2_insert698 (
);

FILL FILL_1__16118_ (
);

FILL FILL_2_BUFX2_insert699 (
);

FILL FILL_3__10639_ (
);

FILL FILL_1__11673_ (
);

FILL FILL_1__11253_ (
);

NOR2X1 _15816_ (
    .A(_6274_),
    .B(_6276_),
    .Y(_6277_)
);

FILL FILL_2__8698_ (
);

FILL SFILL79160x57050 (
);

INVX1 _10951_ (
    .A(_2074_),
    .Y(_2084_)
);

FILL FILL_0__8260_ (
);

FILL FILL_0__10666_ (
);

INVX1 _10531_ (
    .A(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_1852_)
);

FILL FILL_0__10246_ (
);

INVX1 _10111_ (
    .A(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_1633_)
);

FILL FILL_5__13858_ (
);

FILL FILL_5__13438_ (
);

FILL FILL_3__14892_ (
);

FILL FILL_3__14472_ (
);

FILL FILL_5__13018_ (
);

FILL FILL_3__14052_ (
);

OAI21X1 _7738_ (
    .A(_436_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_437_),
    .Y(_393_[22])
);

OAI21X1 _7318_ (
    .A(_217_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .C(_218_),
    .Y(_198_[10])
);

FILL FILL_4__9985_ (
);

FILL FILL_4__9145_ (
);

FILL FILL_2__13885_ (
);

FILL FILL_2__13465_ (
);

FILL FILL111800x61050 (
);

FILL FILL_2__13045_ (
);

FILL SFILL63960x41050 (
);

FILL SFILL94360x32050 (
);

FILL FILL_1__12878_ (
);

FILL FILL_1__12458_ (
);

FILL FILL_1__12038_ (
);

FILL FILL_6_CLKBUF1_insert142 (
);

FILL FILL_3__7982_ (
);

FILL FILL_0__9885_ (
);

FILL FILL_3__7562_ (
);

FILL FILL_0__9465_ (
);

FILL FILL_0__9045_ (
);

OAI21X1 _11736_ (
    .A(_2147_),
    .B(_2160_),
    .C(_2503_),
    .Y(_2833_)
);

AND2X2 _11316_ (
    .A(_2432_),
    .B(_2434_),
    .Y(_2435_)
);

FILL FILL_6_CLKBUF1_insert147 (
);

FILL FILL_5__7488_ (
);

FILL SFILL79160x12050 (
);

FILL FILL_5__7068_ (
);

FILL FILL_4__16264_ (
);

FILL FILL_3__15677_ (
);

FILL FILL_3__15257_ (
);

FILL FILL_1__16291_ (
);

FILL FILL_3__10392_ (
);

FILL FILL_0__15284_ (
);

FILL SFILL84360x75050 (
);

FILL FILL_1__8841_ (
);

FILL SFILL79160x2050 (
);

FILL FILL_1__8001_ (
);

FILL FILL_2__15611_ (
);

FILL FILL_3__8767_ (
);

FILL FILL_3__8347_ (
);

FILL FILL_1__14604_ (
);

OAI21X1 _7491_ (
    .A(_312_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .C(_313_),
    .Y(_263_[25])
);

OAI21X1 _7071_ (
    .A(_93_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .C(_94_),
    .Y(_68_[13])
);

FILL FILL_4__12184_ (
);

FILL FILL_5__9634_ (
);

FILL FILL_3__11597_ (
);

FILL FILL_5__9214_ (
);

FILL FILL_3__11177_ (
);

INVX1 _16354_ (
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_6790_)
);

FILL FILL_0__16069_ (
);

FILL FILL_5__11924_ (
);

FILL FILL_1__9626_ (
);

FILL FILL_5__11504_ (
);

FILL FILL_1__9206_ (
);

FILL SFILL84360x30050 (
);

FILL FILL_4__7631_ (
);

FILL FILL_4__10917_ (
);

FILL FILL_4__7211_ (
);

FILL FILL_2__11951_ (
);

FILL FILL_5__14396_ (
);

FILL FILL_2__11531_ (
);

FILL FILL_2__11111_ (
);

OAI21X1 _8696_ (
    .A(_976_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .C(_977_),
    .Y(_913_[0])
);

FILL FILL_1__15809_ (
);

NAND2X1 _8276_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_715_)
);

FILL FILL_1__10944_ (
);

FILL FILL_4__13389_ (
);

FILL FILL_1__10524_ (
);

FILL FILL_1__10104_ (
);

FILL FILL_0__7951_ (
);

FILL FILL_2__7969_ (
);

BUFX2 BUFX2_insert380 (
    .A(_3196_),
    .Y(_3196__bF$buf0)
);

FILL FILL_2__7549_ (
);

BUFX2 BUFX2_insert381 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf7 )
);

FILL FILL_0__7111_ (
);

BUFX2 BUFX2_insert382 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf6 )
);

BUFX2 BUFX2_insert383 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf5 )
);

BUFX2 BUFX2_insert384 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf4 )
);

BUFX2 BUFX2_insert385 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf3 )
);

FILL FILL_4__14750_ (
);

BUFX2 BUFX2_insert386 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf2 )
);

FILL FILL_4__14330_ (
);

FILL SFILL3720x75050 (
);

BUFX2 BUFX2_insert387 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf1 )
);

BUFX2 BUFX2_insert388 (
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf0 )
);

DFFSR _12694_ (
    .Q(\datapath_1.Data [31]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3425_[31])
);

BUFX2 BUFX2_insert389 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf4 )
);

NAND3X1 _12274_ (
    .A(_3242_),
    .B(_3243_),
    .C(_3244_),
    .Y(\datapath_1.alu_1.ALUInB [14])
);

FILL FILL_2__8910_ (
);

FILL FILL_5__12709_ (
);

FILL FILL_3__13743_ (
);

FILL SFILL43960x82050 (
);

FILL FILL_3__13323_ (
);

FILL FILL_4__8836_ (
);

FILL SFILL69080x17050 (
);

FILL FILL_2__12736_ (
);

FILL FILL_0__13770_ (
);

FILL FILL_2__12316_ (
);

FILL FILL_0__13350_ (
);

FILL FILL_1__11729_ (
);

FILL FILL_1__11309_ (
);

FILL SFILL78680x81050 (
);

FILL FILL_0__8736_ (
);

FILL FILL_5__16122_ (
);

FILL FILL_0__8316_ (
);

FILL FILL_4__15955_ (
);

FILL FILL_4__15535_ (
);

FILL SFILL114520x11050 (
);

FILL FILL_4__15115_ (
);

AOI22X1 _13899_ (
    .A(_4038__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [9]),
    .C(\datapath_1.regfile_1.regOut[18] [9]),
    .D(_4135_),
    .Y(_4402_)
);

FILL FILL_4__10670_ (
);

OAI22X1 _13479_ (
    .A(_3989_),
    .B(_3949_),
    .C(_3983__bF$buf2),
    .D(_3988_),
    .Y(_3990_)
);

FILL FILL_4__10250_ (
);

DFFSR _13059_ (
    .Q(_2_[12]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3620_[12])
);

FILL FILL_3__14948_ (
);

FILL SFILL3720x30050 (
);

FILL FILL_1__15982_ (
);

FILL FILL_3__14528_ (
);

FILL FILL_1__15562_ (
);

FILL FILL_3__14108_ (
);

FILL FILL_1__15142_ (
);

FILL FILL_5__7700_ (
);

FILL FILL_0__14975_ (
);

INVX1 _14840_ (
    .A(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_5323_)
);

FILL FILL_0__14555_ (
);

FILL FILL_0__14135_ (
);

OAI22X1 _14420_ (
    .A(_4910_),
    .B(_3930__bF$buf1),
    .C(_3920_),
    .D(_4911_),
    .Y(_4912_)
);

NOR2X1 _14000_ (
    .A(_4500_),
    .B(_3971__bF$buf0),
    .Y(_4501_)
);

FILL FILL_3__7618_ (
);

FILL SFILL3640x37050 (
);

FILL FILL_5__12882_ (
);

FILL FILL_5__12462_ (
);

FILL FILL_5__12042_ (
);

FILL SFILL43880x44050 (
);

FILL FILL_4__11875_ (
);

FILL FILL_4__11455_ (
);

FILL FILL_4__11035_ (
);

FILL FILL_1__16347_ (
);

FILL FILL_5__8905_ (
);

FILL FILL_3__10448_ (
);

FILL FILL_3__10028_ (
);

FILL FILL_1__11482_ (
);

FILL FILL_1__11062_ (
);

FILL SFILL108840x62050 (
);

INVX1 _15625_ (
    .A(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_6091_)
);

FILL SFILL38120x17050 (
);

NOR2X1 _15205_ (
    .A(_5680_),
    .B(_5681_),
    .Y(_5682_)
);

FILL SFILL59080x15050 (
);

FILL FILL_0__10895_ (
);

INVX1 _10760_ (
    .A(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_1964_)
);

FILL FILL_2__8087_ (
);

DFFSR _10340_ (
    .Q(\datapath_1.regfile_1.regOut[27] [14]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_1693_[14])
);

FILL FILL_0__10055_ (
);

FILL FILL_4__6902_ (
);

FILL FILL_5__13667_ (
);

FILL FILL_2__10802_ (
);

FILL FILL_5__13247_ (
);

FILL FILL_3__14281_ (
);

OAI21X1 _7967_ (
    .A(_548_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .C(_549_),
    .Y(_523_[13])
);

OAI21X1 _7547_ (
    .A(_329_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .C(_330_),
    .Y(_328_[1])
);

DFFSR _7127_ (
    .Q(\datapath_1.regfile_1.regOut[2] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_68_[1])
);

FILL FILL_4__9794_ (
);

FILL FILL_4__9374_ (
);

FILL FILL_2__13694_ (
);

FILL FILL_2__13274_ (
);

FILL FILL_1__12267_ (
);

FILL FILL_4__13601_ (
);

FILL SFILL59000x13050 (
);

FILL SFILL49080x58050 (
);

FILL FILL_3__7371_ (
);

INVX1 _11965_ (
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3018_)
);

FILL FILL_0__9274_ (
);

OAI21X1 _11545_ (
    .A(_2410_),
    .B(_2344__bF$buf2),
    .C(_2654_),
    .Y(_2655_)
);

FILL FILL_5_CLKBUF1_insert130 (
);

NOR2X1 _11125_ (
    .A(_2242_),
    .B(_2243_),
    .Y(_2244_)
);

FILL FILL_5_CLKBUF1_insert131 (
);

FILL FILL_6__15879_ (
);

FILL FILL_5_CLKBUF1_insert132 (
);

FILL FILL_6__15459_ (
);

FILL FILL_5__7297_ (
);

FILL FILL_5_CLKBUF1_insert133 (
);

FILL FILL_5_CLKBUF1_insert134 (
);

FILL FILL_4__16073_ (
);

FILL FILL_5_CLKBUF1_insert135 (
);

FILL FILL_5_CLKBUF1_insert136 (
);

FILL FILL_5_CLKBUF1_insert137 (
);

FILL FILL_5_CLKBUF1_insert138 (
);

FILL FILL_5_CLKBUF1_insert139 (
);

FILL FILL_0__12621_ (
);

FILL FILL_3__15486_ (
);

FILL FILL_3__15066_ (
);

FILL FILL_0__12201_ (
);

FILL FILL_6_BUFX2_insert920 (
);

FILL FILL_1__7289_ (
);

FILL FILL_2__14899_ (
);

FILL FILL_2__14479_ (
);

FILL SFILL28520x29050 (
);

FILL FILL_2__14059_ (
);

FILL FILL_0__15093_ (
);

FILL FILL_6_BUFX2_insert925 (
);

FILL SFILL33880x42050 (
);

FILL FILL_5__15813_ (
);

FILL FILL_1__8650_ (
);

FILL FILL_1__8230_ (
);

FILL FILL_4__14806_ (
);

FILL FILL_2__15840_ (
);

FILL FILL_3__8996_ (
);

FILL FILL_2__15420_ (
);

FILL SFILL49000x56050 (
);

FILL FILL_3__8576_ (
);

FILL FILL_2__15000_ (
);

FILL FILL_1__14833_ (
);

FILL SFILL49080x13050 (
);

FILL FILL_1__14413_ (
);

FILL FILL_6__11799_ (
);

FILL FILL_6__11379_ (
);

FILL SFILL94440x65050 (
);

FILL FILL_0__13826_ (
);

FILL FILL_0__13406_ (
);

FILL FILL_2__6993_ (
);

FILL FILL_5__9863_ (
);

FILL FILL_5__9023_ (
);

FILL FILL_0__16298_ (
);

NOR3X1 _16163_ (
    .A(_6606_),
    .B(_6594_),
    .C(_6615_),
    .Y(_6616_)
);

FILL FILL_2__10399_ (
);

FILL FILL_1__9855_ (
);

FILL FILL_5__11733_ (
);

FILL FILL_5__11313_ (
);

FILL FILL_1__9015_ (
);

FILL FILL_2__16205_ (
);

FILL FILL_4__7860_ (
);

FILL FILL_4__7440_ (
);

FILL FILL_2__11760_ (
);

FILL FILL_4__10306_ (
);

FILL FILL_2__11340_ (
);

FILL SFILL49000x11050 (
);

FILL FILL_1__15618_ (
);

NAND2X1 _8085_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_608_)
);

FILL FILL_1__10753_ (
);

FILL FILL_0__7760_ (
);

FILL SFILL94440x20050 (
);

FILL FILL_2__7358_ (
);

FILL FILL_0__7340_ (
);

FILL FILL_6__13945_ (
);

FILL SFILL18840x3050 (
);

FILL FILL_6__13105_ (
);

FILL SFILL23800x83050 (
);

FILL SFILL18760x8050 (
);

NAND3X1 _12083_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[24]),
    .C(_3032__bF$buf0),
    .Y(_3108_)
);

FILL FILL_5__12518_ (
);

FILL FILL_3__13972_ (
);

FILL FILL_3__13552_ (
);

FILL FILL_3__13132_ (
);

FILL SFILL8840x82050 (
);

FILL FILL_4__8645_ (
);

FILL FILL_4__8225_ (
);

FILL FILL_5_BUFX2_insert940 (
);

FILL FILL_2__12965_ (
);

FILL FILL_5_BUFX2_insert941 (
);

FILL FILL_5_BUFX2_insert942 (
);

FILL FILL_2__12125_ (
);

FILL FILL_5_BUFX2_insert943 (
);

FILL FILL_5_BUFX2_insert944 (
);

FILL SFILL94360x27050 (
);

FILL FILL_5_BUFX2_insert945 (
);

FILL FILL_5_BUFX2_insert946 (
);

FILL FILL_5_BUFX2_insert947 (
);

FILL FILL_1__11958_ (
);

FILL FILL_5_BUFX2_insert948 (
);

FILL FILL_5_BUFX2_insert949 (
);

FILL FILL_1__11538_ (
);

FILL FILL_1__11118_ (
);

FILL FILL_0__8965_ (
);

FILL FILL_5__16351_ (
);

FILL FILL_6__9932_ (
);

FILL SFILL84440x63050 (
);

FILL FILL_0__8125_ (
);

OAI21X1 _10816_ (
    .A(_2000_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .C(_2001_),
    .Y(_1953_[24])
);

FILL FILL_5__6988_ (
);

FILL SFILL63560x22050 (
);

FILL FILL_4__15764_ (
);

FILL FILL_4__15344_ (
);

NAND2X1 _13288_ (
    .A(_3763_),
    .B(_3772_),
    .Y(_3826_)
);

FILL FILL_2__9924_ (
);

FILL FILL_2__9504_ (
);

FILL FILL_3__14757_ (
);

FILL FILL_1__15791_ (
);

FILL FILL_3__14337_ (
);

FILL FILL_1__15371_ (
);

FILL FILL_0__14784_ (
);

FILL FILL_0__14364_ (
);

FILL FILL111800x11050 (
);

FILL FILL_1__7501_ (
);

FILL FILL_3__7847_ (
);

FILL FILL_3__7427_ (
);

FILL FILL_5__12271_ (
);

OAI21X1 _6991_ (
    .A(_60_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .C(_61_),
    .Y(_3_[29])
);

FILL FILL_4__16129_ (
);

FILL FILL_4__11684_ (
);

FILL FILL_4__11264_ (
);

FILL SFILL13800x81050 (
);

FILL FILL_1__16156_ (
);

FILL FILL_3__10677_ (
);

FILL FILL_5__8714_ (
);

FILL FILL_3__10257_ (
);

FILL FILL_1__11291_ (
);

FILL FILL_0__15989_ (
);

INVX2 _15854_ (
    .A(_5527__bF$buf1),
    .Y(_6314_)
);

FILL FILL_0__15569_ (
);

FILL FILL_0__15149_ (
);

NOR2X1 _15434_ (
    .A(_5904_),
    .B(_5897_),
    .Y(_5905_)
);

NOR3X1 _15014_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5492_),
    .C(_5493_),
    .Y(_5494_)
);

FILL FILL_0__10284_ (
);

FILL FILL_3_BUFX2_insert1020 (
);

FILL FILL_1__8706_ (
);

FILL FILL_3_BUFX2_insert1021 (
);

FILL SFILL84360x25050 (
);

FILL FILL_3_BUFX2_insert1022 (
);

FILL FILL_6__14063_ (
);

FILL FILL_3_BUFX2_insert1023 (
);

FILL FILL_3_BUFX2_insert1024 (
);

FILL FILL_3_BUFX2_insert1025 (
);

FILL FILL_3_BUFX2_insert1026 (
);

FILL FILL_3_BUFX2_insert1027 (
);

FILL FILL_3_BUFX2_insert1028 (
);

FILL FILL_5__13896_ (
);

FILL FILL_3_BUFX2_insert1029 (
);

FILL FILL_5__13476_ (
);

DFFSR _7776_ (
    .Q(\datapath_1.regfile_1.regOut[7] [10]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_393_[10])
);

FILL FILL_3__14090_ (
);

NAND2X1 _7356_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_244_)
);

FILL FILL_4__12889_ (
);

FILL FILL_4__12469_ (
);

FILL FILL_4__12049_ (
);

FILL FILL_2__13083_ (
);

FILL FILL_5__9919_ (
);

FILL FILL_1__12496_ (
);

FILL FILL_1__12076_ (
);

FILL FILL_4__13830_ (
);

NAND3X1 _16219_ (
    .A(_6662_),
    .B(_6663_),
    .C(_6669_),
    .Y(_6670_)
);

FILL FILL_4__13410_ (
);

FILL FILL_3__7180_ (
);

INVX1 _11774_ (
    .A(_2868_),
    .Y(\datapath_1.ALUResult [7])
);

FILL FILL_0__9083_ (
);

FILL FILL_0__11489_ (
);

OAI21X1 _11354_ (
    .A(_2469_),
    .B(_2471_),
    .C(_2468_),
    .Y(_2472_)
);

FILL FILL_0__11069_ (
);

FILL SFILL43960x77050 (
);

FILL FILL_3__12823_ (
);

FILL FILL_3__12403_ (
);

FILL FILL_4_CLKBUF1_insert120 (
);

FILL FILL_4_CLKBUF1_insert121 (
);

FILL FILL_2__11816_ (
);

FILL FILL_4_CLKBUF1_insert122 (
);

FILL FILL_0__12850_ (
);

FILL FILL_0__12430_ (
);

FILL FILL_4_CLKBUF1_insert123 (
);

FILL FILL_3__15295_ (
);

FILL SFILL114680x50 (
);

FILL FILL_0__12010_ (
);

FILL FILL_4_CLKBUF1_insert124 (
);

FILL FILL_4_CLKBUF1_insert125 (
);

FILL FILL_4_CLKBUF1_insert126 (
);

FILL FILL_1__7098_ (
);

FILL FILL_4_CLKBUF1_insert127 (
);

FILL FILL_1__10809_ (
);

FILL FILL_4_CLKBUF1_insert128 (
);

FILL FILL_4_CLKBUF1_insert129 (
);

FILL FILL112360x81050 (
);

FILL FILL_2__14288_ (
);

FILL FILL_5__15622_ (
);

FILL FILL_5__15202_ (
);

FILL FILL_0__7816_ (
);

NAND2X1 _9922_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1548_)
);

NAND2X1 _9502_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1329_)
);

FILL FILL_4__14615_ (
);

NAND2X1 _12979_ (
    .A(vdd),
    .B(\datapath_1.rd2 [9]),
    .Y(_3638_)
);

FILL FILL_3__8385_ (
);

DFFSR _12559_ (
    .Q(ALUOut[24]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3360_[24])
);

FILL SFILL89960x50 (
);

INVX1 _12139_ (
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_3146_)
);

FILL SFILL3720x25050 (
);

FILL FILL_3__13608_ (
);

FILL FILL_1__14642_ (
);

FILL FILL_1__14222_ (
);

FILL FILL_0__13635_ (
);

INVX1 _13920_ (
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_4423_)
);

FILL FILL_0__13215_ (
);

INVX1 _13500_ (
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_4011_)
);

FILL FILL_5__9672_ (
);

FILL FILL_5__9252_ (
);

OAI21X1 _16392_ (
    .A(_6814_),
    .B(gnd),
    .C(_6815_),
    .Y(_6769_[23])
);

FILL FILL_5__16407_ (
);

FILL FILL_5__11962_ (
);

FILL FILL_1__9664_ (
);

FILL FILL_5__11542_ (
);

FILL FILL_1__9244_ (
);

FILL FILL_5__11122_ (
);

FILL SFILL104520x49050 (
);

FILL SFILL43880x39050 (
);

FILL FILL_2__16014_ (
);

FILL FILL_4__10955_ (
);

FILL FILL_4__10535_ (
);

FILL FILL_4__10115_ (
);

FILL FILL_1__15847_ (
);

FILL FILL_1__15427_ (
);

FILL FILL_1__15007_ (
);

FILL FILL_1__10982_ (
);

FILL FILL_1__10562_ (
);

FILL FILL_1__10142_ (
);

OAI22X1 _14705_ (
    .A(_3949_),
    .B(_5190_),
    .C(_5189_),
    .D(_3967__bF$buf0),
    .Y(_5191_)
);

FILL SFILL43480x25050 (
);

FILL FILL112280x43050 (
);

FILL FILL_2__7587_ (
);

BUFX2 BUFX2_insert760 (
    .A(_3924_),
    .Y(_3924__bF$buf3)
);

FILL FILL_2__7167_ (
);

BUFX2 BUFX2_insert761 (
    .A(_3924_),
    .Y(_3924__bF$buf2)
);

BUFX2 BUFX2_insert762 (
    .A(_3924_),
    .Y(_3924__bF$buf1)
);

BUFX2 BUFX2_insert763 (
    .A(_3924_),
    .Y(_3924__bF$buf0)
);

BUFX2 BUFX2_insert764 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf4 )
);

BUFX2 BUFX2_insert765 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf3 )
);

BUFX2 BUFX2_insert766 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf2 )
);

BUFX2 BUFX2_insert767 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf1 )
);

BUFX2 BUFX2_insert768 (
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf0 )
);

BUFX2 BUFX2_insert769 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf7 )
);

FILL FILL_5__12747_ (
);

FILL FILL_3__13781_ (
);

FILL FILL_5__12327_ (
);

FILL FILL_3__13361_ (
);

FILL FILL_4__8874_ (
);

FILL FILL_4__8454_ (
);

FILL FILL_2__12774_ (
);

FILL FILL_2__12354_ (
);

INVX1 _9099_ (
    .A(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_1121_)
);

FILL FILL_1__11767_ (
);

FILL FILL_1__11347_ (
);

FILL FILL_0__8774_ (
);

FILL FILL_5__16160_ (
);

FILL FILL_3__6871_ (
);

FILL FILL_6__9741_ (
);

FILL FILL_0__8354_ (
);

OAI21X1 _10625_ (
    .A(_1893_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .C(_1894_),
    .Y(_1888_[3])
);

DFFSR _10205_ (
    .Q(\datapath_1.regfile_1.regOut[26] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_1628_[7])
);

FILL FILL_4__15993_ (
);

FILL FILL_6__14539_ (
);

FILL FILL_4__15573_ (
);

FILL FILL_6__14119_ (
);

FILL FILL_4__15153_ (
);

INVX1 _13097_ (
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_3696_)
);

FILL FILL_3__14986_ (
);

FILL FILL_2__9733_ (
);

FILL FILL_3__14566_ (
);

FILL FILL_0__11701_ (
);

FILL FILL_3__14146_ (
);

FILL FILL_1__15180_ (
);

FILL FILL_4__9659_ (
);

FILL SFILL54760x78050 (
);

FILL FILL_4__9239_ (
);

FILL FILL_2__13979_ (
);

FILL FILL_2__13559_ (
);

FILL FILL_0__14593_ (
);

FILL FILL_2__13139_ (
);

FILL SFILL33880x37050 (
);

FILL FILL_0__14173_ (
);

FILL FILL_1__7730_ (
);

FILL FILL_1__7310_ (
);

FILL FILL_2__14920_ (
);

FILL FILL_2__14500_ (
);

FILL FILL_0__9979_ (
);

FILL FILL_3__7236_ (
);

FILL FILL_0__9139_ (
);

FILL FILL_5__12080_ (
);

FILL FILL_1__13913_ (
);

FILL FILL_4__16358_ (
);

FILL FILL_6__10879_ (
);

FILL FILL_4__11493_ (
);

FILL FILL_4__11073_ (
);

FILL FILL_0__12906_ (
);

FILL FILL_1__16385_ (
);

FILL FILL_3__10486_ (
);

FILL FILL_5__8523_ (
);

FILL FILL_5__8103_ (
);

FILL FILL_3__10066_ (
);

FILL FILL_0__15798_ (
);

FILL FILL_0__15378_ (
);

OAI22X1 _15663_ (
    .A(_5526__bF$buf3),
    .B(_4706_),
    .C(_4688_),
    .D(_5527__bF$buf4),
    .Y(_6128_)
);

FILL FILL_6__11400_ (
);

AOI21X1 _15243_ (
    .A(_5696_),
    .B(_5718_),
    .C(_5509_),
    .Y(_5719_)
);

FILL FILL_5__10813_ (
);

FILL FILL_1__8515_ (
);

FILL FILL_2__15705_ (
);

FILL FILL_4__6940_ (
);

FILL FILL_5__13285_ (
);

FILL FILL_2__10420_ (
);

FILL FILL_2__10000_ (
);

NAND2X1 _7585_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_356_)
);

NAND2X1 _7165_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_137_)
);

FILL FILL_4__12698_ (
);

FILL FILL_4__12278_ (
);

FILL FILL_3__9802_ (
);

FILL SFILL94440x15050 (
);

FILL FILL_2__6858_ (
);

FILL FILL_0__6840_ (
);

FILL FILL_5__9728_ (
);

FILL SFILL23800x78050 (
);

DFFSR _16448_ (
    .Q(\datapath_1.regfile_1.regOut[0] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_6769_[31])
);

INVX1 _16028_ (
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_6484_)
);

OAI21X1 _11583_ (
    .A(_2689_),
    .B(_2272_),
    .C(_2248_),
    .Y(_2690_)
);

FILL FILL_0__11298_ (
);

OAI21X1 _11163_ (
    .A(_2221_),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .C(_2281_),
    .Y(_2282_)
);

FILL SFILL23880x35050 (
);

FILL SFILL54280x26050 (
);

FILL FILL_3__12632_ (
);

FILL FILL_3__12212_ (
);

FILL FILL_4__7725_ (
);

FILL FILL_4__7305_ (
);

FILL FILL_2__11625_ (
);

FILL FILL_2__11205_ (
);

FILL SFILL39000x49050 (
);

FILL FILL_1__10618_ (
);

FILL FILL_2__14097_ (
);

FILL FILL_5__15851_ (
);

FILL FILL_5__15431_ (
);

FILL FILL_5__15011_ (
);

FILL FILL_0__7625_ (
);

FILL FILL_0__7205_ (
);

NAND2X1 _9731_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1441_)
);

DFFSR _9311_ (
    .Q(\datapath_1.regfile_1.regOut[19] [9]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_1173_[9])
);

FILL FILL_4__14844_ (
);

FILL FILL_4__14424_ (
);

FILL FILL_4__14004_ (
);

INVX1 _12788_ (
    .A(\control_1.op [5]),
    .Y(_3551_)
);

FILL FILL_3__8194_ (
);

NAND2X1 _12368_ (
    .A(MemToReg_bF$buf2),
    .B(\datapath_1.Data [8]),
    .Y(_3311_)
);

FILL FILL_3__13837_ (
);

FILL FILL_1__14871_ (
);

FILL FILL_3__13417_ (
);

FILL FILL_1__14451_ (
);

FILL FILL_1__14031_ (
);

FILL FILL_0__13864_ (
);

FILL FILL_0__13444_ (
);

FILL FILL_0__13024_ (
);

FILL FILL_5__9481_ (
);

FILL FILL_3__6927_ (
);

FILL FILL_5__16216_ (
);

FILL FILL_1__9893_ (
);

FILL FILL_5__11771_ (
);

FILL FILL_1__9473_ (
);

FILL FILL_5__11351_ (
);

FILL FILL_4__15629_ (
);

FILL FILL_4__15209_ (
);

FILL FILL_2__16243_ (
);

FILL FILL_3__9399_ (
);

FILL FILL_4__10764_ (
);

FILL SFILL13800x76050 (
);

FILL FILL_1__15656_ (
);

FILL FILL_1__15236_ (
);

FILL FILL_3_BUFX2_insert0 (
);

FILL FILL_1__10791_ (
);

FILL FILL_3_BUFX2_insert1 (
);

FILL FILL_1__10371_ (
);

FILL FILL_3_BUFX2_insert2 (
);

FILL FILL_3_BUFX2_insert3 (
);

FILL FILL_3_BUFX2_insert4 (
);

OAI22X1 _14934_ (
    .A(_5414_),
    .B(_3936__bF$buf4),
    .C(_3944__bF$buf4),
    .D(_5413_),
    .Y(_5415_)
);

FILL FILL_0__14649_ (
);

FILL FILL_0__14229_ (
);

INVX1 _14514_ (
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_5004_)
);

FILL FILL_3_BUFX2_insert5 (
);

FILL FILL_3_BUFX2_insert6 (
);

FILL FILL_3_BUFX2_insert7 (
);

FILL FILL_3_BUFX2_insert8 (
);

FILL FILL_3_BUFX2_insert9 (
);

FILL SFILL53960x29050 (
);

FILL FILL_5__12976_ (
);

FILL FILL_3__13590_ (
);

FILL FILL_5__12136_ (
);

BUFX2 _6856_ (
    .A(_1_[18]),
    .Y(memoryAddress[18])
);

FILL FILL_3__13170_ (
);

FILL FILL_4__11969_ (
);

FILL FILL_4__8263_ (
);

FILL FILL_4__11549_ (
);

FILL FILL_2__12583_ (
);

FILL FILL_4__11129_ (
);

FILL FILL_2__12163_ (
);

FILL FILL_1__11996_ (
);

FILL FILL_1__11576_ (
);

FILL FILL_1__11156_ (
);

NOR3X1 _15719_ (
    .A(_6182_),
    .B(_6179_),
    .C(_6181_),
    .Y(_6183_)
);

FILL FILL_4__12910_ (
);

FILL SFILL74040x42050 (
);

FILL FILL_0__10989_ (
);

FILL FILL_0__8583_ (
);

DFFSR _10854_ (
    .Q(\datapath_1.regfile_1.regOut[31] [16]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_1953_[16])
);

FILL FILL_0__10569_ (
);

FILL FILL_0__10149_ (
);

NAND2X1 _10434_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1808_)
);

NAND2X1 _10014_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1589_)
);

FILL FILL_3__11903_ (
);

FILL FILL_4__15382_ (
);

FILL FILL_3__14795_ (
);

FILL FILL_0__11930_ (
);

FILL FILL_2__9542_ (
);

FILL FILL_2__9122_ (
);

FILL FILL_3__14375_ (
);

FILL FILL_0__11510_ (
);

FILL SFILL3640x50 (
);

FILL FILL_4__9888_ (
);

FILL FILL_4__9468_ (
);

FILL FILL112360x76050 (
);

FILL FILL_2__13788_ (
);

FILL FILL_2__13368_ (
);

FILL FILL_5__14702_ (
);

FILL FILL_3__7885_ (
);

FILL FILL_0__9788_ (
);

FILL FILL_0__9368_ (
);

FILL FILL_3__7465_ (
);

FILL FILL_3__7045_ (
);

AOI21X1 _11639_ (
    .A(_2502_),
    .B(_2496_),
    .C(_2174_),
    .Y(_2742_)
);

AOI21X1 _11219_ (
    .A(_2111_),
    .B(_2332_),
    .C(_2337_),
    .Y(_2338_)
);

FILL FILL_1__13722_ (
);

FILL FILL_1__13302_ (
);

FILL FILL_4__16167_ (
);

FILL FILL_0__12715_ (
);

FILL FILL_1__16194_ (
);

FILL FILL_5__8752_ (
);

FILL FILL_5__8332_ (
);

FILL FILL_3__10295_ (
);

NAND2X1 _15892_ (
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .B(_5693_),
    .Y(_6351_)
);

FILL FILL_0__15187_ (
);

NAND3X1 _15472_ (
    .A(_5937_),
    .B(_5938_),
    .C(_5941_),
    .Y(_5942_)
);

FILL FILL_5__15907_ (
);

NAND2X1 _15052_ (
    .A(_5465_),
    .B(_5531__bF$buf1),
    .Y(_5532_)
);

FILL SFILL104200x23050 (
);

FILL FILL112360x31050 (
);

FILL FILL_3__16101_ (
);

FILL FILL_1__8744_ (
);

FILL FILL_5__10622_ (
);

FILL FILL_1__8324_ (
);

FILL FILL_2__15934_ (
);

FILL FILL_2__15514_ (
);

FILL SFILL64040x40050 (
);

FILL FILL_5__13094_ (
);

FILL FILL_1__14927_ (
);

FILL FILL_1__14507_ (
);

DFFSR _7394_ (
    .Q(\datapath_1.regfile_1.regOut[4] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_198_[12])
);

FILL FILL_4__12087_ (
);

FILL FILL_3__9611_ (
);

FILL FILL112280x38050 (
);

FILL FILL_5__9537_ (
);

FILL FILL_5__9117_ (
);

NOR2X1 _16257_ (
    .A(_6706_),
    .B(_6704_),
    .Y(_6707_)
);

FILL SFILL24680x34050 (
);

OAI21X1 _11392_ (
    .A(_2168_),
    .B(_2198_),
    .C(_2508_),
    .Y(_2509_)
);

FILL FILL_5__11827_ (
);

FILL FILL_1__9529_ (
);

FILL FILL_3__12861_ (
);

FILL FILL_5__11407_ (
);

FILL FILL_3__12441_ (
);

FILL FILL_1__9109_ (
);

FILL FILL_3__12021_ (
);

FILL FILL_4__7954_ (
);

FILL FILL_4__7114_ (
);

FILL FILL_2__11854_ (
);

FILL FILL_5__14299_ (
);

FILL FILL_2__11434_ (
);

FILL SFILL54040x83050 (
);

FILL FILL_2__11014_ (
);

INVX1 _8599_ (
    .A(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_869_)
);

DFFSR _8179_ (
    .Q(\datapath_1.regfile_1.regOut[10] [29]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_588_[29])
);

FILL FILL_1__10427_ (
);

FILL FILL_1__10007_ (
);

FILL FILL_5__15660_ (
);

FILL FILL_5__15240_ (
);

FILL FILL_0__7854_ (
);

FILL FILL_0__7434_ (
);

DFFSR _9960_ (
    .Q(\datapath_1.regfile_1.regOut[24] [18]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_1498_[18])
);

INVX1 _9540_ (
    .A(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_1354_)
);

INVX1 _9120_ (
    .A(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_1135_)
);

FILL FILL_4__14653_ (
);

FILL FILL_4__14233_ (
);

INVX1 _12597_ (
    .A(\datapath_1.Data [10]),
    .Y(_3444_)
);

OAI21X1 _12177_ (
    .A(_3170_),
    .B(ALUSrcA_bF$buf3),
    .C(_3171_),
    .Y(\datapath_1.alu_1.ALUInA [20])
);

FILL FILL_3__13646_ (
);

FILL FILL_3__13226_ (
);

FILL FILL_1__14680_ (
);

FILL FILL_1__14260_ (
);

FILL FILL_4__8739_ (
);

FILL FILL_0_BUFX2_insert400 (
);

FILL FILL_4__8319_ (
);

FILL FILL_0_BUFX2_insert401 (
);

FILL FILL_0_BUFX2_insert402 (
);

FILL FILL_2__12639_ (
);

FILL FILL_0_BUFX2_insert403 (
);

FILL FILL_0_BUFX2_insert404 (
);

FILL FILL_0__13673_ (
);

FILL FILL_2__12219_ (
);

FILL FILL_0__13253_ (
);

FILL FILL_0_BUFX2_insert405 (
);

FILL FILL_0_BUFX2_insert406 (
);

FILL FILL_0_BUFX2_insert407 (
);

FILL FILL_0_BUFX2_insert408 (
);

FILL FILL_0_BUFX2_insert409 (
);

FILL FILL_5__9290_ (
);

FILL FILL_0__8639_ (
);

FILL FILL_5__16025_ (
);

FILL FILL_0__8219_ (
);

FILL FILL_5__11580_ (
);

FILL FILL_1__9282_ (
);

FILL FILL_5__11160_ (
);

FILL FILL_4__15858_ (
);

FILL FILL_4__15438_ (
);

FILL FILL_4__15018_ (
);

FILL FILL_2__16052_ (
);

FILL FILL_4__10993_ (
);

FILL FILL_4__10573_ (
);

FILL FILL_4__10153_ (
);

FILL FILL_1__15885_ (
);

FILL FILL_1__15465_ (
);

FILL FILL_1__15045_ (
);

FILL FILL_5__7603_ (
);

FILL FILL_1__10180_ (
);

FILL FILL_6__10900_ (
);

FILL FILL_0__14878_ (
);

FILL FILL_0__14458_ (
);

INVX1 _14743_ (
    .A(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_5228_)
);

FILL FILL_0__14038_ (
);

AOI22X1 _14323_ (
    .A(\datapath_1.regfile_1.regOut[11] [18]),
    .B(_3950__bF$buf2),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_4817_)
);

FILL SFILL44040x81050 (
);

FILL FILL_6__13792_ (
);

FILL FILL_6__13372_ (
);

FILL FILL_5__12785_ (
);

FILL FILL_5__12365_ (
);

FILL FILL_4__8492_ (
);

FILL FILL_4__8072_ (
);

FILL FILL_4__11778_ (
);

FILL FILL_4__11358_ (
);

FILL FILL_2__12392_ (
);

FILL FILL_1__11385_ (
);

OAI22X1 _15948_ (
    .A(_5480__bF$buf2),
    .B(_4994_),
    .C(_6405_),
    .D(_5499__bF$buf3),
    .Y(_6406_)
);

NOR2X1 _15528_ (
    .A(_5996_),
    .B(_5993_),
    .Y(_5997_)
);

OAI22X1 _15108_ (
    .A(_5478__bF$buf2),
    .B(_5586_),
    .C(_5552__bF$buf3),
    .D(_4026_),
    .Y(_5587_)
);

FILL FILL_0__10798_ (
);

FILL FILL_0__8392_ (
);

NAND2X1 _10663_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1920_)
);

FILL FILL_0__10378_ (
);

NAND2X1 _10243_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1701_)
);

FILL FILL_3__11712_ (
);

FILL FILL_4__15191_ (
);

FILL FILL_2__10705_ (
);

FILL FILL_2__9771_ (
);

FILL FILL112440x7050 (
);

FILL FILL_2__9351_ (
);

FILL FILL_3__14184_ (
);

FILL FILL_4_BUFX2_insert980 (
);

FILL FILL_4_BUFX2_insert981 (
);

FILL FILL_4__9277_ (
);

FILL FILL_4_BUFX2_insert982 (
);

FILL FILL_4_BUFX2_insert983 (
);

FILL FILL_2__13597_ (
);

FILL FILL_4_BUFX2_insert984 (
);

FILL FILL_4_BUFX2_insert985 (
);

FILL FILL_4_BUFX2_insert986 (
);

FILL FILL_5__14931_ (
);

FILL FILL_4_BUFX2_insert987 (
);

FILL FILL112120x1050 (
);

FILL FILL_4_BUFX2_insert988 (
);

FILL FILL_5__14511_ (
);

FILL FILL_4_BUFX2_insert989 (
);

DFFSR _8811_ (
    .Q(\datapath_1.regfile_1.regOut[15] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_913_[21])
);

FILL FILL112040x6050 (
);

FILL FILL_4__13924_ (
);

FILL FILL_4__13504_ (
);

FILL FILL_3__7694_ (
);

FILL FILL_0__9597_ (
);

AND2X2 _11868_ (
    .A(_2953_),
    .B(_2954_),
    .Y(_2955_)
);

FILL SFILL23800x28050 (
);

AND2X2 _11448_ (
    .A(_2379_),
    .B(_2382_),
    .Y(_2564_)
);

AOI21X1 _11028_ (
    .A(_2125_),
    .B(_2135_),
    .C(_2146_),
    .Y(_2147_)
);

FILL FILL_3__12917_ (
);

FILL FILL_1__13951_ (
);

FILL FILL_1__13531_ (
);

FILL FILL_4__16396_ (
);

FILL FILL_1__13111_ (
);

FILL FILL_6__10497_ (
);

FILL FILL_3__15389_ (
);

FILL FILL_0__12524_ (
);

FILL FILL_0__12104_ (
);

FILL FILL_5__8981_ (
);

FILL SFILL109720x44050 (
);

FILL SFILL74120x75050 (
);

FILL SFILL74200x9050 (
);

FILL FILL_5__8141_ (
);

NAND3X1 _15281_ (
    .A(\datapath_1.regfile_1.regOut[20] [5]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf3),
    .Y(_5756_)
);

FILL FILL_5__15716_ (
);

FILL FILL_3__16330_ (
);

FILL FILL_1__8973_ (
);

FILL FILL_5__10431_ (
);

FILL FILL_5__10011_ (
);

FILL FILL_1__8133_ (
);

FILL FILL_4__14709_ (
);

FILL FILL_2__15743_ (
);

FILL FILL_2__15323_ (
);

FILL FILL_3__8899_ (
);

FILL FILL_3__8479_ (
);

FILL FILL_3__8059_ (
);

FILL FILL_1__14736_ (
);

FILL FILL_1__14316_ (
);

FILL FILL_3__9420_ (
);

FILL FILL_0__13729_ (
);

FILL FILL_0__13309_ (
);

FILL FILL_3__9000_ (
);

FILL FILL_2__6896_ (
);

FILL FILL_5__9766_ (
);

FILL FILL_5__9346_ (
);

NAND3X1 _16066_ (
    .A(_6515_),
    .B(_6516_),
    .C(_6520_),
    .Y(_6521_)
);

FILL SFILL74120x30050 (
);

FILL FILL_1__9758_ (
);

FILL FILL_5__11636_ (
);

FILL FILL_5__11216_ (
);

FILL FILL_1__9338_ (
);

FILL FILL_3__12250_ (
);

FILL FILL_4__7763_ (
);

FILL FILL_2__16108_ (
);

FILL FILL_4__7343_ (
);

FILL FILL_4__10629_ (
);

FILL FILL_2__11663_ (
);

FILL FILL_2__11243_ (
);

FILL FILL_6__7689_ (
);

FILL SFILL13800x26050 (
);

FILL FILL_1__10656_ (
);

FILL FILL_1__10236_ (
);

FILL FILL_0__7243_ (
);

FILL FILL_6__13848_ (
);

FILL FILL_6__13428_ (
);

FILL FILL_4__14882_ (
);

FILL FILL_4__14462_ (
);

FILL FILL_4__14042_ (
);

FILL SFILL64120x73050 (
);

FILL FILL_3__13875_ (
);

FILL FILL_2__8622_ (
);

FILL FILL_2__8202_ (
);

FILL FILL_3__13455_ (
);

FILL FILL_3__13035_ (
);

FILL FILL_4__8968_ (
);

FILL FILL_4__8128_ (
);

FILL FILL_2__12868_ (
);

FILL FILL_2__12448_ (
);

FILL FILL_2__12028_ (
);

FILL FILL_0__13482_ (
);

FILL SFILL68440x81050 (
);

FILL FILL_0__8868_ (
);

FILL FILL_3__6965_ (
);

FILL FILL_5__16254_ (
);

FILL FILL_0__8448_ (
);

FILL FILL_6__9415_ (
);

DFFSR _10719_ (
    .Q(\datapath_1.regfile_1.regOut[30] [9]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_1888_[9])
);

FILL FILL_1__9091_ (
);

FILL FILL_4__15667_ (
);

FILL FILL_4__15247_ (
);

FILL FILL_2__16281_ (
);

FILL FILL_4__10382_ (
);

FILL FILL_2__9407_ (
);

FILL FILL_1__15694_ (
);

FILL FILL_1__15274_ (
);

FILL FILL_5__7832_ (
);

INVX1 _14972_ (
    .A(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_5453_)
);

FILL FILL_0__14687_ (
);

OAI22X1 _14552_ (
    .A(_5040_),
    .B(_3972__bF$buf0),
    .C(_3920_),
    .D(_5039_),
    .Y(_5041_)
);

FILL FILL_0__14267_ (
);

AOI22X1 _14132_ (
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_4630_)
);

FILL FILL112360x26050 (
);

FILL SFILL85080x9050 (
);

FILL FILL_3__15601_ (
);

FILL FILL_1__7824_ (
);

FILL SFILL64040x35050 (
);

FILL FILL_5__12594_ (
);

FILL FILL_5__12174_ (
);

BUFX2 _6894_ (
    .A(_2_[24]),
    .Y(memoryWriteData[24])
);

FILL FILL_4__11587_ (
);

FILL FILL_4__11167_ (
);

FILL FILL_1__16059_ (
);

FILL FILL_5__8617_ (
);

FILL FILL_1__11194_ (
);

FILL SFILL9320x50050 (
);

FILL SFILL83720x8050 (
);

NOR2X1 _15757_ (
    .A(_6219_),
    .B(_6217_),
    .Y(_6220_)
);

NOR2X1 _15337_ (
    .A(_5798_),
    .B(_5810_),
    .Y(_5811_)
);

NOR3X1 _10892_ (
    .A(\aluControl_1.inst [0]),
    .B(_2030_),
    .C(_2032_),
    .Y(_2038_)
);

FILL FILL_0__10187_ (
);

DFFSR _10472_ (
    .Q(\datapath_1.regfile_1.regOut[28] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1758_[18])
);

FILL FILL_5__10907_ (
);

INVX1 _10052_ (
    .A(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_1614_)
);

FILL FILL_1__8609_ (
);

FILL FILL_3__11941_ (
);

FILL FILL_3__11521_ (
);

FILL FILL_3__11101_ (
);

FILL FILL_0__16413_ (
);

FILL SFILL89640x53050 (
);

FILL FILL_5__13799_ (
);

FILL FILL_2__10934_ (
);

FILL FILL_5__13379_ (
);

FILL FILL_2__10514_ (
);

FILL FILL_2__9160_ (
);

INVX1 _7679_ (
    .A(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_398_)
);

DFFSR _7259_ (
    .Q(\datapath_1.regfile_1.regOut[3] [5]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_133_[5])
);

FILL FILL_4__9086_ (
);

FILL FILL_5__14740_ (
);

FILL FILL_5__14320_ (
);

FILL FILL_0__6934_ (
);

INVX1 _8620_ (
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_883_)
);

INVX1 _8200_ (
    .A(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_664_)
);

FILL FILL_1__12399_ (
);

FILL FILL_4__13733_ (
);

FILL FILL_4__13313_ (
);

FILL FILL_3__7083_ (
);

OAI21X1 _11677_ (
    .A(_2182_),
    .B(_2183_),
    .C(_2777_),
    .Y(_2778_)
);

AOI21X1 _11257_ (
    .A(_2370_),
    .B(_2363_),
    .C(_2375_),
    .Y(_2376_)
);

FILL FILL_3__12726_ (
);

FILL FILL_1__13760_ (
);

FILL FILL_3__12306_ (
);

FILL FILL_1__13340_ (
);

FILL FILL_4__7819_ (
);

FILL FILL_2__11719_ (
);

FILL FILL_0__12753_ (
);

FILL FILL_3__15198_ (
);

FILL FILL_0__12333_ (
);

FILL SFILL54040x33050 (
);

FILL FILL_5__8370_ (
);

NAND3X1 _15090_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5468_),
    .C(_5465_),
    .Y(_5569_)
);

FILL FILL_5__15945_ (
);

FILL FILL_5__15525_ (
);

FILL FILL_0__7719_ (
);

FILL FILL_5__15105_ (
);

DFFSR _9825_ (
    .Q(\datapath_1.regfile_1.regOut[23] [11]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1433_[11])
);

OAI21X1 _9405_ (
    .A(_1283_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .C(_1284_),
    .Y(_1238_[23])
);

FILL SFILL79240x82050 (
);

FILL FILL_5__10660_ (
);

FILL FILL_1__8782_ (
);

FILL FILL_5__10240_ (
);

FILL FILL_1__8362_ (
);

FILL FILL_4__14938_ (
);

FILL FILL_2__15972_ (
);

FILL FILL_4__14518_ (
);

FILL FILL_2__15552_ (
);

FILL FILL_2__15132_ (
);

FILL FILL_1__14965_ (
);

FILL FILL_1__14545_ (
);

FILL FILL_1__14125_ (
);

FILL FILL_0__13958_ (
);

INVX1 _13823_ (
    .A(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_4328_)
);

FILL FILL_0__13538_ (
);

INVX1 _13403_ (
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_3915_)
);

FILL FILL_0__13118_ (
);

FILL FILL_5__9995_ (
);

FILL FILL_5__9155_ (
);

FILL FILL_6__12872_ (
);

NAND3X1 _16295_ (
    .A(_6741_),
    .B(_6743_),
    .C(_6742_),
    .Y(_6744_)
);

FILL FILL_1__9987_ (
);

FILL FILL_5__11865_ (
);

FILL FILL_5__11445_ (
);

FILL FILL_1__9147_ (
);

FILL FILL_5__11025_ (
);

FILL FILL_4__7992_ (
);

FILL FILL_2__16337_ (
);

FILL FILL_4__7572_ (
);

FILL FILL_4__10438_ (
);

FILL FILL_2__11892_ (
);

FILL FILL_4__10018_ (
);

FILL FILL_2__11472_ (
);

FILL FILL_2__11052_ (
);

FILL FILL_1__10885_ (
);

FILL FILL_1__10045_ (
);

AOI22X1 _14608_ (
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .B(_4079__bF$buf1),
    .C(_4038__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_5096_)
);

FILL FILL_0__7892_ (
);

FILL FILL_0__7472_ (
);

FILL FILL_0__7052_ (
);

FILL FILL_4__14691_ (
);

FILL FILL_4__14271_ (
);

FILL SFILL53800x2050 (
);

FILL FILL_2__8851_ (
);

FILL SFILL54040x4050 (
);

FILL FILL_3__13684_ (
);

FILL SFILL53720x7050 (
);

FILL FILL_3__13264_ (
);

FILL FILL_2__8011_ (
);

FILL SFILL94280x2050 (
);

FILL FILL_4__8777_ (
);

FILL FILL_4__8357_ (
);

FILL FILL_2__12257_ (
);

FILL FILL_0__13291_ (
);

FILL FILL_5__16063_ (
);

NAND2X1 _10948_ (
    .A(_2064_),
    .B(_2080_),
    .Y(_2081_)
);

FILL FILL_0__8257_ (
);

FILL FILL_6__9224_ (
);

INVX1 _10528_ (
    .A(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_1850_)
);

INVX1 _10108_ (
    .A(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_1631_)
);

FILL FILL_4__15896_ (
);

FILL FILL_1__12611_ (
);

FILL FILL_4__15476_ (
);

FILL FILL_4__15056_ (
);

FILL FILL_2__16090_ (
);

FILL SFILL104440x5050 (
);

FILL FILL_4__10191_ (
);

FILL FILL_2__9636_ (
);

FILL FILL_3__14889_ (
);

FILL FILL_2__9216_ (
);

FILL FILL_3__14469_ (
);

FILL FILL_0__11604_ (
);

FILL FILL_3__14049_ (
);

FILL FILL_1__15083_ (
);

FILL FILL_5__7221_ (
);

FILL FILL_0__14496_ (
);

OAI22X1 _14781_ (
    .A(_3909_),
    .B(_5265_),
    .C(_5264_),
    .D(_3944__bF$buf4),
    .Y(_5266_)
);

INVX1 _14361_ (
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_4854_)
);

FILL FILL_0__14076_ (
);

FILL FILL_3__15830_ (
);

FILL FILL_3__15410_ (
);

FILL FILL_1__7633_ (
);

FILL FILL_1__7213_ (
);

FILL FILL_2__14823_ (
);

FILL FILL_2__14403_ (
);

FILL FILL_3__7979_ (
);

FILL FILL_3__7559_ (
);

FILL FILL_1__13816_ (
);

FILL SFILL74520x39050 (
);

FILL SFILL43880x50 (
);

FILL FILL_4__11396_ (
);

FILL SFILL38760x51050 (
);

FILL SFILL69160x42050 (
);

FILL FILL_3__8500_ (
);

FILL FILL_1__16288_ (
);

FILL FILL_5__8846_ (
);

FILL FILL_3__10389_ (
);

FILL FILL_5__8006_ (
);

OAI22X1 _15986_ (
    .A(_5065_),
    .B(_5501_),
    .C(_5524__bF$buf3),
    .D(_5078_),
    .Y(_6443_)
);

INVX1 _15566_ (
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_6034_)
);

FILL FILL_6__11303_ (
);

NAND3X1 _15146_ (
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf1),
    .Y(_5624_)
);

INVX1 _10281_ (
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_1726_)
);

FILL FILL_1__8838_ (
);

FILL FILL_3__11750_ (
);

FILL FILL_3__11330_ (
);

FILL FILL_2__15608_ (
);

FILL FILL_4__6843_ (
);

FILL SFILL38680x58050 (
);

FILL FILL_0__16222_ (
);

FILL FILL_2__10743_ (
);

FILL FILL_2__10323_ (
);

OAI21X1 _7488_ (
    .A(_310_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .C(_311_),
    .Y(_263_[24])
);

OAI21X1 _7068_ (
    .A(_91_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_92_),
    .Y(_68_[12])
);

FILL FILL_6__7710_ (
);

FILL FILL_4__13962_ (
);

FILL FILL_4__13542_ (
);

FILL SFILL64120x68050 (
);

FILL FILL_4__13122_ (
);

FILL SFILL95000x21050 (
);

NAND3X1 _11486_ (
    .A(_2289_),
    .B(_2446_),
    .C(_2590_),
    .Y(_2600_)
);

NOR2X1 _11066_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2185_)
);

FILL FILL_3__12955_ (
);

FILL FILL_2__7702_ (
);

FILL FILL_3__12115_ (
);

FILL FILL_4__7628_ (
);

FILL FILL_4__7208_ (
);

FILL FILL_2__11948_ (
);

FILL FILL_0__12982_ (
);

FILL FILL_2__11528_ (
);

FILL SFILL68440x76050 (
);

FILL FILL_2__11108_ (
);

FILL FILL_0__12142_ (
);

FILL SFILL89320x3050 (
);

FILL SFILL23800x1050 (
);

FILL SFILL23720x6050 (
);

FILL FILL_5__15754_ (
);

FILL FILL_0__7948_ (
);

FILL FILL_5__15334_ (
);

OAI21X1 _9634_ (
    .A(_1395_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1396_),
    .Y(_1368_[14])
);

FILL FILL_0__7108_ (
);

FILL SFILL59160x40050 (
);

OAI21X1 _9214_ (
    .A(_1176_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .C(_1177_),
    .Y(_1173_[2])
);

FILL FILL_1__8591_ (
);

FILL SFILL63880x9050 (
);

FILL FILL_4__14747_ (
);

FILL FILL_2__15781_ (
);

FILL FILL_4__14327_ (
);

FILL FILL_2__15361_ (
);

FILL FILL_3__8097_ (
);

FILL FILL_2__8907_ (
);

FILL SFILL64120x23050 (
);

FILL SFILL3640x2050 (
);

FILL FILL_1__14774_ (
);

FILL FILL_1__14354_ (
);

FILL FILL_5__6912_ (
);

FILL FILL_0__13767_ (
);

INVX1 _13632_ (
    .A(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_4141_)
);

FILL FILL_0__13347_ (
);

FILL SFILL89320x72050 (
);

AND2X2 _13212_ (
    .A(_3752_),
    .B(_3754_),
    .Y(_3755_)
);

FILL FILL_5__9384_ (
);

FILL FILL_1__6904_ (
);

FILL SFILL113800x77050 (
);

FILL FILL_5__16119_ (
);

FILL FILL_1__9796_ (
);

FILL FILL_5__11674_ (
);

FILL FILL_1__9376_ (
);

FILL FILL_5__11254_ (
);

FILL FILL_2__16146_ (
);

FILL FILL_4__7381_ (
);

FILL FILL_4__10667_ (
);

FILL FILL_4__10247_ (
);

FILL FILL_2__11281_ (
);

FILL FILL_1__15979_ (
);

FILL FILL_1__15559_ (
);

FILL FILL_1__15139_ (
);

FILL FILL_1__10694_ (
);

FILL FILL_2_BUFX2_insert310 (
);

FILL FILL_1__10274_ (
);

FILL FILL_2_BUFX2_insert311 (
);

FILL FILL_2_BUFX2_insert312 (
);

NOR2X1 _14837_ (
    .A(_5319_),
    .B(_3935__bF$buf4),
    .Y(_5320_)
);

FILL FILL_2_BUFX2_insert313 (
);

FILL FILL_2_BUFX2_insert314 (
);

OAI22X1 _14417_ (
    .A(_3916_),
    .B(_4907_),
    .C(_3977__bF$buf2),
    .D(_4908_),
    .Y(_4909_)
);

FILL FILL_2_BUFX2_insert315 (
);

FILL FILL_2_BUFX2_insert316 (
);

FILL FILL_2__7299_ (
);

FILL FILL_2_BUFX2_insert317 (
);

FILL FILL_2_BUFX2_insert318 (
);

FILL FILL_2_BUFX2_insert319 (
);

FILL FILL_4__14080_ (
);

FILL FILL_0__15913_ (
);

FILL FILL_5__12879_ (
);

FILL FILL_5__12459_ (
);

FILL FILL_2__8660_ (
);

FILL FILL_5__12039_ (
);

FILL FILL_2__8240_ (
);

FILL FILL_3__13493_ (
);

FILL FILL_4__8586_ (
);

FILL FILL_2__12486_ (
);

FILL FILL_2__12066_ (
);

FILL FILL_5__13820_ (
);

FILL FILL_5__13400_ (
);

FILL FILL_2_BUFX2_insert1030 (
);

FILL SFILL58840x43050 (
);

FILL FILL_2_BUFX2_insert1031 (
);

FILL SFILL89240x34050 (
);

FILL FILL_2_BUFX2_insert1032 (
);

FILL FILL_1__11899_ (
);

INVX1 _7700_ (
    .A(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_412_)
);

FILL SFILL54120x21050 (
);

FILL FILL_2_BUFX2_insert1033 (
);

FILL FILL_1__11479_ (
);

FILL FILL_2_BUFX2_insert1034 (
);

FILL FILL_1__11059_ (
);

FILL FILL_2_BUFX2_insert1035 (
);

FILL FILL_2_BUFX2_insert1036 (
);

FILL FILL_2_BUFX2_insert1037 (
);

FILL FILL_2_BUFX2_insert1038 (
);

FILL FILL_5__16292_ (
);

FILL FILL_2_BUFX2_insert1039 (
);

FILL FILL_0__8486_ (
);

FILL FILL_0__8066_ (
);

INVX1 _10757_ (
    .A(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_1962_)
);

DFFSR _10337_ (
    .Q(\datapath_1.regfile_1.regOut[27] [11]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1693_[11])
);

FILL FILL_3__11806_ (
);

FILL SFILL18680x54050 (
);

FILL FILL_1__12840_ (
);

FILL FILL_1__12420_ (
);

FILL FILL_4__15285_ (
);

FILL FILL_1__12000_ (
);

FILL FILL_2__9865_ (
);

FILL FILL_3__14698_ (
);

FILL FILL_0__11833_ (
);

FILL FILL_3__14278_ (
);

FILL FILL_0__11413_ (
);

FILL FILL_2__9025_ (
);

FILL FILL_5__7870_ (
);

FILL FILL_5__7450_ (
);

FILL FILL_5__7030_ (
);

OAI22X1 _14590_ (
    .A(_3978_),
    .B(_5077_),
    .C(_3977__bF$buf1),
    .D(_5078_),
    .Y(_5079_)
);

NOR2X1 _14170_ (
    .A(_4667_),
    .B(_4652_),
    .Y(_4668_)
);

FILL FILL_5__14605_ (
);

OAI21X1 _8905_ (
    .A(_1031_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .C(_1032_),
    .Y(_978_[27])
);

FILL FILL_1__7862_ (
);

FILL FILL_1__7442_ (
);

FILL FILL_2__14632_ (
);

FILL FILL_2__14212_ (
);

FILL FILL_3__7368_ (
);

FILL FILL_1__13625_ (
);

FILL FILL_1_BUFX2_insert330 (
);

FILL FILL_1_BUFX2_insert331 (
);

FILL SFILL33880x8050 (
);

FILL FILL_0__12618_ (
);

OAI21X1 _12903_ (
    .A(_3606_),
    .B(vdd),
    .C(_3607_),
    .Y(_3555_[26])
);

FILL FILL_1_BUFX2_insert332 (
);

FILL FILL_1_BUFX2_insert333 (
);

FILL FILL_1_BUFX2_insert334 (
);

FILL FILL_1__16097_ (
);

FILL FILL_1_BUFX2_insert335 (
);

FILL FILL_5__8655_ (
);

FILL FILL_1_BUFX2_insert336 (
);

FILL FILL_5__8235_ (
);

FILL FILL_1_BUFX2_insert337 (
);

FILL FILL_1_BUFX2_insert338 (
);

FILL FILL_6__11952_ (
);

FILL FILL_1_BUFX2_insert339 (
);

FILL FILL_6_BUFX2_insert894 (
);

OAI21X1 _15795_ (
    .A(_4809_),
    .B(_5535__bF$buf1),
    .C(_6256_),
    .Y(_6257_)
);

NOR2X1 _15375_ (
    .A(_4379_),
    .B(_5549__bF$buf2),
    .Y(_5847_)
);

FILL FILL_3__16004_ (
);

FILL FILL_6_BUFX2_insert899 (
);

FILL FILL_5__10945_ (
);

DFFSR _10090_ (
    .Q(\datapath_1.regfile_1.regOut[25] [20]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_1563_[20])
);

FILL FILL_1__8647_ (
);

FILL FILL_5__10525_ (
);

FILL FILL_1__8227_ (
);

FILL FILL_5__10105_ (
);

FILL FILL_2__15837_ (
);

FILL SFILL79240x32050 (
);

FILL FILL_2__15417_ (
);

FILL FILL_0__16451_ (
);

FILL FILL_0__16031_ (
);

FILL FILL_2__10972_ (
);

FILL FILL_2__10552_ (
);

FILL FILL_2__10132_ (
);

OAI21X1 _7297_ (
    .A(_203_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .C(_204_),
    .Y(_198_[3])
);

FILL FILL_3__9934_ (
);

FILL FILL_3__9514_ (
);

FILL FILL_0__6972_ (
);

FILL FILL_4__13771_ (
);

FILL FILL_4__13351_ (
);

INVX1 _11295_ (
    .A(_2413_),
    .Y(_2414_)
);

FILL FILL_2__7931_ (
);

FILL FILL_3__12764_ (
);

FILL FILL_3__12344_ (
);

FILL SFILL69240x75050 (
);

FILL FILL_4__7857_ (
);

FILL FILL_4__7437_ (
);

FILL FILL_2__11757_ (
);

FILL FILL_2__11337_ (
);

FILL FILL_0__12371_ (
);

FILL FILL_6__16150_ (
);

FILL FILL_5__15983_ (
);

FILL FILL_5__15563_ (
);

FILL FILL_0__7757_ (
);

FILL FILL_5__15143_ (
);

FILL FILL_0__7337_ (
);

OAI21X1 _9863_ (
    .A(_1507_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .C(_1508_),
    .Y(_1498_[5])
);

DFFSR _9443_ (
    .Q(\datapath_1.regfile_1.regOut[20] [13]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_1238_[13])
);

NAND2X1 _9023_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1091_)
);

FILL FILL_4__14976_ (
);

FILL FILL_4__14556_ (
);

FILL FILL_4__14136_ (
);

FILL FILL_2__15590_ (
);

FILL FILL_2__15170_ (
);

FILL SFILL109400x13050 (
);

FILL FILL_2__8716_ (
);

FILL FILL_3__13969_ (
);

FILL FILL_3__13549_ (
);

FILL FILL_1__14583_ (
);

FILL FILL_3__13129_ (
);

FILL FILL_1__14163_ (
);

FILL FILL_0__13996_ (
);

NOR2X1 _13861_ (
    .A(_4364_),
    .B(_4361_),
    .Y(_4365_)
);

FILL FILL_0__13576_ (
);

FILL SFILL69240x30050 (
);

INVX1 _13441_ (
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_3953_)
);

FILL FILL_0__13156_ (
);

NAND2X1 _13021_ (
    .A(vdd),
    .B(\datapath_1.rd2 [23]),
    .Y(_3666_)
);

FILL FILL_3__14910_ (
);

FILL FILL_6__12490_ (
);

FILL FILL_6__12070_ (
);

FILL FILL_2__13903_ (
);

FILL FILL_5__16348_ (
);

FILL FILL_5__11483_ (
);

FILL FILL_5__11063_ (
);

FILL FILL_2__16375_ (
);

FILL SFILL99400x62050 (
);

FILL FILL_4__10896_ (
);

FILL FILL_4__7190_ (
);

FILL SFILL38760x46050 (
);

FILL SFILL69160x37050 (
);

FILL FILL_0__9903_ (
);

FILL FILL_4__10056_ (
);

FILL FILL_2__11090_ (
);

FILL FILL_1__15788_ (
);

FILL FILL_1__15368_ (
);

FILL FILL_5__7926_ (
);

FILL FILL_5__7506_ (
);

NOR2X1 _14646_ (
    .A(_5133_),
    .B(_5118_),
    .Y(_5134_)
);

AOI22X1 _14226_ (
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .B(_3942__bF$buf1),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_4722_)
);

FILL SFILL28920x9050 (
);

FILL FILL_0__7090_ (
);

FILL FILL_3__10830_ (
);

FILL FILL_6__13275_ (
);

FILL FILL_3__10410_ (
);

FILL SFILL99320x69050 (
);

FILL FILL_0__15722_ (
);

FILL FILL_0__15302_ (
);

FILL FILL_5__12268_ (
);

OAI21X1 _6988_ (
    .A(_58_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_59_),
    .Y(_3_[28])
);

FILL SFILL3800x50050 (
);

FILL SFILL69080x3050 (
);

FILL FILL_4__8395_ (
);

FILL FILL_2__12295_ (
);

FILL SFILL24040x67050 (
);

FILL FILL_1__11288_ (
);

FILL FILL_4__12622_ (
);

FILL FILL_4__12202_ (
);

DFFSR _10986_ (
    .Q(\control_1.reg_state.dout [2]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_2098_[2])
);

OAI21X1 _10566_ (
    .A(_1874_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .C(_1875_),
    .Y(_1823_[26])
);

OAI21X1 _10146_ (
    .A(_1655_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1656_),
    .Y(_1628_[14])
);

FILL FILL_3__11615_ (
);

FILL FILL_4__15094_ (
);

FILL FILL_2__9674_ (
);

FILL SFILL99320x24050 (
);

FILL FILL_2__9254_ (
);

FILL FILL_0__11642_ (
);

FILL FILL_0__11222_ (
);

FILL FILL_3__14087_ (
);

FILL FILL_5__14834_ (
);

FILL SFILL89400x60050 (
);

FILL FILL_5__14414_ (
);

OAI21X1 _8714_ (
    .A(_924_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_925_),
    .Y(_913_[6])
);

FILL FILL_1__7671_ (
);

FILL FILL_1__7251_ (
);

FILL FILL_4__13827_ (
);

FILL FILL_2__14861_ (
);

FILL FILL_4__13407_ (
);

FILL FILL_2__14441_ (
);

FILL FILL_2__14021_ (
);

FILL FILL_3__7597_ (
);

FILL FILL_3__7177_ (
);

FILL SFILL64120x18050 (
);

FILL FILL_1__13854_ (
);

FILL FILL_1__13434_ (
);

FILL FILL_4__16299_ (
);

FILL FILL_1__13014_ (
);

FILL FILL_0__12847_ (
);

FILL SFILL89320x67050 (
);

OAI21X1 _12712_ (
    .A(_3499_),
    .B(IRWrite_bF$buf0),
    .C(_3500_),
    .Y(_3490_[5])
);

FILL FILL_0__12427_ (
);

FILL FILL_0__12007_ (
);

FILL FILL_5__8884_ (
);

FILL FILL_5__8464_ (
);

FILL FILL_6__16206_ (
);

NAND3X1 _15184_ (
    .A(_5654_),
    .B(_5655_),
    .C(_5660_),
    .Y(_5661_)
);

FILL FILL_5__15619_ (
);

FILL FILL_3__16233_ (
);

NAND2X1 _9919_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1546_)
);

FILL FILL_5__10754_ (
);

FILL FILL_1__8876_ (
);

FILL FILL_1__8456_ (
);

FILL FILL_2__15646_ (
);

FILL FILL_2__15226_ (
);

FILL FILL_4__6881_ (
);

FILL FILL_0__16260_ (
);

FILL FILL_2__10781_ (
);

FILL FILL_2__10361_ (
);

FILL FILL_1__14639_ (
);

FILL FILL_1__14219_ (
);

FILL SFILL84840x50 (
);

FILL FILL_3__9743_ (
);

NOR2X1 _13917_ (
    .A(_4419_),
    .B(_4416_),
    .Y(_4420_)
);

FILL FILL_5__9669_ (
);

FILL FILL_5__9249_ (
);

FILL SFILL89320x22050 (
);

OAI21X1 _16389_ (
    .A(_6812_),
    .B(gnd),
    .C(_6813_),
    .Y(_6769_[22])
);

FILL FILL_6__12126_ (
);

FILL FILL_4__13580_ (
);

FILL FILL_4__13160_ (
);

FILL FILL_5__11959_ (
);

FILL FILL_2__7740_ (
);

FILL FILL_3__12993_ (
);

FILL FILL_5__11539_ (
);

FILL FILL_3__12573_ (
);

FILL FILL_2__7320_ (
);

FILL FILL_5__11119_ (
);

FILL FILL_3__12153_ (
);

FILL SFILL18760x42050 (
);

FILL SFILL49160x33050 (
);

FILL FILL_4__7246_ (
);

FILL FILL_2__11986_ (
);

FILL FILL_2__11566_ (
);

FILL FILL_2__11146_ (
);

FILL FILL_0__12180_ (
);

FILL FILL_5__12900_ (
);

FILL SFILL54120x16050 (
);

FILL FILL_1__10979_ (
);

FILL FILL_1__10559_ (
);

FILL FILL_1__10139_ (
);

FILL FILL_5__15792_ (
);

FILL FILL_5__15372_ (
);

FILL FILL_0__7986_ (
);

FILL FILL_0__7566_ (
);

NAND2X1 _9672_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1422_)
);

NAND2X1 _9252_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1203_)
);

FILL FILL_6__8113_ (
);

FILL SFILL79320x65050 (
);

FILL SFILL18680x49050 (
);

FILL FILL_1__11920_ (
);

FILL FILL_4__14785_ (
);

FILL FILL_4__14365_ (
);

FILL FILL_1__11500_ (
);

FILL FILL_2__8525_ (
);

FILL FILL_0__10913_ (
);

FILL FILL_3__13778_ (
);

FILL FILL_3__13358_ (
);

FILL FILL_2__8105_ (
);

FILL FILL_1__14392_ (
);

FILL FILL_5__6950_ (
);

INVX1 _13670_ (
    .A(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_4178_)
);

FILL FILL_0__13385_ (
);

NAND2X1 _13250_ (
    .A(_3770_),
    .B(_3754_),
    .Y(_3793_)
);

FILL SFILL110120x82050 (
);

FILL FILL_1__6942_ (
);

FILL FILL_4__9812_ (
);

FILL FILL_2__13712_ (
);

FILL FILL_3__6868_ (
);

FILL FILL_5__16157_ (
);

FILL FILL_5__11292_ (
);

FILL FILL_1__12705_ (
);

FILL FILL_2__16184_ (
);

FILL SFILL79320x20050 (
);

FILL FILL_4__10285_ (
);

FILL FILL_1__15597_ (
);

FILL FILL_1__15177_ (
);

FILL FILL_5__7735_ (
);

FILL FILL_5__7315_ (
);

FILL FILL111960x33050 (
);

OAI22X1 _14875_ (
    .A(_5356_),
    .B(_3967__bF$buf3),
    .C(_3978_),
    .D(_5357_),
    .Y(_5358_)
);

FILL SFILL39160x31050 (
);

INVX1 _14455_ (
    .A(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_4946_)
);

AOI21X1 _14035_ (
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .B(_4079__bF$buf0),
    .C(_4534_),
    .Y(_4535_)
);

FILL FILL_3__15924_ (
);

FILL FILL_3__15504_ (
);

FILL FILL_1__7727_ (
);

FILL FILL_1__7307_ (
);

FILL FILL_6__13084_ (
);

FILL FILL_2__14917_ (
);

FILL FILL_0__15951_ (
);

FILL FILL_0__15531_ (
);

FILL FILL_0__15111_ (
);

FILL FILL_5__12497_ (
);

FILL FILL_5__12077_ (
);

FILL FILL_1__11097_ (
);

FILL FILL_4__12851_ (
);

FILL FILL_4__12431_ (
);

FILL FILL_4__12011_ (
);

OAI21X1 _10795_ (
    .A(_1986_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1987_),
    .Y(_1953_[17])
);

OAI21X1 _10375_ (
    .A(_1767_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .C(_1768_),
    .Y(_1758_[5])
);

FILL FILL_3__11844_ (
);

FILL FILL_3__11424_ (
);

FILL FILL_3__11004_ (
);

FILL FILL_4__6937_ (
);

FILL FILL_0__16316_ (
);

FILL FILL_2__10837_ (
);

FILL FILL_2__9483_ (
);

FILL FILL_0__11871_ (
);

FILL FILL_2__10417_ (
);

FILL FILL_0__11451_ (
);

FILL FILL_0__11031_ (
);

FILL FILL_5__14643_ (
);

FILL FILL_0__6837_ (
);

FILL FILL_5__14223_ (
);

DFFSR _8943_ (
    .Q(\datapath_1.regfile_1.regOut[16] [25]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_978_[25])
);

NAND2X1 _8523_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_839_)
);

NAND2X1 _8103_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_620_)
);

FILL FILL_1__7480_ (
);

FILL FILL_1__7060_ (
);

FILL FILL_4__13636_ (
);

FILL FILL_4__13216_ (
);

FILL FILL_2__14670_ (
);

FILL FILL_2__14250_ (
);

FILL SFILL114280x59050 (
);

FILL FILL_3__12629_ (
);

FILL FILL_1__13663_ (
);

FILL FILL_3__12209_ (
);

FILL FILL_1__13243_ (
);

FILL FILL_1_BUFX2_insert710 (
);

FILL FILL_1_BUFX2_insert711 (
);

FILL SFILL69240x25050 (
);

FILL FILL_0__12656_ (
);

FILL FILL_1_BUFX2_insert712 (
);

DFFSR _12941_ (
    .Q(\datapath_1.a [22]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3555_[22])
);

FILL FILL_1_BUFX2_insert713 (
);

NAND2X1 _12521_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [27]),
    .Y(_3414_)
);

FILL FILL_0__12236_ (
);

AOI22X1 _12101_ (
    .A(\datapath_1.ALUResult [28]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3122_)
);

FILL FILL_1_BUFX2_insert714 (
);

FILL FILL_1_BUFX2_insert715 (
);

FILL FILL_1_BUFX2_insert716 (
);

FILL FILL_1_BUFX2_insert717 (
);

FILL FILL_5__8273_ (
);

FILL FILL_1_BUFX2_insert718 (
);

FILL FILL_1_BUFX2_insert719 (
);

FILL FILL_5__15848_ (
);

FILL FILL_5__15428_ (
);

FILL FILL_5__15008_ (
);

NAND2X1 _9728_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1439_)
);

FILL FILL_3__16042_ (
);

FILL FILL_5__10983_ (
);

DFFSR _9308_ (
    .Q(\datapath_1.regfile_1.regOut[19] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1173_[6])
);

FILL FILL_5__10563_ (
);

FILL FILL_1__8265_ (
);

FILL FILL_5__10143_ (
);

FILL FILL_2__15875_ (
);

FILL FILL_2__15455_ (
);

FILL SFILL99400x57050 (
);

FILL FILL_2__15035_ (
);

FILL FILL_2__10170_ (
);

FILL FILL_1__14868_ (
);

FILL FILL_1__14448_ (
);

FILL FILL_1__14028_ (
);

FILL FILL_3__9552_ (
);

FILL FILL_3__9132_ (
);

NOR2X1 _13726_ (
    .A(_4229_),
    .B(_4232_),
    .Y(_4233_)
);

NOR3X1 _13306_ (
    .A(_3781_),
    .B(_3835_),
    .C(_3840_),
    .Y(\datapath_1.regfile_1.regEn [9])
);

FILL FILL_5__9898_ (
);

FILL FILL_5__9478_ (
);

FILL SFILL104360x50050 (
);

FILL SFILL83720x79050 (
);

INVX1 _16198_ (
    .A(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_6650_)
);

FILL FILL_0__14802_ (
);

FILL FILL_5__11768_ (
);

FILL FILL_5__11348_ (
);

FILL FILL_3__12382_ (
);

FILL FILL_4__7475_ (
);

FILL FILL_4__7055_ (
);

FILL FILL_2__11795_ (
);

FILL FILL_2__11375_ (
);

FILL SFILL99400x12050 (
);

FILL FILL_1__10788_ (
);

FILL FILL_1__10368_ (
);

FILL FILL_4__11702_ (
);

FILL FILL_5__15181_ (
);

FILL FILL_0__7375_ (
);

NAND2X1 _9481_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1315_)
);

DFFSR _9061_ (
    .Q(\datapath_1.regfile_1.regOut[17] [15]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1043_[15])
);

FILL FILL_4__14594_ (
);

FILL FILL_4__14174_ (
);

FILL FILL_2__8754_ (
);

FILL FILL_2__8334_ (
);

FILL FILL_3__13587_ (
);

FILL FILL_0__10302_ (
);

FILL FILL_3__13167_ (
);

FILL FILL_5__13914_ (
);

FILL SFILL28760x39050 (
);

FILL FILL_4__9621_ (
);

FILL FILL_4__12907_ (
);

FILL FILL_2__13941_ (
);

FILL FILL_5__16386_ (
);

FILL FILL_2__13521_ (
);

FILL FILL_4_BUFX2_insert225 (
);

FILL FILL_2__13101_ (
);

FILL FILL_4_BUFX2_insert226 (
);

FILL FILL_4_BUFX2_insert227 (
);

FILL FILL_4_BUFX2_insert228 (
);

FILL FILL_4_BUFX2_insert229 (
);

FILL FILL_4__15799_ (
);

FILL FILL_4__15379_ (
);

FILL FILL_1__12514_ (
);

FILL FILL_0__9941_ (
);

FILL SFILL73720x77050 (
);

FILL SFILL89800x24050 (
);

FILL FILL_0__11927_ (
);

FILL FILL_0__9521_ (
);

FILL FILL_2__9539_ (
);

FILL FILL_0__9101_ (
);

FILL FILL_0__11507_ (
);

FILL FILL_2__9119_ (
);

FILL FILL_5__7964_ (
);

FILL FILL_5__7544_ (
);

FILL FILL_5__7124_ (
);

FILL FILL_4__16320_ (
);

FILL FILL_0__14399_ (
);

INVX1 _14684_ (
    .A(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_5171_)
);

NOR2X1 _14264_ (
    .A(_4749_),
    .B(_4759_),
    .Y(_4760_)
);

FILL FILL_3__15733_ (
);

FILL FILL_3__15313_ (
);

FILL FILL_1__7956_ (
);

FILL FILL_1__7116_ (
);

FILL SFILL94280x61050 (
);

FILL FILL_2__14726_ (
);

FILL FILL_0__15760_ (
);

FILL FILL_2__14306_ (
);

FILL FILL_0__15340_ (
);

FILL FILL_1__13719_ (
);

FILL FILL_4__11299_ (
);

FILL FILL_3__8823_ (
);

FILL FILL_3__8403_ (
);

FILL FILL_5__8749_ (
);

FILL SFILL89320x17050 (
);

FILL FILL_5__8329_ (
);

NAND2X1 _15889_ (
    .A(_6342_),
    .B(_6348_),
    .Y(_6349_)
);

FILL FILL_4__12660_ (
);

OAI22X1 _15469_ (
    .A(_5526__bF$buf1),
    .B(_4457_),
    .C(_4460_),
    .D(_5527__bF$buf2),
    .Y(_5939_)
);

NOR2X1 _15049_ (
    .A(_5525_),
    .B(_5528_),
    .Y(_5529_)
);

FILL FILL_4__12240_ (
);

NAND2X1 _10184_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1682_)
);

FILL FILL_5__10619_ (
);

FILL FILL_3__11653_ (
);

FILL SFILL18760x37050 (
);

FILL FILL_3__11233_ (
);

OAI21X1 _16410_ (
    .A(_6826_),
    .B(gnd),
    .C(_6827_),
    .Y(_6769_[29])
);

FILL FILL_0__16125_ (
);

FILL FILL_2__10646_ (
);

FILL FILL_2__9292_ (
);

FILL FILL_0__11680_ (
);

FILL FILL_0__11260_ (
);

FILL FILL_3__9608_ (
);

FILL FILL_3_BUFX2_insert240 (
);

FILL FILL_3_BUFX2_insert241 (
);

FILL FILL_5__14872_ (
);

FILL FILL_3_BUFX2_insert242 (
);

FILL FILL_5__14452_ (
);

FILL FILL_3_BUFX2_insert243 (
);

FILL FILL_3_BUFX2_insert244 (
);

FILL FILL_5__14032_ (
);

FILL FILL_3_BUFX2_insert245 (
);

NAND2X1 _8752_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_951_)
);

NAND2X1 _8332_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_732_)
);

FILL FILL_3_BUFX2_insert246 (
);

FILL FILL_3_BUFX2_insert247 (
);

FILL SFILL33960x12050 (
);

FILL FILL_3_BUFX2_insert248 (
);

FILL FILL_4__13865_ (
);

FILL FILL_3_BUFX2_insert249 (
);

FILL FILL_4__13445_ (
);

FILL FILL_4__13025_ (
);

NAND2X1 _11389_ (
    .A(_2187_),
    .B(_2505_),
    .Y(_2506_)
);

FILL FILL_2__7605_ (
);

FILL FILL_3__12858_ (
);

FILL FILL_3__12438_ (
);

FILL FILL_1__13892_ (
);

FILL FILL_3__12018_ (
);

FILL FILL_1__13472_ (
);

FILL FILL_0__12885_ (
);

NAND2X1 _12750_ (
    .A(IRWrite_bF$buf7),
    .B(memoryOutData[18]),
    .Y(_3526_)
);

FILL FILL_0__12465_ (
);

FILL FILL_0__12045_ (
);

NAND3X1 _12330_ (
    .A(_3284_),
    .B(_3285_),
    .C(_3286_),
    .Y(\datapath_1.alu_1.ALUInB [28])
);

FILL FILL_5__8082_ (
);

FILL FILL_5__15657_ (
);

FILL FILL_5__15237_ (
);

DFFSR _9957_ (
    .Q(\datapath_1.regfile_1.regOut[24] [15]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_1498_[15])
);

FILL FILL_3__16271_ (
);

INVX1 _9537_ (
    .A(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_1352_)
);

FILL FILL_5__10792_ (
);

INVX1 _9117_ (
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_1133_)
);

FILL FILL_5__10372_ (
);

FILL FILL_1__8494_ (
);

FILL FILL_1__8074_ (
);

FILL FILL_2__15684_ (
);

FILL FILL_2__15264_ (
);

FILL FILL_1__14677_ (
);

FILL FILL_1__14257_ (
);

FILL FILL_0_BUFX2_insert370 (
);

FILL FILL111960x28050 (
);

FILL FILL_0_BUFX2_insert371 (
);

FILL FILL_0_BUFX2_insert372 (
);

FILL FILL_3__9781_ (
);

FILL FILL_0_BUFX2_insert373 (
);

FILL FILL_0_BUFX2_insert374 (
);

INVX1 _13955_ (
    .A(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_4457_)
);

FILL FILL_3__9361_ (
);

FILL FILL_0_BUFX2_insert375 (
);

INVX1 _13535_ (
    .A(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_4045_)
);

INVX1 _13115_ (
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_3708_)
);

FILL FILL_0_BUFX2_insert376 (
);

FILL FILL_0_BUFX2_insert377 (
);

FILL FILL_0_BUFX2_insert378 (
);

FILL FILL_5__9287_ (
);

FILL FILL_0_BUFX2_insert379 (
);

FILL FILL_0__14611_ (
);

FILL FILL_5__11997_ (
);

FILL FILL_5__11577_ (
);

FILL FILL_1__9279_ (
);

FILL FILL_5__11157_ (
);

FILL FILL_3__12191_ (
);

FILL SFILL69320x58050 (
);

FILL SFILL69800x20050 (
);

FILL FILL_2__16049_ (
);

FILL SFILL74680x71050 (
);

FILL FILL_2__11184_ (
);

FILL FILL_1__10177_ (
);

FILL FILL_4__11931_ (
);

FILL FILL_4__11511_ (
);

FILL FILL_6__8991_ (
);

FILL FILL_0__7184_ (
);

FILL FILL_2_BUFX2_insert50 (
);

FILL FILL_2_BUFX2_insert51 (
);

INVX1 _9290_ (
    .A(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_1228_)
);

FILL FILL_1__16403_ (
);

FILL FILL_2_BUFX2_insert52 (
);

FILL FILL_3__10924_ (
);

FILL FILL_2_BUFX2_insert53 (
);

FILL FILL_3__10504_ (
);

FILL FILL_2_BUFX2_insert54 (
);

FILL FILL_2_BUFX2_insert55 (
);

FILL FILL_2_BUFX2_insert56 (
);

FILL FILL_2_BUFX2_insert57 (
);

FILL FILL_0__15816_ (
);

FILL FILL_2_BUFX2_insert58 (
);

FILL FILL_2_BUFX2_insert59 (
);

FILL FILL_2__8983_ (
);

FILL FILL_0__10951_ (
);

FILL FILL_2__8143_ (
);

FILL FILL_0__10531_ (
);

FILL FILL_3__13396_ (
);

FILL FILL_0__10111_ (
);

FILL FILL_4__8489_ (
);

FILL FILL_4__8069_ (
);

FILL FILL_2__12389_ (
);

FILL SFILL69320x13050 (
);

FILL FILL_5__13723_ (
);

FILL FILL_5__13303_ (
);

NAND2X1 _7603_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_368_)
);

FILL FILL_1__6980_ (
);

FILL FILL_4__9850_ (
);

FILL FILL_4__12716_ (
);

FILL FILL_4__9010_ (
);

FILL FILL_2__13750_ (
);

FILL FILL_2__13330_ (
);

FILL FILL_5__16195_ (
);

FILL FILL_0__8389_ (
);

FILL FILL_3__11709_ (
);

FILL FILL_1__12743_ (
);

FILL FILL_4__15188_ (
);

FILL FILL_1__12323_ (
);

FILL FILL_2__9768_ (
);

FILL FILL_0__9750_ (
);

FILL FILL_2__9348_ (
);

FILL FILL_0__11736_ (
);

FILL SFILL19240x60050 (
);

OAI21X1 _11601_ (
    .A(_2676_),
    .B(_2258_),
    .C(_2523_),
    .Y(_2707_)
);

FILL FILL_0__11316_ (
);

FILL FILL_6__15935_ (
);

FILL FILL_5__7353_ (
);

OAI22X1 _14493_ (
    .A(_4982_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf3),
    .D(_4983_),
    .Y(_4984_)
);

NAND3X1 _14073_ (
    .A(_4564_),
    .B(_4565_),
    .C(_4572_),
    .Y(_4573_)
);

FILL FILL_5__14928_ (
);

FILL FILL_5__14508_ (
);

FILL FILL_3__15962_ (
);

FILL FILL_3__15542_ (
);

DFFSR _8808_ (
    .Q(\datapath_1.regfile_1.regOut[15] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_913_[18])
);

FILL FILL_3__15122_ (
);

FILL FILL_1__7765_ (
);

FILL FILL_1__7345_ (
);

FILL FILL_2__14955_ (
);

FILL FILL_2__14535_ (
);

FILL FILL_2__14115_ (
);

FILL FILL_1__13948_ (
);

FILL FILL_1__13528_ (
);

FILL FILL_1__13108_ (
);

FILL FILL_3__8632_ (
);

DFFSR _12806_ (
    .Q(\datapath_1.PCJump [17]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3490_[15])
);

FILL FILL_3__8212_ (
);

FILL FILL_5__8978_ (
);

FILL SFILL104360x45050 (
);

FILL FILL_5__8138_ (
);

FILL FILL_6__11855_ (
);

INVX1 _15698_ (
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_6162_)
);

FILL SFILL3000x57050 (
);

OAI21X1 _15278_ (
    .A(_5524__bF$buf2),
    .B(_4236_),
    .C(_5752_),
    .Y(_5753_)
);

FILL FILL_3__16327_ (
);

FILL FILL_5__10428_ (
);

FILL FILL_3__11882_ (
);

FILL FILL_5__10008_ (
);

FILL FILL_3__11462_ (
);

FILL FILL_3__11042_ (
);

FILL FILL_4__6975_ (
);

FILL FILL_0__16354_ (
);

FILL FILL_2__10875_ (
);

FILL FILL_2__10035_ (
);

FILL FILL_1__9911_ (
);

FILL SFILL3400x26050 (
);

FILL FILL_3__9417_ (
);

FILL FILL_5__14681_ (
);

FILL FILL_5__14261_ (
);

FILL FILL_0__6875_ (
);

NAND2X1 _8981_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1063_)
);

FILL FILL112440x51050 (
);

DFFSR _8561_ (
    .Q(\datapath_1.regfile_1.regOut[13] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_783_[27])
);

INVX1 _8141_ (
    .A(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_645_)
);

FILL FILL_4__13674_ (
);

FILL FILL_4__13254_ (
);

INVX2 _11198_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .Y(_2317_)
);

FILL FILL_2__7834_ (
);

FILL FILL_2__7414_ (
);

FILL FILL_3__12247_ (
);

FILL FILL_1__13281_ (
);

FILL FILL_0__12274_ (
);

FILL FILL_6__16053_ (
);

FILL FILL_4__8701_ (
);

FILL FILL_5__15886_ (
);

FILL FILL_2__12601_ (
);

FILL FILL_5__15466_ (
);

FILL FILL_5__15046_ (
);

INVX1 _9766_ (
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_1464_)
);

FILL FILL_3__16080_ (
);

INVX1 _9346_ (
    .A(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_1245_)
);

FILL FILL_5__10181_ (
);

FILL FILL_4__14879_ (
);

FILL FILL_4__14459_ (
);

FILL FILL_4__14039_ (
);

FILL FILL_2__15493_ (
);

FILL FILL_2__15073_ (
);

FILL FILL_0__8601_ (
);

FILL FILL_2__8619_ (
);

FILL FILL_1__14486_ (
);

FILL FILL_1__14066_ (
);

FILL FILL_4__15820_ (
);

FILL FILL_4__15400_ (
);

FILL FILL_3__9590_ (
);

FILL FILL_0__13899_ (
);

INVX1 _13764_ (
    .A(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_4270_)
);

FILL FILL_3__9170_ (
);

FILL FILL_0__13479_ (
);

AND2X2 _13344_ (
    .A(_3864_),
    .B(_3769_),
    .Y(\datapath_1.regfile_1.regEn [23])
);

FILL FILL_3__14813_ (
);

FILL FILL_5__9096_ (
);

FILL FILL_4__9906_ (
);

FILL SFILL94280x56050 (
);

FILL FILL_2__13806_ (
);

FILL FILL_0__14840_ (
);

FILL FILL_0__14420_ (
);

FILL FILL_0__14000_ (
);

FILL FILL_5__11386_ (
);

FILL FILL_1__9088_ (
);

FILL FILL_2__16278_ (
);

FILL FILL_4__7093_ (
);

FILL FILL_4__10799_ (
);

FILL FILL_4__10379_ (
);

FILL FILL_0__9806_ (
);

FILL SFILL94600x68050 (
);

FILL FILL_5__7829_ (
);

INVX1 _14969_ (
    .A(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_5450_)
);

AOI21X1 _14549_ (
    .A(_5017_),
    .B(_5038_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [22])
);

FILL FILL_4__11740_ (
);

NOR2X1 _14129_ (
    .A(_4623_),
    .B(_4626_),
    .Y(_4627_)
);

FILL FILL_4__11320_ (
);

FILL SFILL98920x76050 (
);

FILL FILL_1__16212_ (
);

FILL SFILL79400x48050 (
);

FILL FILL_3__10313_ (
);

NOR2X1 _15910_ (
    .A(_6368_),
    .B(_6361_),
    .Y(_6369_)
);

FILL FILL_0__15625_ (
);

FILL FILL_0__15205_ (
);

FILL SFILL94280x11050 (
);

FILL FILL_0__10760_ (
);

FILL FILL_2__8372_ (
);

FILL SFILL23640x74050 (
);

FILL FILL_2__12198_ (
);

FILL FILL_5__13952_ (
);

FILL FILL_5__13532_ (
);

FILL FILL_5__13112_ (
);

NAND2X1 _7832_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_480_)
);

FILL SFILL8680x73050 (
);

DFFSR _7412_ (
    .Q(\datapath_1.regfile_1.regOut[4] [30]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_198_[30])
);

FILL FILL_4_BUFX2_insert600 (
);

FILL FILL_4_BUFX2_insert601 (
);

FILL FILL_4_BUFX2_insert602 (
);

FILL FILL_4_BUFX2_insert603 (
);

FILL FILL_4__12525_ (
);

FILL FILL_4_BUFX2_insert604 (
);

FILL FILL_4__12105_ (
);

FILL FILL_4_BUFX2_insert605 (
);

FILL FILL_4_BUFX2_insert606 (
);

NAND2X1 _10889_ (
    .A(_2035_),
    .B(_2034_),
    .Y(ALUControl[1])
);

FILL FILL_0__8198_ (
);

FILL FILL_4_BUFX2_insert607 (
);

DFFSR _10469_ (
    .Q(\datapath_1.regfile_1.regOut[28] [15]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_1758_[15])
);

FILL FILL_4_BUFX2_insert608 (
);

INVX1 _10049_ (
    .A(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_1612_)
);

FILL FILL_3__11938_ (
);

FILL FILL_4_BUFX2_insert609 (
);

FILL FILL_1__12972_ (
);

FILL FILL_3__11518_ (
);

FILL FILL_1__12132_ (
);

FILL FILL_2__9997_ (
);

FILL FILL_0__11965_ (
);

INVX1 _11830_ (
    .A(_2919_),
    .Y(\datapath_1.ALUResult [2])
);

FILL FILL_2__9157_ (
);

FILL FILL_0__11545_ (
);

INVX1 _11410_ (
    .A(_2303_),
    .Y(_2527_)
);

FILL FILL_0__11125_ (
);

FILL FILL_5__7582_ (
);

FILL SFILL59960x6050 (
);

FILL FILL_5__7162_ (
);

FILL FILL_5__14737_ (
);

FILL FILL_5__14317_ (
);

FILL FILL_3__15771_ (
);

FILL FILL_3__15351_ (
);

FILL SFILL8600x71050 (
);

INVX1 _8617_ (
    .A(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_881_)
);

FILL FILL_1__7994_ (
);

FILL FILL_1__7574_ (
);

FILL FILL_2__14764_ (
);

FILL FILL_2__14344_ (
);

FILL FILL_1__13757_ (
);

FILL FILL_1__13337_ (
);

FILL FILL_3__8861_ (
);

FILL FILL_3__8441_ (
);

INVX1 _12615_ (
    .A(\datapath_1.Data [16]),
    .Y(_3456_)
);

FILL FILL_3__8021_ (
);

FILL FILL_5__8787_ (
);

FILL FILL_6__16109_ (
);

FILL FILL_5__8367_ (
);

FILL SFILL13640x72050 (
);

NAND2X1 _15087_ (
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .B(_5565__bF$buf0),
    .Y(_5566_)
);

FILL FILL_3__16136_ (
);

FILL FILL_5__10657_ (
);

FILL FILL_1__8779_ (
);

FILL FILL_1__8359_ (
);

FILL FILL_5__10237_ (
);

FILL FILL_3__11691_ (
);

FILL FILL_3__11271_ (
);

FILL FILL_2__15969_ (
);

FILL FILL_2__15549_ (
);

FILL FILL_2__15129_ (
);

FILL FILL_0__16163_ (
);

FILL FILL_2__10684_ (
);

FILL SFILL114440x35050 (
);

FILL FILL_2__10264_ (
);

FILL FILL_1__9720_ (
);

FILL FILL_1__9300_ (
);

FILL FILL_3_BUFX2_insert620 (
);

FILL FILL_3__9646_ (
);

FILL FILL_3__9226_ (
);

FILL FILL_3_BUFX2_insert621 (
);

FILL SFILL109560x5050 (
);

FILL FILL_3_BUFX2_insert622 (
);

FILL FILL_5__14490_ (
);

FILL FILL_3_BUFX2_insert623 (
);

FILL FILL_3_BUFX2_insert624 (
);

FILL FILL_5__14070_ (
);

FILL FILL_1__15903_ (
);

FILL FILL_3_BUFX2_insert625 (
);

DFFSR _8790_ (
    .Q(\datapath_1.regfile_1.regOut[15] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_913_[0])
);

FILL FILL_3_BUFX2_insert626 (
);

INVX1 _8370_ (
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_757_)
);

FILL FILL_3_BUFX2_insert627 (
);

FILL FILL_3_BUFX2_insert628 (
);

FILL FILL_6__12449_ (
);

FILL FILL_3_BUFX2_insert629 (
);

FILL FILL_6__12029_ (
);

FILL FILL_4__13483_ (
);

FILL SFILL13160x65050 (
);

FILL FILL_3__12896_ (
);

FILL FILL_2__7223_ (
);

FILL FILL_3__12476_ (
);

FILL FILL_3__12056_ (
);

FILL FILL_1__13090_ (
);

FILL FILL_4__7989_ (
);

FILL FILL_4__7569_ (
);

FILL FILL_2__11889_ (
);

FILL FILL_2__11469_ (
);

FILL FILL_2__11049_ (
);

FILL FILL_0__12083_ (
);

FILL FILL_4__8510_ (
);

FILL FILL_5__15695_ (
);

FILL FILL_2__12830_ (
);

FILL FILL_2__12410_ (
);

FILL FILL_0__7889_ (
);

FILL FILL_5__15275_ (
);

FILL SFILL74200x50050 (
);

INVX1 _9995_ (
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_1576_)
);

FILL FILL_0__7469_ (
);

FILL FILL_0__7049_ (
);

DFFSR _9575_ (
    .Q(\datapath_1.regfile_1.regOut[21] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_1303_[17])
);

OAI21X1 _9155_ (
    .A(_1157_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1158_),
    .Y(_1108_[25])
);

FILL FILL_1__11823_ (
);

FILL FILL_4__14688_ (
);

FILL FILL_4__14268_ (
);

FILL FILL_1__11403_ (
);

FILL FILL_2__8848_ (
);

FILL FILL_0__8830_ (
);

FILL FILL_0__10816_ (
);

FILL FILL_2__8008_ (
);

FILL FILL_1__14295_ (
);

FILL FILL_5__6853_ (
);

FILL FILL_0_BUFX2_insert750 (
);

FILL FILL_0_BUFX2_insert751 (
);

FILL FILL_0_BUFX2_insert752 (
);

FILL FILL_0_BUFX2_insert753 (
);

INVX1 _13993_ (
    .A(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_4494_)
);

FILL FILL_0_BUFX2_insert754 (
);

FILL FILL_0__13288_ (
);

FILL FILL_0_BUFX2_insert755 (
);

INVX1 _13573_ (
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_4083_)
);

OAI21X1 _13153_ (
    .A(_3732_),
    .B(PCEn_bF$buf4),
    .C(_3733_),
    .Y(_3685_[24])
);

FILL FILL_0_BUFX2_insert756 (
);

FILL FILL_0_BUFX2_insert757 (
);

FILL FILL_3__14622_ (
);

FILL FILL_0_BUFX2_insert758 (
);

FILL FILL_3__14202_ (
);

FILL FILL_0_BUFX2_insert759 (
);

FILL FILL_1__6845_ (
);

FILL FILL_2__13615_ (
);

FILL FILL_5__11195_ (
);

FILL FILL_1__12608_ (
);

FILL FILL_2__16087_ (
);

FILL FILL_4__10188_ (
);

FILL FILL_0__9615_ (
);

FILL FILL_3__7712_ (
);

FILL FILL_4__16414_ (
);

FILL FILL_5__7218_ (
);

FILL FILL_6__10935_ (
);

OAI22X1 _14778_ (
    .A(_5261_),
    .B(_3930__bF$buf2),
    .C(_3966__bF$buf2),
    .D(_5262_),
    .Y(_5263_)
);

AOI22X1 _14358_ (
    .A(\datapath_1.regfile_1.regOut[31] [19]),
    .B(_3995__bF$buf2),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_4851_)
);

FILL FILL_3__15827_ (
);

FILL FILL_3__15407_ (
);

FILL FILL_1__16021_ (
);

FILL FILL_3__10962_ (
);

FILL FILL_3__10542_ (
);

FILL FILL_3__10122_ (
);

FILL FILL_0__15854_ (
);

FILL FILL_0__15434_ (
);

FILL FILL_0__15014_ (
);

FILL FILL_3__8917_ (
);

FILL FILL_5__13761_ (
);

FILL FILL_5__13341_ (
);

FILL FILL112440x46050 (
);

DFFSR _7641_ (
    .Q(\datapath_1.regfile_1.regOut[6] [3]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_328_[3])
);

INVX1 _7221_ (
    .A(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_174_)
);

FILL FILL_4__12754_ (
);

FILL FILL_4__12334_ (
);

INVX1 _10698_ (
    .A(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_1943_)
);

FILL FILL_6__9394_ (
);

INVX1 _10278_ (
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_1724_)
);

FILL FILL_2__6914_ (
);

FILL FILL_3__11747_ (
);

FILL FILL_1__12781_ (
);

FILL FILL_3__11327_ (
);

FILL FILL_1__12361_ (
);

FILL FILL_0__16219_ (
);

FILL FILL_0__11774_ (
);

FILL FILL_2__9386_ (
);

FILL FILL_0__11354_ (
);

FILL FILL_5__14966_ (
);

FILL FILL_5__14546_ (
);

FILL FILL_5__14126_ (
);

FILL FILL_3__15580_ (
);

INVX1 _8846_ (
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_993_)
);

FILL FILL_3__15160_ (
);

DFFSR _8426_ (
    .Q(\datapath_1.regfile_1.regOut[12] [20]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_718_[20])
);

OAI21X1 _8006_ (
    .A(_574_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .C(_575_),
    .Y(_523_[26])
);

FILL FILL_4__13959_ (
);

FILL FILL_2__14993_ (
);

FILL FILL_4__13539_ (
);

FILL FILL_2__14573_ (
);

FILL FILL_4__13119_ (
);

FILL FILL_2__14153_ (
);

FILL FILL_1__13986_ (
);

FILL FILL_1__13566_ (
);

FILL FILL_1__13146_ (
);

FILL FILL_4__14900_ (
);

FILL FILL_0__12979_ (
);

FILL FILL_3__8250_ (
);

INVX1 _12844_ (
    .A(\datapath_1.a [7]),
    .Y(_3568_)
);

FILL FILL_0__12139_ (
);

INVX1 _12424_ (
    .A(ALUOut[27]),
    .Y(_3348_)
);

NAND3X1 _12004_ (
    .A(PCSource_1_bF$buf2),
    .B(\aluControl_1.inst [2]),
    .C(_3034__bF$buf4),
    .Y(_3049_)
);

FILL FILL_5__8596_ (
);

FILL FILL_0__13920_ (
);

FILL FILL_3__16365_ (
);

FILL FILL_0__13500_ (
);

FILL FILL_5__10886_ (
);

FILL FILL_1__8588_ (
);

FILL FILL_5__10046_ (
);

FILL FILL_3__11080_ (
);

FILL FILL_2__15778_ (
);

FILL FILL_2__15358_ (
);

FILL FILL_0__16392_ (
);

FILL FILL_2__10493_ (
);

FILL FILL_5__6909_ (
);

FILL FILL_3__9875_ (
);

INVX1 _13629_ (
    .A(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_4138_)
);

FILL FILL_3__9035_ (
);

FILL FILL_4__10820_ (
);

NOR2X1 _13209_ (
    .A(\datapath_1.a3 [1]),
    .B(_3751_),
    .Y(_3752_)
);

FILL FILL_4__10400_ (
);

FILL FILL_6__7880_ (
);

FILL FILL_1__15712_ (
);

FILL FILL_4__13292_ (
);

FILL SFILL58440x61050 (
);

FILL FILL_0__14705_ (
);

FILL FILL_2__7872_ (
);

FILL FILL_2__7452_ (
);

FILL FILL_2__7032_ (
);

FILL FILL_3__12285_ (
);

FILL SFILL23640x69050 (
);

FILL FILL_4__7798_ (
);

FILL FILL_4__7378_ (
);

FILL FILL_2__11698_ (
);

FILL FILL_2__11278_ (
);

FILL FILL_5__12612_ (
);

FILL SFILL8680x68050 (
);

NAND2X1 _6912_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_9_)
);

FILL FILL_2_BUFX2_insert280 (
);

FILL FILL_2_BUFX2_insert281 (
);

FILL FILL_2_BUFX2_insert282 (
);

FILL FILL_2_BUFX2_insert283 (
);

FILL FILL_2_BUFX2_insert284 (
);

FILL FILL_4__11605_ (
);

FILL FILL_2_BUFX2_insert285 (
);

FILL FILL_2_BUFX2_insert286 (
);

FILL FILL_5__15084_ (
);

FILL FILL_0__7698_ (
);

FILL FILL_2_BUFX2_insert287 (
);

FILL SFILL99000x8050 (
);

OAI21X1 _9384_ (
    .A(_1269_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .C(_1270_),
    .Y(_1238_[16])
);

FILL FILL_2_BUFX2_insert288 (
);

FILL FILL_2_BUFX2_insert289 (
);

FILL FILL_4__14497_ (
);

FILL FILL_1__11632_ (
);

FILL FILL_1__11212_ (
);

FILL FILL_4__14077_ (
);

FILL FILL_2__8657_ (
);

FILL FILL_0__10625_ (
);

OAI21X1 _10910_ (
    .A(_2046_),
    .B(_2052_),
    .C(_2055_),
    .Y(_2056_)
);

FILL FILL_2__8237_ (
);

FILL FILL_0__13097_ (
);

INVX8 _13382_ (
    .A(_3893__bF$buf1),
    .Y(_3894_)
);

FILL FILL_5__13817_ (
);

FILL FILL_3__14851_ (
);

FILL FILL_3__14431_ (
);

FILL FILL_3__14011_ (
);

FILL FILL_4__9524_ (
);

FILL FILL_4__9104_ (
);

FILL SFILL8680x23050 (
);

FILL FILL_2__13844_ (
);

FILL SFILL13720x60050 (
);

FILL FILL_2__13424_ (
);

FILL FILL_5__16289_ (
);

FILL FILL_2__13004_ (
);

FILL FILL_1__12837_ (
);

FILL FILL_1__12417_ (
);

FILL SFILL84200x47050 (
);

FILL FILL_3__7941_ (
);

FILL FILL_0__9424_ (
);

FILL FILL_3__7101_ (
);

FILL FILL_0__9004_ (
);

FILL FILL_5__7867_ (
);

FILL FILL_5__7447_ (
);

FILL FILL_4__16223_ (
);

FILL SFILL13640x67050 (
);

NOR2X1 _14587_ (
    .A(_5072_),
    .B(_5075_),
    .Y(_5076_)
);

OAI22X1 _14167_ (
    .A(_4664_),
    .B(_3982__bF$buf1),
    .C(_3983__bF$buf4),
    .D(_4663_),
    .Y(_4665_)
);

FILL FILL_3__15636_ (
);

FILL SFILL109480x47050 (
);

FILL FILL_3__15216_ (
);

FILL FILL_1__16250_ (
);

FILL FILL_1__7859_ (
);

FILL FILL_1__7439_ (
);

FILL FILL_3__10771_ (
);

FILL SFILL8600x21050 (
);

FILL FILL_2__14629_ (
);

FILL FILL_0__15663_ (
);

FILL FILL_2__14209_ (
);

FILL FILL_0__15243_ (
);

FILL SFILL109080x33050 (
);

FILL FILL_3__8726_ (
);

FILL FILL_5__13990_ (
);

FILL FILL_5__13570_ (
);

FILL SFILL74280x47050 (
);

FILL FILL_5__13150_ (
);

INVX1 _7870_ (
    .A(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_505_)
);

INVX1 _7450_ (
    .A(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_286_)
);

INVX1 _7030_ (
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_131_)
);

FILL FILL_4__12983_ (
);

FILL FILL_4__12143_ (
);

FILL SFILL13640x22050 (
);

DFFSR _10087_ (
    .Q(\datapath_1.regfile_1.regOut[25] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_1563_[17])
);

FILL FILL_3__11976_ (
);

FILL FILL_3__11556_ (
);

FILL FILL_1__12590_ (
);

FILL FILL_3__11136_ (
);

FILL FILL_1__12170_ (
);

FILL FILL_0__16028_ (
);

INVX1 _16313_ (
    .A(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_6762_)
);

FILL FILL_2__10969_ (
);

FILL FILL_2__10549_ (
);

FILL SFILL38840x71050 (
);

FILL FILL_2__10129_ (
);

FILL FILL_0__11583_ (
);

FILL FILL_0__11163_ (
);

FILL FILL_6__15782_ (
);

FILL FILL_6__15362_ (
);

FILL SFILL43800x54050 (
);

FILL FILL_2__11910_ (
);

FILL FILL_5__14775_ (
);

FILL SFILL74200x45050 (
);

FILL FILL_0__6969_ (
);

FILL FILL_5__14355_ (
);

FILL SFILL13560x29050 (
);

OAI21X1 _8655_ (
    .A(_905_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .C(_906_),
    .Y(_848_[29])
);

OAI21X1 _8235_ (
    .A(_686_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_687_),
    .Y(_653_[17])
);

FILL FILL_1__7192_ (
);

FILL FILL_1__10903_ (
);

FILL FILL_4__13768_ (
);

FILL FILL_4__13348_ (
);

FILL FILL_2__14382_ (
);

FILL FILL_2__7928_ (
);

FILL FILL_2__7508_ (
);

FILL FILL_1__13795_ (
);

FILL FILL_1__13375_ (
);

FILL SFILL99480x51050 (
);

FILL FILL_0__12788_ (
);

OAI21X1 _12653_ (
    .A(_3480_),
    .B(vdd),
    .C(_3481_),
    .Y(_3425_[28])
);

FILL FILL_0__12368_ (
);

FILL SFILL64680x59050 (
);

AOI22X1 _12233_ (
    .A(_2_[4]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf0),
    .D(\aluControl_1.inst [2]),
    .Y(_3214_)
);

FILL FILL_3__13702_ (
);

FILL FILL_6__11282_ (
);

FILL FILL_3__16174_ (
);

FILL FILL_5__10695_ (
);

FILL FILL112120x65050 (
);

FILL FILL_5__10275_ (
);

FILL FILL_1__8397_ (
);

FILL FILL_2__15587_ (
);

FILL FILL_2__15167_ (
);

FILL FILL_4__15914_ (
);

FILL FILL_3__9684_ (
);

INVX1 _13858_ (
    .A(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_4362_)
);

FILL FILL_3__9264_ (
);

INVX8 _13438_ (
    .A(_3949_),
    .Y(_3950_)
);

NAND2X1 _13018_ (
    .A(vdd),
    .B(\datapath_1.rd2 [22]),
    .Y(_3664_)
);

FILL FILL_3__14907_ (
);

FILL FILL_1__15941_ (
);

FILL FILL_1__15521_ (
);

FILL FILL_1__15101_ (
);

FILL FILL_0__14934_ (
);

FILL FILL_0__14514_ (
);

FILL FILL_2__7681_ (
);

FILL FILL_3__12094_ (
);

FILL FILL112120x20050 (
);

FILL FILL_4__7187_ (
);

FILL FILL_2__11087_ (
);

FILL FILL_5__12841_ (
);

FILL FILL_5__12421_ (
);

FILL FILL_5__12001_ (
);

FILL FILL_4__11834_ (
);

FILL FILL_4__11414_ (
);

FILL FILL_0__7087_ (
);

DFFSR _9193_ (
    .Q(\datapath_1.regfile_1.regOut[18] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1108_[19])
);

FILL FILL_1__16306_ (
);

FILL FILL_3__10827_ (
);

FILL FILL_3__10407_ (
);

FILL FILL_1__11861_ (
);

FILL FILL_1__11441_ (
);

FILL FILL112040x27050 (
);

FILL FILL_1__11021_ (
);

FILL FILL_0__15719_ (
);

FILL FILL_2__8886_ (
);

FILL FILL_2__8466_ (
);

FILL FILL_3__13299_ (
);

FILL FILL_0__10434_ (
);

FILL FILL_0__10014_ (
);

FILL FILL_5__6891_ (
);

DFFSR _13191_ (
    .Q(\datapath_1.mux_iord.din0 [16]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3685_[16])
);

FILL FILL_5__13626_ (
);

FILL FILL_3__14660_ (
);

FILL FILL_3__14240_ (
);

INVX1 _7926_ (
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_586_)
);

OAI21X1 _7506_ (
    .A(_322_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .C(_323_),
    .Y(_263_[30])
);

FILL FILL_1__6883_ (
);

FILL FILL_4__9753_ (
);

FILL FILL_4__12619_ (
);

FILL FILL_2__13653_ (
);

FILL FILL_2__13233_ (
);

FILL FILL_5__16098_ (
);

FILL FILL_1__12646_ (
);

FILL FILL_1__12226_ (
);

FILL FILL_0__9653_ (
);

FILL FILL_3__7750_ (
);

FILL FILL_3__7330_ (
);

NAND2X1 _11924_ (
    .A(IorD_bF$buf4),
    .B(ALUOut[12]),
    .Y(_2991_)
);

FILL FILL_0__11639_ (
);

FILL FILL_0__9233_ (
);

FILL FILL_0__11219_ (
);

OAI21X1 _11504_ (
    .A(_2605_),
    .B(_2606_),
    .C(_2616_),
    .Y(\datapath_1.ALUResult [25])
);

FILL FILL_6__15838_ (
);

FILL FILL_5__7676_ (
);

FILL FILL_4__16032_ (
);

FILL FILL_6__10553_ (
);

OAI22X1 _14396_ (
    .A(_3983__bF$buf1),
    .B(_4888_),
    .C(_3954__bF$buf0),
    .D(_4887_),
    .Y(_4889_)
);

FILL FILL_3__15865_ (
);

FILL FILL_3__15445_ (
);

FILL FILL_3__15025_ (
);

FILL SFILL39000x6050 (
);

FILL SFILL13720x2050 (
);

FILL FILL_6_BUFX2_insert510 (
);

FILL FILL_3__10580_ (
);

FILL FILL_1__7248_ (
);

FILL FILL_3__10160_ (
);

FILL FILL_2__14858_ (
);

FILL FILL_0__15892_ (
);

FILL FILL_2__14438_ (
);

FILL FILL_2__14018_ (
);

FILL FILL_0__15472_ (
);

FILL FILL_6_BUFX2_insert515 (
);

FILL FILL_0__15052_ (
);

FILL SFILL23720x57050 (
);

FILL FILL_3__8955_ (
);

OAI21X1 _12709_ (
    .A(_3497_),
    .B(IRWrite_bF$buf2),
    .C(_3498_),
    .Y(_3490_[4])
);

FILL FILL_3__8115_ (
);

FILL FILL_6__6960_ (
);

FILL FILL_6__11758_ (
);

FILL FILL_6__11338_ (
);

FILL FILL_4__12372_ (
);

FILL FILL_2__6952_ (
);

FILL FILL_3__11785_ (
);

FILL FILL_5__9402_ (
);

FILL FILL_3__11365_ (
);

FILL FILL_4__6878_ (
);

FILL FILL_0__16257_ (
);

NAND3X1 _16122_ (
    .A(_6570_),
    .B(_6575_),
    .C(_6566_),
    .Y(_6576_)
);

FILL FILL_2__10778_ (
);

FILL FILL_2__10358_ (
);

FILL FILL_0__11392_ (
);

FILL SFILL23720x12050 (
);

FILL FILL_5__14584_ (
);

FILL FILL_5__14164_ (
);

FILL FILL_6__7745_ (
);

OAI21X1 _8884_ (
    .A(_1017_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1018_),
    .Y(_978_[20])
);

OAI21X1 _8464_ (
    .A(_798_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .C(_799_),
    .Y(_783_[8])
);

DFFSR _8044_ (
    .Q(\datapath_1.regfile_1.regOut[9] [22]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_523_[22])
);

FILL FILL_4__13997_ (
);

FILL FILL_4__13577_ (
);

FILL FILL_4__13157_ (
);

FILL SFILL48920x61050 (
);

FILL FILL_2__14191_ (
);

FILL FILL_2__7737_ (
);

FILL FILL_2__7317_ (
);

FILL FILL_6__13904_ (
);

FILL SFILL23640x19050 (
);

FILL FILL_0__12597_ (
);

OAI21X1 _12882_ (
    .A(_3592_),
    .B(vdd),
    .C(_3593_),
    .Y(_3555_[19])
);

OAI21X1 _12462_ (
    .A(_3373_),
    .B(vdd),
    .C(_3374_),
    .Y(_3360_[7])
);

FILL FILL_0__12177_ (
);

NAND3X1 _12042_ (
    .A(_3075_),
    .B(_3076_),
    .C(_3077_),
    .Y(\datapath_1.mux_pcsrc.dout [13])
);

FILL FILL_3__13931_ (
);

FILL FILL_3__13511_ (
);

FILL FILL_4__8604_ (
);

FILL SFILL8680x18050 (
);

FILL FILL_5_BUFX2_insert530 (
);

FILL SFILL13720x55050 (
);

FILL FILL_5__15789_ (
);

FILL FILL_5_BUFX2_insert531 (
);

FILL FILL_5_BUFX2_insert532 (
);

FILL FILL_5__15369_ (
);

FILL FILL_2__12504_ (
);

FILL FILL_5_BUFX2_insert533 (
);

FILL FILL_5_BUFX2_insert534 (
);

NAND2X1 _9669_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1420_)
);

FILL FILL_5_BUFX2_insert535 (
);

NAND2X1 _9249_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1201_)
);

FILL FILL_5_BUFX2_insert536 (
);

FILL FILL_5_BUFX2_insert537 (
);

FILL FILL_5_BUFX2_insert538 (
);

FILL FILL_1__11917_ (
);

FILL FILL_5_BUFX2_insert539 (
);

FILL FILL_2__15396_ (
);

FILL FILL_5__16310_ (
);

FILL FILL_0__8504_ (
);

FILL SFILL13320x41050 (
);

FILL FILL_1__14389_ (
);

FILL FILL_5__6947_ (
);

FILL FILL_4__15723_ (
);

FILL FILL_1_BUFX2_insert1060 (
);

FILL FILL_4__15303_ (
);

FILL FILL_1_BUFX2_insert1061 (
);

FILL FILL_1_BUFX2_insert1062 (
);

FILL FILL_1_BUFX2_insert1063 (
);

FILL FILL_3__9493_ (
);

FILL FILL_1_BUFX2_insert1064 (
);

INVX1 _13667_ (
    .A(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_4175_)
);

NOR2X1 _13247_ (
    .A(\datapath_1.a3 [4]),
    .B(_3789_),
    .Y(_3790_)
);

FILL FILL_1_BUFX2_insert1065 (
);

FILL FILL_1_BUFX2_insert1066 (
);

FILL FILL_3__14716_ (
);

FILL FILL_1_BUFX2_insert1067 (
);

FILL FILL_1_BUFX2_insert1068 (
);

FILL FILL_1__15750_ (
);

FILL FILL_1__15330_ (
);

FILL FILL_1_BUFX2_insert1069 (
);

FILL FILL_1__6939_ (
);

FILL FILL_4__9809_ (
);

FILL SFILL8600x16050 (
);

FILL FILL_2__13709_ (
);

FILL SFILL34600x51050 (
);

FILL FILL_0__14743_ (
);

FILL FILL_0__14323_ (
);

FILL SFILL13720x10050 (
);

FILL FILL_2__7490_ (
);

FILL FILL_5__11289_ (
);

FILL FILL_2__7070_ (
);

FILL FILL_3__7806_ (
);

FILL FILL_5__12650_ (
);

FILL FILL_5__12230_ (
);

INVX1 _6950_ (
    .A(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_34_)
);

FILL FILL_2_BUFX2_insert660 (
);

FILL FILL_2_BUFX2_insert661 (
);

FILL FILL_2_BUFX2_insert662 (
);

FILL FILL_2_BUFX2_insert663 (
);

FILL FILL_2_BUFX2_insert664 (
);

FILL FILL_4__11643_ (
);

FILL FILL_4__11223_ (
);

FILL FILL_2_BUFX2_insert665 (
);

FILL FILL_2_BUFX2_insert666 (
);

FILL FILL_2_BUFX2_insert667 (
);

FILL SFILL13640x17050 (
);

FILL FILL_2_BUFX2_insert668 (
);

FILL FILL_2_BUFX2_insert669 (
);

FILL FILL_1__16115_ (
);

FILL FILL_3__10636_ (
);

FILL FILL_1__11670_ (
);

FILL FILL_1__11250_ (
);

FILL FILL_0__15948_ (
);

FILL FILL_0__15528_ (
);

OAI22X1 _15813_ (
    .A(_5489__bF$buf0),
    .B(_4885_),
    .C(_5527__bF$buf2),
    .D(_4874_),
    .Y(_6274_)
);

FILL FILL_0__15108_ (
);

FILL SFILL38840x66050 (
);

FILL FILL_2__8695_ (
);

FILL FILL_0__10663_ (
);

FILL FILL_2__8275_ (
);

FILL FILL_0__10243_ (
);

FILL FILL_6__14022_ (
);

FILL FILL_5__13855_ (
);

FILL FILL_5__13435_ (
);

FILL FILL_5__13015_ (
);

OAI21X1 _7735_ (
    .A(_434_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_435_),
    .Y(_393_[21])
);

OAI21X1 _7315_ (
    .A(_215_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .C(_216_),
    .Y(_198_[9])
);

FILL FILL_4__9982_ (
);

FILL FILL_4__9142_ (
);

FILL FILL_4__12848_ (
);

FILL FILL_4__12428_ (
);

FILL FILL_2__13882_ (
);

FILL FILL_2__13462_ (
);

FILL FILL_4__12008_ (
);

FILL FILL_2__13042_ (
);

FILL FILL_6__9488_ (
);

FILL FILL112200x53050 (
);

FILL FILL_1__12875_ (
);

FILL SFILL99480x46050 (
);

FILL FILL_1__12455_ (
);

FILL FILL_1__12035_ (
);

FILL FILL_6_CLKBUF1_insert111 (
);

FILL FILL_0__9882_ (
);

FILL FILL_0__9462_ (
);

FILL FILL_0__11868_ (
);

FILL FILL_0__9042_ (
);

FILL FILL_6_CLKBUF1_insert116 (
);

OAI21X1 _11733_ (
    .A(_2387_),
    .B(_2480_),
    .C(_2829_),
    .Y(_2830_)
);

FILL FILL_0__11448_ (
);

FILL FILL_0__11028_ (
);

NAND2X1 _11313_ (
    .A(_2431_),
    .B(_2412_),
    .Y(_2432_)
);

FILL SFILL38840x21050 (
);

FILL FILL_5__7485_ (
);

FILL FILL_5__7065_ (
);

FILL FILL_4__16261_ (
);

FILL FILL_6__10362_ (
);

FILL FILL_3__15674_ (
);

FILL FILL_3__15254_ (
);

FILL SFILL78920x17050 (
);

FILL FILL_1__7477_ (
);

FILL FILL_1__7057_ (
);

FILL FILL_2__14667_ (
);

FILL FILL_2__14247_ (
);

FILL FILL_0__15281_ (
);

FILL FILL_1_BUFX2_insert680 (
);

FILL FILL_3__8764_ (
);

FILL FILL_1_BUFX2_insert681 (
);

FILL FILL_3__8344_ (
);

DFFSR _12938_ (
    .Q(\datapath_1.a [19]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3555_[19])
);

FILL FILL_1_BUFX2_insert682 (
);

NAND2X1 _12518_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [26]),
    .Y(_3412_)
);

FILL FILL_1_BUFX2_insert683 (
);

FILL FILL_1_BUFX2_insert684 (
);

FILL FILL_1_BUFX2_insert685 (
);

FILL FILL_1_BUFX2_insert686 (
);

FILL FILL_1__14601_ (
);

FILL FILL_1_BUFX2_insert687 (
);

FILL FILL_1_BUFX2_insert688 (
);

FILL FILL_1_BUFX2_insert689 (
);

FILL FILL_4__12181_ (
);

FILL FILL_3__16039_ (
);

FILL SFILL33800x47050 (
);

FILL SFILL64200x38050 (
);

FILL FILL_3__11594_ (
);

FILL FILL_5__9631_ (
);

FILL FILL_5__9211_ (
);

FILL FILL_3__11174_ (
);

FILL SFILL28440x50050 (
);

FILL FILL_0__16066_ (
);

INVX1 _16351_ (
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_6788_)
);

FILL FILL_2__10167_ (
);

FILL FILL_5__11921_ (
);

FILL FILL_1__9623_ (
);

FILL FILL_5__11501_ (
);

FILL SFILL89480x44050 (
);

FILL FILL_3__9549_ (
);

FILL FILL_4__10914_ (
);

FILL FILL_3__9129_ (
);

FILL FILL_5__14393_ (
);

FILL FILL_1__15806_ (
);

DFFSR _8693_ (
    .Q(\datapath_1.regfile_1.regOut[14] [31]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_848_[31])
);

NAND2X1 _8273_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_713_)
);

FILL FILL_1__10941_ (
);

FILL FILL_4__13386_ (
);

FILL FILL_1__10521_ (
);

FILL FILL_2__7966_ (
);

BUFX2 BUFX2_insert350 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf1)
);

FILL FILL_2__7546_ (
);

FILL FILL_3__12379_ (
);

BUFX2 BUFX2_insert351 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf0)
);

BUFX2 BUFX2_insert352 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf7 )
);

BUFX2 BUFX2_insert353 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf6 )
);

BUFX2 BUFX2_insert354 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf5 )
);

BUFX2 BUFX2_insert355 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf4 )
);

BUFX2 BUFX2_insert356 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf3 )
);

BUFX2 BUFX2_insert357 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf2 )
);

BUFX2 BUFX2_insert358 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf1 )
);

DFFSR _12691_ (
    .Q(\datapath_1.Data [28]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3425_[28])
);

BUFX2 BUFX2_insert359 (
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf0 )
);

NAND3X1 _12271_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3242_)
);

FILL FILL_5__12706_ (
);

FILL FILL_3__13740_ (
);

FILL FILL_3__13320_ (
);

FILL FILL_4__8833_ (
);

FILL FILL_2__12733_ (
);

FILL FILL_5__15598_ (
);

FILL FILL_5__15178_ (
);

FILL FILL_2__12313_ (
);

FILL FILL_6__8759_ (
);

NAND2X1 _9898_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1532_)
);

NAND2X1 _9478_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1313_)
);

DFFSR _9058_ (
    .Q(\datapath_1.regfile_1.regOut[17] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_1043_[12])
);

FILL FILL_1__11726_ (
);

FILL FILL_1__11306_ (
);

FILL FILL_0__8733_ (
);

FILL FILL_0__8313_ (
);

FILL FILL_1__14198_ (
);

FILL FILL_4__15952_ (
);

FILL FILL_4__15532_ (
);

FILL FILL_4__15112_ (
);

AOI22X1 _13896_ (
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .B(_3942__bF$buf3),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_4399_)
);

AOI21X1 _13476_ (
    .A(_3940_),
    .B(_3987_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [0])
);

DFFSR _13056_ (
    .Q(_2_[9]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_3620_[9])
);

FILL FILL_3__14945_ (
);

FILL FILL_3__14525_ (
);

FILL FILL_3__14105_ (
);

FILL FILL_4__9618_ (
);

FILL FILL_2__13938_ (
);

FILL FILL_0__14972_ (
);

FILL FILL_2__13518_ (
);

FILL FILL_0__14552_ (
);

FILL FILL_0__14132_ (
);

FILL FILL_5__11098_ (
);

FILL SFILL48600x80050 (
);

FILL FILL_0__9938_ (
);

FILL FILL_3__7615_ (
);

FILL FILL_0__9518_ (
);

FILL FILL_4__16317_ (
);

FILL FILL_4__11872_ (
);

FILL SFILL109640x68050 (
);

FILL FILL_4__11452_ (
);

FILL FILL_4__11032_ (
);

FILL FILL_6__8092_ (
);

FILL FILL_1__16344_ (
);

FILL FILL_5__8902_ (
);

FILL FILL_3__10445_ (
);

FILL FILL_3__10025_ (
);

FILL FILL_0__15757_ (
);

FILL FILL_0__15337_ (
);

OAI22X1 _15622_ (
    .A(_5544__bF$buf1),
    .B(_6087_),
    .C(_5545__bF$buf2),
    .D(_4654_),
    .Y(_6088_)
);

NAND3X1 _15202_ (
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf4),
    .Y(_5679_)
);

FILL FILL_0__10892_ (
);

FILL FILL_2__8084_ (
);

FILL FILL_0__10052_ (
);

FILL FILL_5__13664_ (
);

FILL FILL_5__13244_ (
);

OAI21X1 _7964_ (
    .A(_546_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .C(_547_),
    .Y(_523_[12])
);

OAI21X1 _7544_ (
    .A(_391_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .C(_392_),
    .Y(_328_[0])
);

FILL SFILL69080x71050 (
);

NAND2X1 _7124_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_130_)
);

FILL FILL_4__9791_ (
);

FILL FILL_4__9371_ (
);

FILL FILL_4__12657_ (
);

FILL SFILL48920x56050 (
);

FILL FILL_4__12237_ (
);

FILL FILL_2__13691_ (
);

FILL FILL_2__13271_ (
);

FILL FILL_1__12264_ (
);

OAI21X1 _16407_ (
    .A(_6824_),
    .B(gnd),
    .C(_6825_),
    .Y(_6769_[28])
);

FILL FILL_0__9271_ (
);

INVX1 _11962_ (
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3016_)
);

FILL FILL_2__9289_ (
);

FILL FILL_0__11677_ (
);

FILL FILL_0__11257_ (
);

NAND3X1 _11542_ (
    .A(_2220_),
    .B(_2634_),
    .C(_2636_),
    .Y(_2652_)
);

INVX2 _11122_ (
    .A(_2240_),
    .Y(_2241_)
);

FILL FILL_5__7294_ (
);

FILL FILL_4__16070_ (
);

FILL FILL_5__14869_ (
);

FILL FILL_5__14449_ (
);

FILL FILL_5__14029_ (
);

FILL FILL_3__15483_ (
);

FILL FILL_3__15063_ (
);

NAND2X1 _8749_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_949_)
);

NAND2X1 _8329_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_730_)
);

FILL FILL_1__7286_ (
);

FILL FILL_2__14896_ (
);

FILL FILL_2__14476_ (
);

FILL FILL_2__14056_ (
);

FILL FILL_0__15090_ (
);

FILL FILL_5__15810_ (
);

FILL SFILL48920x11050 (
);

FILL FILL_1__13889_ (
);

FILL FILL_1__13469_ (
);

FILL FILL_4__14803_ (
);

FILL FILL_3__8993_ (
);

FILL FILL_3__8573_ (
);

NAND2X1 _12747_ (
    .A(IRWrite_bF$buf5),
    .B(memoryOutData[17]),
    .Y(_3524_)
);

NAND3X1 _12327_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3284_)
);

FILL FILL_1__14830_ (
);

FILL FILL_5__8499_ (
);

FILL FILL_5__8079_ (
);

FILL FILL_1__14410_ (
);

FILL FILL_0__13823_ (
);

FILL FILL_0__13403_ (
);

FILL FILL_3__16268_ (
);

FILL SFILL99560x79050 (
);

FILL FILL_2__6990_ (
);

FILL FILL_5__10789_ (
);

FILL FILL_5__10369_ (
);

FILL FILL_5__9860_ (
);

FILL FILL_5__9020_ (
);

FILL FILL_0__16295_ (
);

OAI22X1 _16160_ (
    .A(_5485__bF$buf0),
    .B(_6612_),
    .C(_5244_),
    .D(_5549__bF$buf1),
    .Y(_6613_)
);

FILL FILL_2__10396_ (
);

FILL FILL_5__11730_ (
);

FILL FILL_1__9852_ (
);

FILL FILL_5__11310_ (
);

FILL FILL_1__9012_ (
);

FILL FILL_2__16202_ (
);

FILL FILL_3__9778_ (
);

FILL FILL_3__9358_ (
);

FILL FILL_4__10303_ (
);

FILL FILL_1__15615_ (
);

FILL FILL_6__7363_ (
);

NAND2X1 _8082_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_606_)
);

FILL SFILL38520x40050 (
);

FILL FILL_1__10750_ (
);

FILL FILL_0__14608_ (
);

FILL FILL_2__7355_ (
);

FILL FILL_3__12188_ (
);

FILL SFILL3560x53050 (
);

NAND3X1 _12080_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [23]),
    .C(_3034__bF$buf2),
    .Y(_3106_)
);

FILL FILL_5__12515_ (
);

FILL SFILL104440x70050 (
);

FILL FILL_4__8642_ (
);

FILL FILL_5_BUFX2_insert910 (
);

FILL FILL_4__11928_ (
);

FILL FILL_4__8222_ (
);

FILL FILL_2__12962_ (
);

FILL FILL_5_BUFX2_insert911 (
);

FILL FILL_4__11508_ (
);

FILL FILL_5_BUFX2_insert912 (
);

FILL FILL_2__12122_ (
);

FILL FILL_5_BUFX2_insert913 (
);

FILL FILL_6__8568_ (
);

FILL FILL_5_BUFX2_insert914 (
);

FILL FILL_6__8148_ (
);

INVX1 _9287_ (
    .A(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_1226_)
);

FILL FILL_5_BUFX2_insert915 (
);

FILL FILL_5_BUFX2_insert916 (
);

FILL FILL112200x48050 (
);

FILL FILL_5_BUFX2_insert917 (
);

FILL FILL_5_BUFX2_insert918 (
);

FILL FILL_1__11955_ (
);

FILL FILL_5_BUFX2_insert919 (
);

FILL FILL_1__11535_ (
);

FILL FILL_1__11115_ (
);

FILL FILL_0__8962_ (
);

FILL FILL_0__10948_ (
);

OAI21X1 _10813_ (
    .A(_1998_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1999_),
    .Y(_1953_[23])
);

FILL FILL_0__8122_ (
);

FILL FILL_0__10528_ (
);

FILL FILL_0__10108_ (
);

FILL SFILL89560x77050 (
);

FILL SFILL38840x16050 (
);

FILL FILL_5__6985_ (
);

FILL FILL_4__15761_ (
);

FILL FILL_4__15341_ (
);

NAND3X1 _13285_ (
    .A(_3821_),
    .B(_3817_),
    .C(_3823_),
    .Y(_3824_)
);

FILL FILL_2__9921_ (
);

FILL FILL_3__14754_ (
);

FILL FILL_2__9501_ (
);

FILL FILL_3__14334_ (
);

FILL SFILL28920x52050 (
);

FILL FILL_1__6977_ (
);

FILL FILL_4__9847_ (
);

FILL FILL_4__9427_ (
);

FILL FILL_4__9007_ (
);

FILL FILL_2__13747_ (
);

FILL SFILL89160x63050 (
);

FILL FILL_2__13327_ (
);

FILL FILL_0__14781_ (
);

FILL FILL_0__14361_ (
);

FILL SFILL64920x4050 (
);

FILL FILL_3__7844_ (
);

FILL FILL_0__9747_ (
);

FILL FILL_3__7424_ (
);

FILL SFILL28840x59050 (
);

FILL FILL_4__16126_ (
);

FILL FILL_4__11681_ (
);

FILL FILL_4__11261_ (
);

FILL FILL_3__15959_ (
);

FILL FILL_3__15539_ (
);

FILL FILL_3__15119_ (
);

FILL FILL_1__16153_ (
);

FILL FILL_3__10674_ (
);

FILL FILL_5__8711_ (
);

FILL FILL_3__10254_ (
);

FILL FILL_0__15986_ (
);

FILL FILL_0__15566_ (
);

NOR3X1 _15851_ (
    .A(_6301_),
    .B(_6288_),
    .C(_6311_),
    .Y(_6312_)
);

FILL FILL_0__15146_ (
);

OAI22X1 _15431_ (
    .A(_4406_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf3),
    .D(_5901_),
    .Y(_5902_)
);

NAND2X1 _15011_ (
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .B(_5490_),
    .Y(_5491_)
);

FILL FILL_0__10281_ (
);

FILL FILL_1__8703_ (
);

FILL FILL_3__8629_ (
);

FILL FILL_3__8209_ (
);

FILL FILL_5__13893_ (
);

FILL FILL_5__13473_ (
);

DFFSR _7773_ (
    .Q(\datapath_1.regfile_1.regOut[7] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_393_[7])
);

NAND2X1 _7353_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_242_)
);

FILL FILL_4__12886_ (
);

FILL SFILL28840x14050 (
);

FILL FILL_4__12466_ (
);

FILL SFILL94360x81050 (
);

FILL FILL_4__12046_ (
);

FILL FILL_2__13080_ (
);

FILL FILL_5__9916_ (
);

FILL FILL_3__11879_ (
);

FILL FILL_3__11459_ (
);

FILL FILL_1__12493_ (
);

FILL FILL_3__11039_ (
);

FILL FILL_1__12073_ (
);

NAND2X1 _16216_ (
    .A(\datapath_1.PCJump [26]),
    .B(_5470_),
    .Y(_6667_)
);

FILL FILL_2__9098_ (
);

FILL FILL_0__9080_ (
);

OAI21X1 _11771_ (
    .A(_2364_),
    .B(_2864_),
    .C(_2865_),
    .Y(_2866_)
);

FILL FILL_0__11486_ (
);

FILL SFILL79160x61050 (
);

AND2X2 _11351_ (
    .A(_2456_),
    .B(_2117_),
    .Y(_2469_)
);

FILL FILL_0__11066_ (
);

FILL FILL_1__9908_ (
);

FILL FILL_6__15685_ (
);

FILL FILL_3__12400_ (
);

FILL FILL_6__15265_ (
);

FILL FILL_2__11813_ (
);

FILL FILL_5__14678_ (
);

FILL FILL_5__14258_ (
);

NAND2X1 _8978_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1061_)
);

FILL FILL_3__15292_ (
);

FILL FILL_6__7839_ (
);

DFFSR _8558_ (
    .Q(\datapath_1.regfile_1.regOut[13] [24]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_783_[24])
);

INVX1 _8138_ (
    .A(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_643_)
);

FILL FILL_1__7095_ (
);

FILL FILL_1__10806_ (
);

FILL SFILL18840x57050 (
);

FILL FILL_2__14285_ (
);

FILL FILL_0__7813_ (
);

FILL FILL_1__13698_ (
);

FILL FILL_1__13278_ (
);

FILL FILL_4__14612_ (
);

NAND2X1 _12976_ (
    .A(vdd),
    .B(\datapath_1.rd2 [8]),
    .Y(_3636_)
);

FILL FILL_3__8382_ (
);

DFFSR _12556_ (
    .Q(ALUOut[21]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3360_[21])
);

INVX1 _12136_ (
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_3144_)
);

FILL FILL_3__13605_ (
);

FILL FILL_6__11185_ (
);

FILL FILL_0__13632_ (
);

FILL FILL_0__13212_ (
);

FILL FILL_3__16077_ (
);

FILL FILL_5__10178_ (
);

FILL FILL_5__16404_ (
);

FILL SFILL18840x12050 (
);

FILL FILL_1__9661_ (
);

FILL FILL_1__9241_ (
);

FILL FILL_4__15817_ (
);

FILL FILL_2__16011_ (
);

FILL FILL_4__10952_ (
);

FILL FILL_3__9167_ (
);

FILL FILL_4__10532_ (
);

FILL FILL_4__10112_ (
);

FILL FILL_1__15844_ (
);

FILL FILL_6__7172_ (
);

FILL FILL_1__15424_ (
);

FILL FILL_1__15004_ (
);

FILL FILL_0__14837_ (
);

NAND3X1 _14702_ (
    .A(_5179_),
    .B(_5180_),
    .C(_5187_),
    .Y(_5188_)
);

FILL FILL_0__14417_ (
);

FILL FILL_2__7584_ (
);

BUFX2 BUFX2_insert730 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf2 )
);

BUFX2 BUFX2_insert731 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf1 )
);

FILL FILL_2__7164_ (
);

BUFX2 BUFX2_insert732 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf0 )
);

BUFX2 BUFX2_insert733 (
    .A(_5500_),
    .Y(_5500__bF$buf3)
);

FILL FILL_6__13751_ (
);

BUFX2 BUFX2_insert734 (
    .A(_5500_),
    .Y(_5500__bF$buf2)
);

FILL FILL_6__13331_ (
);

BUFX2 BUFX2_insert735 (
    .A(_5500_),
    .Y(_5500__bF$buf1)
);

BUFX2 BUFX2_insert736 (
    .A(_5500_),
    .Y(_5500__bF$buf0)
);

BUFX2 BUFX2_insert737 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf4 )
);

BUFX2 BUFX2_insert738 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf3 )
);

BUFX2 BUFX2_insert739 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf2 )
);

FILL FILL_5__12744_ (
);

FILL FILL_5__12324_ (
);

FILL SFILL69080x66050 (
);

FILL FILL_4__8871_ (
);

FILL FILL_4__8451_ (
);

FILL FILL_4__11737_ (
);

FILL FILL_2__12771_ (
);

FILL FILL_4__11317_ (
);

FILL FILL_2__12351_ (
);

FILL FILL_1__16209_ (
);

INVX1 _9096_ (
    .A(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_1119_)
);

FILL FILL_1__11764_ (
);

FILL FILL_1__11344_ (
);

OAI22X1 _15907_ (
    .A(_6365_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf0),
    .D(_4975_),
    .Y(_6366_)
);

FILL FILL_2__8789_ (
);

FILL FILL_0__8771_ (
);

FILL FILL_2__8369_ (
);

FILL FILL_0__10757_ (
);

FILL FILL_0__8351_ (
);

OAI21X1 _10622_ (
    .A(_1891_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1892_),
    .Y(_1888_[2])
);

FILL SFILL114520x60050 (
);

DFFSR _10202_ (
    .Q(\datapath_1.regfile_1.regOut[26] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_1628_[4])
);

FILL SFILL53880x50050 (
);

FILL FILL_4__15990_ (
);

FILL FILL_4__15570_ (
);

FILL FILL_4__15150_ (
);

INVX1 _13094_ (
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_3694_)
);

FILL FILL_5__13949_ (
);

FILL FILL_2__9730_ (
);

FILL FILL_3__14983_ (
);

FILL FILL_5__13529_ (
);

FILL FILL_3__14563_ (
);

FILL FILL_5__13109_ (
);

FILL FILL_3__14143_ (
);

NAND2X1 _7829_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_478_)
);

DFFSR _7409_ (
    .Q(\datapath_1.regfile_1.regOut[4] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_198_[27])
);

FILL FILL_4_BUFX2_insert570 (
);

FILL FILL_4__9656_ (
);

FILL FILL_4_BUFX2_insert571 (
);

FILL FILL_4_BUFX2_insert572 (
);

FILL FILL_4__9236_ (
);

FILL FILL_4_BUFX2_insert573 (
);

FILL FILL_2__13976_ (
);

FILL FILL_2__13556_ (
);

FILL FILL_4_BUFX2_insert574 (
);

FILL FILL_0__14590_ (
);

FILL FILL_4_BUFX2_insert575 (
);

FILL FILL_2__13136_ (
);

FILL FILL_0__14170_ (
);

FILL FILL_4_BUFX2_insert576 (
);

FILL FILL_4_BUFX2_insert577 (
);

FILL FILL_4_BUFX2_insert578 (
);

FILL FILL_4_BUFX2_insert579 (
);

FILL FILL_1__12969_ (
);

FILL FILL_1__12129_ (
);

FILL FILL_0__9976_ (
);

FILL FILL_0__9556_ (
);

FILL FILL_0__9136_ (
);

OAI21X1 _11827_ (
    .A(_2353_),
    .B(_2359_),
    .C(_2916_),
    .Y(_2917_)
);

FILL FILL_3__7233_ (
);

OAI21X1 _11407_ (
    .A(_2523_),
    .B(_2249_),
    .C(_2274_),
    .Y(_2524_)
);

FILL FILL_5__7999_ (
);

FILL FILL_5__7579_ (
);

FILL FILL_1__13910_ (
);

FILL FILL_4__16355_ (
);

FILL FILL_5__7159_ (
);

INVX1 _14299_ (
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_4794_)
);

FILL FILL_4__11490_ (
);

FILL FILL_6__10036_ (
);

FILL FILL_4__11070_ (
);

FILL FILL_0__12903_ (
);

FILL FILL_3__15768_ (
);

FILL FILL_3__15348_ (
);

FILL FILL_1__16382_ (
);

FILL FILL_5__8520_ (
);

FILL FILL_5__8100_ (
);

FILL FILL_3__10063_ (
);

FILL SFILL59080x64050 (
);

FILL FILL_0__15795_ (
);

FILL FILL_0__15375_ (
);

NAND3X1 _15660_ (
    .A(_6117_),
    .B(_6124_),
    .C(_6123_),
    .Y(_6125_)
);

NOR2X1 _15240_ (
    .A(_5715_),
    .B(_5712_),
    .Y(_5716_)
);

FILL SFILL38920x49050 (
);

FILL FILL_5__10810_ (
);

FILL FILL_1__8512_ (
);

FILL FILL_2__15702_ (
);

FILL FILL_3__8858_ (
);

FILL FILL_3__8438_ (
);

FILL FILL_3__8018_ (
);

FILL SFILL3640x41050 (
);

FILL FILL_5__13282_ (
);

FILL FILL_6__6863_ (
);

NAND2X1 _7582_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_354_)
);

NAND2X1 _7162_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_135_)
);

FILL FILL_4__12695_ (
);

FILL FILL_4__12275_ (
);

FILL FILL_2__6855_ (
);

FILL FILL_3__11688_ (
);

FILL FILL_5__9725_ (
);

FILL FILL_3__11268_ (
);

FILL SFILL59000x62050 (
);

DFFSR _16445_ (
    .Q(\datapath_1.regfile_1.regOut[0] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_6769_[28])
);

INVX1 _16025_ (
    .A(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_6481_)
);

INVX1 _11580_ (
    .A(_2687_),
    .Y(\datapath_1.ALUResult [20])
);

FILL FILL_0__11295_ (
);

INVX1 _11160_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .Y(_2279_)
);

FILL SFILL104440x65050 (
);

FILL FILL_3_BUFX2_insert590 (
);

FILL FILL_4__7722_ (
);

FILL FILL_3_BUFX2_insert591 (
);

FILL FILL_4__7302_ (
);

FILL FILL_3_BUFX2_insert592 (
);

FILL FILL_5__14487_ (
);

FILL FILL_3_BUFX2_insert593 (
);

FILL FILL_2__11622_ (
);

FILL FILL_3_BUFX2_insert594 (
);

FILL FILL_5__14067_ (
);

FILL FILL_2__11202_ (
);

FILL FILL_3_BUFX2_insert595 (
);

INVX1 _8787_ (
    .A(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_974_)
);

FILL FILL_3_BUFX2_insert596 (
);

INVX1 _8367_ (
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_755_)
);

FILL FILL_3_BUFX2_insert597 (
);

FILL FILL_3_BUFX2_insert598 (
);

FILL FILL_3_BUFX2_insert599 (
);

FILL FILL_1__10615_ (
);

FILL FILL_2__14094_ (
);

FILL FILL_0__7622_ (
);

FILL FILL_0__7202_ (
);

FILL FILL_1__13087_ (
);

FILL FILL_6__13807_ (
);

FILL FILL_4__14841_ (
);

FILL FILL_4__14421_ (
);

FILL FILL_4__14001_ (
);

FILL SFILL43960x6050 (
);

INVX1 _12785_ (
    .A(\control_1.op [4]),
    .Y(_3549_)
);

FILL FILL_3__8191_ (
);

FILL SFILL49080x62050 (
);

NAND2X1 _12365_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [7]),
    .Y(_3309_)
);

FILL FILL_3__13834_ (
);

FILL FILL_3__13414_ (
);

FILL SFILL28920x47050 (
);

FILL FILL_4__8507_ (
);

FILL FILL_2__12827_ (
);

FILL SFILL104440x20050 (
);

FILL FILL_2__12407_ (
);

FILL FILL_0__13861_ (
);

FILL FILL_0__13441_ (
);

FILL FILL_0__13021_ (
);

FILL FILL_2__15299_ (
);

FILL FILL_5__16213_ (
);

FILL FILL_3__6924_ (
);

FILL FILL_0__8827_ (
);

FILL FILL_1__9890_ (
);

FILL FILL_1__9470_ (
);

FILL FILL_4__15626_ (
);

FILL FILL_4__15206_ (
);

FILL FILL_2__16240_ (
);

FILL FILL_3__9396_ (
);

FILL SFILL49000x60050 (
);

FILL FILL_4__10761_ (
);

FILL FILL_3__14619_ (
);

FILL FILL_1__15653_ (
);

FILL FILL_1__15233_ (
);

FILL FILL_0__14646_ (
);

AOI22X1 _14931_ (
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .B(_4005__bF$buf1),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_5412_)
);

FILL FILL_0__14226_ (
);

AOI22X1 _14511_ (
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .B(_4135_),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_5001_)
);

FILL SFILL58920x50 (
);

FILL FILL_3__7709_ (
);

FILL FILL_5__12973_ (
);

FILL FILL_5__12133_ (
);

BUFX2 _6853_ (
    .A(_1_[15]),
    .Y(memoryAddress[15])
);

FILL FILL_4__11966_ (
);

FILL FILL_4__8260_ (
);

FILL SFILL94360x76050 (
);

FILL FILL_4__11546_ (
);

FILL FILL_2__12580_ (
);

FILL FILL_4__11126_ (
);

FILL FILL_2__12160_ (
);

FILL FILL_6__8186_ (
);

FILL FILL_1__16018_ (
);

FILL FILL_3__10959_ (
);

FILL FILL_3__10539_ (
);

FILL FILL_1__11993_ (
);

FILL FILL_1__11573_ (
);

FILL FILL_3__10119_ (
);

FILL FILL_1__11153_ (
);

INVX1 _15716_ (
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_6180_)
);

FILL FILL_0__8580_ (
);

FILL FILL_2__8598_ (
);

FILL SFILL79160x56050 (
);

FILL FILL_0__10566_ (
);

DFFSR _10851_ (
    .Q(\datapath_1.regfile_1.regOut[31] [13]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_1953_[13])
);

NAND2X1 _10431_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1806_)
);

FILL FILL_0__10146_ (
);

NAND2X1 _10011_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1587_)
);

FILL FILL_3__11900_ (
);

FILL FILL_5__13758_ (
);

FILL SFILL18040x69050 (
);

FILL FILL_5__13338_ (
);

FILL FILL_3__14792_ (
);

FILL FILL_3__14372_ (
);

FILL FILL_6__6919_ (
);

DFFSR _7638_ (
    .Q(\datapath_1.regfile_1.regOut[6] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_328_[0])
);

INVX1 _7218_ (
    .A(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_172_)
);

FILL FILL_4__9885_ (
);

FILL FILL_4__9465_ (
);

FILL FILL_4__9045_ (
);

FILL FILL_2__13785_ (
);

FILL FILL_2__13365_ (
);

FILL FILL_1__12778_ (
);

FILL FILL_1__12358_ (
);

FILL FILL_3__7882_ (
);

FILL FILL_0__9785_ (
);

FILL FILL_3__7462_ (
);

FILL FILL_0__9365_ (
);

FILL FILL_3__7042_ (
);

AOI21X1 _11636_ (
    .A(_2720_),
    .B(_2408_),
    .C(_2458_),
    .Y(_2740_)
);

INVX1 _11216_ (
    .A(ALUControl[2]),
    .Y(_2335_)
);

FILL SFILL79160x11050 (
);

FILL FILL_4__16164_ (
);

FILL FILL_3__15997_ (
);

FILL FILL_0__12712_ (
);

FILL FILL_3__15577_ (
);

FILL FILL_3__15157_ (
);

FILL FILL_1__16191_ (
);

FILL FILL_3__10292_ (
);

FILL FILL_0__15184_ (
);

FILL FILL_5__15904_ (
);

FILL SFILL53960x83050 (
);

FILL SFILL84360x74050 (
);

FILL FILL_1__8741_ (
);

FILL SFILL79080x18050 (
);

FILL FILL_1__8321_ (
);

FILL FILL_2__15931_ (
);

FILL FILL_2__15511_ (
);

FILL FILL_3__8247_ (
);

FILL FILL_5__13091_ (
);

FILL FILL_1__14924_ (
);

FILL FILL_1__14504_ (
);

DFFSR _7391_ (
    .Q(\datapath_1.regfile_1.regOut[4] [9]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_198_[9])
);

FILL FILL_4__12084_ (
);

FILL FILL_0__13917_ (
);

FILL FILL_5__9534_ (
);

FILL FILL_3__11497_ (
);

FILL FILL_5__9114_ (
);

FILL FILL_3__11077_ (
);

FILL FILL_6__12831_ (
);

FILL FILL_0__16389_ (
);

OAI22X1 _16254_ (
    .A(_5526__bF$buf1),
    .B(_5404_),
    .C(_5385_),
    .D(_5527__bF$buf2),
    .Y(_6704_)
);

FILL FILL_5__11824_ (
);

FILL FILL_1__9526_ (
);

FILL FILL_5__11404_ (
);

FILL FILL_1__9106_ (
);

FILL FILL_4__7951_ (
);

FILL SFILL114920x69050 (
);

FILL FILL_4__7111_ (
);

FILL FILL_4__10817_ (
);

FILL FILL_2__11851_ (
);

FILL FILL_5__14296_ (
);

FILL FILL_2__11431_ (
);

FILL FILL_2__11011_ (
);

FILL FILL_1__15709_ (
);

INVX1 _8596_ (
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_867_)
);

DFFSR _8176_ (
    .Q(\datapath_1.regfile_1.regOut[10] [26]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_588_[26])
);

FILL FILL_4__13289_ (
);

FILL FILL_1__10424_ (
);

FILL FILL_1__10004_ (
);

FILL FILL_2__7869_ (
);

FILL FILL_0__7851_ (
);

FILL FILL_2__7449_ (
);

FILL FILL_0__7431_ (
);

FILL FILL_4__14650_ (
);

FILL FILL_4__14230_ (
);

FILL SFILL3720x74050 (
);

INVX1 _12594_ (
    .A(\datapath_1.Data [9]),
    .Y(_3442_)
);

OAI21X1 _12174_ (
    .A(_3168_),
    .B(ALUSrcA_bF$buf1),
    .C(_3169_),
    .Y(\datapath_1.alu_1.ALUInA [19])
);

FILL FILL_5__12609_ (
);

FILL FILL_3__13643_ (
);

FILL SFILL43960x81050 (
);

FILL FILL_3__13223_ (
);

NAND2X1 _6909_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_7_)
);

FILL FILL_4__8736_ (
);

FILL FILL_4__8316_ (
);

FILL SFILL53480x31050 (
);

FILL SFILL69080x16050 (
);

FILL FILL_2__12636_ (
);

FILL FILL_0__13670_ (
);

FILL FILL_2__12216_ (
);

FILL FILL_0__13250_ (
);

FILL FILL_1__11629_ (
);

FILL FILL_1__11209_ (
);

FILL FILL_0__8636_ (
);

FILL FILL_5__16022_ (
);

NAND2X1 _10907_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2050_),
    .Y(_2054_)
);

FILL FILL_0__8216_ (
);

FILL FILL_4__15855_ (
);

FILL FILL_4__15435_ (
);

FILL SFILL114520x10050 (
);

FILL FILL_4__15015_ (
);

INVX1 _13799_ (
    .A(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_4304_)
);

FILL FILL_4__10990_ (
);

FILL FILL_4__10570_ (
);

INVX8 _13379_ (
    .A(_3890_),
    .Y(_3891_)
);

FILL FILL_4__10150_ (
);

FILL FILL_3__14848_ (
);

FILL FILL_1__15882_ (
);

FILL FILL_3__14428_ (
);

FILL FILL_3__14008_ (
);

FILL FILL_1__15462_ (
);

FILL FILL_1__15042_ (
);

FILL FILL_5__7600_ (
);

FILL SFILL59080x59050 (
);

FILL FILL_0__14875_ (
);

FILL FILL_0__14455_ (
);

NAND3X1 _14740_ (
    .A(_5224_),
    .B(_5225_),
    .C(_5223_),
    .Y(_5226_)
);

FILL FILL_0__14035_ (
);

OAI22X1 _14320_ (
    .A(_3947__bF$buf3),
    .B(_4813_),
    .C(_3935__bF$buf2),
    .D(_4812_),
    .Y(_4814_)
);

FILL FILL_3__7938_ (
);

FILL SFILL3640x36050 (
);

FILL FILL_5__12782_ (
);

FILL FILL_5__12362_ (
);

FILL SFILL43880x43050 (
);

FILL FILL_4__11775_ (
);

FILL FILL_4__11355_ (
);

FILL FILL_1__16247_ (
);

FILL FILL_3__10768_ (
);

FILL FILL_1__11382_ (
);

NAND3X1 _15945_ (
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf2),
    .Y(_6403_)
);

INVX1 _15525_ (
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_5994_)
);

INVX1 _15105_ (
    .A(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_5584_)
);

FILL SFILL59080x14050 (
);

FILL FILL_0__10795_ (
);

NAND2X1 _10660_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1918_)
);

FILL FILL_0__10375_ (
);

NAND2X1 _10240_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1699_)
);

FILL FILL_6__14994_ (
);

FILL FILL_6__14574_ (
);

FILL FILL_5__13987_ (
);

FILL FILL_2__10702_ (
);

FILL FILL_5__13567_ (
);

FILL FILL_5__13147_ (
);

INVX1 _7867_ (
    .A(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_503_)
);

FILL FILL_3__14181_ (
);

INVX1 _7447_ (
    .A(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_284_)
);

DFFSR _7027_ (
    .Q(\datapath_1.regfile_1.regOut[1] [29]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_3_[29])
);

FILL FILL_4_BUFX2_insert950 (
);

FILL FILL_4_BUFX2_insert951 (
);

FILL FILL_4__9274_ (
);

FILL FILL_4_BUFX2_insert952 (
);

FILL FILL_4_BUFX2_insert953 (
);

FILL FILL_4_BUFX2_insert954 (
);

FILL FILL_2__13594_ (
);

FILL FILL_4_BUFX2_insert955 (
);

FILL FILL_2__13174_ (
);

FILL FILL_4_BUFX2_insert956 (
);

FILL FILL_4_BUFX2_insert957 (
);

FILL FILL_4_BUFX2_insert958 (
);

FILL FILL_4_BUFX2_insert959 (
);

FILL FILL_1__12587_ (
);

FILL FILL_1__12167_ (
);

FILL FILL_4__13921_ (
);

FILL FILL_4__13501_ (
);

FILL FILL_3__7691_ (
);

FILL FILL_0__9594_ (
);

FILL SFILL49080x57050 (
);

NAND3X1 _11865_ (
    .A(_2950_),
    .B(_2951_),
    .C(_2945_),
    .Y(_2952_)
);

NOR2X1 _11445_ (
    .A(_2148_),
    .B(_2560_),
    .Y(_2561_)
);

NOR2X1 _11025_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2144_)
);

FILL FILL_3__12914_ (
);

FILL FILL_4__16393_ (
);

FILL FILL_5__7197_ (
);

FILL FILL_2__11907_ (
);

FILL FILL_3__15386_ (
);

FILL FILL_0__12521_ (
);

FILL FILL_0__12101_ (
);

FILL FILL_1__7189_ (
);

FILL FILL_2__14799_ (
);

FILL FILL_2__14379_ (
);

FILL SFILL33880x41050 (
);

FILL FILL_5__15713_ (
);

FILL FILL_1__8970_ (
);

FILL FILL_1__8130_ (
);

FILL FILL_4__14706_ (
);

FILL FILL_2__15740_ (
);

FILL FILL_3__8896_ (
);

FILL FILL_2__15320_ (
);

FILL SFILL49000x55050 (
);

FILL FILL_3__8476_ (
);

FILL FILL_3__8056_ (
);

FILL FILL_1__14733_ (
);

FILL FILL_1__14313_ (
);

FILL SFILL94440x64050 (
);

FILL FILL_0__13726_ (
);

FILL FILL_0__13306_ (
);

FILL FILL_2__6893_ (
);

FILL FILL_5__9763_ (
);

FILL FILL_5__9343_ (
);

FILL FILL_0_BUFX2_insert1070 (
);

FILL FILL_0_BUFX2_insert1071 (
);

FILL FILL_0_BUFX2_insert1072 (
);

FILL FILL_0_BUFX2_insert1073 (
);

FILL FILL_0__16198_ (
);

INVX1 _16063_ (
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_6518_)
);

FILL FILL_2__10299_ (
);

FILL SFILL98760x72050 (
);

FILL FILL_1__9755_ (
);

FILL FILL_5__11633_ (
);

FILL FILL_1__9335_ (
);

FILL FILL_5__11213_ (
);

FILL FILL_3_BUFX2_insert970 (
);

FILL FILL_2__16105_ (
);

FILL FILL_4__7760_ (
);

FILL FILL_3_BUFX2_insert971 (
);

FILL FILL_4__7340_ (
);

FILL FILL_3_BUFX2_insert972 (
);

FILL FILL_4__10626_ (
);

FILL FILL_3_BUFX2_insert973 (
);

FILL FILL_2__11660_ (
);

FILL FILL_3_BUFX2_insert974 (
);

FILL FILL_2__11240_ (
);

FILL FILL_3_BUFX2_insert975 (
);

FILL FILL_1__15938_ (
);

FILL SFILL49000x10050 (
);

FILL FILL_1__15518_ (
);

FILL FILL_3_BUFX2_insert976 (
);

FILL FILL_3_BUFX2_insert977 (
);

FILL FILL_3_BUFX2_insert978 (
);

FILL FILL_3_BUFX2_insert979 (
);

FILL FILL_1__10653_ (
);

FILL FILL_4__13098_ (
);

FILL FILL_1__10233_ (
);

FILL FILL_2__7678_ (
);

FILL FILL_0__7240_ (
);

FILL SFILL18840x2050 (
);

FILL SFILL23800x82050 (
);

FILL SFILL18760x7050 (
);

FILL FILL_5__12838_ (
);

FILL FILL_3__13872_ (
);

FILL FILL_5__12418_ (
);

FILL SFILL39480x24050 (
);

FILL FILL_3__13452_ (
);

FILL FILL_3__13032_ (
);

FILL FILL_4__8965_ (
);

FILL FILL_4__8125_ (
);

FILL FILL_2__12865_ (
);

FILL FILL_2__12445_ (
);

FILL FILL_2__12025_ (
);

FILL SFILL63960x35050 (
);

FILL SFILL94360x26050 (
);

FILL FILL_1__11858_ (
);

FILL FILL_1__11438_ (
);

FILL FILL_1__11018_ (
);

FILL FILL_0__8865_ (
);

FILL FILL_5__16251_ (
);

FILL FILL_3__6962_ (
);

FILL FILL_0__8445_ (
);

DFFSR _10716_ (
    .Q(\datapath_1.regfile_1.regOut[30] [6]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1888_[6])
);

FILL FILL_5__6888_ (
);

FILL FILL_4__15664_ (
);

FILL FILL_4__15244_ (
);

DFFSR _13188_ (
    .Q(\datapath_1.mux_iord.din0 [13]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[13])
);

FILL FILL_2__9404_ (
);

FILL FILL_3__14657_ (
);

FILL FILL_1__15691_ (
);

FILL FILL_3__14237_ (
);

FILL FILL_1__15271_ (
);

FILL FILL_0__14684_ (
);

FILL FILL_0__14264_ (
);

FILL FILL_1__7821_ (
);

FILL FILL_3__7747_ (
);

FILL FILL_3__7327_ (
);

FILL FILL_5__12591_ (
);

FILL FILL_5__12171_ (
);

BUFX2 _6891_ (
    .A(_2_[21]),
    .Y(memoryWriteData[21])
);

FILL FILL_4__16449_ (
);

FILL FILL_4__16029_ (
);

FILL FILL_4__11584_ (
);

FILL FILL_4__11164_ (
);

FILL SFILL8760x43050 (
);

FILL FILL_1__16056_ (
);

FILL FILL_3__10997_ (
);

FILL FILL_5__8614_ (
);

FILL FILL_6_BUFX2_insert480 (
);

FILL FILL_3__10577_ (
);

FILL FILL_3__10157_ (
);

FILL FILL_1__11191_ (
);

FILL FILL_6__11911_ (
);

FILL FILL_0__15889_ (
);

OAI22X1 _15754_ (
    .A(_5472__bF$buf2),
    .B(_4774_),
    .C(_4762_),
    .D(_5527__bF$buf3),
    .Y(_6217_)
);

FILL FILL_0__15469_ (
);

OAI22X1 _15334_ (
    .A(_5463__bF$buf0),
    .B(_5807_),
    .C(_5806_),
    .D(_5504__bF$buf4),
    .Y(_5808_)
);

FILL FILL_0__15049_ (
);

FILL FILL_6_BUFX2_insert485 (
);

FILL FILL_0__10184_ (
);

FILL SFILL114600x43050 (
);

FILL FILL_5__10904_ (
);

FILL FILL_1__8606_ (
);

FILL FILL_0__16410_ (
);

FILL FILL_2__10931_ (
);

FILL FILL_5__13796_ (
);

FILL FILL_2__10511_ (
);

FILL FILL_5__13376_ (
);

INVX1 _7676_ (
    .A(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_396_)
);

DFFSR _7256_ (
    .Q(\datapath_1.regfile_1.regOut[3] [2]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_133_[2])
);

FILL FILL_4__12789_ (
);

FILL FILL_4__9083_ (
);

FILL FILL_4__12369_ (
);

FILL FILL_2__6949_ (
);

FILL FILL_0__6931_ (
);

FILL FILL_1__12396_ (
);

FILL FILL_4__13730_ (
);

FILL SFILL3720x69050 (
);

FILL FILL_4__13310_ (
);

INVX1 _16119_ (
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_6573_)
);

FILL FILL_3__7080_ (
);

FILL FILL_0__11389_ (
);

NOR2X1 _11674_ (
    .A(_2775_),
    .B(_2767_),
    .Y(_2776_)
);

INVX1 _11254_ (
    .A(_2137_),
    .Y(_2373_)
);

FILL FILL_3__12723_ (
);

FILL FILL_6__15168_ (
);

FILL FILL_3__12303_ (
);

FILL FILL_4__7816_ (
);

FILL FILL_2__11716_ (
);

FILL FILL_0__12750_ (
);

FILL FILL_3__15195_ (
);

FILL FILL_0__12330_ (
);

FILL FILL_1__10709_ (
);

FILL FILL112360x80050 (
);

FILL FILL_2__14188_ (
);

FILL FILL_5__15942_ (
);

FILL FILL_5__15522_ (
);

FILL FILL_0__7716_ (
);

FILL FILL_5__15102_ (
);

DFFSR _9822_ (
    .Q(\datapath_1.regfile_1.regOut[23] [8]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_1433_[8])
);

OAI21X1 _9402_ (
    .A(_1281_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .C(_1282_),
    .Y(_1238_[22])
);

FILL SFILL74760x36050 (
);

FILL FILL_4__14935_ (
);

FILL FILL_4__14515_ (
);

OAI21X1 _12879_ (
    .A(_3590_),
    .B(vdd),
    .C(_3591_),
    .Y(_3555_[18])
);

OAI21X1 _12459_ (
    .A(_3371_),
    .B(vdd),
    .C(_3372_),
    .Y(_3360_[6])
);

NAND3X1 _12039_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[13]),
    .C(_3032__bF$buf3),
    .Y(_3075_)
);

FILL FILL_3__13928_ (
);

FILL FILL_1__14962_ (
);

FILL FILL_3__13508_ (
);

FILL FILL_1__14542_ (
);

FILL FILL_1__14122_ (
);

FILL SFILL43960x31050 (
);

FILL FILL_6__11088_ (
);

FILL FILL_0__13955_ (
);

INVX1 _13820_ (
    .A(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_4325_)
);

FILL FILL_0__13535_ (
);

NOR2X1 _13400_ (
    .A(_3906_),
    .B(_3911_),
    .Y(_3912_)
);

FILL FILL_0__13115_ (
);

FILL FILL_5__9992_ (
);

FILL FILL_5__9152_ (
);

AOI21X1 _16292_ (
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .B(_5649_),
    .C(_6740_),
    .Y(_6741_)
);

FILL FILL_5__16307_ (
);

FILL FILL_1__9984_ (
);

FILL FILL_5__11862_ (
);

FILL FILL_5__11442_ (
);

FILL FILL_1__9144_ (
);

FILL FILL_5__11022_ (
);

FILL SFILL104520x48050 (
);

FILL SFILL43880x38050 (
);

FILL FILL_2__16334_ (
);

FILL FILL_4__10435_ (
);

FILL FILL_4__10015_ (
);

FILL FILL_1__15747_ (
);

FILL FILL_1__15327_ (
);

FILL FILL_1__10882_ (
);

FILL FILL_1__10042_ (
);

AOI22X1 _14605_ (
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .B(_4005__bF$buf3),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_5093_)
);

FILL FILL112280x42050 (
);

FILL FILL_2__7487_ (
);

FILL FILL_2__7067_ (
);

FILL FILL_6__13654_ (
);

FILL FILL_6__13234_ (
);

FILL FILL_5__12647_ (
);

FILL FILL_3__13681_ (
);

FILL FILL_5__12227_ (
);

FILL FILL_3__13261_ (
);

INVX1 _6947_ (
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_32_)
);

FILL FILL_4__8774_ (
);

FILL FILL_4__8354_ (
);

FILL FILL_2__12254_ (
);

FILL FILL_1__11667_ (
);

FILL FILL_1__11247_ (
);

FILL FILL_5__16060_ (
);

FILL FILL_0__8254_ (
);

NAND3X1 _10945_ (
    .A(_2078_),
    .B(_2077_),
    .C(_2070_),
    .Y(\control_1.next [0])
);

INVX1 _10525_ (
    .A(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_1848_)
);

INVX1 _10105_ (
    .A(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_1629_)
);

FILL FILL_4__15893_ (
);

FILL FILL_4__15473_ (
);

FILL FILL_4__15053_ (
);

FILL FILL_2__9633_ (
);

FILL FILL_3__14886_ (
);

FILL FILL_3__14466_ (
);

FILL FILL_2__9213_ (
);

FILL FILL_0__11601_ (
);

FILL FILL_3__14046_ (
);

FILL FILL_1__15080_ (
);

FILL FILL_4__9979_ (
);

FILL FILL_4__9139_ (
);

FILL FILL_2__13879_ (
);

FILL FILL_2__13459_ (
);

FILL FILL_0__14493_ (
);

FILL FILL_2__13039_ (
);

FILL SFILL33880x36050 (
);

FILL FILL_0__14073_ (
);

FILL FILL_1__7630_ (
);

FILL FILL_1__7210_ (
);

FILL FILL_2__14820_ (
);

FILL FILL_3__7976_ (
);

FILL FILL_0__9879_ (
);

FILL FILL_2__14400_ (
);

FILL FILL_3__7556_ (
);

FILL FILL_0__9039_ (
);

FILL FILL_1__13813_ (
);

FILL FILL_4__16258_ (
);

FILL FILL_4__11393_ (
);

FILL FILL_1__16285_ (
);

FILL FILL_5__8843_ (
);

FILL FILL_3__10386_ (
);

FILL FILL_5__8003_ (
);

NAND3X1 _15983_ (
    .A(_6434_),
    .B(_6435_),
    .C(_6439_),
    .Y(_6440_)
);

FILL FILL_0__15698_ (
);

FILL SFILL49400x19050 (
);

OAI22X1 _15563_ (
    .A(_5478__bF$buf2),
    .B(_4539_),
    .C(_5552__bF$buf3),
    .D(_4559_),
    .Y(_6031_)
);

FILL FILL_0__15278_ (
);

FILL SFILL23880x79050 (
);

NAND3X1 _15143_ (
    .A(_5615_),
    .B(_5616_),
    .C(_5620_),
    .Y(_5621_)
);

FILL FILL_1__8835_ (
);

FILL FILL_2__15605_ (
);

FILL FILL_4__6840_ (
);

FILL SFILL18600x14050 (
);

FILL FILL_2__10320_ (
);

OAI21X1 _7485_ (
    .A(_308_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_309_),
    .Y(_263_[23])
);

OAI21X1 _7065_ (
    .A(_89_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .C(_90_),
    .Y(_68_[11])
);

FILL FILL_4__12598_ (
);

FILL FILL_4__12178_ (
);

FILL FILL_5__9628_ (
);

FILL FILL_5__9208_ (
);

FILL FILL_6__12505_ (
);

FILL SFILL23800x77050 (
);

INVX1 _16348_ (
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .Y(_6786_)
);

FILL FILL_0__11198_ (
);

OAI21X1 _11483_ (
    .A(_2289_),
    .B(_2344__bF$buf0),
    .C(_2596_),
    .Y(_2597_)
);

FILL SFILL84520x50050 (
);

FILL FILL_5__11918_ (
);

INVX1 _11063_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .Y(_2182_)
);

FILL FILL_3__12952_ (
);

FILL FILL_3__12532_ (
);

FILL FILL_3__12112_ (
);

FILL FILL_4__7625_ (
);

FILL FILL_4__7205_ (
);

FILL FILL_2__11945_ (
);

FILL FILL_2__11525_ (
);

FILL FILL_2__11105_ (
);

FILL FILL_1__10938_ (
);

FILL FILL_1__10518_ (
);

FILL FILL_5__15751_ (
);

FILL FILL_0__7945_ (
);

FILL FILL_5__15331_ (
);

FILL FILL_0__7105_ (
);

OAI21X1 _9631_ (
    .A(_1393_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .C(_1394_),
    .Y(_1368_[13])
);

OAI21X1 _9211_ (
    .A(_1174_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .C(_1175_),
    .Y(_1173_[1])
);

FILL FILL_4__14744_ (
);

FILL FILL_4__14324_ (
);

DFFSR _12688_ (
    .Q(\datapath_1.Data [25]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3425_[25])
);

FILL FILL_3__8094_ (
);

NAND3X1 _12268_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [15]),
    .C(_3198__bF$buf3),
    .Y(_3240_)
);

FILL FILL_2__8904_ (
);

FILL FILL_3__13737_ (
);

FILL FILL_3__13317_ (
);

FILL FILL_1__14771_ (
);

FILL FILL_1__14351_ (
);

FILL FILL_0__13764_ (
);

FILL SFILL8840x31050 (
);

FILL FILL_0__13344_ (
);

FILL FILL_5__9381_ (
);

FILL FILL_1__6901_ (
);

FILL FILL_5__16116_ (
);

FILL FILL_1__9793_ (
);

FILL FILL_5__11671_ (
);

FILL FILL_5__11251_ (
);

FILL FILL_1__9373_ (
);

FILL FILL_4__15949_ (
);

FILL FILL_4__15529_ (
);

FILL FILL_4__15109_ (
);

FILL FILL_2__16143_ (
);

FILL FILL_3__9299_ (
);

FILL FILL_4__10664_ (
);

FILL FILL_4__10244_ (
);

FILL SFILL13800x75050 (
);

FILL FILL_1__15976_ (
);

FILL FILL_1__15556_ (
);

FILL FILL_1__15136_ (
);

FILL FILL_1__10691_ (
);

FILL FILL_1__10271_ (
);

FILL FILL_0__14969_ (
);

AOI21X1 _14834_ (
    .A(_5296_),
    .B(_5317_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [28])
);

FILL FILL_0__14549_ (
);

FILL FILL_0__14129_ (
);

AOI22X1 _14414_ (
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .B(_4005__bF$buf0),
    .C(_3885_),
    .D(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_4906_)
);

FILL FILL_2__7296_ (
);

FILL SFILL84360x19050 (
);

FILL FILL_0__15910_ (
);

FILL FILL_5__12876_ (
);

FILL FILL_5__12456_ (
);

FILL FILL_3__13490_ (
);

FILL FILL_5__12036_ (
);

FILL FILL_4__8583_ (
);

FILL FILL_4__11869_ (
);

FILL FILL_4__11449_ (
);

FILL FILL_2__12483_ (
);

FILL FILL_4__11029_ (
);

FILL FILL_2__12063_ (
);

FILL FILL_2_BUFX2_insert1000 (
);

FILL FILL_2_BUFX2_insert1001 (
);

FILL SFILL13800x30050 (
);

FILL FILL_1__11896_ (
);

FILL FILL_2_BUFX2_insert1002 (
);

FILL FILL_2_BUFX2_insert1003 (
);

FILL FILL_1__11476_ (
);

FILL FILL_2_BUFX2_insert1004 (
);

FILL FILL_1__11056_ (
);

FILL FILL_2_BUFX2_insert1005 (
);

NAND2X1 _15619_ (
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .B(_5606_),
    .Y(_6085_)
);

FILL FILL_2_BUFX2_insert1006 (
);

FILL SFILL74040x41050 (
);

FILL FILL_2_BUFX2_insert1007 (
);

FILL FILL_2_BUFX2_insert1008 (
);

FILL FILL_6__9870_ (
);

FILL FILL_0__8483_ (
);

FILL FILL_2_BUFX2_insert1009 (
);

FILL FILL_0__10889_ (
);

FILL FILL_0__8063_ (
);

INVX1 _10754_ (
    .A(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_1960_)
);

DFFSR _10334_ (
    .Q(\datapath_1.regfile_1.regOut[27] [8]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_1693_[8])
);

FILL FILL_0__10049_ (
);

FILL FILL_3__11803_ (
);

FILL FILL_4__15282_ (
);

FILL FILL_2__9862_ (
);

FILL FILL_0__11830_ (
);

FILL FILL_3__14695_ (
);

FILL FILL_3__14275_ (
);

FILL FILL_0__11410_ (
);

FILL FILL_2__9022_ (
);

FILL FILL_4__9788_ (
);

FILL FILL_4__9368_ (
);

FILL FILL112360x75050 (
);

FILL FILL_2__13688_ (
);

FILL FILL_2__13268_ (
);

FILL FILL_5__14602_ (
);

OAI21X1 _8902_ (
    .A(_1029_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1030_),
    .Y(_978_[26])
);

INVX1 _11959_ (
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3014_)
);

FILL FILL_3__7365_ (
);

FILL FILL_0__9268_ (
);

OAI21X1 _11539_ (
    .A(_2649_),
    .B(_2219_),
    .C(_2225_),
    .Y(_2650_)
);

FILL SFILL3720x19050 (
);

AND2X2 _11119_ (
    .A(_2237_),
    .B(_2226_),
    .Y(_2238_)
);

FILL FILL_1__13622_ (
);

FILL FILL_4__16067_ (
);

FILL FILL_1_BUFX2_insert300 (
);

FILL FILL_1_BUFX2_insert301 (
);

FILL FILL_0__12615_ (
);

FILL FILL_1_BUFX2_insert302 (
);

OAI21X1 _12900_ (
    .A(_3604_),
    .B(vdd),
    .C(_3605_),
    .Y(_3555_[25])
);

FILL FILL_1_BUFX2_insert303 (
);

FILL FILL_1_BUFX2_insert304 (
);

FILL FILL_1__16094_ (
);

FILL FILL_1_BUFX2_insert305 (
);

FILL FILL_5__8652_ (
);

FILL FILL_1_BUFX2_insert306 (
);

FILL FILL_5__8232_ (
);

FILL FILL_1_BUFX2_insert307 (
);

FILL FILL_3__10195_ (
);

FILL FILL_1_BUFX2_insert308 (
);

FILL FILL_6_BUFX2_insert863 (
);

FILL FILL_1_BUFX2_insert309 (
);

OAI22X1 _15792_ (
    .A(_6253_),
    .B(_5544__bF$buf0),
    .C(_5499__bF$buf1),
    .D(_4841_),
    .Y(_6254_)
);

NOR2X1 _15372_ (
    .A(_5834_),
    .B(_5844_),
    .Y(_5845_)
);

FILL FILL_0__15087_ (
);

FILL FILL_5__15807_ (
);

FILL FILL112360x30050 (
);

FILL FILL_6_BUFX2_insert868 (
);

FILL FILL_3__16001_ (
);

FILL FILL_5__10942_ (
);

FILL FILL_1__8644_ (
);

FILL FILL_5__10522_ (
);

FILL FILL_1__8224_ (
);

FILL FILL_5__10102_ (
);

FILL FILL_2__15834_ (
);

FILL FILL_2__15414_ (
);

FILL FILL_1__14827_ (
);

FILL FILL_1__14407_ (
);

OAI21X1 _7294_ (
    .A(_201_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_202_),
    .Y(_198_[2])
);

FILL FILL_3__9931_ (
);

FILL FILL_3__9511_ (
);

FILL FILL112280x37050 (
);

FILL FILL_2__6987_ (
);

FILL FILL_5__9857_ (
);

FILL FILL_5__9017_ (
);

INVX1 _16157_ (
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_6610_)
);

OR2X2 _11292_ (
    .A(_2223_),
    .B(_2224_),
    .Y(_2411_)
);

FILL FILL_1__9849_ (
);

FILL FILL_5__11727_ (
);

FILL FILL_3__12761_ (
);

FILL FILL_1__9429_ (
);

FILL FILL_5__11307_ (
);

FILL FILL_1__9009_ (
);

FILL FILL_3__12341_ (
);

FILL FILL_4__7854_ (
);

FILL FILL_4__7434_ (
);

FILL FILL_2__11754_ (
);

FILL FILL_5__14199_ (
);

FILL FILL_2__11334_ (
);

FILL SFILL54040x82050 (
);

NAND2X1 _8499_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_823_)
);

NAND2X1 _8079_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_604_)
);

FILL FILL_1__10747_ (
);

FILL FILL_5__15980_ (
);

FILL FILL_5__15560_ (
);

FILL FILL_0__7754_ (
);

FILL FILL_5__15140_ (
);

FILL FILL_0__7334_ (
);

OAI21X1 _9860_ (
    .A(_1505_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1506_),
    .Y(_1498_[4])
);

DFFSR _9440_ (
    .Q(\datapath_1.regfile_1.regOut[20] [10]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_1238_[10])
);

NAND2X1 _9020_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1089_)
);

FILL FILL_4__14973_ (
);

FILL FILL_4__14553_ (
);

FILL FILL_4__14133_ (
);

NAND2X1 _12497_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [19]),
    .Y(_3398_)
);

AOI22X1 _12077_ (
    .A(\datapath_1.ALUResult [22]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3104_)
);

FILL FILL_2__8713_ (
);

FILL FILL_3__13966_ (
);

FILL FILL_3__13546_ (
);

FILL SFILL68680x23050 (
);

FILL FILL_1__14580_ (
);

FILL FILL_3__13126_ (
);

FILL FILL_1__14160_ (
);

FILL FILL_4__8639_ (
);

FILL FILL_4__8219_ (
);

FILL FILL_5_BUFX2_insert880 (
);

FILL FILL_5_BUFX2_insert881 (
);

FILL FILL_2__12959_ (
);

FILL SFILL94520x47050 (
);

FILL FILL_0__13993_ (
);

FILL FILL_5_BUFX2_insert882 (
);

FILL FILL_5_BUFX2_insert883 (
);

FILL FILL_2__12119_ (
);

FILL FILL_0__13573_ (
);

FILL FILL_0__13153_ (
);

FILL FILL_5_BUFX2_insert884 (
);

FILL FILL_5_BUFX2_insert885 (
);

FILL FILL_5_BUFX2_insert886 (
);

FILL FILL_5_BUFX2_insert887 (
);

FILL FILL_5_BUFX2_insert888 (
);

FILL FILL_5_BUFX2_insert889 (
);

FILL FILL_2__13900_ (
);

FILL FILL_0__8959_ (
);

FILL FILL_5__16345_ (
);

FILL FILL_0__8119_ (
);

FILL FILL_5__11480_ (
);

FILL FILL_5__11060_ (
);

FILL FILL_4__15758_ (
);

FILL FILL_4__15338_ (
);

FILL FILL_2__16372_ (
);

FILL FILL_4__10893_ (
);

FILL FILL_2__9918_ (
);

FILL FILL_4__10053_ (
);

FILL FILL_0__9900_ (
);

FILL FILL_1__15785_ (
);

FILL FILL_1__15365_ (
);

FILL FILL_5__7503_ (
);

FILL FILL_0__14778_ (
);

OAI22X1 _14643_ (
    .A(_5130_),
    .B(_3982__bF$buf0),
    .C(_3983__bF$buf3),
    .D(_5129_),
    .Y(_5131_)
);

FILL FILL_0__14358_ (
);

OAI22X1 _14223_ (
    .A(_4718_),
    .B(_3936__bF$buf2),
    .C(_3967__bF$buf3),
    .D(_4717_),
    .Y(_4719_)
);

FILL FILL_5__12265_ (
);

OAI21X1 _6985_ (
    .A(_56_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_57_),
    .Y(_3_[27])
);

FILL FILL_4__8392_ (
);

FILL FILL_4__11678_ (
);

FILL FILL_4__11258_ (
);

FILL FILL_2__12292_ (
);

FILL SFILL109800x81050 (
);

FILL FILL_5__8708_ (
);

FILL FILL_1__11285_ (
);

OAI22X1 _15848_ (
    .A(_5549__bF$buf0),
    .B(_6308_),
    .C(_5466__bF$buf4),
    .D(_6307_),
    .Y(_6309_)
);

AOI22X1 _15428_ (
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [9]),
    .C(\datapath_1.regfile_1.regOut[5] [9]),
    .D(_5700_),
    .Y(_5899_)
);

NAND3X1 _15008_ (
    .A(_5482_),
    .B(_5487_),
    .C(_5474_),
    .Y(_5488_)
);

OAI21X1 _10983_ (
    .A(_2105_),
    .B(vdd),
    .C(_2106_),
    .Y(_2098_[3])
);

FILL FILL_0__10698_ (
);

FILL FILL_0__10278_ (
);

OAI21X1 _10563_ (
    .A(_1872_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1873_),
    .Y(_1823_[25])
);

OAI21X1 _10143_ (
    .A(_1653_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .C(_1654_),
    .Y(_1628_[13])
);

FILL FILL_6__14897_ (
);

FILL FILL_6__14477_ (
);

FILL FILL_3__11612_ (
);

FILL FILL_4__15091_ (
);

FILL FILL_2__9671_ (
);

FILL FILL112440x6050 (
);

FILL FILL_2__9251_ (
);

FILL FILL_3__14084_ (
);

FILL FILL_4__9597_ (
);

FILL FILL_2__13497_ (
);

FILL FILL_5__14831_ (
);

FILL FILL_5__14411_ (
);

FILL FILL111800x3050 (
);

OAI21X1 _8711_ (
    .A(_922_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .C(_923_),
    .Y(_913_[5])
);

FILL FILL112040x5050 (
);

FILL FILL_4__13824_ (
);

FILL FILL_4__13404_ (
);

FILL FILL_0__9497_ (
);

FILL FILL_3__7594_ (
);

AOI21X1 _11768_ (
    .A(_2561_),
    .B(_2363_),
    .C(_2862_),
    .Y(_2863_)
);

FILL FILL_3__7174_ (
);

FILL SFILL23800x27050 (
);

OAI21X1 _11348_ (
    .A(_2117_),
    .B(_2344__bF$buf0),
    .C(_2465_),
    .Y(_2466_)
);

FILL FILL_1__13851_ (
);

FILL FILL_1__13431_ (
);

FILL FILL_4__16296_ (
);

FILL FILL_1__13011_ (
);

FILL SFILL8840x26050 (
);

FILL FILL_0__12844_ (
);

FILL FILL_0__12424_ (
);

FILL FILL_3__15289_ (
);

FILL FILL_0__12004_ (
);

FILL FILL_5__8881_ (
);

FILL FILL_5__8461_ (
);

FILL SFILL74200x8050 (
);

INVX1 _15181_ (
    .A(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_5658_)
);

FILL FILL_5__15616_ (
);

NAND2X1 _9916_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1544_)
);

FILL FILL_3__16230_ (
);

FILL FILL_5__10751_ (
);

FILL FILL_1__8873_ (
);

FILL FILL_1__8453_ (
);

FILL FILL_4__14609_ (
);

FILL FILL_2__15643_ (
);

FILL FILL_2__15223_ (
);

FILL FILL_3__8379_ (
);

FILL FILL_1__14636_ (
);

FILL FILL_1__14216_ (
);

FILL FILL_3__9740_ (
);

FILL FILL_0__13629_ (
);

INVX1 _13914_ (
    .A(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_4417_)
);

FILL FILL_0__13209_ (
);

FILL FILL_5__9666_ (
);

FILL FILL_5__9246_ (
);

OAI21X1 _16386_ (
    .A(_6810_),
    .B(gnd),
    .C(_6811_),
    .Y(_6769_[21])
);

FILL FILL_5__11956_ (
);

FILL FILL_1__9658_ (
);

FILL FILL_3__12990_ (
);

FILL FILL_5__11536_ (
);

FILL FILL_3__12570_ (
);

FILL FILL_5__11116_ (
);

FILL FILL_1__9238_ (
);

FILL FILL_3__12150_ (
);

FILL FILL_2__16008_ (
);

FILL FILL_4__10949_ (
);

FILL FILL_4__7243_ (
);

FILL FILL_2__11983_ (
);

FILL FILL_4__10529_ (
);

FILL FILL_2__11563_ (
);

FILL FILL_4__10109_ (
);

FILL FILL_2__11143_ (
);

FILL SFILL13800x25050 (
);

FILL FILL_1__10976_ (
);

FILL FILL_1__10556_ (
);

FILL FILL_1__10136_ (
);

FILL FILL_0__7983_ (
);

FILL FILL_0__7563_ (
);

FILL FILL_4__14782_ (
);

FILL FILL_4__14362_ (
);

FILL SFILL64120x72050 (
);

FILL FILL_0__10910_ (
);

FILL FILL_3__13775_ (
);

FILL FILL_2__8522_ (
);

FILL FILL_3__13355_ (
);

FILL FILL_2__8102_ (
);

FILL FILL_4__8868_ (
);

FILL FILL_4__8448_ (
);

FILL FILL_2__12768_ (
);

FILL FILL_2__12348_ (
);

FILL FILL_0__13382_ (
);

FILL SFILL64040x79050 (
);

FILL FILL_0__8768_ (
);

FILL FILL_3__6865_ (
);

FILL FILL_5__16154_ (
);

FILL FILL_0__8348_ (
);

OAI21X1 _10619_ (
    .A(_1889_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1890_),
    .Y(_1888_[1])
);

FILL FILL_4__15987_ (
);

FILL FILL_1__12702_ (
);

FILL FILL_4__15567_ (
);

FILL FILL_4__15147_ (
);

FILL FILL_2__16181_ (
);

FILL FILL_4__10282_ (
);

FILL FILL_2__9727_ (
);

FILL FILL_1__15594_ (
);

FILL FILL_1__15174_ (
);

FILL FILL_5__7732_ (
);

FILL FILL_5__7312_ (
);

FILL FILL_0__14587_ (
);

OAI22X1 _14872_ (
    .A(_3947__bF$buf1),
    .B(_5354_),
    .C(_3966__bF$buf0),
    .D(_5353_),
    .Y(_5355_)
);

INVX1 _14452_ (
    .A(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_4943_)
);

FILL FILL_0__14167_ (
);

AOI22X1 _14032_ (
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .B(_4090_),
    .C(_3948_),
    .D(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_4532_)
);

FILL FILL112360x25050 (
);

FILL FILL_3__15921_ (
);

FILL FILL_3__15501_ (
);

FILL FILL_1__7724_ (
);

FILL FILL_1__7304_ (
);

FILL FILL_2__14914_ (
);

FILL FILL_5__12494_ (
);

FILL SFILL84440x5050 (
);

FILL FILL_5__12074_ (
);

FILL FILL_1__13907_ (
);

FILL FILL_4__11487_ (
);

FILL FILL_4__11067_ (
);

FILL SFILL89240x83050 (
);

FILL FILL_1__16379_ (
);

FILL FILL_5__8517_ (
);

FILL FILL_1__11094_ (
);

FILL FILL_6__11814_ (
);

NOR2X1 _15657_ (
    .A(_4674_),
    .B(_5534__bF$buf4),
    .Y(_6122_)
);

INVX1 _15237_ (
    .A(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_5713_)
);

OAI21X1 _10792_ (
    .A(_1984_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .C(_1985_),
    .Y(_1953_[16])
);

OAI21X1 _10372_ (
    .A(_1765_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .C(_1766_),
    .Y(_1758_[4])
);

FILL FILL_5__10807_ (
);

FILL FILL_1__8509_ (
);

FILL FILL_3__11841_ (
);

FILL FILL_3__11421_ (
);

FILL FILL_3__11001_ (
);

FILL FILL_4__6934_ (
);

FILL FILL_0__16313_ (
);

FILL FILL_2__10834_ (
);

FILL FILL_5__13699_ (
);

FILL SFILL54040x77050 (
);

FILL FILL_5__13279_ (
);

FILL FILL_2__9480_ (
);

FILL FILL_2__10414_ (
);

NAND2X1 _7999_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_571_)
);

NAND2X1 _7579_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_352_)
);

NAND2X1 _7159_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .Y(_197_)
);

FILL FILL_5__14640_ (
);

FILL FILL_5__14220_ (
);

DFFSR _8940_ (
    .Q(\datapath_1.regfile_1.regOut[16] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_978_[22])
);

NAND2X1 _8520_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_837_)
);

NAND2X1 _8100_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_618_)
);

FILL FILL_1__12299_ (
);

FILL FILL_4__13633_ (
);

FILL FILL_4__13213_ (
);

AOI22X1 _11997_ (
    .A(\datapath_1.ALUResult [2]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3044_)
);

OAI21X1 _11577_ (
    .A(_2659_),
    .B(_2670_),
    .C(_2470__bF$buf2),
    .Y(_2685_)
);

NOR2X1 _11157_ (
    .A(\datapath_1.alu_1.ALUInB [20]),
    .B(_2232_),
    .Y(_2276_)
);

FILL FILL_3__12626_ (
);

FILL FILL_1__13660_ (
);

FILL FILL_3__12206_ (
);

FILL FILL_1__13240_ (
);

FILL FILL_4__7719_ (
);

FILL FILL_2__11619_ (
);

FILL FILL_0__12653_ (
);

FILL FILL_3__15098_ (
);

FILL FILL_0__12233_ (
);

FILL SFILL54040x32050 (
);

FILL FILL_5__8270_ (
);

FILL FILL_6__16012_ (
);

FILL FILL_5__15845_ (
);

FILL FILL_5__15425_ (
);

FILL FILL_5__15005_ (
);

FILL FILL_0__7619_ (
);

NAND2X1 _9725_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1437_)
);

DFFSR _9305_ (
    .Q(\datapath_1.regfile_1.regOut[19] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_1173_[3])
);

FILL FILL_5__10980_ (
);

FILL FILL_5__10560_ (
);

FILL FILL_5__10140_ (
);

FILL FILL_1__8262_ (
);

FILL FILL_4__14838_ (
);

FILL FILL_4__14418_ (
);

FILL FILL_2__15872_ (
);

FILL FILL_2__15452_ (
);

FILL FILL_2__15032_ (
);

FILL FILL_3__8188_ (
);

FILL FILL_1__14865_ (
);

FILL FILL_1__14445_ (
);

FILL FILL_1__14025_ (
);

FILL FILL_0__13858_ (
);

FILL FILL_0__13438_ (
);

INVX1 _13723_ (
    .A(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_4230_)
);

OAI21X1 _13303_ (
    .A(\datapath_1.a3 [4]),
    .B(_3837_),
    .C(_3785_),
    .Y(_3838_)
);

FILL FILL_0__13018_ (
);

FILL FILL_5__9895_ (
);

FILL FILL_5__9475_ (
);

FILL SFILL44040x75050 (
);

NOR2X1 _16195_ (
    .A(_6644_),
    .B(_6646_),
    .Y(_6647_)
);

FILL FILL_5__11765_ (
);

FILL FILL_1__9887_ (
);

FILL FILL_1__9467_ (
);

FILL FILL_5__11345_ (
);

FILL FILL_2__16237_ (
);

FILL FILL_4__7892_ (
);

FILL FILL_4__7472_ (
);

FILL FILL_4__7052_ (
);

FILL FILL_4__10758_ (
);

FILL FILL_2__11792_ (
);

FILL FILL_2__11372_ (
);

FILL FILL_1__10785_ (
);

FILL FILL_1__10365_ (
);

NOR2X1 _14928_ (
    .A(_5399_),
    .B(_5409_),
    .Y(_5410_)
);

INVX1 _14508_ (
    .A(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_4998_)
);

FILL SFILL8520x45050 (
);

FILL FILL_0__7372_ (
);

FILL FILL_4__14591_ (
);

FILL FILL_4__14171_ (
);

FILL SFILL44040x30050 (
);

FILL SFILL53800x1050 (
);

FILL FILL_2__8751_ (
);

FILL FILL_2__8331_ (
);

FILL FILL_3__13584_ (
);

FILL FILL_3__13164_ (
);

FILL FILL_4__8257_ (
);

FILL FILL_2__12997_ (
);

FILL FILL_2__12577_ (
);

FILL FILL_2__12157_ (
);

FILL FILL_5__13911_ (
);

FILL FILL_4__12904_ (
);

FILL FILL_5__16383_ (
);

FILL FILL_0__8997_ (
);

FILL FILL_0__8577_ (
);

FILL FILL_6__9544_ (
);

DFFSR _10848_ (
    .Q(\datapath_1.regfile_1.regOut[31] [10]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1953_[10])
);

NAND2X1 _10428_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1804_)
);

NAND2X1 _10008_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1585_)
);

FILL FILL_4__15796_ (
);

FILL FILL_4__15376_ (
);

FILL FILL_1__12511_ (
);

FILL FILL_2__9536_ (
);

FILL FILL_0__11924_ (
);

FILL FILL_3__14789_ (
);

FILL FILL_2__9116_ (
);

FILL FILL_3__14369_ (
);

FILL FILL_0__11504_ (
);

FILL FILL_5__7961_ (
);

FILL SFILL74120x69050 (
);

FILL FILL_5__7121_ (
);

FILL SFILL103800x1050 (
);

FILL FILL_0__14396_ (
);

INVX1 _14681_ (
    .A(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_5168_)
);

AOI22X1 _14261_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [16]),
    .C(\datapath_1.regfile_1.regOut[2] [16]),
    .D(_3998__bF$buf2),
    .Y(_4757_)
);

FILL FILL_3__15730_ (
);

FILL SFILL104040x3050 (
);

FILL FILL_3__15310_ (
);

FILL FILL_1__7953_ (
);

FILL FILL_1__7113_ (
);

FILL FILL_2__14723_ (
);

FILL FILL_2__14303_ (
);

FILL FILL_3__7879_ (
);

FILL FILL_3__7459_ (
);

FILL FILL_3__7039_ (
);

FILL FILL_1__13716_ (
);

FILL FILL_4__11296_ (
);

FILL FILL_0__12709_ (
);

FILL FILL_3__8400_ (
);

FILL FILL_1__16188_ (
);

FILL FILL_5__8746_ (
);

FILL FILL_3__10289_ (
);

FILL FILL_5__8326_ (
);

INVX1 _15886_ (
    .A(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_6346_)
);

NAND3X1 _15466_ (
    .A(_5927_),
    .B(_5935_),
    .C(_5932_),
    .Y(_5936_)
);

FILL SFILL74120x24050 (
);

NAND3X1 _15046_ (
    .A(_5459__bF$buf3),
    .B(_5461_),
    .C(_5465_),
    .Y(_5526_)
);

NAND2X1 _10181_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1680_)
);

FILL FILL_1__8738_ (
);

FILL FILL_5__10616_ (
);

FILL FILL_3__11650_ (
);

FILL FILL_1__8318_ (
);

FILL FILL_3__11230_ (
);

FILL FILL_2__15928_ (
);

FILL FILL_2__15508_ (
);

FILL SFILL99320x73050 (
);

FILL FILL_0__16122_ (
);

FILL FILL_2__10643_ (
);

FILL FILL_5__13088_ (
);

DFFSR _7388_ (
    .Q(\datapath_1.regfile_1.regOut[4] [6]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_198_[6])
);

FILL FILL_3__9605_ (
);

FILL FILL_6__12408_ (
);

FILL FILL_4__13862_ (
);

FILL FILL_4__13442_ (
);

FILL SFILL64120x67050 (
);

FILL FILL_4__13022_ (
);

XNOR2X1 _11386_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2503_)
);

FILL FILL_3__12855_ (
);

FILL FILL_2__7602_ (
);

FILL FILL_3__12435_ (
);

FILL FILL_3__12015_ (
);

FILL FILL_4__7948_ (
);

FILL FILL_4__7108_ (
);

FILL FILL_2__11848_ (
);

FILL SFILL24440x40050 (
);

FILL FILL_0__12882_ (
);

FILL FILL_2__11428_ (
);

FILL FILL_0__12462_ (
);

FILL FILL_2__11008_ (
);

FILL FILL_0__12042_ (
);

FILL SFILL89320x2050 (
);

FILL SFILL23720x5050 (
);

FILL FILL_5__15654_ (
);

FILL FILL_0__7848_ (
);

FILL FILL_5__15234_ (
);

FILL FILL_0__7428_ (
);

DFFSR _9954_ (
    .Q(\datapath_1.regfile_1.regOut[24] [12]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1498_[12])
);

INVX1 _9534_ (
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_1350_)
);

INVX1 _9114_ (
    .A(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_1131_)
);

FILL FILL_1__8491_ (
);

FILL FILL_1__8071_ (
);

FILL FILL_4__14647_ (
);

FILL FILL_2__15681_ (
);

FILL FILL_4__14227_ (
);

FILL FILL_2__15261_ (
);

FILL SFILL3640x1050 (
);

FILL FILL_1__14674_ (
);

FILL FILL_1__14254_ (
);

FILL FILL_0_BUFX2_insert340 (
);

FILL FILL_0_BUFX2_insert341 (
);

FILL FILL_0_BUFX2_insert342 (
);

FILL FILL_0_BUFX2_insert343 (
);

FILL FILL_0__13667_ (
);

FILL FILL_0_BUFX2_insert344 (
);

NAND3X1 _13952_ (
    .A(_4452_),
    .B(_4453_),
    .C(_4451_),
    .Y(_4454_)
);

FILL FILL_0__13247_ (
);

FILL FILL_0_BUFX2_insert345 (
);

NOR2X1 _13532_ (
    .A(_4030_),
    .B(_4042_),
    .Y(_4043_)
);

FILL SFILL89320x71050 (
);

INVX1 _13112_ (
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_3706_)
);

FILL FILL_0_BUFX2_insert346 (
);

FILL FILL_0_BUFX2_insert347 (
);

FILL FILL_0_BUFX2_insert348 (
);

FILL FILL_5__9284_ (
);

FILL FILL_0_BUFX2_insert349 (
);

FILL FILL_5__16019_ (
);

FILL SFILL64040x29050 (
);

FILL FILL_5__11994_ (
);

FILL SFILL49160x82050 (
);

FILL FILL_5__11574_ (
);

FILL FILL_1__9276_ (
);

FILL FILL_5__11154_ (
);

FILL FILL_2__16046_ (
);

FILL FILL_4__10567_ (
);

FILL FILL_4__10147_ (
);

FILL SFILL89240x78050 (
);

FILL FILL_2__11181_ (
);

FILL SFILL54120x65050 (
);

FILL FILL_1__15879_ (
);

FILL FILL_1__15459_ (
);

FILL FILL_1__15039_ (
);

FILL FILL_1__10174_ (
);

NOR2X1 _14737_ (
    .A(_5219_),
    .B(_5222_),
    .Y(_5223_)
);

OAI22X1 _14317_ (
    .A(_4810_),
    .B(_3936__bF$buf3),
    .C(_3905__bF$buf3),
    .D(_4809_),
    .Y(_4811_)
);

FILL SFILL49560x51050 (
);

FILL FILL_0__7181_ (
);

FILL FILL_2_BUFX2_insert20 (
);

FILL FILL_2__7199_ (
);

FILL FILL_2_BUFX2_insert21 (
);

FILL FILL_1__16400_ (
);

FILL FILL_2_BUFX2_insert22 (
);

FILL FILL_3__10921_ (
);

FILL FILL_2_BUFX2_insert23 (
);

FILL FILL_2_BUFX2_insert24 (
);

FILL FILL_3__10501_ (
);

FILL FILL_2_BUFX2_insert25 (
);

FILL FILL_2_BUFX2_insert26 (
);

FILL FILL_0__15813_ (
);

FILL FILL_2_BUFX2_insert27 (
);

FILL FILL_2_BUFX2_insert28 (
);

FILL SFILL89640x47050 (
);

FILL FILL_2_BUFX2_insert29 (
);

FILL FILL_5__12779_ (
);

FILL FILL_2__8980_ (
);

FILL FILL_5__12359_ (
);

FILL FILL_3__13393_ (
);

FILL FILL_2__8140_ (
);

FILL FILL_4__8486_ (
);

FILL FILL_4__8066_ (
);

FILL FILL_2__12386_ (
);

FILL FILL_5__13720_ (
);

FILL FILL_5__13300_ (
);

NAND2X1 _7600_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_366_)
);

FILL FILL_1__11799_ (
);

FILL SFILL54120x20050 (
);

FILL FILL_1__11379_ (
);

FILL FILL_4__12713_ (
);

FILL FILL_5__16192_ (
);

FILL FILL_0__8386_ (
);

FILL FILL_6__9353_ (
);

NAND2X1 _10657_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1916_)
);

NAND2X1 _10237_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1697_)
);

FILL FILL_3__11706_ (
);

FILL FILL_1__12740_ (
);

FILL FILL_4__15185_ (
);

FILL FILL_1__12320_ (
);

FILL FILL_2__9765_ (
);

FILL FILL_3__14598_ (
);

FILL FILL_2__9345_ (
);

FILL FILL_0__11733_ (
);

FILL FILL_3__14178_ (
);

FILL FILL_0__11313_ (
);

FILL SFILL54040x27050 (
);

FILL FILL_5__7350_ (
);

NOR2X1 _14490_ (
    .A(_4977_),
    .B(_4980_),
    .Y(_4981_)
);

INVX1 _14070_ (
    .A(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_4570_)
);

FILL FILL_5__14925_ (
);

FILL FILL_5__14505_ (
);

DFFSR _8805_ (
    .Q(\datapath_1.regfile_1.regOut[15] [15]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_913_[15])
);

FILL SFILL79240x76050 (
);

FILL FILL_1__7762_ (
);

FILL FILL_1__7342_ (
);

FILL FILL_4__13918_ (
);

FILL FILL_2__14952_ (
);

FILL FILL_2__14532_ (
);

FILL FILL_3__7688_ (
);

FILL FILL_2__14112_ (
);

FILL FILL_1__13945_ (
);

FILL FILL_1__13525_ (
);

FILL FILL_1__13105_ (
);

FILL SFILL33960x2050 (
);

FILL SFILL33880x7050 (
);

DFFSR _12803_ (
    .Q(\datapath_1.PCJump [14]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_3490_[12])
);

FILL FILL_0__12518_ (
);

FILL FILL_5__8975_ (
);

FILL FILL_5__8135_ (
);

AOI22X1 _15695_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [16]),
    .C(\datapath_1.regfile_1.regOut[26] [16]),
    .D(_5484_),
    .Y(_6159_)
);

INVX1 _15275_ (
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_5750_)
);

FILL FILL_3__16324_ (
);

FILL FILL_1__8967_ (
);

FILL FILL_5__10425_ (
);

FILL FILL_1__8127_ (
);

FILL FILL_5__10005_ (
);

FILL FILL_2__15737_ (
);

FILL SFILL79240x31050 (
);

FILL FILL_4__6972_ (
);

FILL FILL_2__15317_ (
);

FILL FILL_0__16351_ (
);

FILL FILL_2__10872_ (
);

FILL FILL_2__10452_ (
);

FILL FILL_2__10032_ (
);

INVX1 _7197_ (
    .A(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_158_)
);

FILL FILL111880x44050 (
);

FILL FILL_3__9414_ (
);

FILL FILL_0__6872_ (
);

FILL SFILL109400x57050 (
);

FILL FILL_4__13671_ (
);

FILL FILL_4__13251_ (
);

OAI21X1 _11195_ (
    .A(_2291_),
    .B(_2292_),
    .C(_2313_),
    .Y(_2314_)
);

FILL FILL_2__7831_ (
);

FILL FILL_3__12244_ (
);

FILL FILL_4__7757_ (
);

FILL FILL_4__7337_ (
);

FILL SFILL108520x8050 (
);

FILL FILL_2__11657_ (
);

FILL FILL_2__11237_ (
);

FILL FILL_0__12271_ (
);

FILL FILL_5__15883_ (
);

FILL FILL_5__15463_ (
);

FILL FILL_5__15043_ (
);

INVX1 _9763_ (
    .A(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_1462_)
);

FILL FILL_0__7237_ (
);

FILL FILL_6__8624_ (
);

INVX1 _9343_ (
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_1243_)
);

FILL FILL_4__14876_ (
);

FILL FILL_4__14456_ (
);

FILL FILL_4__14036_ (
);

FILL FILL_2__15490_ (
);

FILL FILL_2__15070_ (
);

FILL FILL_3__13869_ (
);

FILL FILL_2__8616_ (
);

FILL FILL_3__13449_ (
);

FILL FILL_1__14483_ (
);

FILL FILL_3__13029_ (
);

FILL FILL_1__14063_ (
);

FILL FILL_0__13896_ (
);

NOR2X1 _13761_ (
    .A(_4256_),
    .B(_4266_),
    .Y(_4267_)
);

FILL FILL_0__13476_ (
);

OAI21X1 _13341_ (
    .A(_3776_),
    .B(_3789_),
    .C(_3856_),
    .Y(_3862_)
);

FILL FILL_3__14810_ (
);

FILL FILL_5__9093_ (
);

FILL FILL_4__9903_ (
);

FILL FILL_2__13803_ (
);

FILL FILL_3__6959_ (
);

FILL FILL_5__16248_ (
);

FILL FILL_5__11383_ (
);

FILL FILL_1__9085_ (
);

FILL FILL_2__16275_ (
);

FILL FILL_4__10796_ (
);

FILL FILL_4__7090_ (
);

FILL FILL_4__10376_ (
);

FILL SFILL69160x36050 (
);

FILL FILL_0__9803_ (
);

FILL FILL_1__15688_ (
);

FILL FILL_1__15268_ (
);

FILL FILL_5__7826_ (
);

FILL FILL_6__10703_ (
);

INVX1 _14966_ (
    .A(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_5447_)
);

FILL SFILL74120x19050 (
);

NOR2X1 _14546_ (
    .A(_5032_),
    .B(_5035_),
    .Y(_5036_)
);

INVX1 _14126_ (
    .A(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_4624_)
);

FILL SFILL28920x8050 (
);

FILL FILL_1__7818_ (
);

FILL FILL_3__10310_ (
);

FILL SFILL99320x68050 (
);

FILL FILL_0__15622_ (
);

FILL FILL_0__15202_ (
);

FILL FILL_5__12588_ (
);

FILL FILL_5__12168_ (
);

BUFX2 _6888_ (
    .A(_2_[18]),
    .Y(memoryWriteData[18])
);

FILL SFILL69080x2050 (
);

FILL SFILL8760x9050 (
);

FILL FILL_2__12195_ (
);

FILL SFILL104280x61050 (
);

FILL FILL_1__11188_ (
);

FILL FILL_4__12522_ (
);

FILL FILL_4__12102_ (
);

FILL FILL_0__8195_ (
);

NOR2X1 _10886_ (
    .A(_2032_),
    .B(_2019_),
    .Y(_2033_)
);

FILL FILL_6__9162_ (
);

DFFSR _10466_ (
    .Q(\datapath_1.regfile_1.regOut[28] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_1758_[12])
);

INVX1 _10046_ (
    .A(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_1610_)
);

FILL SFILL43160x80050 (
);

FILL FILL_3__11935_ (
);

FILL FILL_3__11515_ (
);

FILL FILL_0__16407_ (
);

FILL FILL_2__10928_ (
);

FILL FILL_2__9994_ (
);

FILL FILL_2__10508_ (
);

FILL FILL_0__11962_ (
);

FILL SFILL99320x23050 (
);

FILL FILL_0__11542_ (
);

FILL FILL_2__9154_ (
);

FILL FILL_0__11122_ (
);

FILL FILL_6__15741_ (
);

FILL FILL_6__15321_ (
);

FILL FILL_5__14734_ (
);

FILL FILL_0__6928_ (
);

FILL FILL_5__14314_ (
);

INVX1 _8614_ (
    .A(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_879_)
);

FILL FILL_1__7991_ (
);

FILL FILL_1__7571_ (
);

FILL FILL_4__13727_ (
);

FILL FILL_4__13307_ (
);

FILL FILL_2__14761_ (
);

FILL FILL_2__14341_ (
);

FILL FILL_3__7497_ (
);

FILL FILL_3__7077_ (
);

FILL SFILL64120x17050 (
);

FILL FILL_1__13754_ (
);

FILL FILL_1__13334_ (
);

FILL FILL_4__16199_ (
);

FILL FILL_0__12747_ (
);

FILL SFILL89320x66050 (
);

INVX1 _12612_ (
    .A(\datapath_1.Data [15]),
    .Y(_3454_)
);

FILL FILL_0__12327_ (
);

FILL FILL_5__8784_ (
);

FILL FILL_5__8364_ (
);

FILL FILL_6__11661_ (
);

FILL FILL_6__11241_ (
);

FILL FILL_5__15939_ (
);

NAND2X1 _15084_ (
    .A(\datapath_1.regfile_1.regOut[25] [1]),
    .B(_5562_),
    .Y(_5563_)
);

FILL FILL_5__15519_ (
);

FILL FILL_3__16133_ (
);

DFFSR _9819_ (
    .Q(\datapath_1.regfile_1.regOut[23] [5]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_1433_[5])
);

FILL FILL_1__8776_ (
);

FILL FILL_5__10654_ (
);

FILL FILL_1__8356_ (
);

FILL FILL_5__10234_ (
);

FILL FILL_2__15966_ (
);

FILL FILL_2__15546_ (
);

FILL FILL_2__15126_ (
);

FILL FILL_0__16160_ (
);

FILL FILL_2__10681_ (
);

FILL FILL_2__10261_ (
);

FILL FILL_1__14959_ (
);

FILL FILL_1__14539_ (
);

FILL FILL_1__14119_ (
);

FILL FILL_3__9643_ (
);

AOI22X1 _13817_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [7]),
    .C(\datapath_1.regfile_1.regOut[6] [7]),
    .D(_4001__bF$buf0),
    .Y(_4322_)
);

FILL FILL_3__9223_ (
);

FILL SFILL33960x61050 (
);

FILL FILL_5__9989_ (
);

FILL FILL_1__15900_ (
);

FILL FILL_5__9149_ (
);

FILL SFILL89320x21050 (
);

AOI22X1 _16289_ (
    .A(_5496_),
    .B(\datapath_1.regfile_1.regOut[11] [31]),
    .C(\datapath_1.regfile_1.regOut[14] [31]),
    .D(_5971_),
    .Y(_6738_)
);

FILL FILL_4__13480_ (
);

FILL FILL_5__11859_ (
);

FILL FILL_3__12893_ (
);

FILL FILL_5__11439_ (
);

FILL FILL_3__12473_ (
);

FILL FILL_5__11019_ (
);

FILL FILL_2__7220_ (
);

FILL FILL_3__12053_ (
);

FILL SFILL18760x41050 (
);

FILL FILL_4__7986_ (
);

FILL FILL_4__7566_ (
);

FILL FILL_2__11886_ (
);

FILL FILL_2__11466_ (
);

FILL FILL_2__11046_ (
);

FILL FILL_0__12080_ (
);

FILL SFILL54120x15050 (
);

FILL FILL_1__10879_ (
);

FILL FILL_1__10039_ (
);

FILL FILL_5__15692_ (
);

FILL FILL_0__7886_ (
);

FILL FILL_5__15272_ (
);

INVX1 _9992_ (
    .A(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_1574_)
);

FILL FILL_0__7466_ (
);

DFFSR _9572_ (
    .Q(\datapath_1.regfile_1.regOut[21] [14]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_1303_[14])
);

FILL FILL_0__7046_ (
);

OAI21X1 _9152_ (
    .A(_1155_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .C(_1156_),
    .Y(_1108_[24])
);

FILL SFILL18680x48050 (
);

FILL FILL_1__11820_ (
);

FILL FILL_4__14685_ (
);

FILL SFILL38680x9050 (
);

FILL FILL_4__14265_ (
);

FILL FILL_1__11400_ (
);

FILL FILL_2__8845_ (
);

FILL FILL_0__10813_ (
);

FILL FILL_3__13678_ (
);

FILL FILL_3__13258_ (
);

FILL FILL_2__8005_ (
);

FILL FILL_1__14292_ (
);

FILL FILL_5__6850_ (
);

FILL FILL_0_BUFX2_insert720 (
);

FILL FILL_0_BUFX2_insert721 (
);

FILL FILL_0_BUFX2_insert722 (
);

FILL FILL_0_BUFX2_insert723 (
);

FILL FILL_0_BUFX2_insert724 (
);

INVX1 _13990_ (
    .A(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_4491_)
);

FILL FILL_0__13285_ (
);

FILL FILL_0_BUFX2_insert725 (
);

AOI22X1 _13570_ (
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .B(_4038__bF$buf1),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_4080_)
);

FILL FILL_0_BUFX2_insert726 (
);

OAI21X1 _13150_ (
    .A(_3730_),
    .B(PCEn_bF$buf7),
    .C(_3731_),
    .Y(_3685_[23])
);

FILL FILL_0_BUFX2_insert727 (
);

FILL FILL_0_BUFX2_insert728 (
);

FILL FILL_0_BUFX2_insert729 (
);

FILL FILL_1__6842_ (
);

FILL FILL_2__13612_ (
);

FILL FILL_5__16057_ (
);

FILL FILL_5__11192_ (
);

FILL FILL_1__12605_ (
);

FILL FILL_2__16084_ (
);

FILL FILL_4__10185_ (
);

FILL FILL_0__9612_ (
);

FILL FILL_1__15497_ (
);

FILL FILL_1__15077_ (
);

FILL FILL_5__7635_ (
);

FILL FILL_5__7215_ (
);

FILL FILL_4__16411_ (
);

FILL FILL_6__10512_ (
);

NAND3X1 _14775_ (
    .A(_5258_),
    .B(_5259_),
    .C(_5257_),
    .Y(_5260_)
);

NAND3X1 _14355_ (
    .A(_4847_),
    .B(_4848_),
    .C(_4846_),
    .Y(_4849_)
);

FILL FILL_3__15824_ (
);

FILL FILL_3__15404_ (
);

FILL FILL_1__7627_ (
);

FILL FILL_1__7207_ (
);

FILL FILL_6_BUFX2_insert101 (
);

FILL SFILL79240x26050 (
);

FILL FILL_2__14817_ (
);

FILL FILL_0__15851_ (
);

FILL FILL_0__15431_ (
);

FILL FILL_0__15011_ (
);

FILL FILL_6_BUFX2_insert106 (
);

FILL FILL_5__12397_ (
);

FILL FILL_3__8914_ (
);

FILL FILL_6__11717_ (
);

FILL FILL_4__12751_ (
);

FILL FILL_4__12331_ (
);

INVX1 _10695_ (
    .A(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_1941_)
);

INVX1 _10275_ (
    .A(\datapath_1.regfile_1.regOut[27] [15]),
    .Y(_1722_)
);

FILL FILL_2__6911_ (
);

FILL FILL_3__11744_ (
);

FILL FILL_3__11324_ (
);

FILL FILL_4__6837_ (
);

FILL FILL_0__16216_ (
);

FILL FILL_2__10317_ (
);

FILL FILL_2__9383_ (
);

FILL FILL_0__11771_ (
);

FILL FILL_0__11351_ (
);

FILL FILL_5__14963_ (
);

FILL FILL_5__14543_ (
);

FILL FILL_5__14123_ (
);

INVX1 _8843_ (
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_991_)
);

DFFSR _8423_ (
    .Q(\datapath_1.regfile_1.regOut[12] [17]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_718_[17])
);

OAI21X1 _8003_ (
    .A(_572_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .C(_573_),
    .Y(_523_[25])
);

FILL FILL_1__7380_ (
);

FILL FILL_4__13956_ (
);

FILL FILL_2__14990_ (
);

FILL FILL_4__13536_ (
);

FILL FILL_2__14570_ (
);

FILL FILL_4__13116_ (
);

FILL FILL_2__14150_ (
);

FILL FILL_1__13983_ (
);

FILL FILL_3__12529_ (
);

FILL FILL_3__12109_ (
);

FILL FILL_1__13563_ (
);

FILL FILL_1__13143_ (
);

FILL FILL_0__12976_ (
);

FILL SFILL69240x24050 (
);

INVX1 _12841_ (
    .A(\datapath_1.a [6]),
    .Y(_3566_)
);

FILL FILL_0__12136_ (
);

INVX1 _12421_ (
    .A(ALUOut[26]),
    .Y(_3346_)
);

AOI22X1 _12001_ (
    .A(\datapath_1.ALUResult [3]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3047_)
);

FILL FILL_5__8593_ (
);

FILL FILL_5__15748_ (
);

FILL FILL_5__15328_ (
);

FILL FILL_3__16362_ (
);

OAI21X1 _9628_ (
    .A(_1391_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .C(_1392_),
    .Y(_1368_[12])
);

OAI21X1 _9208_ (
    .A(_1236_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1237_),
    .Y(_1173_[0])
);

FILL FILL_5__10883_ (
);

FILL FILL_1__8585_ (
);

FILL FILL_5__10043_ (
);

FILL FILL_2__15775_ (
);

FILL FILL_2__15355_ (
);

FILL SFILL83800x71050 (
);

FILL SFILL99400x56050 (
);

FILL FILL_2__10490_ (
);

FILL FILL_1__14768_ (
);

FILL FILL_1__14348_ (
);

FILL FILL_5__6906_ (
);

FILL FILL_3__9872_ (
);

INVX8 _13626_ (
    .A(_3972__bF$buf0),
    .Y(_4135_)
);

FILL FILL_3__9032_ (
);

DFFSR _13206_ (
    .Q(\datapath_1.PCJump [31]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[31])
);

FILL FILL_5__9798_ (
);

FILL FILL_5__9378_ (
);

OAI22X1 _16098_ (
    .A(_5526__bF$buf0),
    .B(_5206_),
    .C(_5184_),
    .D(_5527__bF$buf0),
    .Y(_6552_)
);

FILL FILL_0__14702_ (
);

FILL FILL_5__11668_ (
);

FILL FILL_5__11248_ (
);

FILL FILL_3__12282_ (
);

FILL FILL_4__7375_ (
);

FILL FILL_2__11695_ (
);

FILL FILL_2__11275_ (
);

FILL SFILL99400x11050 (
);

FILL FILL_1__10688_ (
);

FILL FILL_2_BUFX2_insert250 (
);

FILL FILL_2_BUFX2_insert251 (
);

FILL FILL_1__10268_ (
);

FILL FILL_2_BUFX2_insert252 (
);

FILL FILL_2_BUFX2_insert253 (
);

FILL FILL_2_BUFX2_insert254 (
);

FILL FILL_4__11602_ (
);

FILL FILL_2_BUFX2_insert255 (
);

FILL FILL_0__7695_ (
);

FILL FILL_5__15081_ (
);

FILL FILL_2_BUFX2_insert256 (
);

FILL FILL_2_BUFX2_insert257 (
);

OAI21X1 _9381_ (
    .A(_1267_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .C(_1268_),
    .Y(_1238_[15])
);

FILL FILL_2_BUFX2_insert258 (
);

FILL FILL_6__8242_ (
);

FILL FILL_2_BUFX2_insert259 (
);

FILL FILL_4__14494_ (
);

FILL FILL_4__14074_ (
);

FILL FILL_0__15907_ (
);

FILL SFILL99320x18050 (
);

FILL FILL_2__8654_ (
);

FILL FILL_3__13487_ (
);

FILL FILL_2__8234_ (
);

FILL FILL_0__10622_ (
);

FILL FILL_0__13094_ (
);

FILL FILL_5__13814_ (
);

FILL SFILL59160x29050 (
);

FILL FILL_4__9941_ (
);

FILL FILL_4__9521_ (
);

FILL FILL_4__9101_ (
);

FILL FILL_2__13841_ (
);

FILL FILL_2__13421_ (
);

FILL FILL_3__6997_ (
);

FILL FILL_5__16286_ (
);

FILL FILL_2__13001_ (
);

FILL FILL_6__9027_ (
);

FILL FILL_4__15699_ (
);

FILL FILL_1__12834_ (
);

FILL FILL_1__12414_ (
);

FILL FILL_4__15279_ (
);

FILL FILL_2__9859_ (
);

FILL FILL_0__9421_ (
);

FILL FILL_0__11827_ (
);

FILL FILL_2__9019_ (
);

FILL FILL_0__9001_ (
);

FILL FILL_0__11407_ (
);

FILL FILL_5__7864_ (
);

FILL FILL_5__7444_ (
);

FILL FILL_4__16220_ (
);

INVX1 _14584_ (
    .A(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_5073_)
);

FILL FILL_0__14299_ (
);

OAI22X1 _14164_ (
    .A(_3978_),
    .B(_4660_),
    .C(_3977__bF$buf3),
    .D(_4661_),
    .Y(_4662_)
);

FILL FILL_3__15633_ (
);

FILL FILL_3__15213_ (
);

FILL SFILL14040x59050 (
);

FILL FILL_1__7856_ (
);

FILL FILL_1__7436_ (
);

FILL SFILL94280x60050 (
);

FILL FILL_2__14626_ (
);

FILL FILL_0__15660_ (
);

FILL FILL_2__14206_ (
);

FILL FILL_0__15240_ (
);

FILL FILL_1__13619_ (
);

FILL FILL_1_BUFX2_insert270 (
);

FILL FILL_4__11199_ (
);

FILL FILL_1_BUFX2_insert271 (
);

FILL FILL_3__8723_ (
);

FILL FILL_1_BUFX2_insert272 (
);

FILL FILL_1_BUFX2_insert273 (
);

FILL SFILL33960x56050 (
);

FILL FILL_1_BUFX2_insert274 (
);

FILL FILL_1_BUFX2_insert275 (
);

FILL FILL_5__8649_ (
);

FILL FILL_1_BUFX2_insert276 (
);

FILL FILL_5__8229_ (
);

FILL FILL_1_BUFX2_insert277 (
);

FILL FILL_1_BUFX2_insert278 (
);

FILL FILL_1_BUFX2_insert279 (
);

NAND3X1 _15789_ (
    .A(\datapath_1.regfile_1.regOut[4] [18]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf4),
    .Y(_6251_)
);

FILL FILL_4__12980_ (
);

OAI22X1 _15369_ (
    .A(_5463__bF$buf1),
    .B(_4336_),
    .C(_4340_),
    .D(_5504__bF$buf3),
    .Y(_5842_)
);

FILL FILL_4__12140_ (
);

FILL FILL_5__10939_ (
);

DFFSR _10084_ (
    .Q(\datapath_1.regfile_1.regOut[25] [14]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_1563_[14])
);

FILL FILL_3__11973_ (
);

FILL FILL_5__10519_ (
);

FILL FILL_3__11553_ (
);

FILL SFILL18760x36050 (
);

FILL FILL_3__11133_ (
);

FILL FILL_0__16025_ (
);

INVX1 _16310_ (
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_6759_)
);

FILL FILL_2__10966_ (
);

FILL FILL_2__10546_ (
);

FILL FILL_2__10126_ (
);

FILL FILL_0__11580_ (
);

FILL FILL_0__11160_ (
);

FILL FILL_3__9928_ (
);

FILL FILL_3__9508_ (
);

FILL FILL_5__14772_ (
);

FILL FILL_0__6966_ (
);

FILL FILL_5__14352_ (
);

OAI21X1 _8652_ (
    .A(_903_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .C(_904_),
    .Y(_848_[28])
);

OAI21X1 _8232_ (
    .A(_684_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_685_),
    .Y(_653_[16])
);

FILL SFILL33960x11050 (
);

FILL FILL_1__10900_ (
);

FILL FILL_4__13765_ (
);

FILL FILL_4__13345_ (
);

OAI21X1 _11289_ (
    .A(_2376_),
    .B(_2383_),
    .C(_2407_),
    .Y(_2408_)
);

FILL FILL_3__12758_ (
);

FILL FILL_2__7505_ (
);

FILL FILL_1__13792_ (
);

FILL FILL_3__12338_ (
);

FILL FILL_1__13372_ (
);

FILL FILL_0__12785_ (
);

OAI21X1 _12650_ (
    .A(_3478_),
    .B(vdd),
    .C(_3479_),
    .Y(_3425_[27])
);

FILL FILL_0__12365_ (
);

NAND3X1 _12230_ (
    .A(_3209_),
    .B(_3210_),
    .C(_3211_),
    .Y(\datapath_1.alu_1.ALUInB [3])
);

FILL FILL_5__15977_ (
);

FILL FILL_5__15557_ (
);

FILL FILL_5__15137_ (
);

FILL FILL_6__8718_ (
);

OAI21X1 _9857_ (
    .A(_1503_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1504_),
    .Y(_1498_[3])
);

FILL FILL_3__16171_ (
);

DFFSR _9437_ (
    .Q(\datapath_1.regfile_1.regOut[20] [7]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_1238_[7])
);

FILL FILL_5__10692_ (
);

NAND2X1 _9017_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1087_)
);

FILL FILL_1__8394_ (
);

FILL FILL_5__10272_ (
);

FILL FILL_2__15584_ (
);

FILL SFILL79320x14050 (
);

FILL FILL_2__15164_ (
);

FILL FILL_1__14997_ (
);

FILL FILL_1__14577_ (
);

FILL FILL_1__14157_ (
);

FILL FILL_4__15911_ (
);

FILL FILL111960x27050 (
);

FILL FILL_3__9681_ (
);

INVX1 _13855_ (
    .A(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_4359_)
);

FILL FILL_3__9261_ (
);

NAND3X1 _13435_ (
    .A(_3898_),
    .B(_3903_),
    .C(_3888_),
    .Y(_3947_)
);

NAND2X1 _13015_ (
    .A(vdd),
    .B(\datapath_1.rd2 [21]),
    .Y(_3662_)
);

FILL FILL_3__14904_ (
);

FILL FILL_6__12484_ (
);

FILL SFILL29240x61050 (
);

FILL FILL_0__14931_ (
);

FILL FILL_0__14511_ (
);

FILL FILL_5__11897_ (
);

FILL FILL_1__9599_ (
);

FILL FILL_5__11477_ (
);

FILL FILL_5__11057_ (
);

FILL FILL_3__12091_ (
);

FILL FILL_2__16369_ (
);

FILL SFILL53720x72050 (
);

FILL FILL_4__7184_ (
);

FILL FILL_2__11084_ (
);

FILL FILL_1__10497_ (
);

FILL FILL_4__11831_ (
);

FILL FILL_4__11411_ (
);

FILL FILL_0__7084_ (
);

DFFSR _9190_ (
    .Q(\datapath_1.regfile_1.regOut[18] [16]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_1108_[16])
);

FILL FILL_1__16303_ (
);

FILL FILL_3__10824_ (
);

FILL FILL_6__13689_ (
);

FILL FILL_3__10404_ (
);

FILL FILL_0__15716_ (
);

FILL FILL_2__8883_ (
);

FILL FILL_2__8463_ (
);

FILL FILL_3__13296_ (
);

FILL FILL_0__10431_ (
);

FILL FILL_0__10011_ (
);

FILL FILL_4__8389_ (
);

FILL FILL_2__12289_ (
);

FILL SFILL69320x12050 (
);

FILL FILL_5__13623_ (
);

DFFSR _7923_ (
    .Q(\datapath_1.regfile_1.regOut[8] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_458_[29])
);

OAI21X1 _7503_ (
    .A(_320_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_321_),
    .Y(_263_[29])
);

FILL FILL_1__6880_ (
);

FILL FILL_4__9750_ (
);

FILL FILL_4__12616_ (
);

FILL FILL_2__13650_ (
);

FILL FILL_2__13230_ (
);

FILL FILL_5__16095_ (
);

FILL FILL_3__11609_ (
);

FILL FILL_1__12643_ (
);

FILL FILL_4__15088_ (
);

FILL FILL_1__12223_ (
);

FILL SFILL69240x19050 (
);

FILL FILL_2__9668_ (
);

FILL FILL_0__9650_ (
);

FILL FILL_0__9230_ (
);

FILL FILL_2__9248_ (
);

NAND2X1 _11921_ (
    .A(IorD_bF$buf4),
    .B(ALUOut[11]),
    .Y(_2989_)
);

FILL FILL_0__11636_ (
);

FILL FILL_0__11216_ (
);

OAI21X1 _11501_ (
    .A(_2296_),
    .B(_2305_),
    .C(_2462__bF$buf2),
    .Y(_2614_)
);

FILL FILL_5__7673_ (
);

FILL FILL_5__7253_ (
);

OAI22X1 _14393_ (
    .A(_3947__bF$buf0),
    .B(_4885_),
    .C(_3909_),
    .D(_4884_),
    .Y(_4886_)
);

FILL FILL_6__10130_ (
);

FILL FILL_5__14828_ (
);

FILL FILL_5__14408_ (
);

FILL FILL_3__15862_ (
);

FILL FILL_3__15442_ (
);

OAI21X1 _8708_ (
    .A(_920_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .C(_921_),
    .Y(_913_[4])
);

FILL FILL_3__15022_ (
);

FILL FILL_1__7245_ (
);

FILL FILL_2__14855_ (
);

FILL FILL_2__14435_ (
);

FILL FILL_2__14015_ (
);

FILL FILL_1__13848_ (
);

FILL FILL_1__13428_ (
);

FILL FILL_1__13008_ (
);

FILL FILL_3__8952_ (
);

FILL FILL_3__8532_ (
);

OAI21X1 _12706_ (
    .A(_3495_),
    .B(IRWrite_bF$buf1),
    .C(_3496_),
    .Y(_3490_[3])
);

FILL FILL_3__8112_ (
);

FILL FILL_5__8878_ (
);

FILL SFILL104360x44050 (
);

FILL FILL_5__8458_ (
);

NAND2X1 _15598_ (
    .A(_6060_),
    .B(_6064_),
    .Y(_6065_)
);

AOI22X1 _15178_ (
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .B(_5606_),
    .C(_5570__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_5655_)
);

FILL FILL_3__16227_ (
);

FILL FILL_5__10748_ (
);

FILL SFILL3800x39050 (
);

FILL FILL_3__11782_ (
);

FILL FILL_3__11362_ (
);

FILL FILL_4__6875_ (
);

FILL FILL_0__16254_ (
);

FILL FILL_2__10775_ (
);

FILL FILL_1__9811_ (
);

FILL FILL_3__9737_ (
);

FILL FILL_5__14581_ (
);

FILL FILL_5__14161_ (
);

OAI21X1 _8881_ (
    .A(_1015_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1016_),
    .Y(_978_[19])
);

FILL FILL112440x50050 (
);

OAI21X1 _8461_ (
    .A(_796_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .C(_797_),
    .Y(_783_[7])
);

FILL FILL_6__7322_ (
);

DFFSR _8041_ (
    .Q(\datapath_1.regfile_1.regOut[9] [19]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_523_[19])
);

FILL FILL_4__13994_ (
);

FILL FILL_4__13574_ (
);

FILL FILL_4__13154_ (
);

NOR2X1 _11098_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2217_)
);

FILL FILL_2__7734_ (
);

FILL FILL_3__12987_ (
);

FILL FILL_3__12567_ (
);

FILL FILL_2__7314_ (
);

FILL FILL_3__12147_ (
);

FILL FILL_0__12594_ (
);

FILL SFILL89400x49050 (
);

FILL FILL_0__12174_ (
);

FILL FILL_4__8601_ (
);

FILL FILL_5_BUFX2_insert500 (
);

FILL FILL_5_BUFX2_insert501 (
);

FILL FILL_5__15786_ (
);

FILL FILL_5__15366_ (
);

FILL FILL_2__12501_ (
);

FILL FILL_5_BUFX2_insert502 (
);

FILL FILL_5_BUFX2_insert503 (
);

FILL FILL_5_BUFX2_insert504 (
);

NAND2X1 _9666_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1418_)
);

FILL FILL_5_BUFX2_insert505 (
);

NAND2X1 _9246_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1199_)
);

FILL FILL_5_BUFX2_insert506 (
);

FILL FILL_5_BUFX2_insert507 (
);

FILL FILL_5_BUFX2_insert508 (
);

FILL FILL_1__11914_ (
);

FILL FILL_4__14779_ (
);

FILL FILL_4__14359_ (
);

FILL FILL_5_BUFX2_insert509 (
);

FILL FILL_2__15393_ (
);

FILL FILL_0__8501_ (
);

FILL FILL_0__10907_ (
);

FILL FILL_2__8519_ (
);

FILL FILL_1__14386_ (
);

FILL FILL_5__6944_ (
);

FILL FILL_4__15720_ (
);

FILL FILL_1_BUFX2_insert1030 (
);

FILL FILL_4__15300_ (
);

FILL FILL_1_BUFX2_insert1031 (
);

FILL FILL_1_BUFX2_insert1032 (
);

FILL FILL_0__13799_ (
);

FILL FILL_1_BUFX2_insert1033 (
);

FILL FILL_3__9490_ (
);

NOR2X1 _13664_ (
    .A(_4171_),
    .B(_4156_),
    .Y(_4172_)
);

FILL FILL_1_BUFX2_insert1034 (
);

FILL FILL_0__13379_ (
);

OR2X2 _13244_ (
    .A(_3765_),
    .B(_3786_),
    .Y(_3787_)
);

FILL FILL_1_BUFX2_insert1035 (
);

FILL FILL_1_BUFX2_insert1036 (
);

FILL FILL_1_BUFX2_insert1037 (
);

FILL FILL_3__14713_ (
);

FILL FILL_1_BUFX2_insert1038 (
);

FILL FILL_1_BUFX2_insert1039 (
);

FILL FILL_1__6936_ (
);

FILL FILL_4__9806_ (
);

FILL SFILL94280x55050 (
);

FILL FILL_2__13706_ (
);

FILL FILL_0__14740_ (
);

FILL FILL_0__14320_ (
);

FILL FILL_5__11286_ (
);

FILL SFILL33640x30050 (
);

FILL FILL_2__16178_ (
);

FILL FILL_4__10699_ (
);

FILL FILL_4__10279_ (
);

FILL FILL_3__7803_ (
);

FILL FILL_5__7729_ (
);

FILL FILL_5__7309_ (
);

FILL FILL_2_BUFX2_insert630 (
);

FILL FILL_2_BUFX2_insert631 (
);

FILL FILL_2_BUFX2_insert632 (
);

FILL FILL_2_BUFX2_insert633 (
);

NAND3X1 _14869_ (
    .A(_5350_),
    .B(_5351_),
    .C(_5349_),
    .Y(_5352_)
);

FILL FILL_2_BUFX2_insert634 (
);

NOR2X1 _14449_ (
    .A(_4930_),
    .B(_4940_),
    .Y(_4941_)
);

FILL FILL_4__11640_ (
);

FILL FILL_2_BUFX2_insert635 (
);

INVX1 _14029_ (
    .A(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_4529_)
);

FILL FILL_4__11220_ (
);

FILL FILL_2_BUFX2_insert636 (
);

FILL FILL_3__15918_ (
);

FILL FILL_2_BUFX2_insert637 (
);

FILL FILL_2_BUFX2_insert638 (
);

FILL FILL_1__16112_ (
);

FILL FILL_2_BUFX2_insert639 (
);

FILL SFILL79400x47050 (
);

FILL FILL_3__10633_ (
);

FILL FILL_0__15945_ (
);

FILL FILL_0__15525_ (
);

NAND2X1 _15810_ (
    .A(_6271_),
    .B(_6265_),
    .Y(_6272_)
);

FILL FILL_0__15105_ (
);

FILL SFILL94280x10050 (
);

FILL FILL_0__10660_ (
);

FILL FILL_2__8272_ (
);

FILL FILL_0__10240_ (
);

FILL FILL_4__8198_ (
);

FILL SFILL79000x33050 (
);

FILL FILL_2__12098_ (
);

FILL FILL_5__13852_ (
);

FILL FILL_5__13432_ (
);

FILL FILL_5__13012_ (
);

OAI21X1 _7732_ (
    .A(_432_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_433_),
    .Y(_393_[20])
);

OAI21X1 _7312_ (
    .A(_213_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .C(_214_),
    .Y(_198_[8])
);

FILL FILL_4__12845_ (
);

FILL FILL_4__12425_ (
);

FILL FILL_4__12005_ (
);

OAI21X1 _10789_ (
    .A(_1982_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .C(_1983_),
    .Y(_1953_[15])
);

FILL FILL_0__8098_ (
);

OAI21X1 _10369_ (
    .A(_1763_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1764_),
    .Y(_1758_[3])
);

FILL FILL_3__11838_ (
);

FILL FILL_1__12872_ (
);

FILL FILL_3__11418_ (
);

FILL FILL_1__12452_ (
);

FILL FILL_1__12032_ (
);

FILL SFILL84280x53050 (
);

FILL FILL_2__9897_ (
);

FILL FILL_0__11865_ (
);

FILL FILL_2__9477_ (
);

FILL FILL_0__11445_ (
);

AND2X2 _11730_ (
    .A(_2826_),
    .B(_2168_),
    .Y(_2827_)
);

FILL FILL_0__11025_ (
);

INVX1 _11310_ (
    .A(_2229_),
    .Y(_2429_)
);

FILL FILL_6__15644_ (
);

FILL FILL_5__7482_ (
);

FILL FILL_6__15224_ (
);

FILL FILL_5__7062_ (
);

FILL SFILL39240x13050 (
);

FILL FILL_5__14637_ (
);

FILL FILL_3__15671_ (
);

FILL FILL_5__14217_ (
);

FILL FILL_3__15251_ (
);

DFFSR _8937_ (
    .Q(\datapath_1.regfile_1.regOut[16] [19]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_978_[19])
);

NAND2X1 _8517_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_835_)
);

FILL FILL_1__7474_ (
);

FILL FILL_1__7054_ (
);

FILL SFILL114440x79050 (
);

FILL FILL_2__14664_ (
);

FILL FILL_2__14244_ (
);

FILL FILL_3_BUFX2_insert90 (
);

FILL FILL_3_BUFX2_insert91 (
);

FILL FILL_1__13657_ (
);

FILL FILL_1__13237_ (
);

FILL FILL_3_BUFX2_insert92 (
);

FILL FILL_3_BUFX2_insert93 (
);

FILL SFILL94200x5050 (
);

FILL FILL_3_BUFX2_insert94 (
);

FILL FILL_3_BUFX2_insert95 (
);

FILL SFILL84200x51050 (
);

FILL FILL_3_BUFX2_insert96 (
);

FILL FILL_1_BUFX2_insert650 (
);

FILL FILL_1_BUFX2_insert651 (
);

FILL FILL_3__8761_ (
);

FILL FILL_3_BUFX2_insert97 (
);

FILL FILL_1_BUFX2_insert652 (
);

FILL FILL_3_BUFX2_insert98 (
);

DFFSR _12935_ (
    .Q(\datapath_1.a [16]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3555_[16])
);

FILL FILL_3__8341_ (
);

FILL FILL_1_BUFX2_insert653 (
);

NAND2X1 _12515_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [25]),
    .Y(_3410_)
);

FILL FILL_3_BUFX2_insert99 (
);

FILL FILL_1_BUFX2_insert654 (
);

FILL FILL_1_BUFX2_insert655 (
);

FILL FILL_1_BUFX2_insert656 (
);

FILL FILL_5__8267_ (
);

FILL FILL_1_BUFX2_insert657 (
);

FILL FILL_1_BUFX2_insert658 (
);

FILL FILL_1_BUFX2_insert659 (
);

FILL FILL_6__11564_ (
);

FILL FILL_6__11144_ (
);

FILL SFILL13640x71050 (
);

FILL SFILL29240x56050 (
);

FILL FILL_3__16036_ (
);

FILL SFILL109480x51050 (
);

FILL FILL_5__10977_ (
);

FILL FILL_5__10557_ (
);

FILL FILL_5__10137_ (
);

FILL FILL_3__11591_ (
);

FILL FILL_1__8259_ (
);

FILL FILL_3__11171_ (
);

FILL FILL_2__15869_ (
);

FILL FILL_2__15449_ (
);

FILL FILL_2__15029_ (
);

FILL FILL_0__16063_ (
);

FILL FILL_2__10164_ (
);

FILL FILL_1__9620_ (
);

FILL FILL_3__9546_ (
);

FILL FILL_4__10911_ (
);

FILL FILL_3__9126_ (
);

FILL FILL_5__14390_ (
);

DFFSR _8690_ (
    .Q(\datapath_1.regfile_1.regOut[14] [28]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_848_[28])
);

FILL FILL_1__15803_ (
);

NAND2X1 _8270_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_711_)
);

FILL FILL_4__13383_ (
);

FILL FILL_2__7963_ (
);

BUFX2 BUFX2_insert320 (
    .A(_5480_),
    .Y(_5480__bF$buf0)
);

FILL FILL_2__7543_ (
);

FILL FILL_3__12376_ (
);

BUFX2 BUFX2_insert321 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf7 )
);

FILL FILL_2__7123_ (
);

BUFX2 BUFX2_insert322 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf6 )
);

BUFX2 BUFX2_insert323 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf5 )
);

BUFX2 BUFX2_insert324 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf4 )
);

FILL FILL_4__7889_ (
);

FILL FILL_6__13710_ (
);

BUFX2 BUFX2_insert325 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf3 )
);

FILL FILL_4__7469_ (
);

BUFX2 BUFX2_insert326 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf2 )
);

FILL FILL_4__7049_ (
);

BUFX2 BUFX2_insert327 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf1 )
);

FILL FILL_2__11789_ (
);

BUFX2 BUFX2_insert328 (
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf0 )
);

FILL FILL_2__11369_ (
);

BUFX2 BUFX2_insert329 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf4 )
);

FILL FILL_5__12703_ (
);

FILL FILL_4__8830_ (
);

FILL FILL_2__12730_ (
);

FILL FILL_5__15595_ (
);

FILL FILL_5__15175_ (
);

FILL FILL_2__12310_ (
);

NAND2X1 _9895_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1530_)
);

FILL FILL_0__7369_ (
);

NAND2X1 _9475_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1311_)
);

DFFSR _9055_ (
    .Q(\datapath_1.regfile_1.regOut[17] [9]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_1043_[9])
);

FILL FILL_4__14588_ (
);

FILL FILL_1__11723_ (
);

FILL FILL_4__14168_ (
);

FILL FILL_1__11303_ (
);

FILL FILL_0__8730_ (
);

FILL FILL_2__8748_ (
);

FILL FILL_2__8328_ (
);

FILL FILL_0__8310_ (
);

FILL FILL_1__14195_ (
);

OAI22X1 _13893_ (
    .A(_4394_),
    .B(_3893__bF$buf3),
    .C(_3944__bF$buf1),
    .D(_4395_),
    .Y(_4396_)
);

NOR2X1 _13473_ (
    .A(_3984_),
    .B(_3979_),
    .Y(_3985_)
);

DFFSR _13053_ (
    .Q(_2_[6]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3620_[6])
);

FILL FILL_5__13908_ (
);

FILL FILL_3__14942_ (
);

FILL FILL_3__14522_ (
);

FILL FILL_3__14102_ (
);

FILL FILL_4__9615_ (
);

FILL FILL_2__13935_ (
);

FILL FILL_2__13515_ (
);

FILL FILL_5__11095_ (
);

FILL FILL_1__12508_ (
);

FILL FILL_0__9935_ (
);

FILL FILL_3__7612_ (
);

FILL FILL_0__9515_ (
);

FILL SFILL104360x39050 (
);

FILL FILL_5__7958_ (
);

FILL FILL_5__7118_ (
);

FILL FILL_4__16314_ (
);

OAI22X1 _14678_ (
    .A(_3947__bF$buf2),
    .B(_5163_),
    .C(_3977__bF$buf0),
    .D(_5164_),
    .Y(_5165_)
);

INVX1 _14258_ (
    .A(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_4754_)
);

FILL FILL_3__15727_ (
);

FILL FILL_3__15307_ (
);

FILL FILL_1__16341_ (
);

FILL FILL112040x76050 (
);

FILL FILL_3__10442_ (
);

FILL FILL_3__10022_ (
);

FILL FILL_0__15754_ (
);

FILL FILL_0__15334_ (
);

FILL FILL_2__8081_ (
);

FILL FILL_5__13661_ (
);

FILL FILL_5__13241_ (
);

FILL FILL112440x45050 (
);

OAI21X1 _7961_ (
    .A(_544_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_545_),
    .Y(_523_[11])
);

DFFSR _7541_ (
    .Q(\datapath_1.regfile_1.regOut[5] [31]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_263_[31])
);

NAND2X1 _7121_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_128_)
);

FILL FILL_4__12654_ (
);

FILL FILL_4__12234_ (
);

DFFSR _10598_ (
    .Q(\datapath_1.regfile_1.regOut[29] [16]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_1823_[16])
);

NAND2X1 _10178_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1678_)
);

FILL FILL_3__11647_ (
);

FILL FILL_3__11227_ (
);

FILL FILL_1__12261_ (
);

FILL FILL112040x31050 (
);

FILL FILL_0__16119_ (
);

OAI21X1 _16404_ (
    .A(_6822_),
    .B(gnd),
    .C(_6823_),
    .Y(_6769_[27])
);

FILL FILL_2__9286_ (
);

FILL FILL_0__11674_ (
);

FILL FILL_0__11254_ (
);

FILL FILL_5__7291_ (
);

FILL FILL_5__14866_ (
);

FILL FILL_5__14446_ (
);

FILL FILL_5__14026_ (
);

FILL FILL_3__15480_ (
);

FILL FILL_3__15060_ (
);

NAND2X1 _8746_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_947_)
);

NAND2X1 _8326_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_728_)
);

FILL FILL_4__13859_ (
);

FILL FILL_4__13439_ (
);

FILL FILL_2__14893_ (
);

FILL FILL_2__14473_ (
);

FILL FILL_4__13019_ (
);

FILL FILL_2__14053_ (
);

FILL FILL_1__13886_ (
);

FILL FILL_1__13466_ (
);

FILL FILL_1__13046_ (
);

FILL FILL_4__14800_ (
);

FILL FILL_3__8990_ (
);

FILL FILL_0__12879_ (
);

FILL FILL_3__8570_ (
);

NAND2X1 _12744_ (
    .A(IRWrite_bF$buf5),
    .B(memoryOutData[16]),
    .Y(_3522_)
);

FILL FILL_0__12459_ (
);

FILL FILL_0__12039_ (
);

NAND3X1 _12324_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf1),
    .Y(_3282_)
);

FILL FILL_5__8496_ (
);

FILL FILL_5__8076_ (
);

FILL FILL_0__13820_ (
);

FILL FILL_0__13400_ (
);

FILL FILL_3__16265_ (
);

FILL FILL_5__10786_ (
);

FILL FILL_1__8488_ (
);

FILL FILL_5__10366_ (
);

FILL FILL_1__8068_ (
);

FILL FILL_2__15678_ (
);

FILL FILL_2__15258_ (
);

FILL FILL_0__16292_ (
);

FILL FILL_2__10393_ (
);

FILL SFILL23720x61050 (
);

FILL FILL_3__9775_ (
);

FILL FILL_3__9355_ (
);

NOR2X1 _13949_ (
    .A(_4447_),
    .B(_4450_),
    .Y(_4451_)
);

INVX8 _13529_ (
    .A(_3966__bF$buf1),
    .Y(_4040_)
);

FILL FILL_4__10300_ (
);

INVX1 _13109_ (
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_3704_)
);

FILL SFILL34600x4050 (
);

FILL FILL_1__15612_ (
);

FILL FILL_6__12578_ (
);

FILL FILL_0__14605_ (
);

FILL SFILL4360x59050 (
);

FILL SFILL3720x50 (
);

FILL FILL_2__7352_ (
);

FILL FILL_3__12185_ (
);

FILL FILL_4__7698_ (
);

FILL FILL_2__11598_ (
);

FILL FILL_2__11178_ (
);

FILL FILL_5__12512_ (
);

FILL SFILL8680x67050 (
);

FILL FILL_4__11925_ (
);

FILL FILL_4__11505_ (
);

FILL SFILL23240x54050 (
);

FILL FILL_0__7598_ (
);

FILL FILL_0__7178_ (
);

INVX1 _9284_ (
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_1224_)
);

FILL FILL_3__10918_ (
);

FILL FILL_1__11952_ (
);

FILL FILL_4__14397_ (
);

FILL FILL_1__11532_ (
);

FILL FILL_1__11112_ (
);

FILL SFILL84280x48050 (
);

FILL FILL_2__8977_ (
);

FILL FILL_0__10945_ (
);

OAI21X1 _10810_ (
    .A(_1996_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .C(_1997_),
    .Y(_1953_[22])
);

FILL FILL_2__8137_ (
);

FILL FILL_0__10525_ (
);

FILL SFILL109160x70050 (
);

FILL FILL_0__10105_ (
);

FILL FILL_5__6982_ (
);

FILL SFILL23640x23050 (
);

NAND2X1 _13282_ (
    .A(_3750_),
    .B(_3820_),
    .Y(_3821_)
);

FILL FILL_5__13717_ (
);

FILL FILL_3__14751_ (
);

FILL FILL_3__14331_ (
);

FILL FILL_1__6974_ (
);

FILL FILL_4__9424_ (
);

FILL FILL_4__9004_ (
);

FILL SFILL8680x22050 (
);

FILL FILL_2__13744_ (
);

FILL SFILL84680x17050 (
);

FILL FILL_2__13324_ (
);

FILL FILL_5__16189_ (
);

FILL SFILL44120x50050 (
);

FILL FILL_1__12737_ (
);

FILL FILL_1__12317_ (
);

FILL FILL_0__9744_ (
);

FILL FILL_3__7841_ (
);

FILL FILL_3__7421_ (
);

FILL FILL_5__7347_ (
);

FILL FILL_4__16123_ (
);

FILL SFILL13640x66050 (
);

INVX1 _14487_ (
    .A(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_4978_)
);

INVX1 _14067_ (
    .A(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_4567_)
);

FILL FILL_3__15956_ (
);

FILL FILL_3__15536_ (
);

FILL SFILL109480x46050 (
);

FILL FILL_3__15116_ (
);

FILL FILL_1__16150_ (
);

FILL FILL_1__7759_ (
);

FILL FILL_3__10671_ (
);

FILL FILL_1__7339_ (
);

FILL FILL_3__10251_ (
);

FILL SFILL8600x20050 (
);

FILL FILL_2__14949_ (
);

FILL FILL_0__15983_ (
);

FILL FILL_2__14529_ (
);

FILL FILL_0__15563_ (
);

FILL FILL_2__14109_ (
);

FILL FILL_0__15143_ (
);

FILL SFILL114440x29050 (
);

FILL FILL_1__8700_ (
);

FILL FILL_3__8626_ (
);

FILL FILL_3__8206_ (
);

FILL FILL_5__13890_ (
);

FILL FILL_5__13470_ (
);

FILL SFILL74280x46050 (
);

DFFSR _7770_ (
    .Q(\datapath_1.regfile_1.regOut[7] [4]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_393_[4])
);

NAND2X1 _7350_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_240_)
);

FILL FILL_4__12883_ (
);

FILL FILL_4__12463_ (
);

FILL FILL_4__12043_ (
);

FILL SFILL13640x21050 (
);

FILL FILL_3__11876_ (
);

FILL FILL_5__9913_ (
);

FILL FILL_3__11456_ (
);

FILL FILL_1__12490_ (
);

FILL FILL_3__11036_ (
);

FILL FILL_1__12070_ (
);

FILL FILL_4__6969_ (
);

FILL FILL_0__16348_ (
);

OAI22X1 _16213_ (
    .A(_5335_),
    .B(_5539__bF$buf3),
    .C(_5503__bF$buf3),
    .D(_5346_),
    .Y(_6664_)
);

FILL FILL_2__10449_ (
);

FILL SFILL38840x70050 (
);

FILL FILL_2__10029_ (
);

FILL FILL_0__11483_ (
);

FILL FILL_2__9095_ (
);

FILL FILL_0__11063_ (
);

FILL FILL_1__9905_ (
);

FILL FILL_2__11810_ (
);

FILL FILL_5__14675_ (
);

FILL SFILL74200x44050 (
);

FILL FILL_5__14255_ (
);

FILL FILL_0__6869_ (
);

NAND2X1 _8975_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1059_)
);

DFFSR _8555_ (
    .Q(\datapath_1.regfile_1.regOut[13] [21]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_783_[21])
);

INVX1 _8135_ (
    .A(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_641_)
);

FILL FILL_1__7092_ (
);

FILL FILL_4__13668_ (
);

FILL FILL_1__10803_ (
);

FILL FILL_4__13248_ (
);

FILL FILL_2__14282_ (
);

FILL FILL_0__7810_ (
);

FILL FILL_2__7828_ (
);

FILL FILL_1__13695_ (
);

FILL FILL_1__13275_ (
);

FILL SFILL99480x50050 (
);

NAND2X1 _12973_ (
    .A(vdd),
    .B(\datapath_1.rd2 [7]),
    .Y(_3634_)
);

DFFSR _12553_ (
    .Q(ALUOut[18]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[18])
);

FILL FILL_0__12268_ (
);

INVX1 _12133_ (
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_3142_)
);

FILL FILL_3__13602_ (
);

FILL FILL_3__16074_ (
);

FILL FILL112120x64050 (
);

FILL FILL_5__10175_ (
);

FILL FILL_2__15487_ (
);

FILL FILL_2__15067_ (
);

FILL FILL_5__16401_ (
);

FILL FILL_4__15814_ (
);

FILL FILL_3__9164_ (
);

OAI22X1 _13758_ (
    .A(_3884__bF$buf1),
    .B(_4262_),
    .C(_3977__bF$buf1),
    .D(_4263_),
    .Y(_4264_)
);

NOR2X1 _13338_ (
    .A(_3860_),
    .B(_3858_),
    .Y(\datapath_1.regfile_1.regEn [21])
);

FILL FILL_3__14807_ (
);

FILL FILL_1__15841_ (
);

FILL FILL_1__15421_ (
);

FILL FILL_1__15001_ (
);

FILL FILL_6__12387_ (
);

FILL FILL_0__14834_ (
);

FILL FILL_0__14414_ (
);

BUFX2 BUFX2_insert700 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf1 )
);

FILL FILL_2__7581_ (
);

FILL FILL_2__7161_ (
);

BUFX2 BUFX2_insert701 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf0 )
);

FILL SFILL64200x42050 (
);

BUFX2 BUFX2_insert702 (
    .A(_3034_),
    .Y(_3034__bF$buf4)
);

BUFX2 BUFX2_insert703 (
    .A(_3034_),
    .Y(_3034__bF$buf3)
);

BUFX2 BUFX2_insert704 (
    .A(_3034_),
    .Y(_3034__bF$buf2)
);

BUFX2 BUFX2_insert705 (
    .A(_3034_),
    .Y(_3034__bF$buf1)
);

BUFX2 BUFX2_insert706 (
    .A(_3034_),
    .Y(_3034__bF$buf0)
);

FILL FILL_4__7087_ (
);

BUFX2 BUFX2_insert707 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf4 )
);

BUFX2 BUFX2_insert708 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf3 )
);

BUFX2 BUFX2_insert709 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf2 )
);

FILL FILL_5__12741_ (
);

FILL FILL_5__12321_ (
);

FILL FILL_4__11734_ (
);

FILL FILL_4__11314_ (
);

FILL FILL_1__16206_ (
);

INVX1 _9093_ (
    .A(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_1117_)
);

FILL FILL_1__11761_ (
);

FILL FILL_3__10307_ (
);

FILL FILL_1__11341_ (
);

AOI22X1 _15904_ (
    .A(_5565__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [21]),
    .C(\datapath_1.regfile_1.regOut[5] [21]),
    .D(_5700_),
    .Y(_6363_)
);

FILL FILL_0__15619_ (
);

FILL FILL_2__8786_ (
);

FILL FILL_0__10754_ (
);

FILL FILL_2__8366_ (
);

FILL FILL_6__14953_ (
);

FILL FILL_6__14533_ (
);

INVX1 _13091_ (
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_3692_)
);

FILL FILL_5__13946_ (
);

FILL FILL_3__14980_ (
);

FILL FILL_5__13526_ (
);

FILL FILL_3__14560_ (
);

FILL FILL_5__13106_ (
);

FILL FILL_3__14140_ (
);

NAND2X1 _7826_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_476_)
);

DFFSR _7406_ (
    .Q(\datapath_1.regfile_1.regOut[4] [24]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_198_[24])
);

FILL FILL_4_BUFX2_insert540 (
);

FILL FILL_4__9653_ (
);

FILL FILL_4_BUFX2_insert541 (
);

FILL FILL_4_BUFX2_insert542 (
);

FILL FILL_4__9233_ (
);

FILL FILL_4__12519_ (
);

FILL FILL_4_BUFX2_insert543 (
);

FILL FILL_2__13973_ (
);

FILL FILL_4_BUFX2_insert544 (
);

FILL FILL_2__13553_ (
);

FILL FILL_2__13133_ (
);

FILL FILL_4_BUFX2_insert545 (
);

FILL FILL_6__9999_ (
);

FILL FILL_4_BUFX2_insert546 (
);

FILL FILL_4_BUFX2_insert547 (
);

FILL FILL_4_BUFX2_insert548 (
);

FILL FILL_4_BUFX2_insert549 (
);

FILL FILL_1__12966_ (
);

FILL FILL_1__12126_ (
);

FILL SFILL115320x21050 (
);

FILL FILL_0__11959_ (
);

FILL FILL_0__9553_ (
);

FILL FILL_3__7230_ (
);

FILL FILL_0__9133_ (
);

AOI22X1 _11824_ (
    .A(_2478_),
    .B(_2353_),
    .C(_2352_),
    .D(_2341__bF$buf3),
    .Y(_2914_)
);

FILL FILL_0__11539_ (
);

NOR2X1 _11404_ (
    .A(_2262_),
    .B(_2520_),
    .Y(_2521_)
);

FILL FILL_0__11119_ (
);

FILL FILL_5__7996_ (
);

FILL FILL_5__7576_ (
);

FILL SFILL58920x62050 (
);

FILL FILL_4__16352_ (
);

OAI22X1 _14296_ (
    .A(_4789_),
    .B(_3884__bF$buf3),
    .C(_3881_),
    .D(_4790_),
    .Y(_4791_)
);

FILL FILL_3__15765_ (
);

FILL FILL_0__12900_ (
);

FILL FILL_3__15345_ (
);

FILL SFILL39000x5050 (
);

FILL FILL_1__7988_ (
);

FILL FILL_1__7568_ (
);

FILL SFILL13720x1050 (
);

FILL FILL_3__10060_ (
);

FILL FILL_2__14758_ (
);

FILL FILL_2__14338_ (
);

FILL FILL_0__15792_ (
);

FILL FILL_0__15372_ (
);

FILL SFILL13640x6050 (
);

FILL SFILL23720x56050 (
);

FILL FILL_3__8855_ (
);

FILL FILL_3__8015_ (
);

INVX1 _12609_ (
    .A(\datapath_1.Data [14]),
    .Y(_3452_)
);

FILL FILL_4__12272_ (
);

FILL FILL_2__6852_ (
);

FILL FILL_5__9722_ (
);

FILL FILL_3__11685_ (
);

FILL FILL_3__11265_ (
);

FILL FILL_0__16157_ (
);

DFFSR _16442_ (
    .Q(\datapath_1.regfile_1.regOut[0] [25]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_6769_[25])
);

NOR3X1 _16022_ (
    .A(_5515__bF$buf1),
    .B(_5098_),
    .C(_5521__bF$buf0),
    .Y(_6478_)
);

FILL FILL_2__10678_ (
);

FILL FILL_2__10258_ (
);

FILL FILL_0__11292_ (
);

FILL FILL_6__15071_ (
);

FILL FILL_3_BUFX2_insert560 (
);

FILL SFILL109560x79050 (
);

FILL FILL_3_BUFX2_insert561 (
);

FILL SFILL23720x11050 (
);

FILL FILL_3_BUFX2_insert562 (
);

FILL FILL_3_BUFX2_insert563 (
);

FILL FILL_5__14484_ (
);

FILL FILL_5__14064_ (
);

FILL FILL_3_BUFX2_insert564 (
);

FILL FILL_3_BUFX2_insert565 (
);

INVX1 _8784_ (
    .A(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_972_)
);

FILL FILL_3_BUFX2_insert566 (
);

INVX1 _8364_ (
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_753_)
);

FILL FILL_3_BUFX2_insert567 (
);

FILL FILL_3_BUFX2_insert568 (
);

FILL FILL_3_BUFX2_insert569 (
);

FILL FILL_4__13897_ (
);

FILL FILL_4__13477_ (
);

FILL SFILL48920x60050 (
);

FILL FILL_2__14091_ (
);

FILL FILL_2__7637_ (
);

FILL FILL_2__7217_ (
);

FILL FILL_1__13084_ (
);

INVX1 _12782_ (
    .A(\control_1.op [3]),
    .Y(_3547_)
);

FILL FILL_0__12497_ (
);

NAND2X1 _12362_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [6]),
    .Y(_3307_)
);

FILL FILL_0__12077_ (
);

FILL FILL_3__13831_ (
);

FILL FILL_3__13411_ (
);

FILL FILL_4__8504_ (
);

FILL SFILL8680x17050 (
);

FILL SFILL13720x54050 (
);

FILL FILL_5__15689_ (
);

FILL FILL_2__12824_ (
);

FILL SFILL44120x45050 (
);

FILL FILL_2__12404_ (
);

FILL FILL_5__15269_ (
);

INVX1 _9989_ (
    .A(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_1572_)
);

DFFSR _9569_ (
    .Q(\datapath_1.regfile_1.regOut[21] [11]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_1303_[11])
);

FILL SFILL109560x34050 (
);

OAI21X1 _9149_ (
    .A(_1153_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1154_),
    .Y(_1108_[23])
);

FILL FILL_1__11817_ (
);

FILL FILL_2__15296_ (
);

FILL FILL_5__16210_ (
);

FILL FILL_3__6921_ (
);

FILL FILL_0__8824_ (
);

FILL FILL_0__8404_ (
);

FILL FILL_1__14289_ (
);

FILL FILL_5__6847_ (
);

FILL FILL_0_BUFX2_insert690 (
);

FILL FILL_4__15623_ (
);

FILL FILL_0_BUFX2_insert691 (
);

FILL FILL_4__15203_ (
);

FILL FILL_0_BUFX2_insert692 (
);

FILL FILL_0_BUFX2_insert693 (
);

FILL FILL_0_BUFX2_insert694 (
);

NAND3X1 _13987_ (
    .A(_4477_),
    .B(_4480_),
    .C(_4487_),
    .Y(_4488_)
);

FILL FILL_3__9393_ (
);

FILL FILL_0_BUFX2_insert695 (
);

NOR2X1 _13567_ (
    .A(_4073_),
    .B(_4076_),
    .Y(_4077_)
);

OAI21X1 _13147_ (
    .A(_3728_),
    .B(PCEn_bF$buf7),
    .C(_3729_),
    .Y(_3685_[22])
);

FILL FILL_0_BUFX2_insert696 (
);

FILL FILL_0_BUFX2_insert697 (
);

FILL FILL_3__14616_ (
);

FILL FILL_0_BUFX2_insert698 (
);

FILL FILL_1__15650_ (
);

FILL FILL_0_BUFX2_insert699 (
);

FILL FILL_1__15230_ (
);

FILL FILL_1__6839_ (
);

FILL SFILL8600x15050 (
);

FILL FILL_2__13609_ (
);

FILL FILL_0__14643_ (
);

FILL FILL_0__14223_ (
);

FILL FILL_5__11189_ (
);

FILL FILL_0__9609_ (
);

FILL FILL_3__7706_ (
);

FILL FILL_5__12970_ (
);

FILL FILL_5__12130_ (
);

BUFX2 _6850_ (
    .A(_1_[12]),
    .Y(memoryAddress[12])
);

FILL FILL_4__16408_ (
);

FILL FILL_4__11963_ (
);

FILL FILL_4__11543_ (
);

FILL FILL_4__11123_ (
);

FILL SFILL13640x16050 (
);

FILL FILL_1__16015_ (
);

FILL FILL_3__10956_ (
);

FILL FILL_3__10536_ (
);

FILL FILL_1__11990_ (
);

FILL FILL_3__10116_ (
);

FILL FILL_1__11570_ (
);

FILL FILL_1__11150_ (
);

FILL FILL_0__15848_ (
);

OAI22X1 _15713_ (
    .A(_4714_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf2),
    .D(_6176_),
    .Y(_6177_)
);

FILL FILL_0__15428_ (
);

FILL FILL_0__15008_ (
);

FILL SFILL38840x65050 (
);

FILL FILL_0__10983_ (
);

FILL FILL_2__8595_ (
);

FILL FILL_0__10563_ (
);

FILL FILL_0__10143_ (
);

FILL FILL_5__13755_ (
);

FILL FILL_5__13335_ (
);

INVX1 _7635_ (
    .A(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_389_)
);

INVX1 _7215_ (
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_170_)
);

FILL FILL_4__9882_ (
);

FILL FILL_4__9462_ (
);

FILL FILL_4__12748_ (
);

FILL FILL_4__9042_ (
);

FILL FILL_2__13782_ (
);

FILL FILL_4__12328_ (
);

FILL FILL_2__13362_ (
);

FILL FILL_2__6908_ (
);

FILL FILL112200x52050 (
);

FILL FILL_1__12775_ (
);

FILL FILL_1__12355_ (
);

FILL FILL_0__9782_ (
);

FILL FILL_0__11768_ (
);

FILL FILL_0__9362_ (
);

FILL FILL_0__11348_ (
);

OAI21X1 _11633_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .C(_2620_),
    .Y(_2737_)
);

OAI21X1 _11213_ (
    .A(_2112_),
    .B(\datapath_1.alu_1.ALUInB [30]),
    .C(_2331_),
    .Y(_2332_)
);

FILL SFILL38840x20050 (
);

FILL FILL_6__15127_ (
);

FILL FILL_4__16161_ (
);

FILL FILL_6__10682_ (
);

FILL FILL_3__15994_ (
);

FILL FILL_3__15574_ (
);

FILL FILL_3__15154_ (
);

FILL FILL112120x59050 (
);

FILL FILL_1__7377_ (
);

FILL SFILL64280x39050 (
);

FILL FILL_2__14987_ (
);

FILL FILL_2__14567_ (
);

FILL FILL_2__14147_ (
);

FILL FILL_0__15181_ (
);

FILL FILL_5__15901_ (
);

FILL FILL_3__8244_ (
);

INVX1 _12838_ (
    .A(\datapath_1.a [5]),
    .Y(_3564_)
);

INVX1 _12418_ (
    .A(ALUOut[25]),
    .Y(_3344_)
);

FILL FILL_1__14921_ (
);

FILL SFILL28840x63050 (
);

FILL FILL_1__14501_ (
);

FILL FILL_6__11047_ (
);

FILL FILL_4__12081_ (
);

FILL FILL_0__13914_ (
);

FILL FILL_3__16359_ (
);

FILL SFILL33800x46050 (
);

FILL SFILL64200x37050 (
);

FILL FILL_5__9531_ (
);

FILL FILL_3__11494_ (
);

FILL FILL_5__9111_ (
);

FILL FILL_3__11074_ (
);

FILL FILL112120x14050 (
);

FILL FILL_0__16386_ (
);

NAND3X1 _16251_ (
    .A(_6695_),
    .B(_6700_),
    .C(_6699_),
    .Y(_6701_)
);

FILL FILL_2__10487_ (
);

FILL FILL_2__10067_ (
);

FILL FILL_5__11821_ (
);

FILL FILL_1__9523_ (
);

FILL FILL_5__11401_ (
);

FILL FILL_1__9103_ (
);

FILL FILL_3__9869_ (
);

FILL FILL_4__10814_ (
);

FILL FILL_3__9029_ (
);

FILL FILL_5__14293_ (
);

FILL FILL_1__15706_ (
);

INVX1 _8593_ (
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_865_)
);

DFFSR _8173_ (
    .Q(\datapath_1.regfile_1.regOut[10] [23]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_588_[23])
);

FILL FILL_1__10421_ (
);

FILL FILL_4__13286_ (
);

FILL FILL_1__10001_ (
);

FILL FILL_2__7866_ (
);

FILL FILL_3__12699_ (
);

FILL FILL_2__7446_ (
);

FILL FILL_3__12279_ (
);

FILL FILL_6__13613_ (
);

INVX1 _12591_ (
    .A(\datapath_1.Data [8]),
    .Y(_3440_)
);

OAI21X1 _12171_ (
    .A(_3166_),
    .B(ALUSrcA_bF$buf1),
    .C(_3167_),
    .Y(\datapath_1.alu_1.ALUInA [18])
);

FILL FILL_5__12606_ (
);

FILL FILL_3__13640_ (
);

FILL FILL_3__13220_ (
);

NAND2X1 _6906_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_5_)
);

FILL FILL_4__8733_ (
);

FILL FILL_4__8313_ (
);

FILL FILL_2__12633_ (
);

FILL FILL_5__15498_ (
);

FILL FILL_2__12213_ (
);

FILL FILL_5__15078_ (
);

OAI21X1 _9798_ (
    .A(_1484_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1485_),
    .Y(_1433_[26])
);

OAI21X1 _9378_ (
    .A(_1265_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1266_),
    .Y(_1238_[14])
);

FILL FILL_1__11626_ (
);

FILL SFILL43960x50 (
);

FILL FILL_1__11206_ (
);

FILL SFILL18840x61050 (
);

FILL FILL_0__8633_ (
);

NOR2X1 _10904_ (
    .A(_2047_),
    .B(_2051_),
    .Y(Branch)
);

FILL FILL_0__10619_ (
);

FILL FILL_0__8213_ (
);

FILL FILL_1__14098_ (
);

FILL FILL_4__15852_ (
);

FILL FILL_4__15432_ (
);

FILL FILL_4__15012_ (
);

NOR2X1 _13796_ (
    .A(_4300_),
    .B(_4297_),
    .Y(_4301_)
);

NOR2X1 _13376_ (
    .A(\datapath_1.PCJump [21]),
    .B(_3887_),
    .Y(_3888_)
);

FILL FILL_3__14845_ (
);

FILL FILL_3__14425_ (
);

FILL FILL_3__14005_ (
);

FILL FILL_4__9938_ (
);

FILL FILL_4__9518_ (
);

FILL FILL_2__13838_ (
);

FILL FILL_0__14872_ (
);

FILL FILL_2__13418_ (
);

FILL FILL_0__14452_ (
);

FILL FILL_0__14032_ (
);

FILL FILL_3__7935_ (
);

FILL FILL_0__9418_ (
);

FILL FILL_4__16217_ (
);

FILL FILL_4__11772_ (
);

FILL FILL_4__11352_ (
);

FILL FILL_1__16244_ (
);

FILL FILL_3__10765_ (
);

FILL FILL_0__15657_ (
);

NAND3X1 _15942_ (
    .A(_6397_),
    .B(_6399_),
    .C(_6396_),
    .Y(_6400_)
);

FILL FILL_0__15237_ (
);

NOR2X1 _15522_ (
    .A(_5989_),
    .B(_5990_),
    .Y(_5991_)
);

NAND3X1 _15102_ (
    .A(_5575_),
    .B(_5580_),
    .C(_5578_),
    .Y(_5581_)
);

FILL FILL_0__10792_ (
);

FILL FILL_0__10372_ (
);

FILL FILL_5__13984_ (
);

FILL FILL_5__13564_ (
);

FILL FILL_5__13144_ (
);

INVX1 _7864_ (
    .A(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_501_)
);

INVX1 _7444_ (
    .A(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_282_)
);

DFFSR _7024_ (
    .Q(\datapath_1.regfile_1.regOut[1] [26]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_3_[26])
);

FILL FILL_4_BUFX2_insert920 (
);

FILL FILL_4_BUFX2_insert921 (
);

FILL FILL_4__9271_ (
);

FILL FILL_4__12977_ (
);

FILL FILL_4_BUFX2_insert922 (
);

FILL FILL_4_BUFX2_insert923 (
);

FILL SFILL48920x55050 (
);

FILL FILL_2__13591_ (
);

FILL FILL_4__12137_ (
);

FILL FILL_4_BUFX2_insert924 (
);

FILL FILL_2__13171_ (
);

FILL FILL_4_BUFX2_insert925 (
);

FILL FILL_4_BUFX2_insert926 (
);

FILL FILL_4_BUFX2_insert927 (
);

FILL FILL_4_BUFX2_insert928 (
);

FILL FILL_4_BUFX2_insert929 (
);

FILL FILL_1__12584_ (
);

FILL FILL_1__12164_ (
);

NOR2X1 _16307_ (
    .A(_6753_),
    .B(_6755_),
    .Y(_6756_)
);

FILL FILL_0__11997_ (
);

FILL FILL_0__9591_ (
);

FILL FILL_0__9171_ (
);

NAND2X1 _11862_ (
    .A(_2627_),
    .B(_2948_),
    .Y(_2949_)
);

FILL FILL_0__11577_ (
);

XNOR2X1 _11442_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2558_)
);

FILL FILL_0__11157_ (
);

AND2X2 _11022_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2141_)
);

FILL FILL_3__12911_ (
);

FILL FILL_4__16390_ (
);

FILL FILL_5__7194_ (
);

FILL SFILL13720x49050 (
);

FILL FILL_2__11904_ (
);

FILL FILL_5__14769_ (
);

FILL FILL_5__14349_ (
);

FILL FILL_3__15383_ (
);

FILL SFILL109560x29050 (
);

OAI21X1 _8649_ (
    .A(_901_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_902_),
    .Y(_848_[27])
);

OAI21X1 _8229_ (
    .A(_682_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .C(_683_),
    .Y(_653_[15])
);

FILL FILL_1__7186_ (
);

FILL FILL_2__14796_ (
);

FILL FILL_2__14376_ (
);

FILL FILL_5__15710_ (
);

FILL SFILL48920x10050 (
);

FILL FILL_1__13789_ (
);

FILL FILL_1__13369_ (
);

FILL FILL_4__14703_ (
);

FILL FILL_3__8893_ (
);

FILL FILL_3__8473_ (
);

OAI21X1 _12647_ (
    .A(_3476_),
    .B(vdd),
    .C(_3477_),
    .Y(_3425_[26])
);

NAND3X1 _12227_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3209_)
);

FILL FILL_5__8399_ (
);

FILL FILL_1__14730_ (
);

FILL FILL_1__14310_ (
);

FILL FILL_0__13723_ (
);

FILL FILL_0__13303_ (
);

FILL FILL_3__16168_ (
);

FILL FILL_2__6890_ (
);

FILL FILL_5__10689_ (
);

FILL FILL_5__9760_ (
);

FILL FILL_5__10269_ (
);

FILL FILL_5__9340_ (
);

FILL FILL_0_BUFX2_insert1040 (
);

FILL FILL_0_BUFX2_insert1041 (
);

FILL FILL_0_BUFX2_insert1042 (
);

FILL FILL_0_BUFX2_insert1043 (
);

FILL FILL_0__16195_ (
);

FILL FILL_0_BUFX2_insert1044 (
);

AOI22X1 _16060_ (
    .A(\datapath_1.regfile_1.regOut[1] [25]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_6515_)
);

FILL FILL_0_BUFX2_insert1045 (
);

FILL FILL_2__10296_ (
);

FILL FILL_0_BUFX2_insert1046 (
);

FILL FILL_0_BUFX2_insert1047 (
);

FILL FILL_0_BUFX2_insert1048 (
);

FILL FILL_1__9752_ (
);

FILL FILL_0_BUFX2_insert1049 (
);

FILL FILL_5__11630_ (
);

FILL FILL_5__11210_ (
);

FILL FILL_4__15908_ (
);

FILL FILL_3__9678_ (
);

FILL FILL_2__16102_ (
);

FILL FILL_3_BUFX2_insert940 (
);

FILL FILL_3__9258_ (
);

FILL FILL_3_BUFX2_insert941 (
);

FILL FILL_4__10623_ (
);

FILL FILL_3_BUFX2_insert942 (
);

FILL FILL_3_BUFX2_insert943 (
);

FILL FILL_3_BUFX2_insert944 (
);

FILL FILL_1__15935_ (
);

FILL FILL_3_BUFX2_insert945 (
);

FILL FILL_1__15515_ (
);

FILL FILL_3_BUFX2_insert946 (
);

FILL FILL_3_BUFX2_insert947 (
);

FILL FILL_3_BUFX2_insert948 (
);

FILL SFILL38040x77050 (
);

FILL FILL_3_BUFX2_insert949 (
);

FILL FILL_1__10650_ (
);

FILL FILL_1__10230_ (
);

FILL FILL_4__13095_ (
);

FILL FILL_0__14928_ (
);

FILL FILL_0__14508_ (
);

FILL FILL_2__7675_ (
);

FILL FILL_3__12088_ (
);

FILL SFILL3560x52050 (
);

FILL FILL_5__12835_ (
);

FILL FILL_5__12415_ (
);

FILL FILL_4__8962_ (
);

FILL FILL_4__8122_ (
);

FILL FILL_4__11828_ (
);

FILL FILL_2__12862_ (
);

FILL FILL_4__11408_ (
);

FILL FILL_2__12442_ (
);

FILL FILL_2__12022_ (
);

FILL FILL_6__8888_ (
);

DFFSR _9187_ (
    .Q(\datapath_1.regfile_1.regOut[18] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_1108_[13])
);

FILL FILL112200x47050 (
);

FILL FILL_1__11855_ (
);

FILL FILL_1__11435_ (
);

FILL FILL_1__11015_ (
);

FILL FILL_0__8862_ (
);

FILL FILL_0__8442_ (
);

FILL SFILL24600x43050 (
);

DFFSR _10713_ (
    .Q(\datapath_1.regfile_1.regOut[30] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_1888_[3])
);

FILL FILL_0__10428_ (
);

FILL FILL_0__10008_ (
);

FILL FILL_5__6885_ (
);

FILL FILL_4__15661_ (
);

FILL FILL_4__15241_ (
);

DFFSR _13185_ (
    .Q(\datapath_1.mux_iord.din0 [10]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3685_[10])
);

FILL FILL_2__9401_ (
);

FILL FILL_3__14654_ (
);

FILL FILL_3__14234_ (
);

FILL SFILL28920x51050 (
);

FILL FILL_1__6877_ (
);

FILL FILL_4__9747_ (
);

FILL FILL_2__13647_ (
);

FILL FILL_2__13227_ (
);

FILL FILL_0__14681_ (
);

FILL FILL_0__14261_ (
);

FILL SFILL83880x10050 (
);

FILL FILL_3__7744_ (
);

FILL FILL_0__9647_ (
);

FILL FILL_0__9227_ (
);

FILL FILL_3__7324_ (
);

NAND2X1 _11918_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[10]),
    .Y(_2987_)
);

FILL SFILL3480x14050 (
);

FILL FILL_4__16026_ (
);

FILL FILL_4__11581_ (
);

FILL FILL_4__11161_ (
);

FILL FILL_3__15859_ (
);

FILL FILL_3__15439_ (
);

FILL FILL_3__15019_ (
);

FILL FILL_1__16053_ (
);

FILL FILL_3__10994_ (
);

FILL FILL_3__10574_ (
);

FILL FILL_5__8611_ (
);

FILL FILL_3__10154_ (
);

FILL FILL_0__15886_ (
);

FILL SFILL28440x44050 (
);

FILL FILL_6_BUFX2_insert454 (
);

INVX1 _15751_ (
    .A(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_6214_)
);

FILL FILL_0__15466_ (
);

OAI22X1 _15331_ (
    .A(_5804_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf1),
    .D(_4260_),
    .Y(_5805_)
);

FILL FILL_0__15046_ (
);

FILL FILL_0__10181_ (
);

FILL FILL_6_BUFX2_insert459 (
);

FILL FILL_5__10901_ (
);

FILL FILL_1__8603_ (
);

FILL FILL_6__14380_ (
);

FILL SFILL89480x38050 (
);

FILL FILL_3__8529_ (
);

FILL FILL_3__8109_ (
);

FILL FILL_5__13793_ (
);

FILL FILL_5__13373_ (
);

INVX1 _7673_ (
    .A(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_394_)
);

OAI21X1 _7253_ (
    .A(_194_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .C(_195_),
    .Y(_133_[31])
);

FILL SFILL115160x5050 (
);

FILL FILL_4__12786_ (
);

FILL FILL_4__9080_ (
);

FILL SFILL28840x13050 (
);

FILL FILL_4__12366_ (
);

FILL SFILL94360x80050 (
);

FILL FILL_2__6946_ (
);

FILL FILL_3__11779_ (
);

FILL FILL_3__11359_ (
);

FILL FILL_1__12393_ (
);

NOR2X1 _16116_ (
    .A(_6569_),
    .B(_6567_),
    .Y(_6570_)
);

FILL FILL_0__11386_ (
);

AND2X2 _11671_ (
    .A(_2758_),
    .B(_2752_),
    .Y(_2773_)
);

NOR2X1 _11251_ (
    .A(_2366_),
    .B(_2369_),
    .Y(_2370_)
);

FILL FILL_1__9808_ (
);

FILL FILL_3__12720_ (
);

FILL FILL_3__12300_ (
);

FILL FILL_4__7813_ (
);

FILL FILL_5__14998_ (
);

FILL FILL_5__14578_ (
);

FILL FILL_2__11713_ (
);

FILL FILL_5__14158_ (
);

FILL FILL_3__15192_ (
);

OAI21X1 _8878_ (
    .A(_1013_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .C(_1014_),
    .Y(_978_[18])
);

OAI21X1 _8458_ (
    .A(_794_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .C(_795_),
    .Y(_783_[6])
);

DFFSR _8038_ (
    .Q(\datapath_1.regfile_1.regOut[9] [16]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_523_[16])
);

FILL FILL_1__10706_ (
);

FILL SFILL18840x56050 (
);

FILL FILL_2__14185_ (
);

FILL FILL_0__7713_ (
);

FILL FILL_1__13598_ (
);

FILL FILL_4__14932_ (
);

FILL FILL_4__14512_ (
);

OAI21X1 _12876_ (
    .A(_3588_),
    .B(vdd),
    .C(_3589_),
    .Y(_3555_[17])
);

OAI21X1 _12456_ (
    .A(_3369_),
    .B(vdd),
    .C(_3370_),
    .Y(_3360_[5])
);

NAND3X1 _12036_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [12]),
    .C(_3034__bF$buf3),
    .Y(_3073_)
);

FILL FILL_3__13925_ (
);

FILL FILL_3__13505_ (
);

FILL FILL_5_BUFX2_insert470 (
);

FILL FILL_5_BUFX2_insert471 (
);

FILL FILL_2__12918_ (
);

FILL FILL_5_BUFX2_insert472 (
);

FILL FILL_0__13952_ (
);

FILL FILL_5_BUFX2_insert473 (
);

FILL FILL_0__13532_ (
);

FILL FILL_3__16397_ (
);

FILL FILL_0__13112_ (
);

FILL FILL_5_BUFX2_insert474 (
);

FILL FILL_5_BUFX2_insert475 (
);

FILL FILL_5__10498_ (
);

FILL FILL_5_BUFX2_insert476 (
);

FILL FILL_5_BUFX2_insert477 (
);

FILL FILL_5_BUFX2_insert478 (
);

FILL FILL_5_BUFX2_insert479 (
);

FILL FILL_5__16304_ (
);

FILL SFILL18840x11050 (
);

FILL FILL_1__9981_ (
);

FILL FILL_1__9141_ (
);

FILL FILL_4__15717_ (
);

FILL FILL_2__16331_ (
);

FILL FILL_3__9487_ (
);

FILL FILL_4__10432_ (
);

FILL FILL_4__10012_ (
);

FILL FILL_6__7492_ (
);

FILL FILL_1__15744_ (
);

FILL FILL_1__15324_ (
);

FILL FILL_0__14737_ (
);

INVX1 _14602_ (
    .A(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_5090_)
);

FILL FILL_0__14317_ (
);

FILL FILL_2__7484_ (
);

FILL FILL_2__7064_ (
);

FILL FILL_5__12644_ (
);

FILL FILL_5__12224_ (
);

INVX1 _6944_ (
    .A(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_30_)
);

FILL SFILL69080x65050 (
);

FILL FILL_4__8771_ (
);

FILL FILL_4__8351_ (
);

FILL FILL_4__11637_ (
);

FILL FILL_4__11217_ (
);

FILL FILL_2__12251_ (
);

FILL FILL_6__8697_ (
);

FILL FILL_1__16109_ (
);

FILL FILL_1__11664_ (
);

FILL FILL_1__11244_ (
);

INVX1 _15807_ (
    .A(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_6269_)
);

NOR2X1 _10942_ (
    .A(_2075_),
    .B(_2074_),
    .Y(_2076_)
);

FILL FILL_0__8251_ (
);

FILL FILL_2__8269_ (
);

FILL FILL_0__10657_ (
);

INVX1 _10522_ (
    .A(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_1846_)
);

FILL FILL_0__10237_ (
);

INVX1 _10102_ (
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_1691_)
);

FILL FILL_6__14856_ (
);

FILL FILL_4__15890_ (
);

FILL FILL_6__14436_ (
);

FILL FILL_4__15470_ (
);

FILL FILL_4__15050_ (
);

FILL FILL_5__13849_ (
);

FILL FILL_5__13429_ (
);

FILL FILL_3__14883_ (
);

FILL FILL_2__9630_ (
);

FILL FILL_3__14463_ (
);

FILL FILL_5__13009_ (
);

FILL FILL_2__9210_ (
);

FILL FILL_3__14043_ (
);

OAI21X1 _7729_ (
    .A(_430_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_431_),
    .Y(_393_[19])
);

OAI21X1 _7309_ (
    .A(_211_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_212_),
    .Y(_198_[7])
);

FILL FILL_4__9976_ (
);

FILL FILL_4__9556_ (
);

FILL FILL_4__9136_ (
);

FILL FILL_2__13876_ (
);

FILL FILL_2__13456_ (
);

FILL FILL_0__14490_ (
);

FILL FILL_2__13036_ (
);

FILL FILL_0__14070_ (
);

FILL SFILL84920x50 (
);

FILL FILL_1__12869_ (
);

FILL FILL_1__12449_ (
);

FILL FILL_1__12029_ (
);

FILL FILL_3__7973_ (
);

FILL FILL_0__9876_ (
);

FILL FILL_3__7553_ (
);

FILL FILL_0__9036_ (
);

NAND3X1 _11727_ (
    .A(_2822_),
    .B(_2824_),
    .C(_2819_),
    .Y(\datapath_1.ALUResult [10])
);

INVX1 _11307_ (
    .A(_2425_),
    .Y(_2426_)
);

FILL FILL_5__7479_ (
);

FILL FILL_1__13810_ (
);

FILL FILL_4__16255_ (
);

FILL FILL_5__7059_ (
);

FILL FILL_6__10776_ (
);

INVX1 _14199_ (
    .A(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_4696_)
);

FILL FILL_4__11390_ (
);

FILL FILL_3__15668_ (
);

FILL FILL_3__15248_ (
);

FILL FILL_1__16282_ (
);

FILL FILL_5__8840_ (
);

FILL FILL_3__10383_ (
);

FILL FILL_5__8000_ (
);

FILL SFILL59080x63050 (
);

OAI22X1 _15980_ (
    .A(_5530__bF$buf2),
    .B(_6436_),
    .C(_5552__bF$buf0),
    .D(_5062_),
    .Y(_6437_)
);

FILL FILL_0__15695_ (
);

NAND2X1 _15560_ (
    .A(_6023_),
    .B(_6027_),
    .Y(_6028_)
);

FILL FILL_0__15275_ (
);

INVX1 _15140_ (
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_5618_)
);

FILL SFILL38920x48050 (
);

FILL FILL_1__8832_ (
);

FILL FILL_2__15602_ (
);

FILL FILL_3__8758_ (
);

FILL FILL_3__8338_ (
);

FILL SFILL3640x40050 (
);

OAI21X1 _7482_ (
    .A(_306_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_307_),
    .Y(_263_[22])
);

OAI21X1 _7062_ (
    .A(_87_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_88_),
    .Y(_68_[10])
);

FILL FILL_4__12595_ (
);

FILL FILL_4__12175_ (
);

FILL FILL_5__9625_ (
);

FILL FILL_3__11588_ (
);

FILL FILL_3__11168_ (
);

INVX1 _16345_ (
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_6784_)
);

FILL FILL_0__11195_ (
);

NAND3X1 _11480_ (
    .A(_2288_),
    .B(_2309_),
    .C(_2578_),
    .Y(_2594_)
);

FILL FILL_5__11915_ (
);

NOR2X1 _11060_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2179_)
);

FILL FILL_1__9617_ (
);

FILL SFILL104440x64050 (
);

FILL FILL_4__7622_ (
);

FILL FILL_4__10908_ (
);

FILL FILL_4__7202_ (
);

FILL FILL_2__11942_ (
);

FILL FILL_5__14387_ (
);

FILL FILL_2__11522_ (
);

FILL FILL_6__7968_ (
);

FILL FILL_2__11102_ (
);

DFFSR _8687_ (
    .Q(\datapath_1.regfile_1.regOut[14] [25]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_848_[25])
);

NAND2X1 _8267_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_709_)
);

FILL SFILL44680x3050 (
);

FILL FILL_1__10935_ (
);

FILL FILL_1__10515_ (
);

FILL FILL_0__7942_ (
);

BUFX2 BUFX2_insert290 (
    .A(_5539_),
    .Y(_5539__bF$buf0)
);

FILL FILL_0__7102_ (
);

BUFX2 BUFX2_insert291 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf7 )
);

BUFX2 BUFX2_insert292 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf6 )
);

BUFX2 BUFX2_insert293 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf5 )
);

BUFX2 BUFX2_insert294 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf4 )
);

BUFX2 BUFX2_insert295 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf3 )
);

FILL FILL_4__14741_ (
);

BUFX2 BUFX2_insert296 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf2 )
);

FILL FILL_4__14321_ (
);

FILL SFILL69240x9050 (
);

BUFX2 BUFX2_insert297 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf1 )
);

BUFX2 BUFX2_insert298 (
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf0 )
);

FILL SFILL43960x5050 (
);

DFFSR _12685_ (
    .Q(\datapath_1.Data [22]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3425_[22])
);

BUFX2 BUFX2_insert299 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf4 )
);

FILL FILL_3__8091_ (
);

FILL SFILL49080x61050 (
);

AOI22X1 _12265_ (
    .A(_2_[12]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [12]),
    .Y(_3238_)
);

FILL FILL_2__8901_ (
);

FILL FILL_3__13734_ (
);

FILL FILL_3__13314_ (
);

FILL SFILL28920x46050 (
);

FILL FILL_4__8827_ (
);

FILL FILL_2__12727_ (
);

FILL FILL_0__13761_ (
);

FILL FILL_2__12307_ (
);

FILL FILL_0__13341_ (
);

FILL FILL_2__15199_ (
);

FILL FILL_0__8727_ (
);

FILL FILL_5__16113_ (
);

FILL FILL_1__9790_ (
);

FILL FILL_1__9370_ (
);

FILL FILL_4__15946_ (
);

FILL FILL_4__15526_ (
);

FILL FILL_4__15106_ (
);

FILL FILL_2__16140_ (
);

FILL SFILL73960x41050 (
);

FILL SFILL89560x26050 (
);

FILL FILL_3__9296_ (
);

FILL FILL_4__10661_ (
);

FILL FILL_4__10241_ (
);

FILL FILL_3__14939_ (
);

FILL FILL_1__15973_ (
);

FILL FILL_3__14519_ (
);

FILL FILL_1__15553_ (
);

FILL FILL_1__15133_ (
);

FILL FILL_0__14966_ (
);

NOR2X1 _14831_ (
    .A(_5311_),
    .B(_5314_),
    .Y(_5315_)
);

FILL FILL_0__14546_ (
);

FILL FILL_0__14126_ (
);

NOR2X1 _14411_ (
    .A(_4899_),
    .B(_4902_),
    .Y(_4903_)
);

FILL FILL_2__7293_ (
);

FILL FILL_3__7609_ (
);

FILL FILL_5__12873_ (
);

FILL SFILL28040x25050 (
);

FILL FILL_5__12453_ (
);

FILL FILL_5__12033_ (
);

FILL FILL_4__8580_ (
);

FILL FILL_4__11866_ (
);

FILL SFILL94360x75050 (
);

FILL FILL_4__11446_ (
);

FILL FILL_2__12480_ (
);

FILL FILL_4__11026_ (
);

FILL FILL_2__12060_ (
);

FILL FILL_1__16338_ (
);

FILL FILL_1__11893_ (
);

FILL FILL_3__10439_ (
);

FILL FILL_3__10019_ (
);

FILL FILL_1__11473_ (
);

FILL FILL_1__11053_ (
);

AOI22X1 _15616_ (
    .A(\datapath_1.regfile_1.regOut[3] [14]),
    .B(_5494_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_6082_)
);

FILL SFILL58200x57050 (
);

FILL FILL_0__8480_ (
);

FILL FILL_0__10886_ (
);

FILL FILL_2__8498_ (
);

FILL SFILL79160x55050 (
);

FILL FILL_2__8078_ (
);

INVX1 _10751_ (
    .A(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_1958_)
);

FILL FILL_0__8060_ (
);

FILL FILL_0__10046_ (
);

DFFSR _10331_ (
    .Q(\datapath_1.regfile_1.regOut[27] [5]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_1693_[5])
);

FILL FILL_3__11800_ (
);

FILL FILL_5__13658_ (
);

FILL FILL_5__13238_ (
);

FILL FILL_3__14692_ (
);

FILL FILL_3__14272_ (
);

OAI21X1 _7958_ (
    .A(_542_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .C(_543_),
    .Y(_523_[10])
);

DFFSR _7538_ (
    .Q(\datapath_1.regfile_1.regOut[5] [28]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_263_[28])
);

NAND2X1 _7118_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_126_)
);

FILL FILL_4__9785_ (
);

FILL FILL_4__9365_ (
);

FILL FILL_2__13685_ (
);

FILL FILL_2__13265_ (
);

FILL FILL_1__12258_ (
);

FILL FILL_0__9685_ (
);

INVX1 _11956_ (
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3012_)
);

FILL FILL_0__9265_ (
);

FILL FILL_3__7362_ (
);

AOI21X1 _11536_ (
    .A(_2407_),
    .B(_2565_),
    .C(_2421_),
    .Y(_2647_)
);

NOR2X1 _11116_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .B(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2235_)
);

FILL FILL_5__7288_ (
);

FILL SFILL79160x10050 (
);

FILL FILL_4__16064_ (
);

FILL FILL_6__10165_ (
);

FILL SFILL39320x3050 (
);

FILL FILL111720x66050 (
);

FILL FILL_3__15897_ (
);

FILL FILL_0__12612_ (
);

FILL FILL_3__15477_ (
);

FILL FILL_3__15057_ (
);

FILL FILL_1__16091_ (
);

FILL FILL_3__10192_ (
);

FILL FILL_6_BUFX2_insert833 (
);

FILL FILL_0__15084_ (
);

FILL FILL_5__15804_ (
);

FILL SFILL53960x82050 (
);

FILL SFILL84360x73050 (
);

FILL FILL_6_BUFX2_insert838 (
);

FILL FILL_1__8641_ (
);

FILL FILL_1__8221_ (
);

FILL FILL_2__15831_ (
);

FILL FILL_2__15411_ (
);

FILL FILL_3__8987_ (
);

FILL FILL_3__8567_ (
);

FILL FILL_3__8147_ (
);

FILL FILL_1__14824_ (
);

FILL FILL_1__14404_ (
);

OAI21X1 _7291_ (
    .A(_199_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .C(_200_),
    .Y(_198_[1])
);

FILL FILL_0__13817_ (
);

FILL FILL_2__6984_ (
);

FILL FILL111720x21050 (
);

FILL FILL_5__9854_ (
);

FILL FILL_3__11397_ (
);

FILL FILL_5__9014_ (
);

FILL FILL_0__16289_ (
);

OAI22X1 _16154_ (
    .A(_5233_),
    .B(_5539__bF$buf0),
    .C(_5526__bF$buf4),
    .D(_5269_),
    .Y(_6607_)
);

FILL FILL_1__9846_ (
);

FILL FILL_5__11724_ (
);

FILL FILL_1__9426_ (
);

FILL FILL_5__11304_ (
);

FILL FILL_1__9006_ (
);

FILL FILL_4__7851_ (
);

FILL FILL_4__7431_ (
);

FILL FILL_2__11751_ (
);

FILL FILL_5__14196_ (
);

FILL FILL_2__11331_ (
);

NAND2X1 _8496_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_821_)
);

FILL FILL_1__15609_ (
);

NAND2X1 _8076_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_602_)
);

FILL FILL_1__10744_ (
);

FILL FILL_1__10324_ (
);

FILL FILL_0__7751_ (
);

FILL FILL_2__7349_ (
);

FILL FILL_0__7331_ (
);

FILL SFILL114520x54050 (
);

FILL FILL_4__14970_ (
);

FILL FILL_4__14550_ (
);

FILL FILL_4__14130_ (
);

FILL SFILL3720x73050 (
);

NAND2X1 _12494_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [18]),
    .Y(_3396_)
);

NAND3X1 _12074_ (
    .A(_3099_),
    .B(_3100_),
    .C(_3101_),
    .Y(\datapath_1.mux_pcsrc.dout [21])
);

FILL FILL_5__12509_ (
);

FILL FILL_3__13963_ (
);

FILL FILL_2__8710_ (
);

FILL FILL_3__13543_ (
);

FILL FILL_3__13123_ (
);

FILL FILL_4__8636_ (
);

FILL FILL_4__8216_ (
);

FILL FILL_5_BUFX2_insert850 (
);

FILL SFILL69080x15050 (
);

FILL FILL_5_BUFX2_insert851 (
);

FILL FILL_2__12956_ (
);

FILL FILL_5_BUFX2_insert852 (
);

FILL FILL_0__13990_ (
);

FILL FILL_5_BUFX2_insert853 (
);

FILL FILL_2__12116_ (
);

FILL FILL_0__13570_ (
);

FILL FILL_5_BUFX2_insert854 (
);

FILL FILL_0__13150_ (
);

FILL FILL_5_BUFX2_insert855 (
);

FILL FILL_5_BUFX2_insert856 (
);

FILL FILL_5_BUFX2_insert857 (
);

FILL FILL_1__11949_ (
);

FILL FILL_5_BUFX2_insert858 (
);

FILL FILL_5_BUFX2_insert859 (
);

FILL FILL_1__11529_ (
);

FILL FILL_1__11109_ (
);

FILL FILL_5__16342_ (
);

FILL FILL_0__8956_ (
);

OAI21X1 _10807_ (
    .A(_1994_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1995_),
    .Y(_1953_[21])
);

FILL FILL_0__8116_ (
);

FILL FILL_6__9503_ (
);

FILL FILL_5__6979_ (
);

FILL FILL_4__15755_ (
);

FILL FILL_4__15335_ (
);

FILL FILL_4__10890_ (
);

INVX1 _13699_ (
    .A(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_4206_)
);

OR2X2 _13279_ (
    .A(_3796_),
    .B(_3818_),
    .Y(_3819_)
);

FILL FILL_2__9915_ (
);

FILL FILL_4__10050_ (
);

FILL FILL_3__14748_ (
);

FILL FILL_1__15782_ (
);

FILL FILL_3__14328_ (
);

FILL FILL_1__15362_ (
);

FILL FILL_5__7500_ (
);

FILL SFILL59080x58050 (
);

FILL FILL_0__14775_ (
);

OAI22X1 _14640_ (
    .A(_3978_),
    .B(_5126_),
    .C(_3977__bF$buf4),
    .D(_5127_),
    .Y(_5128_)
);

FILL FILL_0__14355_ (
);

OAI22X1 _14220_ (
    .A(_4714_),
    .B(_3910_),
    .C(_3935__bF$buf4),
    .D(_4715_),
    .Y(_4716_)
);

FILL FILL_3__7838_ (
);

FILL FILL_3__7418_ (
);

FILL SFILL49480x5050 (
);

FILL SFILL3640x35050 (
);

FILL FILL_5__12262_ (
);

OAI21X1 _6982_ (
    .A(_54_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_55_),
    .Y(_3_[26])
);

FILL FILL_2_BUFX2_insert980 (
);

FILL FILL_2_BUFX2_insert981 (
);

FILL SFILL104520x52050 (
);

FILL FILL_2_BUFX2_insert982 (
);

FILL SFILL43880x42050 (
);

FILL FILL_2_BUFX2_insert983 (
);

FILL FILL_2_BUFX2_insert984 (
);

FILL FILL_4__11675_ (
);

FILL FILL_2_BUFX2_insert985 (
);

FILL FILL_4__11255_ (
);

FILL FILL_2_BUFX2_insert986 (
);

FILL FILL_2_BUFX2_insert987 (
);

FILL SFILL48840x2050 (
);

FILL FILL_2_BUFX2_insert988 (
);

FILL FILL_2_BUFX2_insert989 (
);

FILL FILL_1__16147_ (
);

FILL FILL_5__8705_ (
);

FILL FILL_3__10668_ (
);

FILL SFILL49080x4050 (
);

FILL FILL_3__10248_ (
);

FILL SFILL59000x56050 (
);

FILL FILL_1__11282_ (
);

OAI22X1 _15845_ (
    .A(_5534__bF$buf1),
    .B(_4888_),
    .C(_5532__bF$buf3),
    .D(_6305_),
    .Y(_6306_)
);

NOR2X1 _15425_ (
    .A(_5894_),
    .B(_5895_),
    .Y(_5896_)
);

NAND3X1 _15005_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5462_),
    .C(_5461_),
    .Y(_5485_)
);

FILL SFILL59080x13050 (
);

OAI21X1 _10980_ (
    .A(_2103_),
    .B(vdd),
    .C(_2104_),
    .Y(_2098_[2])
);

FILL FILL_0__10695_ (
);

FILL FILL_0__10275_ (
);

OAI21X1 _10560_ (
    .A(_1870_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .C(_1871_),
    .Y(_1823_[24])
);

OAI21X1 _10140_ (
    .A(_1651_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1652_),
    .Y(_1628_[12])
);

FILL SFILL104440x59050 (
);

FILL FILL_5__13887_ (
);

FILL FILL_5__13467_ (
);

DFFSR _7767_ (
    .Q(\datapath_1.regfile_1.regOut[7] [1]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_393_[1])
);

FILL FILL_3__14081_ (
);

NAND2X1 _7347_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_238_)
);

FILL FILL_4__9594_ (
);

FILL FILL_2__13494_ (
);

FILL FILL_1__12487_ (
);

FILL FILL_1__12067_ (
);

FILL FILL_4__13821_ (
);

FILL FILL_4__13401_ (
);

FILL SFILL28120x58050 (
);

FILL FILL_3__7591_ (
);

FILL FILL_0__9494_ (
);

FILL SFILL49080x56050 (
);

FILL FILL_3__7171_ (
);

AOI22X1 _11765_ (
    .A(_2136_),
    .B(_2481__bF$buf0),
    .C(_2620_),
    .D(_2373_),
    .Y(_2860_)
);

OAI21X1 _11345_ (
    .A(_2461_),
    .B(_2116_),
    .C(_2462__bF$buf2),
    .Y(_2463_)
);

FILL FILL_6__15679_ (
);

FILL FILL_5__7097_ (
);

FILL FILL_4__16293_ (
);

FILL FILL_2__11807_ (
);

FILL FILL_0__12841_ (
);

FILL FILL_0__12421_ (
);

FILL FILL_3__15286_ (
);

FILL FILL_0__12001_ (
);

FILL FILL_1__7089_ (
);

FILL FILL_2__14699_ (
);

FILL FILL_2__14279_ (
);

FILL FILL_5__15613_ (
);

FILL FILL_0__7807_ (
);

NAND2X1 _9913_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1542_)
);

FILL FILL_1__8870_ (
);

FILL FILL_1__8450_ (
);

FILL FILL_4__14606_ (
);

FILL FILL_2__15640_ (
);

FILL FILL_2__15220_ (
);

FILL SFILL49000x54050 (
);

FILL FILL_3__8376_ (
);

FILL FILL_1__14633_ (
);

FILL SFILL49080x11050 (
);

FILL FILL_1__14213_ (
);

FILL FILL_6__11599_ (
);

FILL SFILL94440x63050 (
);

FILL FILL_0__13626_ (
);

INVX1 _13911_ (
    .A(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_4414_)
);

FILL FILL_5__9663_ (
);

FILL FILL_5__9243_ (
);

FILL FILL_6__12960_ (
);

OAI21X1 _16383_ (
    .A(_6808_),
    .B(gnd),
    .C(_6809_),
    .Y(_6769_[20])
);

FILL FILL_0__16098_ (
);

FILL SFILL23880x83050 (
);

FILL FILL_5__11953_ (
);

FILL FILL_1__9655_ (
);

FILL FILL_5__11533_ (
);

FILL FILL_5__11113_ (
);

FILL FILL_1__9235_ (
);

FILL FILL_2__16005_ (
);

FILL FILL_4__10946_ (
);

FILL FILL_4__7240_ (
);

FILL FILL_2__11980_ (
);

FILL FILL_4__10526_ (
);

FILL FILL_2__11560_ (
);

FILL FILL_4__10106_ (
);

FILL FILL_2__11140_ (
);

FILL FILL_6__7586_ (
);

FILL FILL_1__15838_ (
);

FILL FILL_1__15418_ (
);

FILL FILL_1__10973_ (
);

FILL FILL_1__10553_ (
);

FILL FILL_1__10133_ (
);

FILL FILL_2__7998_ (
);

FILL FILL_0__7980_ (
);

BUFX2 BUFX2_insert670 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf0 )
);

FILL FILL_0__7560_ (
);

FILL FILL_2__7578_ (
);

BUFX2 BUFX2_insert671 (
    .A(_5544_),
    .Y(_5544__bF$buf3)
);

FILL FILL_2__7158_ (
);

BUFX2 BUFX2_insert672 (
    .A(_5544_),
    .Y(_5544__bF$buf2)
);

BUFX2 BUFX2_insert673 (
    .A(_5544_),
    .Y(_5544__bF$buf1)
);

BUFX2 BUFX2_insert674 (
    .A(_5544_),
    .Y(_5544__bF$buf0)
);

BUFX2 BUFX2_insert675 (
    .A(_4051_),
    .Y(_4051__bF$buf3)
);

FILL SFILL18840x1050 (
);

BUFX2 BUFX2_insert676 (
    .A(_4051_),
    .Y(_4051__bF$buf2)
);

FILL SFILL23800x81050 (
);

BUFX2 BUFX2_insert677 (
    .A(_4051_),
    .Y(_4051__bF$buf1)
);

BUFX2 BUFX2_insert678 (
    .A(_4051_),
    .Y(_4051__bF$buf0)
);

BUFX2 BUFX2_insert679 (
    .A(_5485_),
    .Y(_5485__bF$buf4)
);

FILL SFILL18520x25050 (
);

FILL SFILL18760x6050 (
);

FILL FILL_5__12738_ (
);

FILL FILL_3__13772_ (
);

FILL FILL_5__12318_ (
);

FILL FILL_3__13352_ (
);

FILL FILL_4__8865_ (
);

FILL SFILL8840x80050 (
);

FILL FILL_4__8445_ (
);

FILL FILL_2__12765_ (
);

FILL FILL_2__12345_ (
);

FILL SFILL79560x19050 (
);

FILL SFILL39000x52050 (
);

FILL SFILL94360x25050 (
);

FILL FILL_1__11758_ (
);

FILL FILL_1__11338_ (
);

FILL FILL_0__8765_ (
);

FILL FILL_3__6862_ (
);

FILL FILL_5__16151_ (
);

FILL FILL_0__8345_ (
);

FILL SFILL84440x61050 (
);

OAI21X1 _10616_ (
    .A(_1951_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1952_),
    .Y(_1888_[0])
);

FILL FILL_4__15984_ (
);

FILL FILL_4__15564_ (
);

FILL FILL_4__15144_ (
);

INVX1 _13088_ (
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_3690_)
);

FILL FILL_3__14977_ (
);

FILL FILL_2__9724_ (
);

FILL FILL_3__14557_ (
);

FILL FILL_3__14137_ (
);

FILL FILL_1__15591_ (
);

FILL FILL_1__15171_ (
);

FILL FILL_0__14584_ (
);

FILL FILL_0__14164_ (
);

FILL SFILL53960x77050 (
);

FILL FILL_1__7721_ (
);

FILL FILL_1__7301_ (
);

FILL FILL_2__14911_ (
);

FILL FILL_3__7227_ (
);

FILL FILL_5__12491_ (
);

FILL FILL_5__12071_ (
);

FILL FILL_1__13904_ (
);

FILL FILL_4__16349_ (
);

FILL FILL_4__11484_ (
);

FILL FILL_4__11064_ (
);

FILL FILL_1__16376_ (
);

FILL FILL_3__10897_ (
);

FILL FILL_5__8514_ (
);

FILL FILL_3__10057_ (
);

FILL FILL_1__11091_ (
);

FILL FILL_0__15789_ (
);

NOR2X1 _15654_ (
    .A(_6118_),
    .B(_5549__bF$buf2),
    .Y(_6119_)
);

FILL FILL_0__15369_ (
);

AOI21X1 _15234_ (
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .B(_5567_),
    .C(_5709_),
    .Y(_5710_)
);

FILL SFILL114600x42050 (
);

FILL FILL_5__10804_ (
);

FILL SFILL53960x32050 (
);

FILL FILL_1__8506_ (
);

FILL SFILL84360x23050 (
);

FILL FILL_6__14283_ (
);

FILL FILL_4__6931_ (
);

FILL FILL_0__16310_ (
);

FILL FILL_2__10831_ (
);

FILL FILL_5__13696_ (
);

FILL FILL_5__13276_ (
);

FILL FILL_2__10411_ (
);

NAND2X1 _7996_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_569_)
);

NAND2X1 _7576_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_350_)
);

DFFSR _7156_ (
    .Q(\datapath_1.regfile_1.regOut[2] [30]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_68_[30])
);

FILL FILL_4__12269_ (
);

FILL FILL_2__6849_ (
);

FILL FILL_5__9719_ (
);

FILL SFILL53880x39050 (
);

FILL FILL_1__12296_ (
);

FILL FILL_4__13630_ (
);

DFFSR _16439_ (
    .Q(\datapath_1.regfile_1.regOut[0] [22]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_6769_[22])
);

FILL SFILL3720x68050 (
);

FILL FILL_4__13210_ (
);

NOR2X1 _16019_ (
    .A(_6472_),
    .B(_6474_),
    .Y(_6475_)
);

NAND3X1 _11994_ (
    .A(_3039_),
    .B(_3040_),
    .C(_3041_),
    .Y(\datapath_1.mux_pcsrc.dout [1])
);

OAI21X1 _11574_ (
    .A(_2670_),
    .B(_2344__bF$buf2),
    .C(_2681_),
    .Y(_2682_)
);

FILL FILL_0__11289_ (
);

NOR2X1 _11154_ (
    .A(\datapath_1.alu_1.ALUInB [19]),
    .B(_2242_),
    .Y(_2273_)
);

FILL SFILL43960x75050 (
);

FILL FILL_3__12623_ (
);

FILL FILL_3__12203_ (
);

FILL FILL_4__7716_ (
);

FILL FILL_2__11616_ (
);

FILL FILL_0__12650_ (
);

FILL FILL_0__12230_ (
);

FILL FILL_3__15095_ (
);

FILL FILL_2__14088_ (
);

FILL FILL_5__15842_ (
);

FILL FILL_5__15422_ (
);

FILL FILL_0__7616_ (
);

FILL FILL_5__15002_ (
);

NAND2X1 _9722_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1435_)
);

DFFSR _9302_ (
    .Q(\datapath_1.regfile_1.regOut[19] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1173_[0])
);

FILL FILL_4__14835_ (
);

FILL FILL_4__14415_ (
);

INVX1 _12779_ (
    .A(\control_1.op [2]),
    .Y(_3545_)
);

FILL FILL_3__8185_ (
);

NAND2X1 _12359_ (
    .A(MemToReg_bF$buf6),
    .B(\datapath_1.Data [5]),
    .Y(_3305_)
);

FILL SFILL3720x23050 (
);

FILL FILL_3__13828_ (
);

FILL FILL_1__14862_ (
);

FILL FILL_3__13408_ (
);

FILL FILL_1__14442_ (
);

FILL FILL_1__14022_ (
);

FILL SFILL104600x40050 (
);

FILL SFILL43960x30050 (
);

FILL FILL_0__13855_ (
);

FILL FILL_0__13435_ (
);

INVX1 _13720_ (
    .A(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_4227_)
);

OR2X2 _13300_ (
    .A(_3796_),
    .B(_3835_),
    .Y(_3836_)
);

FILL FILL_0__13015_ (
);

FILL FILL_5__9892_ (
);

FILL FILL_5__9472_ (
);

OAI21X1 _16192_ (
    .A(_5526__bF$buf2),
    .B(_5313_),
    .C(_6643_),
    .Y(_6644_)
);

FILL FILL_5__16207_ (
);

FILL FILL_3__6918_ (
);

FILL FILL_1__9884_ (
);

FILL FILL_5__11762_ (
);

FILL FILL_1__9464_ (
);

FILL FILL_5__11342_ (
);

FILL FILL_1__9044_ (
);

FILL SFILL104520x47050 (
);

FILL FILL_2__16234_ (
);

FILL FILL_4__10755_ (
);

FILL FILL_1__15647_ (
);

FILL FILL_1__15227_ (
);

FILL FILL_1__10782_ (
);

FILL FILL_1__10362_ (
);

AOI22X1 _14925_ (
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .B(_4154_),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_5407_)
);

INVX1 _14505_ (
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_4995_)
);

FILL FILL112280x41050 (
);

FILL FILL_5__12967_ (
);

FILL FILL_5__12127_ (
);

FILL FILL_3__13581_ (
);

BUFX2 _6847_ (
    .A(_1_[9]),
    .Y(memoryAddress[9])
);

FILL FILL_3__13161_ (
);

FILL FILL_4__8254_ (
);

FILL FILL_2__12994_ (
);

FILL FILL_2__12574_ (
);

FILL FILL_2__12154_ (
);

FILL FILL_1__11987_ (
);

FILL FILL_1__11567_ (
);

FILL FILL_1__11147_ (
);

FILL FILL_4__12901_ (
);

FILL FILL_0__8994_ (
);

FILL FILL_5__16380_ (
);

FILL FILL_0__8574_ (
);

DFFSR _10845_ (
    .Q(\datapath_1.regfile_1.regOut[31] [7]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1953_[7])
);

FILL FILL_6__9121_ (
);

NAND2X1 _10425_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1802_)
);

NAND2X1 _10005_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1583_)
);

FILL FILL_6__14759_ (
);

FILL FILL_4__15793_ (
);

FILL FILL_6__14339_ (
);

FILL FILL_4__15373_ (
);

FILL FILL_2__9533_ (
);

FILL FILL_0__11921_ (
);

FILL FILL_3__14786_ (
);

FILL FILL_2__9113_ (
);

FILL FILL_3__14366_ (
);

FILL FILL_0__11501_ (
);

FILL FILL_6__15700_ (
);

FILL FILL_4__9879_ (
);

FILL FILL_4__9039_ (
);

FILL FILL_2__13779_ (
);

FILL FILL_2__13359_ (
);

FILL FILL_0__14393_ (
);

FILL SFILL33880x35050 (
);

FILL FILL_1__7950_ (
);

FILL FILL_1__7110_ (
);

FILL FILL_2__14720_ (
);

FILL FILL_3__7876_ (
);

FILL FILL_0__9779_ (
);

FILL FILL_2__14300_ (
);

FILL FILL_0__9359_ (
);

FILL FILL_3__7456_ (
);

FILL FILL_3__7036_ (
);

FILL FILL_1__13713_ (
);

FILL FILL_4__16158_ (
);

FILL FILL_6__10259_ (
);

FILL SFILL94440x58050 (
);

FILL FILL_4__11293_ (
);

FILL FILL_0__12706_ (
);

FILL FILL_1__16185_ (
);

FILL SFILL33000x50050 (
);

FILL FILL_5__8743_ (
);

FILL FILL_5__8323_ (
);

FILL FILL_3__10286_ (
);

INVX1 _15883_ (
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_6343_)
);

FILL FILL_6__11620_ (
);

FILL FILL_0__15598_ (
);

FILL FILL_0__15178_ (
);

FILL FILL_6__11200_ (
);

OAI22X1 _15463_ (
    .A(_5530__bF$buf1),
    .B(_4466_),
    .C(_5532__bF$buf2),
    .D(_4448_),
    .Y(_5933_)
);

FILL SFILL23880x78050 (
);

NAND3X1 _15043_ (
    .A(_5459__bF$buf1),
    .B(_5471__bF$buf3),
    .C(_5476_),
    .Y(_5523_)
);

FILL FILL_1__8735_ (
);

FILL FILL_1__8315_ (
);

FILL FILL_2__15925_ (
);

FILL FILL_2__15505_ (
);

FILL FILL_2__10640_ (
);

FILL FILL_5__13085_ (
);

FILL FILL_1__14918_ (
);

DFFSR _7385_ (
    .Q(\datapath_1.regfile_1.regOut[4] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_198_[3])
);

FILL FILL_4__12498_ (
);

FILL FILL_4__12078_ (
);

FILL FILL_3__9602_ (
);

FILL SFILL94440x13050 (
);

FILL FILL_5__9528_ (
);

FILL FILL_5__9108_ (
);

FILL SFILL23800x76050 (
);

OAI22X1 _16248_ (
    .A(_5365_),
    .B(_5545__bF$buf2),
    .C(_5480__bF$buf2),
    .D(_5364_),
    .Y(_6698_)
);

OAI21X1 _11383_ (
    .A(_2136_),
    .B(_2137_),
    .C(_2156_),
    .Y(_2500_)
);

FILL FILL_0__11098_ (
);

FILL FILL_5__11818_ (
);

FILL FILL_3__12852_ (
);

FILL FILL_3__12432_ (
);

FILL FILL_3__12012_ (
);

FILL SFILL8840x75050 (
);

FILL FILL_4__7945_ (
);

FILL FILL_4__7105_ (
);

FILL FILL111800x49050 (
);

FILL FILL_2__11845_ (
);

FILL FILL_2__11425_ (
);

FILL SFILL63960x29050 (
);

FILL FILL_2__11005_ (
);

FILL SFILL23400x62050 (
);

FILL SFILL39000x47050 (
);

FILL FILL_1__10418_ (
);

FILL FILL_5__15651_ (
);

FILL FILL_0__7845_ (
);

FILL FILL_5__15231_ (
);

FILL SFILL84440x56050 (
);

FILL FILL_0__7425_ (
);

DFFSR _9951_ (
    .Q(\datapath_1.regfile_1.regOut[24] [9]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_1498_[9])
);

INVX1 _9531_ (
    .A(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_1348_)
);

INVX1 _9111_ (
    .A(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_1129_)
);

FILL FILL_4__14644_ (
);

FILL FILL_4__14224_ (
);

INVX1 _12588_ (
    .A(\datapath_1.Data [7]),
    .Y(_3438_)
);

OAI21X1 _12168_ (
    .A(_3164_),
    .B(ALUSrcA_bF$buf1),
    .C(_3165_),
    .Y(\datapath_1.alu_1.ALUInA [17])
);

FILL SFILL13880x76050 (
);

FILL FILL_3__13637_ (
);

FILL FILL_3__13217_ (
);

FILL FILL_1__14671_ (
);

FILL FILL_1__14251_ (
);

FILL FILL_0_BUFX2_insert310 (
);

FILL FILL_0_BUFX2_insert311 (
);

FILL FILL_0_BUFX2_insert312 (
);

FILL FILL_0_BUFX2_insert313 (
);

FILL FILL_0__13664_ (
);

FILL FILL_0_BUFX2_insert314 (
);

FILL FILL_0__13244_ (
);

FILL FILL_0_BUFX2_insert315 (
);

FILL FILL_0_BUFX2_insert316 (
);

FILL FILL_0_BUFX2_insert317 (
);

FILL FILL_0_BUFX2_insert318 (
);

FILL FILL_0_BUFX2_insert319 (
);

FILL FILL_5__9281_ (
);

FILL FILL_5__16016_ (
);

FILL FILL_5__11991_ (
);

FILL FILL_5__11571_ (
);

FILL FILL_1__9273_ (
);

FILL FILL_5__11151_ (
);

FILL FILL_4__15849_ (
);

FILL FILL_4__15429_ (
);

FILL FILL_4__15009_ (
);

FILL FILL_2__16043_ (
);

FILL FILL_4__10564_ (
);

FILL SFILL8760x37050 (
);

FILL FILL_4__10144_ (
);

FILL FILL_1__15876_ (
);

FILL FILL_1__15456_ (
);

FILL FILL_1__15036_ (
);

FILL FILL_1__10171_ (
);

FILL FILL_0__14869_ (
);

INVX1 _14734_ (
    .A(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_5220_)
);

FILL FILL_0__14449_ (
);

FILL FILL_0__14029_ (
);

AOI22X1 _14314_ (
    .A(\datapath_1.regfile_1.regOut[6] [18]),
    .B(_4001__bF$buf2),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_4808_)
);

FILL FILL_2__7196_ (
);

FILL SFILL114600x37050 (
);

FILL SFILL53960x27050 (
);

FILL FILL_0__15810_ (
);

FILL FILL_5__12776_ (
);

FILL FILL_5__12356_ (
);

FILL FILL_3__13390_ (
);

FILL SFILL49000x50 (
);

FILL SFILL74440x54050 (
);

FILL FILL_4__8483_ (
);

FILL FILL_4__8063_ (
);

FILL FILL_4__11769_ (
);

FILL FILL_4__11349_ (
);

FILL FILL_2__12383_ (
);

FILL FILL_1__11796_ (
);

FILL FILL_1__11376_ (
);

AOI22X1 _15939_ (
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .B(_5571_),
    .C(_5570__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_6397_)
);

FILL FILL_4__12710_ (
);

NAND3X1 _15519_ (
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .B(_5471__bF$buf3),
    .C(_5531__bF$buf2),
    .Y(_5988_)
);

FILL FILL_0__10789_ (
);

FILL FILL_0__8383_ (
);

FILL FILL_0__10369_ (
);

NAND2X1 _10654_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1914_)
);

NAND2X1 _10234_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1695_)
);

FILL FILL_3__11703_ (
);

FILL FILL_4__15182_ (
);

FILL FILL_2__9762_ (
);

FILL FILL_3__14595_ (
);

FILL FILL_0__11730_ (
);

FILL FILL_2__9342_ (
);

FILL FILL_3__14175_ (
);

FILL FILL_0__11310_ (
);

FILL FILL_4_BUFX2_insert890 (
);

FILL FILL_4_BUFX2_insert891 (
);

FILL FILL_4_BUFX2_insert892 (
);

FILL FILL_4__9268_ (
);

FILL FILL_4_BUFX2_insert893 (
);

FILL FILL112360x74050 (
);

FILL FILL_4_BUFX2_insert894 (
);

FILL FILL_2__13588_ (
);

FILL FILL_4_BUFX2_insert895 (
);

FILL FILL_2__13168_ (
);

FILL FILL_4_BUFX2_insert896 (
);

FILL FILL_4_BUFX2_insert897 (
);

FILL FILL_5__14922_ (
);

FILL FILL_4_BUFX2_insert898 (
);

FILL FILL_5__14502_ (
);

FILL FILL_4_BUFX2_insert899 (
);

DFFSR _8802_ (
    .Q(\datapath_1.regfile_1.regOut[15] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_913_[12])
);

FILL FILL_4__13915_ (
);

FILL FILL_3__7685_ (
);

NAND3X1 _11859_ (
    .A(_2868_),
    .B(_2790_),
    .C(_2816_),
    .Y(_2946_)
);

FILL FILL_0__9168_ (
);

AOI21X1 _11439_ (
    .A(_2554_),
    .B(_2549_),
    .C(_2445_),
    .Y(_2555_)
);

FILL SFILL3720x18050 (
);

AND2X2 _11019_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2138_)
);

FILL FILL_3__12908_ (
);

FILL FILL_1__13942_ (
);

FILL FILL_4__16387_ (
);

FILL FILL_1__13522_ (
);

FILL FILL_1__13102_ (
);

DFFSR _12800_ (
    .Q(\datapath_1.PCJump [11]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3490_[9])
);

FILL FILL_0__12515_ (
);

FILL FILL_5__8972_ (
);

FILL FILL_5__8132_ (
);

OAI22X1 _15692_ (
    .A(_4743_),
    .B(_5535__bF$buf0),
    .C(_5569_),
    .D(_4717_),
    .Y(_6156_)
);

NOR2X1 _15272_ (
    .A(_5744_),
    .B(_5746_),
    .Y(_5747_)
);

FILL FILL_5__15707_ (
);

FILL FILL_3__16321_ (
);

FILL FILL_1__8964_ (
);

FILL FILL_5__10422_ (
);

FILL FILL_1__8124_ (
);

FILL FILL_5__10002_ (
);

FILL FILL_2__15734_ (
);

FILL FILL_2__15314_ (
);

FILL FILL_1__14727_ (
);

INVX1 _7194_ (
    .A(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_156_)
);

FILL FILL_1__14307_ (
);

FILL FILL_3__9411_ (
);

FILL FILL112280x36050 (
);

FILL FILL_2__6887_ (
);

FILL FILL_5__9757_ (
);

FILL FILL_5__9337_ (
);

FILL FILL_6__12634_ (
);

OAI22X1 _16057_ (
    .A(_5472__bF$buf0),
    .B(_5161_),
    .C(_5160_),
    .D(_5552__bF$buf1),
    .Y(_6512_)
);

INVX1 _11192_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .Y(_2311_)
);

FILL FILL_5__11627_ (
);

FILL FILL_1__9749_ (
);

FILL FILL_3__12661_ (
);

FILL FILL_5__11207_ (
);

FILL FILL_3__12241_ (
);

FILL FILL_4__7754_ (
);

FILL FILL_4__7334_ (
);

FILL FILL_2__11654_ (
);

FILL FILL_2__11234_ (
);

FILL FILL_5__14099_ (
);

FILL SFILL54040x81050 (
);

OAI21X1 _8399_ (
    .A(_775_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .C(_776_),
    .Y(_718_[29])
);

FILL FILL_1__10647_ (
);

FILL FILL_5__15880_ (
);

FILL FILL_5__15460_ (
);

FILL FILL_5__15040_ (
);

INVX1 _9760_ (
    .A(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_1460_)
);

FILL FILL_0__7234_ (
);

FILL FILL_6__8201_ (
);

INVX1 _9340_ (
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_1241_)
);

FILL FILL_4__14873_ (
);

FILL FILL_4__14453_ (
);

FILL FILL_4__14033_ (
);

INVX1 _12397_ (
    .A(ALUOut[18]),
    .Y(_3330_)
);

FILL FILL_3__13866_ (
);

FILL FILL_2__8613_ (
);

FILL FILL_3__13446_ (
);

FILL FILL_1__14480_ (
);

FILL FILL_3__13026_ (
);

FILL FILL_1__14060_ (
);

FILL FILL_4__8959_ (
);

FILL FILL_4__8119_ (
);

FILL FILL_2__12859_ (
);

FILL FILL_2__12439_ (
);

FILL FILL_0__13893_ (
);

FILL FILL_2__12019_ (
);

FILL FILL_0__13473_ (
);

FILL FILL_5__9090_ (
);

FILL FILL_4__9900_ (
);

FILL FILL_2__13800_ (
);

FILL FILL_3__6956_ (
);

FILL FILL_0__8859_ (
);

FILL FILL_5__16245_ (
);

FILL FILL_0__8439_ (
);

FILL FILL_0__8019_ (
);

FILL FILL_5__11380_ (
);

FILL FILL_1__9082_ (
);

FILL FILL_4__15658_ (
);

FILL FILL_4__15238_ (
);

FILL FILL_2__16272_ (
);

FILL FILL_4__10793_ (
);

FILL FILL_4__10373_ (
);

FILL FILL_0__9800_ (
);

FILL FILL_1__15685_ (
);

FILL FILL_1__15265_ (
);

FILL FILL_5__7823_ (
);

NOR2X1 _14963_ (
    .A(_5440_),
    .B(_5443_),
    .Y(_5444_)
);

FILL FILL_0__14678_ (
);

FILL FILL_0__14258_ (
);

INVX1 _14543_ (
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_5033_)
);

INVX1 _14123_ (
    .A(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_4621_)
);

FILL FILL_1__7815_ (
);

FILL FILL_6__13592_ (
);

FILL FILL_5__12585_ (
);

FILL FILL_5__12165_ (
);

BUFX2 _6885_ (
    .A(_2_[15]),
    .Y(memoryWriteData[15])
);

FILL FILL_4__11998_ (
);

FILL FILL_4__11578_ (
);

FILL FILL_4__11158_ (
);

FILL FILL_2__12192_ (
);

FILL FILL_5__8608_ (
);

FILL FILL_1__11185_ (
);

NOR3X1 _15748_ (
    .A(_5515__bF$buf0),
    .B(_6210_),
    .C(_5521__bF$buf2),
    .Y(_6211_)
);

OAI22X1 _15328_ (
    .A(_4270_),
    .B(_5548__bF$buf2),
    .C(_5489__bF$buf1),
    .D(_5801_),
    .Y(_5802_)
);

FILL FILL_0__8192_ (
);

INVX1 _10883_ (
    .A(\aluControl_1.inst [1]),
    .Y(_2030_)
);

FILL FILL_0__10178_ (
);

DFFSR _10463_ (
    .Q(\datapath_1.regfile_1.regOut[28] [9]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_1758_[9])
);

FILL SFILL23880x28050 (
);

INVX1 _10043_ (
    .A(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_1608_)
);

FILL FILL_3__11932_ (
);

FILL FILL_3__11512_ (
);

FILL FILL_0__16404_ (
);

FILL FILL_2__10925_ (
);

FILL FILL_2__9991_ (
);

FILL FILL_2__10505_ (
);

FILL FILL112440x5050 (
);

FILL FILL_2__9151_ (
);

FILL FILL_4__9497_ (
);

FILL FILL_2__13397_ (
);

FILL FILL_5__14731_ (
);

FILL FILL_0__6925_ (
);

FILL FILL_5__14311_ (
);

INVX1 _8611_ (
    .A(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_877_)
);

FILL FILL_4__13724_ (
);

FILL FILL_4__13304_ (
);

FILL FILL_0__9397_ (
);

FILL FILL_3__7494_ (
);

FILL FILL_3__7074_ (
);

NAND2X1 _11668_ (
    .A(_2178_),
    .B(_2481__bF$buf3),
    .Y(_2770_)
);

XOR2X1 _11248_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2367_)
);

FILL FILL_3__12717_ (
);

FILL FILL_1__13751_ (
);

FILL FILL_1__13331_ (
);

FILL FILL_4__16196_ (
);

FILL FILL_0__12744_ (
);

FILL FILL_3__15189_ (
);

FILL FILL_0__12324_ (
);

FILL FILL_5__8781_ (
);

FILL FILL_5__8361_ (
);

FILL SFILL74120x73050 (
);

FILL SFILL74200x7050 (
);

FILL FILL_5__15936_ (
);

INVX2 _15081_ (
    .A(_5526__bF$buf3),
    .Y(_5560_)
);

FILL FILL_5__15516_ (
);

FILL FILL_3__16130_ (
);

DFFSR _9816_ (
    .Q(\datapath_1.regfile_1.regOut[23] [2]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_1433_[2])
);

FILL FILL_1__8773_ (
);

FILL FILL_5__10651_ (
);

FILL SFILL8440x11050 (
);

FILL FILL_1__8353_ (
);

FILL FILL_5__10231_ (
);

FILL FILL_4__14929_ (
);

FILL FILL_4__14509_ (
);

FILL FILL_2__15963_ (
);

FILL FILL_2__15543_ (
);

FILL FILL_2__15123_ (
);

FILL FILL_3__8699_ (
);

FILL SFILL13800x69050 (
);

FILL FILL_1__14956_ (
);

FILL FILL_1__14536_ (
);

FILL FILL_1__14116_ (
);

FILL FILL_3__9640_ (
);

FILL FILL_0__13949_ (
);

NOR2X1 _13814_ (
    .A(_4318_),
    .B(_4315_),
    .Y(_4319_)
);

FILL FILL_3__9220_ (
);

FILL FILL_0__13529_ (
);

FILL FILL_0__13109_ (
);

FILL FILL_5__9986_ (
);

FILL FILL_5__9146_ (
);

FILL FILL_6__12443_ (
);

NAND2X1 _16286_ (
    .A(_6734_),
    .B(_6733_),
    .Y(_6735_)
);

FILL FILL_5__11856_ (
);

FILL FILL_1__9978_ (
);

FILL FILL_3__12890_ (
);

FILL FILL_5__11436_ (
);

FILL FILL_3__12470_ (
);

FILL FILL_1__9138_ (
);

FILL FILL_5__11016_ (
);

FILL FILL_3__12050_ (
);

FILL FILL_4__7983_ (
);

FILL FILL_2__16328_ (
);

FILL FILL_4__7563_ (
);

FILL FILL_4__10429_ (
);

FILL FILL_2__11883_ (
);

FILL FILL_4__10009_ (
);

FILL FILL_2__11463_ (
);

FILL FILL_2__11043_ (
);

FILL FILL_6__7069_ (
);

FILL SFILL13800x24050 (
);

FILL FILL_1__10876_ (
);

FILL FILL_1__10036_ (
);

FILL FILL_0__7883_ (
);

FILL FILL_0__7463_ (
);

FILL FILL_0__7043_ (
);

FILL FILL_6__13648_ (
);

FILL FILL_4__14682_ (
);

FILL FILL_4__14262_ (
);

FILL SFILL64120x71050 (
);

FILL FILL_2__8842_ (
);

FILL FILL_3__13675_ (
);

FILL FILL_0__10810_ (
);

FILL FILL_3__13255_ (
);

FILL FILL_2__8002_ (
);

FILL FILL_4__8768_ (
);

FILL FILL_4__8348_ (
);

FILL FILL112360x69050 (
);

FILL FILL_2__12248_ (
);

FILL FILL_0__13282_ (
);

FILL SFILL64040x78050 (
);

FILL FILL_5__16054_ (
);

INVX1 _10939_ (
    .A(\control_1.op [4]),
    .Y(_2073_)
);

FILL FILL_0__8248_ (
);

INVX1 _10519_ (
    .A(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_1844_)
);

FILL FILL_4__15887_ (
);

FILL FILL_1__12602_ (
);

FILL FILL_4__15467_ (
);

FILL FILL_4__15047_ (
);

FILL FILL_2__16081_ (
);

FILL FILL_4__10182_ (
);

FILL FILL_2__9627_ (
);

FILL FILL_2__9207_ (
);

FILL FILL_1__15494_ (
);

FILL FILL_1__15074_ (
);

FILL FILL_5__7632_ (
);

FILL FILL_5__7212_ (
);

FILL FILL_0__14487_ (
);

NOR2X1 _14772_ (
    .A(_5253_),
    .B(_5256_),
    .Y(_5257_)
);

FILL FILL_0__14067_ (
);

NOR2X1 _14352_ (
    .A(_4845_),
    .B(_4842_),
    .Y(_4846_)
);

FILL FILL_3__15821_ (
);

FILL SFILL85080x7050 (
);

FILL FILL_3__15401_ (
);

FILL FILL_1__7624_ (
);

FILL FILL_1__7204_ (
);

FILL FILL_2__14814_ (
);

FILL SFILL64040x33050 (
);

FILL FILL_5__12394_ (
);

FILL FILL_1__13807_ (
);

FILL FILL_4__11387_ (
);

FILL FILL_3__8911_ (
);

FILL SFILL89240x82050 (
);

FILL FILL_1__16279_ (
);

FILL FILL_5__8837_ (
);

NAND2X1 _15977_ (
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .B(_5494_),
    .Y(_6434_)
);

OAI21X1 _15557_ (
    .A(_4557_),
    .B(_5535__bF$buf2),
    .C(_6024_),
    .Y(_6025_)
);

NAND2X1 _15137_ (
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .B(_5494_),
    .Y(_5615_)
);

INVX1 _10692_ (
    .A(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_1939_)
);

INVX1 _10272_ (
    .A(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_1720_)
);

FILL FILL_5__10707_ (
);

FILL FILL_1__8829_ (
);

FILL FILL_3__11741_ (
);

FILL FILL_6__14186_ (
);

FILL FILL_3__11321_ (
);

FILL FILL_0__16213_ (
);

FILL FILL_5__13599_ (
);

FILL SFILL54040x76050 (
);

FILL FILL_2__10314_ (
);

FILL FILL_2__9380_ (
);

DFFSR _7899_ (
    .Q(\datapath_1.regfile_1.regOut[8] [5]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_458_[5])
);

OAI21X1 _7479_ (
    .A(_304_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_305_),
    .Y(_263_[21])
);

OAI21X1 _7059_ (
    .A(_85_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .C(_86_),
    .Y(_68_[9])
);

FILL FILL_5__14960_ (
);

FILL FILL_5__14540_ (
);

FILL FILL_5__14120_ (
);

INVX1 _8840_ (
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_989_)
);

DFFSR _8420_ (
    .Q(\datapath_1.regfile_1.regOut[12] [14]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_718_[14])
);

OAI21X1 _8000_ (
    .A(_570_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_571_),
    .Y(_523_[24])
);

FILL FILL_1__12199_ (
);

FILL FILL_4__13953_ (
);

FILL FILL_4__13533_ (
);

FILL FILL_4__13113_ (
);

NAND2X1 _11897_ (
    .A(IorD_bF$buf2),
    .B(ALUOut[3]),
    .Y(_2973_)
);

OAI21X1 _11477_ (
    .A(_2591_),
    .B(_2287_),
    .C(_2438_),
    .Y(_2592_)
);

OAI21X1 _11057_ (
    .A(_2147_),
    .B(_2160_),
    .C(_2175_),
    .Y(_2176_)
);

FILL FILL_3__12526_ (
);

FILL FILL_1__13980_ (
);

FILL FILL_3__12106_ (
);

FILL FILL_1__13560_ (
);

FILL FILL_1__13140_ (
);

FILL FILL_4__7619_ (
);

FILL FILL_2__11939_ (
);

FILL FILL_0__12973_ (
);

FILL FILL_2__11519_ (
);

FILL FILL_0__12133_ (
);

FILL FILL_5__8590_ (
);

FILL FILL_5__15745_ (
);

FILL FILL_0__7939_ (
);

FILL FILL_5__15325_ (
);

OAI21X1 _9625_ (
    .A(_1389_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1390_),
    .Y(_1368_[11])
);

FILL FILL_5__10880_ (
);

DFFSR _9205_ (
    .Q(\datapath_1.regfile_1.regOut[18] [31]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_1108_[31])
);

FILL SFILL79240x80050 (
);

FILL FILL_1__8582_ (
);

FILL FILL_5__10040_ (
);

FILL FILL_4__14738_ (
);

FILL FILL_4__14318_ (
);

FILL FILL_2__15772_ (
);

FILL FILL_2__15352_ (
);

FILL FILL_3__8088_ (
);

FILL FILL_1__14765_ (
);

FILL FILL_1__14345_ (
);

FILL FILL_5__6903_ (
);

FILL FILL_0__13758_ (
);

FILL FILL_0__13338_ (
);

INVX1 _13623_ (
    .A(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_4132_)
);

DFFSR _13203_ (
    .Q(\datapath_1.PCJump [28]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3685_[28])
);

FILL FILL_5__9795_ (
);

FILL FILL_5__9375_ (
);

FILL SFILL44040x74050 (
);

NAND3X1 _16095_ (
    .A(_6542_),
    .B(_6548_),
    .C(_6547_),
    .Y(_6549_)
);

FILL FILL_1__9787_ (
);

FILL FILL_5__11665_ (
);

FILL FILL_1__9367_ (
);

FILL FILL_5__11245_ (
);

FILL FILL_2__16137_ (
);

FILL FILL_4__7372_ (
);

FILL FILL_4__10658_ (
);

FILL FILL_4__10238_ (
);

FILL FILL_2__11692_ (
);

FILL FILL_2__11272_ (
);

FILL FILL_1__10685_ (
);

FILL FILL_1__10265_ (
);

INVX1 _14828_ (
    .A(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_5312_)
);

INVX1 _14408_ (
    .A(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_4900_)
);

FILL FILL_2_BUFX2_insert225 (
);

FILL SFILL8520x44050 (
);

FILL FILL_2_BUFX2_insert226 (
);

FILL FILL_0__7692_ (
);

FILL FILL_2_BUFX2_insert227 (
);

FILL FILL_2_BUFX2_insert228 (
);

FILL FILL_2_BUFX2_insert229 (
);

FILL FILL_4__14491_ (
);

FILL FILL_6__13037_ (
);

FILL FILL_4__14071_ (
);

FILL FILL_0__15904_ (
);

FILL FILL_2__8651_ (
);

FILL FILL_2__8231_ (
);

FILL FILL_3__13484_ (
);

FILL FILL_4__8997_ (
);

FILL FILL_4__8577_ (
);

FILL FILL_2__12897_ (
);

FILL FILL_2__12477_ (
);

FILL FILL_2__12057_ (
);

FILL FILL_0__13091_ (
);

FILL FILL_5__13811_ (
);

FILL FILL_3__6994_ (
);

FILL FILL_5__16283_ (
);

FILL FILL_0__8897_ (
);

FILL FILL_0__8477_ (
);

INVX1 _10748_ (
    .A(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_1956_)
);

FILL FILL_0__8057_ (
);

DFFSR _10328_ (
    .Q(\datapath_1.regfile_1.regOut[27] [2]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_1693_[2])
);

FILL FILL_4__15696_ (
);

FILL FILL_1__12831_ (
);

FILL FILL_1__12411_ (
);

FILL FILL_4__15276_ (
);

FILL FILL_2__9856_ (
);

FILL FILL_0__11824_ (
);

FILL FILL_3__14689_ (
);

FILL FILL_2__9016_ (
);

FILL FILL_3__14269_ (
);

FILL FILL_0__11404_ (
);

FILL SFILL104360x8050 (
);

FILL FILL_5__7861_ (
);

FILL FILL_6__15603_ (
);

FILL SFILL74120x68050 (
);

FILL FILL_5__7441_ (
);

INVX1 _14581_ (
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_5070_)
);

FILL FILL_0__14296_ (
);

NOR2X1 _14161_ (
    .A(_4655_),
    .B(_4658_),
    .Y(_4659_)
);

FILL FILL_3__15630_ (
);

FILL FILL_3__15210_ (
);

FILL FILL_1__7853_ (
);

FILL FILL_1__7433_ (
);

FILL FILL_2__14623_ (
);

FILL FILL_2__14203_ (
);

FILL FILL_3__7359_ (
);

FILL FILL_1__13616_ (
);

FILL FILL_1_BUFX2_insert240 (
);

FILL FILL_4__11196_ (
);

FILL FILL_3__8720_ (
);

FILL FILL_1_BUFX2_insert241 (
);

FILL SFILL69160x40050 (
);

FILL FILL_0__12609_ (
);

FILL FILL_1_BUFX2_insert242 (
);

FILL FILL_1_BUFX2_insert243 (
);

FILL FILL_1_BUFX2_insert244 (
);

FILL FILL_1__16088_ (
);

FILL FILL_1_BUFX2_insert245 (
);

FILL FILL_1_BUFX2_insert246 (
);

FILL FILL_5__8646_ (
);

FILL FILL_3__10189_ (
);

FILL FILL_5__8226_ (
);

FILL FILL_1_BUFX2_insert247 (
);

FILL FILL_1_BUFX2_insert248 (
);

FILL FILL_1_BUFX2_insert249 (
);

NOR2X1 _15786_ (
    .A(_6247_),
    .B(_6239_),
    .Y(_6248_)
);

FILL FILL_6__11523_ (
);

OAI22X1 _15366_ (
    .A(_5837_),
    .B(_5548__bF$buf3),
    .C(_5489__bF$buf2),
    .D(_5838_),
    .Y(_5839_)
);

FILL FILL_6__11103_ (
);

FILL SFILL74120x23050 (
);

FILL FILL_3__16415_ (
);

FILL FILL_5__10936_ (
);

DFFSR _10081_ (
    .Q(\datapath_1.regfile_1.regOut[25] [11]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_1563_[11])
);

FILL FILL_1__8638_ (
);

FILL FILL_3__11970_ (
);

FILL FILL_5__10516_ (
);

FILL FILL_1__8218_ (
);

FILL FILL_3__11550_ (
);

FILL FILL_3__11130_ (
);

FILL FILL_2__15828_ (
);

FILL FILL_2__15408_ (
);

FILL FILL_0__16022_ (
);

FILL FILL_2__10963_ (
);

FILL FILL_2__10543_ (
);

FILL FILL_2__10123_ (
);

OAI21X1 _7288_ (
    .A(_261_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_262_),
    .Y(_198_[0])
);

FILL FILL_3__9925_ (
);

FILL FILL_3__9505_ (
);

FILL SFILL59160x83050 (
);

FILL FILL_0__6963_ (
);

FILL SFILL38280x42050 (
);

FILL FILL_4__13762_ (
);

FILL FILL_4__13342_ (
);

FILL SFILL64120x66050 (
);

AOI21X1 _11286_ (
    .A(_2178_),
    .B(_2404_),
    .C(_2402_),
    .Y(_2405_)
);

FILL FILL_2__7502_ (
);

FILL FILL_3__12755_ (
);

FILL FILL_3__12335_ (
);

FILL FILL_4__7848_ (
);

FILL FILL_4__7428_ (
);

FILL FILL_2__11748_ (
);

FILL FILL_0__12782_ (
);

FILL FILL_2__11328_ (
);

FILL FILL_0__12362_ (
);

FILL SFILL89320x1050 (
);

FILL SFILL89240x6050 (
);

FILL FILL_5__15974_ (
);

FILL FILL_5__15554_ (
);

FILL FILL_0__7748_ (
);

FILL FILL_5__15134_ (
);

FILL FILL_0__7328_ (
);

OAI21X1 _9854_ (
    .A(_1501_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .C(_1502_),
    .Y(_1498_[2])
);

DFFSR _9434_ (
    .Q(\datapath_1.regfile_1.regOut[20] [4]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_1238_[4])
);

NAND2X1 _9014_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1085_)
);

FILL FILL_1__8391_ (
);

FILL FILL_4__14967_ (
);

FILL FILL_4__14547_ (
);

FILL FILL_4__14127_ (
);

FILL FILL_2__15581_ (
);

FILL FILL_2__15161_ (
);

FILL FILL_2__8707_ (
);

FILL SFILL64120x21050 (
);

FILL FILL_1__14994_ (
);

FILL FILL_1__14574_ (
);

FILL FILL_1__14154_ (
);

FILL FILL_0__13987_ (
);

NAND3X1 _13852_ (
    .A(_4352_),
    .B(_4355_),
    .C(_4351_),
    .Y(_4356_)
);

FILL FILL_0__13567_ (
);

NAND3X1 _13432_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3883_),
    .C(_3919_),
    .Y(_3944_)
);

FILL FILL_0__13147_ (
);

FILL SFILL89320x70050 (
);

FILL FILL112360x19050 (
);

NAND2X1 _13012_ (
    .A(vdd),
    .B(\datapath_1.rd2 [20]),
    .Y(_3660_)
);

FILL FILL_3__14901_ (
);

FILL FILL_5__16339_ (
);

FILL SFILL64040x28050 (
);

FILL FILL_5__11894_ (
);

FILL FILL_5__11474_ (
);

FILL FILL_1__9596_ (
);

FILL FILL_5__11054_ (
);

FILL FILL_2__16366_ (
);

FILL FILL_4__7181_ (
);

FILL FILL_4__10887_ (
);

FILL FILL_4__10047_ (
);

FILL FILL_2__11081_ (
);

FILL SFILL54120x64050 (
);

FILL FILL_1__15779_ (
);

FILL FILL_1__15359_ (
);

FILL FILL_1__10494_ (
);

NOR2X1 _14637_ (
    .A(_5124_),
    .B(_5121_),
    .Y(_5125_)
);

AOI21X1 _14217_ (
    .A(_4713_),
    .B(_4692_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [15])
);

FILL FILL_2__7099_ (
);

FILL FILL_0__7081_ (
);

FILL FILL_1__16300_ (
);

FILL FILL_3__10821_ (
);

FILL FILL_3__10401_ (
);

FILL FILL_0__15713_ (
);

FILL FILL_2__8880_ (
);

FILL FILL_2__8460_ (
);

FILL FILL_5__12259_ (
);

FILL FILL_3__13293_ (
);

OAI21X1 _6979_ (
    .A(_52_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_53_),
    .Y(_3_[25])
);

FILL FILL_4__8386_ (
);

FILL FILL_2__12286_ (
);

FILL FILL_5__13620_ (
);

DFFSR _7920_ (
    .Q(\datapath_1.regfile_1.regOut[8] [26]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_458_[26])
);

FILL SFILL89240x32050 (
);

OAI21X1 _7500_ (
    .A(_318_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .C(_319_),
    .Y(_263_[28])
);

FILL FILL_1__11699_ (
);

FILL FILL_1__11279_ (
);

FILL FILL_4__12613_ (
);

FILL FILL_5__16092_ (
);

OAI21X1 _10977_ (
    .A(_2101_),
    .B(vdd),
    .C(_2102_),
    .Y(_2098_[1])
);

FILL FILL_6__9673_ (
);

OAI21X1 _10557_ (
    .A(_1868_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1869_),
    .Y(_1823_[23])
);

OAI21X1 _10137_ (
    .A(_1649_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1650_),
    .Y(_1628_[11])
);

FILL FILL_3__11606_ (
);

FILL SFILL18680x52050 (
);

FILL FILL_1__12640_ (
);

FILL FILL_1__12220_ (
);

FILL FILL_4__15085_ (
);

FILL FILL_2__9665_ (
);

FILL FILL_3__14498_ (
);

FILL FILL_0__11633_ (
);

FILL FILL_2__9245_ (
);

FILL FILL_0__11213_ (
);

FILL FILL_3__14078_ (
);

FILL FILL_5__7670_ (
);

FILL FILL_5__7250_ (
);

NAND3X1 _14390_ (
    .A(_4881_),
    .B(_4882_),
    .C(_4880_),
    .Y(_4883_)
);

FILL FILL_5__14825_ (
);

FILL FILL_5__14405_ (
);

OAI21X1 _8705_ (
    .A(_918_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_919_),
    .Y(_913_[3])
);

FILL SFILL79240x75050 (
);

FILL FILL_1__7242_ (
);

FILL FILL_4__13818_ (
);

FILL SFILL58360x34050 (
);

FILL FILL_2__14852_ (
);

FILL FILL_2__14432_ (
);

FILL FILL_3__7588_ (
);

FILL FILL_2__14012_ (
);

FILL FILL_3__7168_ (
);

FILL FILL_1__13845_ (
);

FILL FILL_1__13425_ (
);

FILL SFILL58920x8050 (
);

FILL FILL_1__13005_ (
);

FILL SFILL33960x1050 (
);

FILL FILL_0__12838_ (
);

FILL SFILL33880x6050 (
);

OAI21X1 _12703_ (
    .A(_3493_),
    .B(IRWrite_bF$buf2),
    .C(_3494_),
    .Y(_3490_[2])
);

FILL FILL_0__12418_ (
);

FILL FILL_5__8875_ (
);

FILL SFILL44040x69050 (
);

FILL FILL_5__8455_ (
);

OAI21X1 _15595_ (
    .A(_4601_),
    .B(_5535__bF$buf3),
    .C(_6061_),
    .Y(_6062_)
);

AOI22X1 _15175_ (
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .B(_5567_),
    .C(_5565__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_5652_)
);

FILL FILL_3__16224_ (
);

FILL FILL_5__10745_ (
);

FILL FILL_1__8867_ (
);

FILL FILL_1__8447_ (
);

FILL FILL_5__10325_ (
);

FILL FILL_2__15637_ (
);

FILL SFILL79240x30050 (
);

FILL FILL_2__15217_ (
);

FILL FILL_4__6872_ (
);

FILL FILL_0__16251_ (
);

FILL FILL_2__10772_ (
);

NAND2X1 _7097_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_112_)
);

FILL FILL_3__9734_ (
);

NOR2X1 _13908_ (
    .A(_4410_),
    .B(_4400_),
    .Y(_4411_)
);

FILL SFILL8520x39050 (
);

FILL SFILL109400x56050 (
);

FILL FILL_4__13991_ (
);

FILL FILL_4__13571_ (
);

FILL SFILL44040x24050 (
);

FILL FILL_4__13151_ (
);

AOI21X1 _11095_ (
    .A(_2211_),
    .B(_2177_),
    .C(_2213_),
    .Y(_2214_)
);

FILL FILL_3__12984_ (
);

FILL FILL_2__7731_ (
);

FILL FILL_2__7311_ (
);

FILL FILL_3__12144_ (
);

FILL SFILL69240x73050 (
);

FILL FILL_4__7237_ (
);

FILL FILL_2__11977_ (
);

FILL FILL_2__11557_ (
);

FILL FILL_0__12591_ (
);

FILL FILL_2__11137_ (
);

FILL FILL_0__12171_ (
);

FILL FILL_6__16370_ (
);

FILL SFILL114680x76050 (
);

FILL SFILL88440x28050 (
);

FILL FILL_5__15783_ (
);

FILL FILL_5__15363_ (
);

FILL FILL_0__7977_ (
);

FILL FILL_0__7557_ (
);

NAND2X1 _9663_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1416_)
);

NAND2X1 _9243_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1197_)
);

FILL FILL_1__11911_ (
);

FILL FILL_4__14776_ (
);

FILL FILL_4__14356_ (
);

FILL FILL_2__15390_ (
);

FILL SFILL109400x11050 (
);

FILL FILL_0__10904_ (
);

FILL FILL_3__13769_ (
);

FILL FILL_2__8516_ (
);

FILL FILL_3__13349_ (
);

FILL FILL_1__14383_ (
);

FILL FILL_5__6941_ (
);

FILL FILL_1_BUFX2_insert1000 (
);

FILL FILL_1_BUFX2_insert1001 (
);

FILL FILL_1_BUFX2_insert1002 (
);

FILL FILL_1_BUFX2_insert1003 (
);

FILL FILL_0__13796_ (
);

OAI22X1 _13661_ (
    .A(_4167_),
    .B(_3936__bF$buf0),
    .C(_3978_),
    .D(_4168_),
    .Y(_4169_)
);

FILL FILL_0__13376_ (
);

FILL FILL_1_BUFX2_insert1004 (
);

NOR2X1 _13241_ (
    .A(_3776_),
    .B(_3783_),
    .Y(_3784_)
);

FILL FILL_1_BUFX2_insert1005 (
);

FILL FILL_1_BUFX2_insert1006 (
);

FILL FILL_3__14710_ (
);

FILL FILL_1_BUFX2_insert1007 (
);

FILL FILL_1_BUFX2_insert1008 (
);

FILL FILL_1_BUFX2_insert1009 (
);

FILL FILL_1__6933_ (
);

FILL FILL_4__9803_ (
);

FILL FILL_6__12290_ (
);

FILL FILL_2__13703_ (
);

FILL FILL_3__6859_ (
);

FILL FILL_5__16148_ (
);

FILL FILL_5__11283_ (
);

FILL FILL_2__16175_ (
);

FILL SFILL99400x60050 (
);

FILL FILL_4__10696_ (
);

FILL FILL_4__10276_ (
);

FILL SFILL69160x35050 (
);

FILL FILL_3__7800_ (
);

FILL FILL_1__15588_ (
);

FILL FILL_1__15168_ (
);

FILL FILL_5__7726_ (
);

FILL FILL_5__7306_ (
);

FILL FILL_2_BUFX2_insert600 (
);

FILL FILL_2_BUFX2_insert601 (
);

FILL FILL_2_BUFX2_insert602 (
);

FILL FILL_2_BUFX2_insert603 (
);

NOR2X1 _14866_ (
    .A(_5345_),
    .B(_5348_),
    .Y(_5349_)
);

FILL SFILL74120x18050 (
);

FILL FILL_2_BUFX2_insert604 (
);

AOI22X1 _14446_ (
    .A(_3891__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [20]),
    .C(\datapath_1.regfile_1.regOut[8] [20]),
    .D(_4090_),
    .Y(_4938_)
);

FILL FILL_2_BUFX2_insert605 (
);

INVX1 _14026_ (
    .A(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_4526_)
);

FILL SFILL28920x7050 (
);

FILL FILL_3__15915_ (
);

FILL FILL_2_BUFX2_insert606 (
);

FILL FILL_2_BUFX2_insert607 (
);

FILL FILL_2_BUFX2_insert608 (
);

FILL FILL_2_BUFX2_insert609 (
);

FILL FILL_1__7718_ (
);

FILL FILL_6__13495_ (
);

FILL FILL_3__10630_ (
);

FILL FILL_2__14908_ (
);

FILL SFILL99320x67050 (
);

FILL FILL_0__15942_ (
);

FILL FILL_0__15522_ (
);

FILL FILL_0__15102_ (
);

FILL FILL_5__12488_ (
);

FILL FILL_5__12068_ (
);

FILL SFILL8840x3050 (
);

FILL SFILL69080x1050 (
);

FILL FILL_4__8195_ (
);

FILL SFILL8760x8050 (
);

FILL SFILL59160x78050 (
);

FILL FILL_2__12095_ (
);

FILL FILL_1__11088_ (
);

FILL FILL_4__12842_ (
);

FILL FILL_4__12422_ (
);

FILL FILL_4__12002_ (
);

OAI21X1 _10786_ (
    .A(_1980_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .C(_1981_),
    .Y(_1953_[14])
);

FILL FILL_0__8095_ (
);

OAI21X1 _10366_ (
    .A(_1761_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .C(_1762_),
    .Y(_1758_[2])
);

FILL FILL_3__11835_ (
);

FILL FILL_3__11415_ (
);

FILL FILL_4__6928_ (
);

FILL FILL_0__16307_ (
);

FILL FILL_2__10828_ (
);

FILL FILL_2__9894_ (
);

FILL FILL_2__10408_ (
);

FILL FILL_2__9474_ (
);

FILL FILL_0__11862_ (
);

FILL FILL_0__11442_ (
);

FILL FILL_0__11022_ (
);

FILL FILL_5__14634_ (
);

FILL FILL_5__14214_ (
);

DFFSR _8934_ (
    .Q(\datapath_1.regfile_1.regOut[16] [16]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_978_[16])
);

FILL SFILL59160x33050 (
);

NAND2X1 _8514_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_833_)
);

FILL FILL_1__7891_ (
);

FILL FILL_1__7471_ (
);

FILL FILL_1__7051_ (
);

FILL FILL_4__13627_ (
);

FILL FILL_4__13207_ (
);

FILL FILL_2__14661_ (
);

FILL FILL_2__14241_ (
);

FILL FILL_3_BUFX2_insert60 (
);

FILL FILL_1__13654_ (
);

FILL FILL_3_BUFX2_insert61 (
);

FILL FILL_1__13234_ (
);

FILL FILL_3_BUFX2_insert62 (
);

FILL FILL_4__16099_ (
);

FILL FILL_3_BUFX2_insert63 (
);

FILL FILL_3_BUFX2_insert64 (
);

FILL FILL_3_BUFX2_insert65 (
);

FILL FILL_1_BUFX2_insert620 (
);

FILL FILL_3_BUFX2_insert66 (
);

FILL FILL_1_BUFX2_insert621 (
);

FILL FILL_3_BUFX2_insert67 (
);

FILL FILL_0__12647_ (
);

FILL FILL_1_BUFX2_insert622 (
);

FILL FILL_3_BUFX2_insert68 (
);

DFFSR _12932_ (
    .Q(\datapath_1.a [13]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_3555_[13])
);

FILL SFILL73720x80050 (
);

NAND2X1 _12512_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [24]),
    .Y(_3408_)
);

FILL FILL_1_BUFX2_insert623 (
);

FILL FILL_3_BUFX2_insert69 (
);

FILL FILL_0__12227_ (
);

FILL SFILL28680x49050 (
);

FILL FILL_1_BUFX2_insert624 (
);

FILL FILL_1_BUFX2_insert625 (
);

FILL FILL_1_BUFX2_insert626 (
);

FILL FILL_1_BUFX2_insert627 (
);

FILL FILL_5__8264_ (
);

FILL FILL_1_BUFX2_insert628 (
);

FILL FILL_1_BUFX2_insert629 (
);

FILL FILL_5__15839_ (
);

FILL FILL_5__15419_ (
);

FILL FILL_3__16033_ (
);

NAND2X1 _9719_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .Y(_1497_)
);

FILL SFILL49160x76050 (
);

FILL FILL_5__10974_ (
);

FILL FILL_5__10554_ (
);

FILL FILL_1__8256_ (
);

FILL FILL_5__10134_ (
);

FILL FILL_2__15866_ (
);

FILL FILL_2__15446_ (
);

FILL FILL_2__15026_ (
);

FILL FILL_0__16060_ (
);

FILL FILL_2__10581_ (
);

FILL SFILL54120x59050 (
);

FILL FILL_2__10161_ (
);

FILL FILL_1__14859_ (
);

FILL FILL_1__14439_ (
);

FILL FILL_1__14019_ (
);

FILL FILL_3__9543_ (
);

FILL FILL_3__9123_ (
);

AOI21X1 _13717_ (
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .B(_4090_),
    .C(_4223_),
    .Y(_4224_)
);

FILL FILL_5__9889_ (
);

FILL FILL_1__15800_ (
);

FILL FILL_5__9469_ (
);

FILL FILL_6__12346_ (
);

FILL FILL_4__13380_ (
);

NOR2X1 _16189_ (
    .A(_6638_),
    .B(_6640_),
    .Y(_6641_)
);

FILL FILL_2__7960_ (
);

FILL FILL_5__11759_ (
);

FILL FILL_5__11339_ (
);

FILL FILL_3__12373_ (
);

FILL FILL_2__7120_ (
);

FILL SFILL18760x40050 (
);

FILL FILL_4__7886_ (
);

FILL FILL_4__7466_ (
);

FILL FILL_4__7046_ (
);

FILL FILL_2__11786_ (
);

FILL FILL_2__11366_ (
);

FILL FILL_5__12700_ (
);

FILL SFILL54120x14050 (
);

FILL FILL_1__10779_ (
);

FILL FILL_1__10359_ (
);

FILL FILL_5__15592_ (
);

FILL FILL_5__15172_ (
);

NAND2X1 _9892_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1528_)
);

FILL FILL_0__7366_ (
);

NAND2X1 _9472_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1309_)
);

DFFSR _9052_ (
    .Q(\datapath_1.regfile_1.regOut[17] [6]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1043_[6])
);

FILL SFILL79320x63050 (
);

FILL SFILL18680x47050 (
);

FILL FILL_4__14585_ (
);

FILL FILL_1__11720_ (
);

FILL FILL_4__14165_ (
);

FILL FILL_1__11300_ (
);

FILL FILL_3__13998_ (
);

FILL FILL_2__8745_ (
);

FILL FILL_3__13578_ (
);

FILL FILL_2__8325_ (
);

FILL FILL111960x76050 (
);

FILL FILL_3__13158_ (
);

FILL FILL_1__14192_ (
);

FILL FILL_6__14912_ (
);

OAI22X1 _13890_ (
    .A(_4392_),
    .B(_3983__bF$buf1),
    .C(_3920_),
    .D(_4391_),
    .Y(_4393_)
);

NAND3X1 _13470_ (
    .A(_3898_),
    .B(_3880_),
    .C(_3883_),
    .Y(_3982_)
);

DFFSR _13050_ (
    .Q(_2_[3]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_3620_[3])
);

FILL FILL_5__13905_ (
);

FILL FILL_4__9612_ (
);

FILL FILL_2__13932_ (
);

FILL FILL_5__16377_ (
);

FILL FILL_2__13512_ (
);

FILL FILL_5__11092_ (
);

FILL FILL_1__12505_ (
);

FILL FILL_0__9932_ (
);

FILL FILL_0__9512_ (
);

FILL FILL_0__11918_ (
);

FILL FILL_1__15397_ (
);

FILL FILL_5__7955_ (
);

FILL FILL_5__7115_ (
);

FILL FILL_4__16311_ (
);

FILL FILL111960x31050 (
);

FILL FILL_6__10832_ (
);

OAI22X1 _14675_ (
    .A(_5160_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf0),
    .D(_5161_),
    .Y(_5162_)
);

INVX1 _14255_ (
    .A(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_4751_)
);

FILL FILL_3__15724_ (
);

FILL FILL_3__15304_ (
);

FILL FILL_1__7947_ (
);

FILL FILL_1__7107_ (
);

FILL SFILL79240x25050 (
);

FILL FILL_2__14717_ (
);

FILL FILL_0__15751_ (
);

FILL FILL_0__15331_ (
);

FILL FILL_5__12297_ (
);

FILL FILL111880x38050 (
);

FILL SFILL69320x61050 (
);

FILL SFILL44040x19050 (
);

FILL FILL_4__12651_ (
);

FILL FILL_4__12231_ (
);

FILL FILL_6__9291_ (
);

DFFSR _10595_ (
    .Q(\datapath_1.regfile_1.regOut[29] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1823_[13])
);

NAND2X1 _10175_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1676_)
);

FILL FILL_3__11644_ (
);

FILL FILL_3__11224_ (
);

FILL FILL_0__16116_ (
);

OAI21X1 _16401_ (
    .A(_6820_),
    .B(gnd),
    .C(_6821_),
    .Y(_6769_[26])
);

FILL FILL_2__10637_ (
);

FILL FILL_2__9283_ (
);

FILL FILL_0__11671_ (
);

FILL FILL_0__11251_ (
);

FILL FILL_6__15030_ (
);

FILL FILL_5__14863_ (
);

FILL FILL_5__14443_ (
);

FILL FILL_5__14023_ (
);

NAND2X1 _8743_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_945_)
);

NAND2X1 _8323_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_726_)
);

FILL FILL_4__13856_ (
);

FILL FILL_4__13436_ (
);

FILL FILL_2__14890_ (
);

FILL FILL_2__14470_ (
);

FILL FILL_4__13016_ (
);

FILL FILL_2__14050_ (
);

FILL FILL_3__12849_ (
);

FILL FILL_1__13883_ (
);

FILL FILL_3__12429_ (
);

FILL FILL_1__13463_ (
);

FILL FILL_3__12009_ (
);

FILL FILL_1__13043_ (
);

FILL FILL_0__12876_ (
);

NAND2X1 _12741_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[15]),
    .Y(_3520_)
);

FILL FILL_0__12456_ (
);

FILL FILL_0__12036_ (
);

AOI22X1 _12321_ (
    .A(_2_[26]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3280_)
);

FILL FILL_5__8493_ (
);

FILL FILL_5__8073_ (
);

FILL SFILL93720x34050 (
);

FILL FILL_5__15648_ (
);

FILL FILL_5__15228_ (
);

DFFSR _9948_ (
    .Q(\datapath_1.regfile_1.regOut[24] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_1498_[6])
);

FILL FILL_3__16262_ (
);

INVX1 _9528_ (
    .A(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_1346_)
);

FILL FILL_5__10783_ (
);

INVX1 _9108_ (
    .A(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_1127_)
);

FILL FILL_1__8485_ (
);

FILL FILL_5__10363_ (
);

FILL FILL_1__8065_ (
);

FILL FILL_2__15675_ (
);

FILL FILL_2__15255_ (
);

FILL SFILL99400x55050 (
);

FILL FILL_2__10390_ (
);

FILL FILL_1__14668_ (
);

FILL FILL_1__14248_ (
);

FILL FILL_0_BUFX2_insert280 (
);

FILL FILL_0_BUFX2_insert281 (
);

FILL FILL_0_BUFX2_insert282 (
);

FILL FILL_3__9772_ (
);

FILL FILL_0_BUFX2_insert283 (
);

FILL FILL_3__9352_ (
);

FILL FILL_0_BUFX2_insert284 (
);

INVX1 _13946_ (
    .A(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_4448_)
);

FILL FILL_0_BUFX2_insert285 (
);

NOR2X1 _13526_ (
    .A(_4036_),
    .B(_4033_),
    .Y(_4037_)
);

FILL FILL_0_BUFX2_insert286 (
);

INVX1 _13106_ (
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_3702_)
);

FILL FILL_0_BUFX2_insert287 (
);

FILL FILL_0_BUFX2_insert288 (
);

FILL FILL_5__9278_ (
);

FILL FILL_0_BUFX2_insert289 (
);

FILL SFILL83720x77050 (
);

FILL FILL_0__14602_ (
);

FILL FILL_5__11988_ (
);

FILL FILL_5__11568_ (
);

FILL FILL_5__11148_ (
);

FILL FILL_3__12182_ (
);

FILL FILL_4__7695_ (
);

FILL SFILL59640x35050 (
);

FILL FILL_2__11595_ (
);

FILL FILL_2__11175_ (
);

FILL SFILL99400x10050 (
);

FILL FILL_1__10168_ (
);

FILL FILL_4__11922_ (
);

FILL FILL_4__11502_ (
);

FILL FILL_0__7595_ (
);

FILL FILL_0__7175_ (
);

INVX1 _9281_ (
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_1222_)
);

FILL FILL_3__10915_ (
);

FILL FILL_4__14394_ (
);

FILL FILL_0__15807_ (
);

FILL FILL_2__8974_ (
);

FILL SFILL99320x17050 (
);

FILL FILL_0__10942_ (
);

FILL FILL_3__13387_ (
);

FILL FILL_0__10522_ (
);

FILL FILL_2__8134_ (
);

FILL FILL_0__10102_ (
);

FILL FILL_5__13714_ (
);

FILL SFILL28760x37050 (
);

FILL SFILL59160x28050 (
);

FILL FILL_1__6971_ (
);

FILL FILL_4__9421_ (
);

FILL FILL_4__12707_ (
);

FILL FILL_4__9001_ (
);

FILL FILL_2__13741_ (
);

FILL FILL_2__13321_ (
);

FILL FILL_5__16186_ (
);

FILL FILL_3__6897_ (
);

FILL FILL_6__9767_ (
);

FILL FILL_1__12734_ (
);

FILL FILL_4__15599_ (
);

FILL FILL_4__15179_ (
);

FILL FILL_1__12314_ (
);

FILL FILL_0__9741_ (
);

FILL FILL_2__9759_ (
);

FILL FILL_2__9339_ (
);

FILL FILL_0__11727_ (
);

FILL FILL_0__11307_ (
);

FILL FILL_6__15506_ (
);

FILL FILL_5__7764_ (
);

FILL FILL_5__7344_ (
);

FILL FILL_4__16120_ (
);

FILL FILL_6__10641_ (
);

FILL FILL_0__14199_ (
);

INVX1 _14484_ (
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_4975_)
);

AOI22X1 _14064_ (
    .A(_4129_),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .C(\datapath_1.regfile_1.regOut[6] [12]),
    .D(_4001__bF$buf2),
    .Y(_4564_)
);

FILL FILL_5__14919_ (
);

FILL FILL_3__15953_ (
);

FILL FILL_3__15533_ (
);

FILL FILL_3__15113_ (
);

FILL FILL_1__7756_ (
);

FILL FILL_1__7336_ (
);

FILL FILL_2__14946_ (
);

FILL FILL_0__15980_ (
);

FILL FILL_2__14526_ (
);

FILL FILL_0__15560_ (
);

FILL FILL_2__14106_ (
);

FILL FILL_0__15140_ (
);

FILL SFILL89720x29050 (
);

FILL FILL_1__13939_ (
);

FILL FILL_1__13519_ (
);

FILL FILL_4__11099_ (
);

FILL FILL_3__8623_ (
);

FILL FILL_3__8203_ (
);

FILL FILL_5__8969_ (
);

FILL SFILL89320x15050 (
);

FILL FILL_5__8129_ (
);

FILL SFILL69160x50 (
);

NAND3X1 _15689_ (
    .A(_6149_),
    .B(_6153_),
    .C(_6145_),
    .Y(_6154_)
);

FILL FILL_4__12880_ (
);

FILL FILL_4__12460_ (
);

FILL FILL_6__11006_ (
);

OAI22X1 _15269_ (
    .A(_5743_),
    .B(_5545__bF$buf3),
    .C(_5569_),
    .D(_4207_),
    .Y(_5744_)
);

FILL FILL_4__12040_ (
);

FILL FILL_3__16318_ (
);

FILL FILL_5__9910_ (
);

FILL FILL_3__11873_ (
);

FILL FILL_5__10419_ (
);

FILL FILL_3__11453_ (
);

FILL SFILL18760x35050 (
);

FILL FILL_3__11033_ (
);

FILL FILL_4__6966_ (
);

FILL FILL_0__16345_ (
);

NAND3X1 _16210_ (
    .A(_6655_),
    .B(_6656_),
    .C(_6660_),
    .Y(_6661_)
);

FILL FILL_2__10446_ (
);

FILL FILL_2__9092_ (
);

FILL FILL_2__10026_ (
);

FILL FILL_0__11480_ (
);

FILL FILL_0__11060_ (
);

FILL FILL_1__9902_ (
);

FILL FILL_3__9408_ (
);

FILL FILL_5__14672_ (
);

FILL FILL_5__14252_ (
);

FILL FILL_0__6866_ (
);

NAND2X1 _8972_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1057_)
);

DFFSR _8552_ (
    .Q(\datapath_1.regfile_1.regOut[13] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_783_[18])
);

INVX1 _8132_ (
    .A(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_639_)
);

FILL SFILL33960x10050 (
);

FILL FILL_4__13665_ (
);

FILL FILL_1__10800_ (
);

FILL FILL_4__13245_ (
);

OAI21X1 _11189_ (
    .A(_2296_),
    .B(_2305_),
    .C(_2307_),
    .Y(_2308_)
);

FILL FILL_2__7825_ (
);

FILL FILL_3__12658_ (
);

FILL FILL_3__12238_ (
);

FILL FILL_1__13692_ (
);

FILL FILL_1__13272_ (
);

NAND2X1 _12970_ (
    .A(vdd),
    .B(\datapath_1.rd2 [6]),
    .Y(_3632_)
);

DFFSR _12550_ (
    .Q(ALUOut[15]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3360_[15])
);

FILL FILL_0__12265_ (
);

INVX1 _12130_ (
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_3140_)
);

FILL FILL_5__15877_ (
);

FILL FILL_5__15457_ (
);

FILL FILL_5__15037_ (
);

FILL FILL_3__16071_ (
);

INVX1 _9757_ (
    .A(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_1458_)
);

INVX1 _9337_ (
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_1239_)
);

FILL FILL_5__10172_ (
);

FILL FILL_2__15484_ (
);

FILL SFILL114440x83050 (
);

FILL FILL_2__15064_ (
);

FILL FILL_1__14897_ (
);

FILL FILL_1__14477_ (
);

FILL FILL_1__14057_ (
);

FILL FILL_4__15811_ (
);

OAI22X1 _13755_ (
    .A(_4260_),
    .B(_3949_),
    .C(_3983__bF$buf3),
    .D(_4259_),
    .Y(_4261_)
);

FILL FILL_3__9161_ (
);

INVX1 _13335_ (
    .A(_3769_),
    .Y(_3858_)
);

FILL FILL_3__14804_ (
);

FILL FILL_5__9087_ (
);

FILL FILL_0__14831_ (
);

FILL FILL_0__14411_ (
);

FILL FILL_5__11797_ (
);

FILL FILL_1__9499_ (
);

FILL FILL_5__11377_ (
);

FILL FILL_1__9079_ (
);

FILL FILL_2__16269_ (
);

FILL SFILL69320x56050 (
);

FILL FILL_4__7084_ (
);

FILL FILL_1__10397_ (
);

FILL FILL_4__11731_ (
);

FILL FILL_4__11311_ (
);

FILL FILL_6__8371_ (
);

INVX1 _9090_ (
    .A(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_1115_)
);

FILL FILL_1__16203_ (
);

FILL FILL_3__10304_ (
);

NOR2X1 _15901_ (
    .A(_6358_),
    .B(_6359_),
    .Y(_6360_)
);

FILL FILL_0__15616_ (
);

FILL FILL_2__8783_ (
);

FILL FILL_0__10751_ (
);

FILL FILL_2__8363_ (
);

FILL FILL_2__12189_ (
);

FILL FILL_5__13943_ (
);

FILL FILL_5__13523_ (
);

FILL FILL_5__13103_ (
);

NAND2X1 _7823_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_474_)
);

DFFSR _7403_ (
    .Q(\datapath_1.regfile_1.regOut[4] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_198_[21])
);

FILL FILL_4_BUFX2_insert510 (
);

FILL FILL_4_BUFX2_insert511 (
);

FILL FILL_4__9650_ (
);

FILL FILL_4__9230_ (
);

FILL FILL_4_BUFX2_insert512 (
);

FILL FILL_4__12516_ (
);

FILL FILL_4_BUFX2_insert513 (
);

FILL FILL_2__13970_ (
);

FILL FILL_4_BUFX2_insert514 (
);

FILL FILL_2__13550_ (
);

FILL FILL_4_BUFX2_insert515 (
);

FILL FILL_2__13130_ (
);

FILL FILL_4_BUFX2_insert516 (
);

FILL FILL_0__8189_ (
);

FILL FILL_6__9156_ (
);

FILL FILL_4_BUFX2_insert517 (
);

FILL FILL_4_BUFX2_insert518 (
);

FILL FILL_4_BUFX2_insert519 (
);

FILL FILL_3__11929_ (
);

FILL FILL_1__12963_ (
);

FILL FILL_3__11509_ (
);

FILL FILL_1__12123_ (
);

FILL FILL_2__9988_ (
);

FILL SFILL69240x18050 (
);

FILL FILL_0__9550_ (
);

FILL FILL_0__11956_ (
);

FILL FILL_2__9148_ (
);

FILL FILL_0__9130_ (
);

OAI21X1 _11821_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(_2126_),
    .C(_2492_),
    .Y(_2911_)
);

FILL FILL_0__11536_ (
);

FILL FILL_0__11116_ (
);

OAI21X1 _11401_ (
    .A(_2167_),
    .B(_2513_),
    .C(_2517_),
    .Y(_2518_)
);

FILL FILL_5__7993_ (
);

FILL FILL_5__7573_ (
);

OAI22X1 _14293_ (
    .A(_4786_),
    .B(_3893__bF$buf0),
    .C(_3916_),
    .D(_4787_),
    .Y(_4788_)
);

FILL FILL_5__14728_ (
);

FILL FILL_5__14308_ (
);

FILL FILL_3__15762_ (
);

FILL FILL_3__15342_ (
);

INVX1 _8608_ (
    .A(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_875_)
);

FILL FILL_1__7985_ (
);

FILL FILL_1__7565_ (
);

FILL SFILL7800x70050 (
);

FILL FILL_2__14755_ (
);

FILL FILL_2__14335_ (
);

FILL FILL_1__13748_ (
);

FILL FILL_1__13328_ (
);

FILL FILL_3__8852_ (
);

INVX1 _12606_ (
    .A(\datapath_1.Data [13]),
    .Y(_3450_)
);

FILL FILL_3__8012_ (
);

FILL FILL_5__8778_ (
);

FILL SFILL104360x43050 (
);

FILL FILL_5__8358_ (
);

OAI22X1 _15498_ (
    .A(_5489__bF$buf2),
    .B(_4507_),
    .C(_5527__bF$buf0),
    .D(_4478_),
    .Y(_5967_)
);

INVX1 _15078_ (
    .A(_5534__bF$buf3),
    .Y(_5557_)
);

FILL FILL_3__16127_ (
);

FILL FILL_5__10648_ (
);

FILL FILL_3__11682_ (
);

FILL FILL_3__11262_ (
);

FILL FILL_0__16154_ (
);

FILL FILL_2__10675_ (
);

FILL FILL_2__10255_ (
);

FILL FILL_3__9637_ (
);

FILL FILL_3_BUFX2_insert530 (
);

FILL FILL_3__9217_ (
);

FILL FILL_3_BUFX2_insert531 (
);

FILL FILL_3_BUFX2_insert532 (
);

FILL FILL_5__14481_ (
);

FILL FILL_3_BUFX2_insert533 (
);

FILL FILL_3_BUFX2_insert534 (
);

FILL FILL_5__14061_ (
);

FILL FILL_3_BUFX2_insert535 (
);

INVX1 _8781_ (
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_970_)
);

FILL FILL_3_BUFX2_insert536 (
);

INVX1 _8361_ (
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_751_)
);

FILL FILL_3_BUFX2_insert537 (
);

FILL FILL_3_BUFX2_insert538 (
);

FILL FILL_3_BUFX2_insert539 (
);

FILL FILL_4__13894_ (
);

FILL FILL_4__13474_ (
);

FILL FILL_3__12887_ (
);

FILL FILL_2__7634_ (
);

FILL FILL_3__12467_ (
);

FILL FILL_2__7214_ (
);

FILL FILL_3__12047_ (
);

FILL FILL_1__13081_ (
);

FILL FILL_0__12494_ (
);

FILL SFILL89400x48050 (
);

FILL FILL_0__12074_ (
);

FILL FILL_6__16273_ (
);

FILL FILL_4__8501_ (
);

FILL FILL_5__15686_ (
);

FILL FILL_2__12401_ (
);

FILL FILL_5__15266_ (
);

FILL FILL_6__8847_ (
);

INVX1 _9986_ (
    .A(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_1570_)
);

DFFSR _9566_ (
    .Q(\datapath_1.regfile_1.regOut[21] [8]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_1303_[8])
);

FILL SFILL49240x59050 (
);

OAI21X1 _9146_ (
    .A(_1151_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1152_),
    .Y(_1108_[22])
);

FILL FILL_1__11814_ (
);

FILL FILL_4__14679_ (
);

FILL FILL_4__14259_ (
);

FILL FILL_2__15293_ (
);

FILL FILL_2__8839_ (
);

FILL FILL_0__10807_ (
);

FILL FILL_0__8401_ (
);

FILL FILL_1__14286_ (
);

FILL FILL_5__6844_ (
);

FILL FILL_0_BUFX2_insert660 (
);

FILL FILL_4__15620_ (
);

FILL FILL_0_BUFX2_insert661 (
);

FILL FILL_4__15200_ (
);

FILL FILL_0_BUFX2_insert662 (
);

FILL FILL_0_BUFX2_insert663 (
);

INVX1 _13984_ (
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_4485_)
);

FILL FILL_3__9390_ (
);

FILL FILL_0_BUFX2_insert664 (
);

FILL FILL_0__13699_ (
);

FILL FILL_0__13279_ (
);

INVX1 _13564_ (
    .A(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_4074_)
);

FILL FILL_0_BUFX2_insert665 (
);

OAI21X1 _13144_ (
    .A(_3726_),
    .B(PCEn_bF$buf4),
    .C(_3727_),
    .Y(_3685_[21])
);

FILL FILL_0_BUFX2_insert666 (
);

FILL FILL_0_BUFX2_insert667 (
);

FILL FILL_3__14613_ (
);

FILL FILL_0_BUFX2_insert668 (
);

FILL FILL_0_BUFX2_insert669 (
);

FILL FILL_1__6836_ (
);

FILL SFILL94280x54050 (
);

FILL FILL_6__12193_ (
);

FILL FILL_2__13606_ (
);

FILL FILL_0__14640_ (
);

FILL FILL_0__14220_ (
);

FILL FILL_5__11186_ (
);

FILL FILL_2__16078_ (
);

FILL FILL_4__10179_ (
);

FILL FILL_3__7703_ (
);

FILL FILL_0__9606_ (
);

FILL SFILL73720x25050 (
);

FILL FILL_5__7629_ (
);

FILL FILL_4__16405_ (
);

FILL FILL_5__7209_ (
);

FILL FILL_4__11960_ (
);

INVX1 _14769_ (
    .A(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_5254_)
);

INVX1 _14349_ (
    .A(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_4843_)
);

FILL FILL_4__11540_ (
);

FILL FILL_4__11120_ (
);

FILL FILL_3__15818_ (
);

FILL FILL_1__16012_ (
);

FILL FILL_3__10953_ (
);

FILL FILL_3__10533_ (
);

FILL FILL_6__13398_ (
);

FILL FILL_3__10113_ (
);

FILL FILL_0__15845_ (
);

INVX1 _15710_ (
    .A(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_6174_)
);

FILL FILL_0__15425_ (
);

FILL FILL_0__15005_ (
);

FILL FILL_2__8592_ (
);

FILL FILL_0__10980_ (
);

FILL FILL_0__10560_ (
);

FILL FILL_0__10140_ (
);

FILL FILL_4__8098_ (
);

FILL FILL_3__8908_ (
);

FILL FILL_5__13752_ (
);

FILL FILL_5__13332_ (
);

INVX1 _7632_ (
    .A(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_387_)
);

FILL SFILL8680x71050 (
);

INVX1 _7212_ (
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_168_)
);

FILL FILL_4__12745_ (
);

FILL FILL_4__12325_ (
);

INVX1 _10689_ (
    .A(\datapath_1.regfile_1.regOut[30] [25]),
    .Y(_1937_)
);

INVX1 _10269_ (
    .A(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_1718_)
);

FILL FILL_2__6905_ (
);

FILL FILL_3__11738_ (
);

FILL FILL_1__12772_ (
);

FILL FILL_3__11318_ (
);

FILL FILL_1__12352_ (
);

FILL FILL_2__9797_ (
);

FILL FILL_2__9377_ (
);

FILL FILL_0__11765_ (
);

FILL FILL_0__11345_ (
);

NAND2X1 _11630_ (
    .A(_2720_),
    .B(_2676_),
    .Y(_2734_)
);

OAI21X1 _11210_ (
    .A(_2319_),
    .B(_2320_),
    .C(_2328_),
    .Y(_2329_)
);

FILL FILL_5__14957_ (
);

FILL FILL_3__15991_ (
);

FILL FILL_5__14537_ (
);

FILL FILL_3__15571_ (
);

FILL FILL_5__14117_ (
);

FILL FILL_3__15151_ (
);

INVX1 _8837_ (
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_987_)
);

DFFSR _8417_ (
    .Q(\datapath_1.regfile_1.regOut[12] [11]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_718_[11])
);

FILL SFILL23960x48050 (
);

FILL FILL_1__7374_ (
);

FILL FILL_2__14984_ (
);

FILL SFILL114440x78050 (
);

FILL FILL_2__14564_ (
);

FILL FILL_2__14144_ (
);

FILL FILL_1__13977_ (
);

FILL FILL_1__13557_ (
);

FILL FILL_1__13137_ (
);

FILL SFILL94200x4050 (
);

FILL FILL_3__8661_ (
);

INVX1 _12835_ (
    .A(\datapath_1.a [4]),
    .Y(_3562_)
);

FILL FILL_3__8241_ (
);

INVX1 _12415_ (
    .A(ALUOut[24]),
    .Y(_3342_)
);

FILL FILL_5__8587_ (
);

FILL FILL_6__16329_ (
);

FILL SFILL13640x70050 (
);

FILL FILL_0__13911_ (
);

FILL FILL_3__16356_ (
);

FILL SFILL109480x50050 (
);

FILL FILL_1__8999_ (
);

FILL FILL_5__10877_ (
);

FILL FILL_1__8579_ (
);

FILL FILL_5__10037_ (
);

FILL FILL_3__11491_ (
);

FILL FILL_3__11071_ (
);

FILL FILL_2__15769_ (
);

FILL FILL_2__15349_ (
);

FILL FILL_0__16383_ (
);

FILL SFILL114440x33050 (
);

FILL FILL_2__10064_ (
);

FILL FILL_1__9940_ (
);

FILL FILL_1__9520_ (
);

FILL FILL_1__9100_ (
);

FILL FILL_3__9866_ (
);

FILL FILL_4__10811_ (
);

FILL FILL_3__9026_ (
);

FILL FILL_5__14290_ (
);

FILL SFILL74280x50050 (
);

INVX1 _8590_ (
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_863_)
);

FILL FILL_1__15703_ (
);

FILL FILL_6__7451_ (
);

DFFSR _8170_ (
    .Q(\datapath_1.regfile_1.regOut[10] [20]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_588_[20])
);

FILL FILL_6__12249_ (
);

FILL FILL_4__13283_ (
);

FILL FILL_2__7863_ (
);

FILL FILL_3__12696_ (
);

FILL FILL_2__7443_ (
);

FILL FILL_3__12276_ (
);

FILL FILL_4__7369_ (
);

FILL FILL_2__11689_ (
);

FILL FILL_2__11269_ (
);

FILL FILL_5__12603_ (
);

NAND2X1 _6903_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .Y(_67_)
);

FILL FILL_4__8730_ (
);

FILL FILL_4__8310_ (
);

FILL FILL_2__12630_ (
);

FILL FILL_5__15495_ (
);

FILL FILL_0__7689_ (
);

FILL FILL_5__15075_ (
);

FILL FILL_2__12210_ (
);

OAI21X1 _9795_ (
    .A(_1482_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1483_),
    .Y(_1433_[25])
);

FILL SFILL29160x17050 (
);

OAI21X1 _9375_ (
    .A(_1263_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1264_),
    .Y(_1238_[13])
);

FILL FILL_4__14488_ (
);

FILL FILL_1__11623_ (
);

FILL FILL_4__14068_ (
);

FILL FILL_1__11203_ (
);

FILL FILL_0__8630_ (
);

FILL FILL_2__8648_ (
);

FILL FILL_2__8228_ (
);

NOR2X1 _10901_ (
    .A(_2047_),
    .B(_2049_),
    .Y(BranchNe)
);

FILL FILL_0__10616_ (
);

FILL FILL_0__8210_ (
);

FILL FILL_1__14095_ (
);

FILL FILL_6__14815_ (
);

INVX1 _13793_ (
    .A(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_4298_)
);

FILL FILL_0__13088_ (
);

INVX8 _13373_ (
    .A(_3884__bF$buf2),
    .Y(_3885_)
);

FILL FILL_5__13808_ (
);

FILL SFILL64680x62050 (
);

FILL FILL_3__14842_ (
);

FILL FILL_3__14422_ (
);

FILL FILL_3__14002_ (
);

FILL FILL_4__9935_ (
);

FILL FILL_4__9515_ (
);

FILL FILL_2__13835_ (
);

FILL FILL_2__13415_ (
);

FILL FILL_1__12828_ (
);

FILL FILL_1__12408_ (
);

CLKBUF1 CLKBUF1_insert210 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert211 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert212 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert213 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf11)
);

FILL FILL_3__7932_ (
);

CLKBUF1 CLKBUF1_insert214 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf10)
);

FILL FILL_0__9415_ (
);

CLKBUF1 CLKBUF1_insert215 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert216 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert217 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf7)
);

FILL SFILL104360x38050 (
);

CLKBUF1 CLKBUF1_insert218 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf6)
);

FILL FILL_5__7858_ (
);

FILL FILL_5__7438_ (
);

CLKBUF1 CLKBUF1_insert219 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf5)
);

FILL FILL_4__16214_ (
);

NAND3X1 _14998_ (
    .A(_5459__bF$buf1),
    .B(_5477_),
    .C(_5476_),
    .Y(_5478_)
);

FILL FILL_6__10315_ (
);

OAI22X1 _14578_ (
    .A(_5065_),
    .B(_3890_),
    .C(_3960_),
    .D(_5066_),
    .Y(_5067_)
);

INVX1 _14158_ (
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_4656_)
);

FILL FILL_3__15627_ (
);

FILL SFILL64200x3050 (
);

FILL FILL_3__15207_ (
);

FILL FILL_1__16241_ (
);

FILL FILL112040x75050 (
);

FILL FILL_3__10762_ (
);

FILL FILL_0__15654_ (
);

FILL FILL_0__15234_ (
);

FILL FILL_3__8717_ (
);

FILL FILL_5__13981_ (
);

FILL FILL_5__13561_ (
);

FILL FILL_5__13141_ (
);

FILL FILL112440x44050 (
);

INVX1 _7861_ (
    .A(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_499_)
);

INVX1 _7441_ (
    .A(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_280_)
);

DFFSR _7021_ (
    .Q(\datapath_1.regfile_1.regOut[1] [23]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_3_[23])
);

FILL FILL_4__12974_ (
);

FILL FILL_4__12134_ (
);

INVX1 _10498_ (
    .A(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_1830_)
);

FILL SFILL114520x9050 (
);

DFFSR _10078_ (
    .Q(\datapath_1.regfile_1.regOut[25] [8]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1563_[8])
);

FILL SFILL33720x62050 (
);

FILL FILL_3__11967_ (
);

FILL FILL_3__11547_ (
);

FILL FILL_1__12581_ (
);

FILL FILL_3__11127_ (
);

FILL FILL_1__12161_ (
);

FILL FILL112040x30050 (
);

FILL FILL_0__16019_ (
);

OAI21X1 _16304_ (
    .A(_5441_),
    .B(_5535__bF$buf3),
    .C(_6752_),
    .Y(_6753_)
);

FILL FILL_0__11994_ (
);

FILL SFILL73800x58050 (
);

FILL FILL_0__11574_ (
);

FILL FILL_0__11154_ (
);

FILL FILL_5__7191_ (
);

FILL FILL_2__11901_ (
);

FILL FILL_5__14766_ (
);

FILL FILL_5__14346_ (
);

FILL FILL_3__15380_ (
);

FILL FILL_6__7927_ (
);

OAI21X1 _8646_ (
    .A(_899_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_900_),
    .Y(_848_[26])
);

OAI21X1 _8226_ (
    .A(_680_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .C(_681_),
    .Y(_653_[14])
);

FILL FILL_1__7183_ (
);

FILL FILL_4__13759_ (
);

FILL FILL_4__13339_ (
);

FILL FILL_2__14793_ (
);

FILL FILL_2__14373_ (
);

FILL FILL_1__13786_ (
);

FILL FILL_1__13366_ (
);

FILL FILL_4__14700_ (
);

FILL FILL_3__8890_ (
);

FILL FILL_0__12779_ (
);

FILL FILL_3__8470_ (
);

OAI21X1 _12644_ (
    .A(_3474_),
    .B(vdd),
    .C(_3475_),
    .Y(_3425_[25])
);

FILL FILL_0__12359_ (
);

NAND3X1 _12224_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [2]),
    .C(_3198__bF$buf4),
    .Y(_3207_)
);

FILL FILL_5__8396_ (
);

FILL SFILL94280x49050 (
);

FILL FILL_0__13720_ (
);

FILL FILL_0__13300_ (
);

FILL FILL_3__16165_ (
);

FILL FILL_5__10686_ (
);

FILL FILL_1__8388_ (
);

FILL FILL_5__10266_ (
);

FILL FILL_2__15998_ (
);

FILL FILL_0_BUFX2_insert1010 (
);

FILL FILL_0_BUFX2_insert1011 (
);

FILL FILL_2__15578_ (
);

FILL FILL_0_BUFX2_insert1012 (
);

FILL FILL_2__15158_ (
);

FILL FILL_0__16192_ (
);

FILL FILL_0_BUFX2_insert1013 (
);

FILL FILL_0_BUFX2_insert1014 (
);

FILL FILL_0_BUFX2_insert1015 (
);

FILL FILL_2__10293_ (
);

FILL FILL_0_BUFX2_insert1016 (
);

FILL FILL_0_BUFX2_insert1017 (
);

FILL FILL_0_BUFX2_insert1018 (
);

FILL FILL_0_BUFX2_insert1019 (
);

FILL FILL_4__15905_ (
);

FILL FILL_3_BUFX2_insert910 (
);

FILL FILL_3__9675_ (
);

INVX1 _13849_ (
    .A(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_4353_)
);

FILL FILL_3__9255_ (
);

FILL FILL_3_BUFX2_insert911 (
);

NAND3X1 _13429_ (
    .A(_3898_),
    .B(_3904_),
    .C(_3903_),
    .Y(_3941_)
);

FILL FILL_4__10620_ (
);

FILL FILL_3_BUFX2_insert912 (
);

NAND2X1 _13009_ (
    .A(vdd),
    .B(\datapath_1.rd2 [19]),
    .Y(_3658_)
);

FILL FILL_3_BUFX2_insert913 (
);

FILL FILL_3_BUFX2_insert914 (
);

FILL FILL_1__15932_ (
);

FILL FILL_3_BUFX2_insert915 (
);

FILL FILL_3_BUFX2_insert916 (
);

FILL FILL_1__15512_ (
);

FILL FILL_3_BUFX2_insert917 (
);

FILL FILL_3_BUFX2_insert918 (
);

FILL FILL_6__12898_ (
);

FILL FILL_3_BUFX2_insert919 (
);

FILL FILL_4__13092_ (
);

FILL FILL_0__14925_ (
);

FILL FILL_0__14505_ (
);

FILL FILL_2__7672_ (
);

FILL FILL_2__7252_ (
);

FILL FILL_3__12085_ (
);

FILL FILL_4__7598_ (
);

FILL FILL_4__7178_ (
);

FILL FILL_2__11498_ (
);

FILL FILL_2__11078_ (
);

FILL FILL_5__12832_ (
);

FILL FILL_5__12412_ (
);

FILL SFILL94600x16050 (
);

FILL FILL_4__11825_ (
);

FILL SFILL109560x83050 (
);

FILL FILL_4__11405_ (
);

FILL FILL_0__7498_ (
);

FILL FILL_0__7078_ (
);

DFFSR _9184_ (
    .Q(\datapath_1.regfile_1.regOut[18] [10]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_1108_[10])
);

FILL FILL_3__10818_ (
);

FILL FILL_1__11852_ (
);

FILL FILL_4__14297_ (
);

FILL FILL_1__11432_ (
);

FILL FILL_1__11012_ (
);

FILL SFILL84280x47050 (
);

FILL FILL_2__8877_ (
);

FILL FILL_2__8457_ (
);

DFFSR _10710_ (
    .Q(\datapath_1.regfile_1.regOut[30] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1888_[0])
);

FILL FILL_0__10425_ (
);

FILL FILL_0__10005_ (
);

FILL FILL_5__6882_ (
);

DFFSR _13182_ (
    .Q(\datapath_1.mux_iord.din0 [7]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3685_[7])
);

FILL FILL_5__13617_ (
);

FILL FILL_3__14651_ (
);

FILL SFILL8600x64050 (
);

DFFSR _7917_ (
    .Q(\datapath_1.regfile_1.regOut[8] [23]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_458_[23])
);

FILL FILL_3__14231_ (
);

FILL FILL_1__6874_ (
);

FILL FILL_4__9744_ (
);

FILL SFILL8680x21050 (
);

FILL FILL_2__13644_ (
);

FILL FILL_2__13224_ (
);

FILL FILL_5__16089_ (
);

FILL FILL_1__12637_ (
);

FILL FILL_1__12217_ (
);

FILL SFILL84200x45050 (
);

FILL SFILL23560x29050 (
);

FILL FILL_3__7741_ (
);

FILL FILL_0__9644_ (
);

FILL FILL_0__9224_ (
);

FILL FILL_3__7321_ (
);

NAND2X1 _11915_ (
    .A(IorD_bF$buf4),
    .B(ALUOut[9]),
    .Y(_2985_)
);

FILL FILL_5__7247_ (
);

FILL FILL_4__16023_ (
);

FILL FILL_6__10124_ (
);

NOR2X1 _14387_ (
    .A(_4879_),
    .B(_4876_),
    .Y(_4880_)
);

FILL FILL_3__15856_ (
);

FILL FILL_3__15436_ (
);

FILL SFILL109480x45050 (
);

FILL FILL_3__15016_ (
);

FILL FILL_1__16050_ (
);

FILL FILL_3__10991_ (
);

FILL FILL_3__10571_ (
);

FILL FILL_1__7239_ (
);

FILL FILL_3__10151_ (
);

FILL FILL_2__14849_ (
);

FILL FILL_0__15883_ (
);

FILL FILL_2__14429_ (
);

FILL FILL_6_BUFX2_insert423 (
);

FILL FILL_2__14009_ (
);

FILL FILL_0__15463_ (
);

FILL FILL_0__15043_ (
);

FILL SFILL114440x28050 (
);

FILL FILL_6_BUFX2_insert428 (
);

FILL FILL_1__8600_ (
);

FILL FILL_3__8526_ (
);

FILL FILL_3__8106_ (
);

FILL FILL_5__13790_ (
);

FILL FILL_5__13370_ (
);

FILL SFILL74280x45050 (
);

INVX1 _7670_ (
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .Y(_456_)
);

OAI21X1 _7250_ (
    .A(_192_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_193_),
    .Y(_133_[30])
);

FILL FILL_4__12783_ (
);

FILL FILL_4__12363_ (
);

FILL SFILL13640x20050 (
);

FILL FILL_2__6943_ (
);

FILL FILL_5__9813_ (
);

FILL FILL_3__11776_ (
);

FILL FILL_3__11356_ (
);

FILL FILL_1__12390_ (
);

FILL FILL_4__6869_ (
);

FILL FILL_0__16248_ (
);

OAI22X1 _16113_ (
    .A(_5221_),
    .B(_5518__bF$buf3),
    .C(_5478__bF$buf1),
    .D(_5213_),
    .Y(_6567_)
);

FILL FILL_2__10769_ (
);

FILL FILL_0__11383_ (
);

FILL FILL_1__9805_ (
);

FILL FILL_6__15582_ (
);

FILL FILL_4__7810_ (
);

FILL FILL_5__14995_ (
);

FILL FILL_5__14575_ (
);

FILL FILL_2__11710_ (
);

FILL FILL_5__14155_ (
);

FILL SFILL13560x27050 (
);

OAI21X1 _8875_ (
    .A(_1011_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .C(_1012_),
    .Y(_978_[17])
);

OAI21X1 _8455_ (
    .A(_792_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_793_),
    .Y(_783_[5])
);

DFFSR _8035_ (
    .Q(\datapath_1.regfile_1.regOut[9] [13]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_523_[13])
);

FILL FILL_4__13988_ (
);

FILL FILL_1__10703_ (
);

FILL FILL_4__13568_ (
);

FILL FILL_4__13148_ (
);

FILL FILL_2__14182_ (
);

FILL FILL_2__7728_ (
);

FILL FILL_0__7710_ (
);

FILL FILL_2__7308_ (
);

FILL FILL_1__13595_ (
);

FILL FILL_0__12588_ (
);

OAI21X1 _12873_ (
    .A(_3586_),
    .B(vdd),
    .C(_3587_),
    .Y(_3555_[16])
);

OAI21X1 _12453_ (
    .A(_3367_),
    .B(vdd),
    .C(_3368_),
    .Y(_3360_[4])
);

FILL FILL_0__12168_ (
);

AOI22X1 _12033_ (
    .A(\datapath_1.ALUResult [11]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3071_)
);

FILL FILL_3__13922_ (
);

FILL FILL_3__13502_ (
);

FILL FILL_5_BUFX2_insert440 (
);

FILL FILL_2__12915_ (
);

FILL FILL_5_BUFX2_insert441 (
);

FILL FILL_5_BUFX2_insert442 (
);

FILL FILL_5_BUFX2_insert443 (
);

FILL FILL_3__16394_ (
);

FILL FILL_5_BUFX2_insert444 (
);

FILL FILL_5_BUFX2_insert445 (
);

FILL FILL_5__10495_ (
);

FILL FILL_5_BUFX2_insert446 (
);

FILL FILL112120x63050 (
);

FILL FILL_1__8197_ (
);

FILL FILL_5_BUFX2_insert447 (
);

FILL FILL_1__11908_ (
);

FILL FILL_5_BUFX2_insert448 (
);

FILL FILL_5_BUFX2_insert449 (
);

FILL FILL_2__15387_ (
);

FILL FILL_5__16301_ (
);

FILL FILL_0__8915_ (
);

FILL FILL_5__6938_ (
);

FILL FILL_4__15714_ (
);

FILL FILL_3__9484_ (
);

OAI22X1 _13658_ (
    .A(_4165_),
    .B(_3902__bF$buf0),
    .C(_3983__bF$buf4),
    .D(_4164_),
    .Y(_4166_)
);

NAND2X1 _13238_ (
    .A(_3780_),
    .B(_3769_),
    .Y(_3781_)
);

FILL FILL_3__14707_ (
);

FILL FILL_1__15741_ (
);

FILL SFILL43720x14050 (
);

FILL FILL_1__15321_ (
);

FILL FILL_0__14734_ (
);

FILL FILL_0__14314_ (
);

FILL FILL_2__7481_ (
);

FILL FILL_2__7061_ (
);

FILL FILL_5__12641_ (
);

FILL FILL112440x39050 (
);

FILL FILL_5__12221_ (
);

INVX1 _6941_ (
    .A(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_28_)
);

FILL FILL_2_BUFX2_insert570 (
);

FILL FILL_2_BUFX2_insert571 (
);

FILL FILL_2_BUFX2_insert572 (
);

FILL FILL_2_BUFX2_insert573 (
);

FILL FILL_4__11634_ (
);

FILL FILL_2_BUFX2_insert574 (
);

FILL FILL_2_BUFX2_insert575 (
);

FILL FILL_4__11214_ (
);

FILL FILL_2_BUFX2_insert576 (
);

FILL FILL_2_BUFX2_insert577 (
);

FILL FILL_2_BUFX2_insert578 (
);

FILL FILL_1__16106_ (
);

FILL FILL_2_BUFX2_insert579 (
);

FILL FILL_3__10627_ (
);

FILL FILL_1__11661_ (
);

FILL FILL_1__11241_ (
);

FILL FILL112040x25050 (
);

FILL FILL_0__15939_ (
);

FILL FILL_0__15519_ (
);

INVX1 _15804_ (
    .A(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_6266_)
);

FILL FILL_2__8266_ (
);

FILL FILL_0__10654_ (
);

FILL FILL_3__13099_ (
);

FILL FILL_0__10234_ (
);

FILL FILL_5__13846_ (
);

FILL FILL_3__14880_ (
);

FILL FILL_5__13426_ (
);

FILL FILL_3__14460_ (
);

FILL FILL_5__13006_ (
);

FILL FILL_3__14040_ (
);

OAI21X1 _7726_ (
    .A(_428_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_429_),
    .Y(_393_[18])
);

OAI21X1 _7306_ (
    .A(_209_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_210_),
    .Y(_198_[6])
);

FILL FILL_4__9553_ (
);

FILL FILL_4__9133_ (
);

FILL FILL_4__12839_ (
);

FILL FILL_2__13873_ (
);

FILL FILL_4__12419_ (
);

FILL FILL_2__13453_ (
);

FILL FILL_2__13033_ (
);

FILL FILL_1__12866_ (
);

FILL FILL_1__12446_ (
);

FILL FILL_1__12026_ (
);

FILL FILL_3__7970_ (
);

FILL FILL_0__9873_ (
);

FILL FILL_0__11859_ (
);

FILL FILL_3__7550_ (
);

FILL FILL_0__9033_ (
);

FILL FILL_0__11439_ (
);

AOI21X1 _11724_ (
    .A(_2810_),
    .B(_2620_),
    .C(_2821_),
    .Y(_2822_)
);

FILL FILL_0__11019_ (
);

OAI21X1 _11304_ (
    .A(_2252_),
    .B(_2253_),
    .C(_2250_),
    .Y(_2423_)
);

FILL FILL_5__7476_ (
);

FILL FILL_5__7056_ (
);

FILL FILL_4__16252_ (
);

AOI22X1 _14196_ (
    .A(_3891__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [15]),
    .C(\datapath_1.regfile_1.regOut[8] [15]),
    .D(_4090_),
    .Y(_4693_)
);

FILL FILL_3__15665_ (
);

FILL FILL_3__15245_ (
);

FILL SFILL39000x4050 (
);

FILL FILL_1__7888_ (
);

FILL FILL_1__7468_ (
);

FILL FILL_3__10380_ (
);

FILL FILL_1__7048_ (
);

FILL FILL_2__14658_ (
);

FILL FILL_2__14238_ (
);

FILL FILL_0__15692_ (
);

FILL FILL_0__15272_ (
);

FILL SFILL13640x5050 (
);

FILL SFILL23720x55050 (
);

FILL FILL_1_BUFX2_insert590 (
);

FILL FILL_1_BUFX2_insert591 (
);

FILL FILL_3__8755_ (
);

FILL FILL_3__8335_ (
);

FILL FILL_1_BUFX2_insert592 (
);

DFFSR _12929_ (
    .Q(\datapath_1.a [10]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_3555_[10])
);

NAND2X1 _12509_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [23]),
    .Y(_3406_)
);

FILL FILL_1_BUFX2_insert593 (
);

FILL FILL_1_BUFX2_insert594 (
);

FILL FILL_1_BUFX2_insert595 (
);

FILL FILL_1_BUFX2_insert596 (
);

FILL FILL_1_BUFX2_insert597 (
);

FILL FILL_1_BUFX2_insert598 (
);

FILL FILL_6__11978_ (
);

FILL FILL_1_BUFX2_insert599 (
);

FILL FILL_6__11558_ (
);

FILL FILL_4__12592_ (
);

FILL FILL_4__12172_ (
);

FILL FILL_5__9622_ (
);

FILL FILL_3__11585_ (
);

FILL FILL_3__11165_ (
);

INVX1 _16342_ (
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .Y(_6782_)
);

FILL FILL_0__16057_ (
);

FILL FILL_2__10998_ (
);

FILL FILL_2__10578_ (
);

FILL FILL_2__10158_ (
);

FILL FILL_0__11192_ (
);

FILL FILL_5__11912_ (
);

FILL FILL_1__9614_ (
);

FILL SFILL109560x78050 (
);

FILL FILL_4__10905_ (
);

FILL SFILL23720x10050 (
);

FILL FILL_5__14384_ (
);

DFFSR _8684_ (
    .Q(\datapath_1.regfile_1.regOut[14] [22]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_848_[22])
);

FILL FILL_6__7545_ (
);

FILL FILL_6__7125_ (
);

NAND2X1 _8264_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_707_)
);

FILL FILL_1__10932_ (
);

FILL FILL_4__13797_ (
);

FILL FILL_1__10512_ (
);

FILL FILL_4__13377_ (
);

FILL FILL_2__7957_ (
);

BUFX2 BUFX2_insert260 (
    .A(_2344_),
    .Y(_2344__bF$buf3)
);

FILL FILL_2__7117_ (
);

BUFX2 BUFX2_insert261 (
    .A(_2344_),
    .Y(_2344__bF$buf2)
);

BUFX2 BUFX2_insert262 (
    .A(_2344_),
    .Y(_2344__bF$buf1)
);

BUFX2 BUFX2_insert263 (
    .A(_2344_),
    .Y(_2344__bF$buf0)
);

BUFX2 BUFX2_insert264 (
    .A(_5504_),
    .Y(_5504__bF$buf4)
);

BUFX2 BUFX2_insert265 (
    .A(_5504_),
    .Y(_5504__bF$buf3)
);

BUFX2 BUFX2_insert266 (
    .A(_5504_),
    .Y(_5504__bF$buf2)
);

BUFX2 BUFX2_insert267 (
    .A(_5504_),
    .Y(_5504__bF$buf1)
);

BUFX2 BUFX2_insert268 (
    .A(_5504_),
    .Y(_5504__bF$buf0)
);

DFFSR _12682_ (
    .Q(\datapath_1.Data [19]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3425_[19])
);

FILL FILL_0__12397_ (
);

BUFX2 BUFX2_insert269 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf7 )
);

NAND3X1 _12262_ (
    .A(_3233_),
    .B(_3234_),
    .C(_3235_),
    .Y(\datapath_1.alu_1.ALUInB [11])
);

FILL SFILL8600x59050 (
);

FILL FILL_3__13731_ (
);

FILL FILL_3__13311_ (
);

FILL FILL_6__16176_ (
);

FILL FILL_4__8824_ (
);

FILL FILL_4__8404_ (
);

FILL SFILL8680x16050 (
);

FILL SFILL13720x53050 (
);

FILL FILL_2__12724_ (
);

FILL FILL_5__15589_ (
);

FILL FILL_5__15169_ (
);

FILL FILL_2__12304_ (
);

FILL SFILL88600x41050 (
);

NAND2X1 _9889_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1526_)
);

NAND2X1 _9469_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1307_)
);

DFFSR _9049_ (
    .Q(\datapath_1.regfile_1.regOut[17] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_1043_[3])
);

FILL FILL_1__11717_ (
);

FILL FILL_2__15196_ (
);

FILL FILL_5__16110_ (
);

FILL FILL_0__8724_ (
);

FILL FILL_1__14189_ (
);

FILL FILL_4__15943_ (
);

FILL FILL_4__15523_ (
);

FILL FILL_4__15103_ (
);

FILL FILL_3__9293_ (
);

AOI21X1 _13887_ (
    .A(_4367_),
    .B(_4390_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [8])
);

OAI22X1 _13467_ (
    .A(_3978_),
    .B(_3975_),
    .C(_3977__bF$buf4),
    .D(_3976_),
    .Y(_3979_)
);

DFFSR _13047_ (
    .Q(_2_[0]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3620_[0])
);

FILL FILL_3__14936_ (
);

FILL FILL_1__15970_ (
);

FILL FILL_3__14516_ (
);

FILL FILL_1__15550_ (
);

FILL FILL_1__15130_ (
);

FILL FILL_4__9609_ (
);

FILL SFILL8600x14050 (
);

FILL FILL_6__12096_ (
);

FILL FILL_2__13929_ (
);

FILL FILL_0__14963_ (
);

FILL FILL_2__13509_ (
);

FILL FILL_0__14543_ (
);

FILL FILL_0__14123_ (
);

FILL FILL_2__7290_ (
);

FILL FILL_5__11089_ (
);

FILL FILL_0__9929_ (
);

FILL FILL_0__9509_ (
);

FILL FILL_3__7606_ (
);

FILL FILL_5__12870_ (
);

FILL FILL_5__12450_ (
);

FILL FILL_5__12030_ (
);

FILL FILL_4__16308_ (
);

FILL FILL_4__11863_ (
);

FILL FILL_4__11443_ (
);

FILL FILL_4__11023_ (
);

FILL SFILL13640x15050 (
);

FILL FILL_1__16335_ (
);

FILL FILL_3__10436_ (
);

FILL FILL_1__11890_ (
);

FILL FILL_3__10016_ (
);

FILL FILL_1__11470_ (
);

FILL FILL_1__11050_ (
);

FILL FILL_0__15748_ (
);

FILL FILL_0__15328_ (
);

INVX1 _15613_ (
    .A(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_6079_)
);

FILL SFILL38840x64050 (
);

FILL FILL_0__10883_ (
);

FILL FILL_2__8495_ (
);

FILL FILL_2__8075_ (
);

FILL FILL_0__10043_ (
);

FILL FILL_6__14242_ (
);

FILL SFILL43800x47050 (
);

FILL SFILL74200x38050 (
);

FILL FILL_5__13655_ (
);

FILL FILL_5__13235_ (
);

OAI21X1 _7955_ (
    .A(_540_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .C(_541_),
    .Y(_523_[9])
);

DFFSR _7535_ (
    .Q(\datapath_1.regfile_1.regOut[5] [25]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_263_[25])
);

NAND2X1 _7115_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_124_)
);

FILL FILL_4__9782_ (
);

FILL FILL_4__9362_ (
);

FILL FILL_4__12648_ (
);

FILL FILL_2__13682_ (
);

FILL FILL_4__12228_ (
);

FILL FILL_2__13262_ (
);

FILL FILL112200x51050 (
);

FILL FILL_1__12255_ (
);

FILL FILL_0__9682_ (
);

INVX1 _11953_ (
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3010_)
);

FILL FILL_0__9262_ (
);

FILL FILL_0__11668_ (
);

FILL SFILL3480x63050 (
);

FILL FILL_0__11248_ (
);

AOI21X1 _11533_ (
    .A(_2428_),
    .B(_2643_),
    .C(_2413_),
    .Y(_2644_)
);

INVX1 _11113_ (
    .A(\datapath_1.alu_1.ALUInA [20]),
    .Y(_2232_)
);

FILL FILL_4__16061_ (
);

FILL FILL_3__15894_ (
);

FILL FILL_3__15474_ (
);

FILL FILL_3__15054_ (
);

FILL SFILL78920x15050 (
);

FILL FILL112120x58050 (
);

FILL FILL_1__7697_ (
);

FILL FILL_6_BUFX2_insert802 (
);

FILL FILL_2__14887_ (
);

FILL FILL_2__14467_ (
);

FILL FILL_2__14047_ (
);

FILL FILL_0__15081_ (
);

FILL FILL_5__15801_ (
);

FILL FILL_6_BUFX2_insert807 (
);

FILL FILL_3__8984_ (
);

NAND2X1 _12738_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[14]),
    .Y(_3518_)
);

FILL FILL_3__8144_ (
);

NAND3X1 _12318_ (
    .A(_3275_),
    .B(_3276_),
    .C(_3277_),
    .Y(\datapath_1.alu_1.ALUInB [25])
);

FILL FILL_1__14821_ (
);

FILL FILL_1__14401_ (
);

FILL FILL_0__13814_ (
);

FILL FILL_3__16259_ (
);

FILL FILL_2__6981_ (
);

FILL SFILL33800x45050 (
);

FILL FILL_5__9851_ (
);

FILL SFILL64200x36050 (
);

FILL FILL_3__11394_ (
);

FILL FILL_5__9011_ (
);

FILL FILL112120x13050 (
);

FILL FILL_0__16286_ (
);

OAI22X1 _16151_ (
    .A(_6603_),
    .B(_5545__bF$buf3),
    .C(_5466__bF$buf1),
    .D(_5262_),
    .Y(_6604_)
);

FILL FILL_2__10387_ (
);

FILL FILL_5__11721_ (
);

FILL FILL_1__9423_ (
);

FILL FILL_5__11301_ (
);

FILL FILL_1__9003_ (
);

FILL SFILL68520x44050 (
);

FILL FILL_3__9769_ (
);

FILL FILL_3__9349_ (
);

FILL FILL_5__14193_ (
);

NAND2X1 _8493_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_819_)
);

FILL FILL_1__15606_ (
);

NAND2X1 _8073_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_600_)
);

FILL SFILL58600x80050 (
);

FILL SFILL113960x47050 (
);

FILL FILL_1__10321_ (
);

FILL FILL_3__12599_ (
);

FILL FILL_2__7346_ (
);

FILL FILL_3__12179_ (
);

NAND2X1 _12491_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [17]),
    .Y(_3394_)
);

NAND3X1 _12071_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[21]),
    .C(_3032__bF$buf0),
    .Y(_3099_)
);

FILL FILL_5__12506_ (
);

FILL FILL_3__13960_ (
);

FILL FILL_3__13540_ (
);

FILL FILL_3__13120_ (
);

FILL FILL_4__8633_ (
);

FILL FILL_4__11919_ (
);

FILL FILL_5_BUFX2_insert820 (
);

FILL FILL_4__8213_ (
);

FILL FILL_2__12953_ (
);

FILL FILL_5_BUFX2_insert821 (
);

FILL FILL_5__15398_ (
);

FILL FILL_2__12533_ (
);

FILL FILL_5_BUFX2_insert822 (
);

FILL FILL_5_BUFX2_insert823 (
);

FILL FILL_2__12113_ (
);

DFFSR _9698_ (
    .Q(\datapath_1.regfile_1.regOut[22] [12]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_1368_[12])
);

FILL FILL_5_BUFX2_insert824 (
);

INVX1 _9278_ (
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_1220_)
);

FILL FILL_5_BUFX2_insert825 (
);

FILL FILL_5_BUFX2_insert826 (
);

FILL FILL_5_BUFX2_insert827 (
);

FILL FILL_5_BUFX2_insert828 (
);

FILL FILL_1__11946_ (
);

FILL FILL_5_BUFX2_insert829 (
);

FILL FILL_1__11526_ (
);

FILL FILL_1__11106_ (
);

FILL FILL_0__8953_ (
);

FILL FILL_0__10939_ (
);

FILL FILL_0__8533_ (
);

FILL FILL_0__10519_ (
);

FILL FILL_0__8113_ (
);

OAI21X1 _10804_ (
    .A(_1992_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1993_),
    .Y(_1953_[20])
);

FILL FILL_5__6976_ (
);

FILL FILL_6__14718_ (
);

FILL FILL_4__15752_ (
);

FILL FILL_4__15332_ (
);

FILL SFILL54200x34050 (
);

OAI22X1 _13696_ (
    .A(_4201_),
    .B(_3893__bF$buf0),
    .C(_3966__bF$buf2),
    .D(_4202_),
    .Y(_4203_)
);

NOR2X1 _13276_ (
    .A(_3781_),
    .B(_3816_),
    .Y(\datapath_1.regfile_1.regEn [3])
);

FILL FILL_2__9912_ (
);

FILL FILL_3__14745_ (
);

FILL FILL_3__14325_ (
);

FILL FILL_1__6968_ (
);

FILL FILL_4__9418_ (
);

FILL FILL_2__13738_ (
);

FILL FILL_2__13318_ (
);

FILL FILL_0__14772_ (
);

FILL FILL_0__14352_ (
);

FILL FILL_0__9738_ (
);

FILL FILL_3__7835_ (
);

FILL FILL_3__7415_ (
);

FILL FILL_2_BUFX2_insert950 (
);

FILL FILL_2_BUFX2_insert951 (
);

FILL FILL_4__16117_ (
);

FILL FILL_2_BUFX2_insert952 (
);

FILL FILL_2_BUFX2_insert953 (
);

FILL FILL_2_BUFX2_insert954 (
);

FILL FILL_4__11672_ (
);

FILL FILL_2_BUFX2_insert955 (
);

FILL FILL_4__11252_ (
);

FILL FILL_2_BUFX2_insert956 (
);

FILL FILL_2_BUFX2_insert957 (
);

FILL FILL_2_BUFX2_insert958 (
);

FILL FILL_1__16144_ (
);

FILL FILL_2_BUFX2_insert959 (
);

FILL FILL_3__10665_ (
);

FILL FILL_5__8702_ (
);

FILL FILL_3__10245_ (
);

FILL FILL_0__15977_ (
);

FILL FILL_0__15557_ (
);

OAI22X1 _15842_ (
    .A(_5463__bF$buf2),
    .B(_4861_),
    .C(_4864_),
    .D(_5495__bF$buf3),
    .Y(_6303_)
);

FILL FILL_0__15137_ (
);

INVX1 _15422_ (
    .A(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_5893_)
);

AOI22X1 _15002_ (
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [0]),
    .C(\datapath_1.regfile_1.regOut[30] [0]),
    .D(_5481_),
    .Y(_5482_)
);

FILL FILL_0__10692_ (
);

FILL FILL_0__10272_ (
);

FILL FILL_5__13884_ (
);

FILL FILL_5__13464_ (
);

FILL FILL_5__13044_ (
);

NAND2X1 _7764_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_455_)
);

NAND2X1 _7344_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_236_)
);

FILL FILL_4__9591_ (
);

FILL FILL_4__12877_ (
);

FILL FILL_4__9171_ (
);

FILL FILL_4__12457_ (
);

FILL SFILL48920x54050 (
);

FILL FILL_4__12037_ (
);

FILL FILL_2__13491_ (
);

FILL SFILL13320x79050 (
);

FILL SFILL109640x21050 (
);

FILL FILL_5__9907_ (
);

FILL FILL_1__12484_ (
);

FILL FILL_1__12064_ (
);

INVX1 _16207_ (
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_6658_)
);

FILL FILL_0__11897_ (
);

FILL FILL_0__9491_ (
);

FILL FILL_2__9089_ (
);

OR2X2 _11762_ (
    .A(_2856_),
    .B(_2337_),
    .Y(_2857_)
);

FILL FILL_0__11477_ (
);

NAND3X1 _11342_ (
    .A(_2349_),
    .B(_2460_),
    .C(_2339_),
    .Y(\datapath_1.ALUResult [31])
);

FILL FILL_0__11057_ (
);

FILL SFILL48520x40050 (
);

FILL SFILL38840x50 (
);

FILL FILL_5__7094_ (
);

FILL FILL_4__16290_ (
);

FILL SFILL13720x48050 (
);

FILL FILL_2__11804_ (
);

FILL FILL_5__14669_ (
);

FILL FILL_5__14249_ (
);

NAND2X1 _8969_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1055_)
);

FILL FILL_3__15283_ (
);

DFFSR _8549_ (
    .Q(\datapath_1.regfile_1.regOut[13] [15]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_783_[15])
);

INVX1 _8129_ (
    .A(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_637_)
);

FILL FILL_1__7086_ (
);

FILL FILL_2__14696_ (
);

FILL FILL_2__14276_ (
);

FILL FILL_5__15610_ (
);

FILL FILL_0__7804_ (
);

NAND2X1 _9910_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1540_)
);

FILL FILL_1__13689_ (
);

FILL FILL_1__13269_ (
);

FILL FILL_4__14603_ (
);

FILL FILL_1_BUFX2_insert970 (
);

FILL FILL_1_BUFX2_insert971 (
);

FILL FILL_3__8373_ (
);

FILL FILL_1_BUFX2_insert972 (
);

NAND2X1 _12967_ (
    .A(vdd),
    .B(\datapath_1.rd2 [5]),
    .Y(_3630_)
);

FILL FILL_1_BUFX2_insert973 (
);

DFFSR _12547_ (
    .Q(ALUOut[12]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3360_[12])
);

FILL FILL_1_BUFX2_insert974 (
);

INVX1 _12127_ (
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_3138_)
);

FILL FILL_1_BUFX2_insert975 (
);

FILL FILL_1_BUFX2_insert976 (
);

FILL FILL_1__14630_ (
);

FILL FILL_1_BUFX2_insert977 (
);

FILL FILL_1__14210_ (
);

FILL FILL_1_BUFX2_insert978 (
);

FILL FILL_1_BUFX2_insert979 (
);

FILL FILL_0__13623_ (
);

FILL FILL_3__16068_ (
);

FILL FILL_5__9660_ (
);

FILL FILL_5__10169_ (
);

FILL FILL_5__9240_ (
);

FILL FILL_0__16095_ (
);

OAI21X1 _16380_ (
    .A(_6806_),
    .B(gnd),
    .C(_6807_),
    .Y(_6769_[19])
);

FILL FILL_2__10196_ (
);

FILL FILL_5__11950_ (
);

FILL FILL_1__9652_ (
);

FILL FILL_5__11530_ (
);

FILL FILL_1__9232_ (
);

FILL FILL_5__11110_ (
);

FILL FILL_4__15808_ (
);

FILL FILL_3__9998_ (
);

FILL FILL_2__16002_ (
);

FILL FILL_4__10943_ (
);

FILL FILL_3__9158_ (
);

FILL FILL_4__10523_ (
);

FILL FILL_4__10103_ (
);

FILL FILL_1__15835_ (
);

FILL FILL_1__15415_ (
);

FILL FILL_1__10970_ (
);

FILL FILL_1__10550_ (
);

FILL FILL_1__10130_ (
);

FILL FILL_0__14828_ (
);

FILL FILL_0__14408_ (
);

FILL SFILL38840x59050 (
);

FILL FILL_2__7995_ (
);

FILL FILL_2__7575_ (
);

BUFX2 BUFX2_insert640 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf1 )
);

BUFX2 BUFX2_insert641 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf0 )
);

BUFX2 BUFX2_insert642 (
    .A(_3936_),
    .Y(_3936__bF$buf4)
);

BUFX2 BUFX2_insert643 (
    .A(_3936_),
    .Y(_3936__bF$buf3)
);

BUFX2 BUFX2_insert644 (
    .A(_3936_),
    .Y(_3936__bF$buf2)
);

BUFX2 BUFX2_insert645 (
    .A(_3936_),
    .Y(_3936__bF$buf1)
);

BUFX2 BUFX2_insert646 (
    .A(_3936_),
    .Y(_3936__bF$buf0)
);

BUFX2 BUFX2_insert647 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf4)
);

BUFX2 BUFX2_insert648 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf3)
);

BUFX2 BUFX2_insert649 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf2)
);

FILL SFILL3560x51050 (
);

FILL FILL_5__12735_ (
);

FILL FILL_5__12315_ (
);

FILL FILL_4__8862_ (
);

FILL FILL_4__8442_ (
);

FILL FILL_4__11728_ (
);

FILL FILL_2__12762_ (
);

FILL FILL_4__11308_ (
);

FILL FILL_2__12342_ (
);

INVX1 _9087_ (
    .A(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_1113_)
);

FILL FILL112200x46050 (
);

FILL FILL_1__11755_ (
);

FILL FILL_1__11335_ (
);

FILL FILL_0__8762_ (
);

FILL SFILL3480x58050 (
);

FILL FILL_0__10748_ (
);

FILL FILL_0__8342_ (
);

DFFSR _10613_ (
    .Q(\datapath_1.regfile_1.regOut[29] [31]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_1823_[31])
);

FILL SFILL38840x14050 (
);

FILL FILL_4__15981_ (
);

FILL FILL_4__15561_ (
);

FILL FILL_4__15141_ (
);

INVX1 _13085_ (
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_3688_)
);

FILL FILL_3__14974_ (
);

FILL FILL_2__9721_ (
);

FILL FILL_3__14554_ (
);

FILL FILL_2__9301_ (
);

FILL FILL_3__14134_ (
);

FILL FILL_4_BUFX2_insert480 (
);

FILL FILL_4_BUFX2_insert481 (
);

FILL FILL_4__9647_ (
);

FILL FILL_4__9227_ (
);

FILL FILL_4_BUFX2_insert482 (
);

FILL FILL_4_BUFX2_insert483 (
);

FILL FILL_2__13967_ (
);

FILL FILL_2__13547_ (
);

FILL FILL_4_BUFX2_insert484 (
);

FILL FILL_0__14581_ (
);

FILL FILL_2__13127_ (
);

FILL FILL_4_BUFX2_insert485 (
);

FILL FILL_0__14161_ (
);

FILL FILL_4_BUFX2_insert486 (
);

FILL FILL_4_BUFX2_insert487 (
);

FILL FILL_4_BUFX2_insert488 (
);

FILL FILL_4_BUFX2_insert489 (
);

FILL FILL_0__9547_ (
);

FILL FILL_0__9127_ (
);

FILL FILL_3__7224_ (
);

OAI21X1 _11818_ (
    .A(_2124_),
    .B(_2907_),
    .C(_2908_),
    .Y(_2909_)
);

FILL SFILL28840x57050 (
);

FILL FILL_1__13901_ (
);

FILL FILL_4__16346_ (
);

FILL FILL_4__11481_ (
);

FILL FILL_4__11061_ (
);

FILL FILL_3__15759_ (
);

FILL FILL_3__15339_ (
);

FILL FILL_1__16373_ (
);

FILL FILL_3__10894_ (
);

FILL FILL_5__8511_ (
);

FILL FILL_3__10054_ (
);

FILL FILL_0__15786_ (
);

FILL SFILL28440x43050 (
);

FILL FILL_0__15366_ (
);

AOI21X1 _15651_ (
    .A(_6095_),
    .B(_6116_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [14])
);

NAND2X1 _15231_ (
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .B(_5649_),
    .Y(_5707_)
);

FILL FILL_5__10801_ (
);

FILL FILL_1__8503_ (
);

FILL SFILL115000x34050 (
);

FILL FILL_3__8849_ (
);

FILL FILL_3__8009_ (
);

FILL FILL_5__13693_ (
);

FILL FILL_5__13273_ (
);

NAND2X1 _7993_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_567_)
);

NAND2X1 _7573_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_348_)
);

DFFSR _7153_ (
    .Q(\datapath_1.regfile_1.regOut[2] [27]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_68_[27])
);

FILL FILL_4__12266_ (
);

FILL FILL_2__6846_ (
);

FILL FILL_3__11679_ (
);

FILL FILL_3__11259_ (
);

FILL FILL_1__12293_ (
);

DFFSR _16436_ (
    .Q(\datapath_1.regfile_1.regOut[0] [19]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_6769_[19])
);

OAI22X1 _16016_ (
    .A(_6471_),
    .B(_5545__bF$buf1),
    .C(_5569_),
    .D(_5119_),
    .Y(_6472_)
);

NAND3X1 _11991_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[1]),
    .C(_3032__bF$buf1),
    .Y(_3039_)
);

NAND2X1 _11571_ (
    .A(_2462__bF$buf1),
    .B(_2671_),
    .Y(_2679_)
);

FILL FILL_0__11286_ (
);

NAND2X1 _11151_ (
    .A(_2269_),
    .B(_2265_),
    .Y(_2270_)
);

FILL FILL_3__12620_ (
);

FILL FILL_6__15485_ (
);

FILL FILL_3__12200_ (
);

FILL FILL_4__7713_ (
);

FILL FILL_5__14898_ (
);

FILL FILL_5__14478_ (
);

FILL FILL_2__11613_ (
);

FILL FILL_5__14058_ (
);

INVX1 _8778_ (
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_968_)
);

FILL FILL_3__15092_ (
);

INVX1 _8358_ (
    .A(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_749_)
);

FILL SFILL18840x55050 (
);

FILL FILL_2__14085_ (
);

FILL FILL_0__7613_ (
);

FILL FILL_1__13498_ (
);

FILL FILL_4__14832_ (
);

FILL FILL_4__14412_ (
);

INVX1 _12776_ (
    .A(\control_1.op [1]),
    .Y(_3543_)
);

FILL FILL_3__8182_ (
);

NAND2X1 _12356_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [4]),
    .Y(_3303_)
);

FILL FILL_3__13825_ (
);

FILL FILL_3__13405_ (
);

FILL FILL_0__13852_ (
);

FILL FILL_0__13432_ (
);

FILL FILL_3__16297_ (
);

FILL FILL_0__13012_ (
);

FILL FILL_5__10398_ (
);

FILL FILL_5__16204_ (
);

FILL FILL_3__6915_ (
);

FILL SFILL18840x10050 (
);

FILL FILL_1__9881_ (
);

FILL FILL_1__9041_ (
);

FILL SFILL79080x21050 (
);

FILL FILL_4__15617_ (
);

FILL FILL_2__16231_ (
);

FILL FILL_3__9387_ (
);

FILL FILL_4__10752_ (
);

FILL FILL_1__15644_ (
);

FILL FILL_1__15224_ (
);

FILL FILL_0__14637_ (
);

INVX1 _14922_ (
    .A(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_5404_)
);

FILL FILL_0__14217_ (
);

INVX1 _14502_ (
    .A(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_4992_)
);

FILL FILL_6__13971_ (
);

FILL FILL_6__13551_ (
);

FILL FILL_5__12964_ (
);

FILL FILL_5__12124_ (
);

BUFX2 _6844_ (
    .A(_1_[6]),
    .Y(memoryAddress[6])
);

FILL SFILL69080x64050 (
);

FILL FILL_4__8251_ (
);

FILL FILL_4__11957_ (
);

FILL SFILL48920x49050 (
);

FILL SFILL99320x4050 (
);

FILL FILL_2__12991_ (
);

FILL FILL_4__11537_ (
);

FILL FILL_2__12571_ (
);

FILL FILL_4__11117_ (
);

FILL FILL_2__12151_ (
);

FILL SFILL109640x16050 (
);

FILL FILL_1__16009_ (
);

FILL FILL_1__11984_ (
);

FILL FILL_1__11564_ (
);

FILL FILL_1__11144_ (
);

INVX1 _15707_ (
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_6171_)
);

FILL FILL_0__8991_ (
);

FILL FILL_2__8589_ (
);

FILL FILL_0__10977_ (
);

FILL FILL_0__8571_ (
);

FILL FILL_0__10557_ (
);

DFFSR _10842_ (
    .Q(\datapath_1.regfile_1.regOut[31] [4]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_1953_[4])
);

FILL SFILL48520x35050 (
);

NAND2X1 _10422_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1800_)
);

FILL FILL_0__10137_ (
);

NAND2X1 _10002_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1581_)
);

FILL FILL_4__15790_ (
);

FILL FILL_4__15370_ (
);

FILL FILL_5__13749_ (
);

FILL FILL_5__13329_ (
);

FILL FILL_2__9530_ (
);

FILL FILL_3__14783_ (
);

FILL FILL_3__14363_ (
);

FILL FILL_2__9110_ (
);

INVX1 _7629_ (
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_385_)
);

INVX1 _7209_ (
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_166_)
);

FILL FILL_4__9876_ (
);

FILL FILL_4__9036_ (
);

FILL FILL_2__13776_ (
);

FILL FILL_2__13356_ (
);

FILL FILL_0__14390_ (
);

FILL FILL_1__12769_ (
);

FILL FILL_1__12349_ (
);

FILL FILL_0__9776_ (
);

FILL FILL_3__7873_ (
);

FILL FILL_0__9356_ (
);

FILL FILL_3__7453_ (
);

OAI21X1 _11627_ (
    .A(_2730_),
    .B(_2731_),
    .C(_2727_),
    .Y(_2732_)
);

FILL FILL_3__7033_ (
);

AOI21X1 _11207_ (
    .A(_2316_),
    .B(_2304_),
    .C(_2325_),
    .Y(_2326_)
);

FILL FILL_5__7799_ (
);

FILL FILL_5__7379_ (
);

FILL FILL_1__13710_ (
);

FILL FILL_4__16155_ (
);

INVX1 _14099_ (
    .A(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_4598_)
);

FILL FILL_4__11290_ (
);

FILL FILL_3__15988_ (
);

FILL FILL_0__12703_ (
);

FILL FILL_3__15568_ (
);

FILL FILL_3__15148_ (
);

FILL FILL_1__16182_ (
);

FILL FILL_5__8740_ (
);

FILL FILL_5__8320_ (
);

FILL FILL_3__10283_ (
);

INVX1 _15880_ (
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_6340_)
);

FILL FILL_0__15595_ (
);

FILL FILL_0__15175_ (
);

NOR3X1 _15460_ (
    .A(_5929_),
    .B(_5509_),
    .C(_5688_),
    .Y(_5930_)
);

OAI21X1 _15040_ (
    .A(_5519_),
    .B(\datapath_1.PCJump_27_bF$buf4 ),
    .C(_5518__bF$buf2),
    .Y(_5520_)
);

FILL SFILL38920x47050 (
);

FILL FILL_1__8732_ (
);

FILL FILL_1__8312_ (
);

FILL FILL_2__15922_ (
);

FILL FILL_2__15502_ (
);

FILL FILL_3__8658_ (
);

FILL FILL_3__8238_ (
);

FILL FILL_5__13082_ (
);

FILL FILL_1__14915_ (
);

DFFSR _7382_ (
    .Q(\datapath_1.regfile_1.regOut[4] [0]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_198_[0])
);

FILL FILL_4__12495_ (
);

FILL FILL_4__12075_ (
);

FILL FILL_0__13908_ (
);

FILL FILL_5__9525_ (
);

FILL FILL_3__11488_ (
);

FILL FILL_5__9105_ (
);

FILL FILL_3__11068_ (
);

FILL SFILL59000x60050 (
);

NAND2X1 _16245_ (
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .B(_5570__bF$buf1),
    .Y(_6695_)
);

FILL SFILL3560x46050 (
);

INVX1 _11380_ (
    .A(_2140_),
    .Y(_2497_)
);

FILL FILL_0__11095_ (
);

FILL FILL_1__9937_ (
);

FILL FILL_5__11815_ (
);

FILL FILL_1__9517_ (
);

FILL SFILL104440x63050 (
);

FILL FILL_4__7942_ (
);

FILL FILL_4__7102_ (
);

FILL FILL_4__10808_ (
);

FILL FILL_2__11842_ (
);

FILL FILL_5__14287_ (
);

FILL FILL_2__11422_ (
);

FILL FILL_2__11002_ (
);

INVX1 _8587_ (
    .A(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_861_)
);

DFFSR _8167_ (
    .Q(\datapath_1.regfile_1.regOut[10] [17]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_588_[17])
);

FILL FILL_1__10835_ (
);

FILL FILL_1__10415_ (
);

FILL FILL_0__7842_ (
);

FILL FILL_0__7422_ (
);

FILL FILL_4__14641_ (
);

FILL FILL_4__14221_ (
);

FILL SFILL69240x8050 (
);

INVX1 _12585_ (
    .A(\datapath_1.Data [6]),
    .Y(_3436_)
);

FILL SFILL49080x60050 (
);

OAI21X1 _12165_ (
    .A(_3162_),
    .B(ALUSrcA_bF$buf2),
    .C(_3163_),
    .Y(\datapath_1.alu_1.ALUInA [16])
);

FILL FILL_3__13634_ (
);

FILL FILL_3__13214_ (
);

FILL FILL_4__8727_ (
);

FILL FILL_2__12627_ (
);

FILL FILL_0__13661_ (
);

FILL FILL_2__12207_ (
);

FILL FILL_0__13241_ (
);

FILL FILL_2__15099_ (
);

FILL FILL_5__16013_ (
);

FILL FILL_0__8627_ (
);

FILL FILL_0__8207_ (
);

FILL FILL_1__9270_ (
);

FILL FILL_4__15846_ (
);

FILL FILL_4__15426_ (
);

FILL FILL_4__15006_ (
);

FILL FILL_2__16040_ (
);

FILL FILL_4__10981_ (
);

FILL FILL_4__10561_ (
);

FILL FILL_4__10141_ (
);

FILL FILL_3__14839_ (
);

FILL FILL_3__14419_ (
);

FILL FILL_1__15873_ (
);

FILL FILL_1__15453_ (
);

FILL FILL_1__15033_ (
);

FILL FILL_0__14866_ (
);

INVX1 _14731_ (
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_5217_)
);

FILL FILL_0__14446_ (
);

FILL FILL_0__14026_ (
);

NOR2X1 _14311_ (
    .A(_4793_),
    .B(_4805_),
    .Y(_4806_)
);

FILL SFILL89160x11050 (
);

FILL FILL_2__7193_ (
);

CLKBUF1 CLKBUF1_insert180 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert181 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert182 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert183 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf41)
);

FILL FILL_3__7929_ (
);

CLKBUF1 CLKBUF1_insert184 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf40)
);

FILL FILL_3__7509_ (
);

CLKBUF1 CLKBUF1_insert185 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf39)
);

FILL FILL_5__12773_ (
);

CLKBUF1 CLKBUF1_insert186 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert187 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf37)
);

FILL FILL_5__12353_ (
);

CLKBUF1 CLKBUF1_insert188 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert189 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf35)
);

FILL FILL_4__8480_ (
);

FILL SFILL63960x83050 (
);

FILL FILL_4__11766_ (
);

FILL FILL_4__8060_ (
);

FILL SFILL94360x74050 (
);

FILL FILL_4__11346_ (
);

FILL FILL_2__12380_ (
);

FILL FILL_1__16238_ (
);

FILL FILL_3__10759_ (
);

FILL FILL_1__11793_ (
);

FILL FILL_1__11373_ (
);

NAND3X1 _15936_ (
    .A(_6392_),
    .B(_6393_),
    .C(_6391_),
    .Y(_6394_)
);

INVX1 _15516_ (
    .A(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_5985_)
);

FILL FILL_0__8380_ (
);

FILL FILL_2__8398_ (
);

FILL FILL_0__10786_ (
);

FILL SFILL79160x54050 (
);

NAND2X1 _10651_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1912_)
);

FILL FILL_0__10366_ (
);

NAND2X1 _10231_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .Y(_1757_)
);

FILL FILL_3__11700_ (
);

FILL FILL_6__14145_ (
);

FILL FILL_5__13978_ (
);

FILL FILL_5__13558_ (
);

FILL FILL_3__14592_ (
);

FILL FILL_5__13138_ (
);

FILL FILL_3__14172_ (
);

INVX1 _7858_ (
    .A(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_497_)
);

INVX1 _7438_ (
    .A(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_278_)
);

FILL FILL_4_BUFX2_insert860 (
);

DFFSR _7018_ (
    .Q(\datapath_1.regfile_1.regOut[1] [20]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_3_[20])
);

FILL FILL_4__9685_ (
);

FILL FILL_4_BUFX2_insert861 (
);

FILL FILL_4_BUFX2_insert862 (
);

FILL FILL_4__9265_ (
);

FILL FILL_4_BUFX2_insert863 (
);

FILL FILL_2__13585_ (
);

FILL FILL_4_BUFX2_insert864 (
);

FILL FILL_2__13165_ (
);

FILL FILL_4_BUFX2_insert865 (
);

FILL FILL_4_BUFX2_insert866 (
);

FILL FILL_4_BUFX2_insert867 (
);

FILL FILL_4_BUFX2_insert868 (
);

FILL FILL_4_BUFX2_insert869 (
);

FILL FILL_1__12998_ (
);

FILL FILL_1__12578_ (
);

FILL FILL_1__12158_ (
);

FILL FILL_4__13912_ (
);

FILL FILL_3__7682_ (
);

FILL FILL_0__9165_ (
);

OR2X2 _11856_ (
    .A(_2661_),
    .B(_2662_),
    .Y(_2943_)
);

INVX2 _11436_ (
    .A(_2431_),
    .Y(_2552_)
);

OAI21X1 _11016_ (
    .A(_2131_),
    .B(_2127_),
    .C(_2134_),
    .Y(_2135_)
);

FILL FILL_3__12905_ (
);

FILL FILL_4__16384_ (
);

FILL FILL_5__7188_ (
);

FILL FILL111720x65050 (
);

FILL FILL_3__15797_ (
);

FILL FILL_3__15377_ (
);

FILL FILL_0__12512_ (
);

FILL FILL_5__15704_ (
);

FILL SFILL53960x81050 (
);

FILL FILL_1__8961_ (
);

FILL SFILL79080x16050 (
);

FILL FILL_1__8121_ (
);

FILL FILL_2__15731_ (
);

FILL FILL_2__15311_ (
);

FILL FILL_3__8887_ (
);

FILL FILL_3__8467_ (
);

FILL FILL_1__14724_ (
);

INVX1 _7191_ (
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_154_)
);

FILL FILL_1__14304_ (
);

FILL FILL_0__13717_ (
);

FILL FILL_2__6884_ (
);

FILL FILL_5__9754_ (
);

FILL FILL_5__9334_ (
);

FILL FILL_3__11297_ (
);

FILL SFILL78360x6050 (
);

FILL FILL_0__16189_ (
);

INVX1 _16054_ (
    .A(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_6509_)
);

FILL FILL_1__9746_ (
);

FILL FILL_5__11624_ (
);

FILL FILL_5__11204_ (
);

FILL SFILL53480x74050 (
);

FILL FILL_3_BUFX2_insert880 (
);

FILL FILL_4__7751_ (
);

FILL FILL_4__7331_ (
);

FILL FILL_3_BUFX2_insert881 (
);

FILL FILL_3_BUFX2_insert882 (
);

FILL FILL_4__10617_ (
);

FILL FILL_3_BUFX2_insert883 (
);

FILL FILL_2__11651_ (
);

FILL FILL_3_BUFX2_insert884 (
);

FILL FILL_2__11231_ (
);

FILL FILL_5__14096_ (
);

FILL FILL_1__15929_ (
);

FILL FILL_3_BUFX2_insert885 (
);

OAI21X1 _8396_ (
    .A(_773_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .C(_774_),
    .Y(_718_[28])
);

FILL FILL_3_BUFX2_insert886 (
);

FILL FILL_1__15509_ (
);

FILL FILL_3_BUFX2_insert887 (
);

FILL FILL_3_BUFX2_insert888 (
);

FILL FILL_3_BUFX2_insert889 (
);

FILL FILL_1__10644_ (
);

FILL FILL_4__13089_ (
);

FILL FILL_0__7231_ (
);

FILL FILL_2__7249_ (
);

FILL SFILL114520x53050 (
);

FILL FILL_4__14870_ (
);

FILL FILL_4__14450_ (
);

FILL FILL_4__14030_ (
);

INVX1 _12394_ (
    .A(ALUOut[17]),
    .Y(_3328_)
);

FILL FILL_5__12829_ (
);

FILL FILL_3__13863_ (
);

FILL FILL_5__12409_ (
);

FILL FILL_2__8610_ (
);

FILL FILL_3__13443_ (
);

FILL FILL_3__13023_ (
);

FILL SFILL74360x70050 (
);

FILL FILL_4__8956_ (
);

FILL FILL_4__8116_ (
);

FILL SFILL69080x14050 (
);

FILL FILL_2__12856_ (
);

FILL FILL_2__12436_ (
);

FILL FILL_0__13890_ (
);

FILL FILL_2__12016_ (
);

FILL FILL_0__13470_ (
);

FILL FILL_1__11849_ (
);

FILL FILL_1__11429_ (
);

FILL FILL_1__11009_ (
);

FILL SFILL3640x79050 (
);

FILL FILL_5__16242_ (
);

FILL FILL_0__8856_ (
);

FILL FILL_3__6953_ (
);

INVX1 _10707_ (
    .A(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_1949_)
);

FILL FILL_0__8016_ (
);

FILL FILL_5__6879_ (
);

FILL FILL_4__15655_ (
);

FILL FILL_4__15235_ (
);

INVX1 _13599_ (
    .A(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_4108_)
);

FILL FILL_4__10790_ (
);

FILL FILL_4__10370_ (
);

DFFSR _13179_ (
    .Q(\datapath_1.mux_iord.din0 [4]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3685_[4])
);

FILL FILL_3__14648_ (
);

FILL FILL_1__15682_ (
);

FILL FILL_3__14228_ (
);

FILL FILL_1__15262_ (
);

FILL FILL_5__7820_ (
);

INVX1 _14960_ (
    .A(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_5441_)
);

FILL FILL_0__14675_ (
);

FILL FILL_0__14255_ (
);

INVX1 _14540_ (
    .A(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_5030_)
);

NAND3X1 _14120_ (
    .A(_4608_),
    .B(_4611_),
    .C(_4618_),
    .Y(_4619_)
);

FILL FILL_1__7812_ (
);

FILL FILL_3__7738_ (
);

FILL FILL_3__7318_ (
);

FILL SFILL3640x34050 (
);

FILL FILL_5__12582_ (
);

FILL FILL_5__12162_ (
);

BUFX2 _6882_ (
    .A(_2_[12]),
    .Y(memoryWriteData[12])
);

FILL SFILL104520x51050 (
);

FILL SFILL43880x41050 (
);

FILL FILL_4__11995_ (
);

FILL FILL_4__11575_ (
);

FILL FILL_4__11155_ (
);

FILL FILL_1__16047_ (
);

FILL FILL_3__10988_ (
);

FILL FILL_3__10568_ (
);

FILL FILL_5__8605_ (
);

FILL SFILL49080x3050 (
);

FILL FILL_3__10148_ (
);

FILL SFILL59000x55050 (
);

FILL FILL_1__11182_ (
);

FILL FILL_6_BUFX2_insert393 (
);

NAND3X1 _15745_ (
    .A(_6205_),
    .B(_6207_),
    .C(_6206_),
    .Y(_6208_)
);

NAND3X1 _15325_ (
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5799_)
);

FILL SFILL59080x12050 (
);

FILL FILL_6_BUFX2_insert398 (
);

NOR2X1 _10880_ (
    .A(_2027_),
    .B(_2026_),
    .Y(_2028_)
);

FILL FILL_0__10175_ (
);

DFFSR _10460_ (
    .Q(\datapath_1.regfile_1.regOut[28] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_1758_[6])
);

INVX1 _10040_ (
    .A(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_1606_)
);

FILL FILL_6__14794_ (
);

FILL SFILL104440x58050 (
);

FILL FILL_0__16401_ (
);

FILL FILL_2__10922_ (
);

FILL FILL_5__13787_ (
);

FILL FILL_5__13367_ (
);

FILL FILL_2__10502_ (
);

DFFSR _7667_ (
    .Q(\datapath_1.regfile_1.regOut[6] [29]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_328_[29])
);

OAI21X1 _7247_ (
    .A(_190_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .C(_191_),
    .Y(_133_[29])
);

FILL FILL_4__9494_ (
);

FILL SFILL108760x66050 (
);

FILL FILL_2__13394_ (
);

FILL FILL_0__6922_ (
);

FILL FILL_1__12387_ (
);

FILL FILL_4__13721_ (
);

FILL FILL_4__13301_ (
);

FILL SFILL59000x10050 (
);

FILL FILL_0__9394_ (
);

FILL FILL_3__7491_ (
);

FILL SFILL49080x55050 (
);

FILL FILL_3__7071_ (
);

NOR3X1 _11665_ (
    .A(_2337_),
    .B(_2744_),
    .C(_2766_),
    .Y(_2767_)
);

XOR2X1 _11245_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2364_)
);

FILL FILL_3__12714_ (
);

FILL FILL_4__16193_ (
);

FILL FILL_4__7807_ (
);

FILL FILL_2__11707_ (
);

FILL FILL_0__12741_ (
);

FILL FILL_3__15186_ (
);

FILL FILL_0__12321_ (
);

FILL FILL_2__14599_ (
);

FILL FILL_2__14179_ (
);

FILL FILL_5__15933_ (
);

FILL FILL_5__15513_ (
);

FILL FILL_0__7707_ (
);

OAI21X1 _9813_ (
    .A(_1494_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .C(_1495_),
    .Y(_1433_[31])
);

FILL FILL_1__8770_ (
);

FILL FILL_1__8350_ (
);

FILL FILL_4__14926_ (
);

FILL FILL_2__15960_ (
);

FILL FILL_4__14506_ (
);

FILL FILL_2__15540_ (
);

FILL FILL_3__8696_ (
);

FILL FILL_2__15120_ (
);

FILL SFILL49000x53050 (
);

FILL FILL_3__8276_ (
);

FILL FILL_3__13919_ (
);

FILL FILL_1__14953_ (
);

FILL FILL_1__14533_ (
);

FILL SFILL49080x10050 (
);

FILL FILL_1__14113_ (
);

FILL SFILL94440x62050 (
);

FILL FILL_0__13946_ (
);

INVX1 _13811_ (
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_4316_)
);

FILL FILL_0__13526_ (
);

FILL FILL_0__13106_ (
);

FILL FILL_5__9983_ (
);

FILL FILL_5__9143_ (
);

AOI21X1 _16283_ (
    .A(_6709_),
    .B(_6732_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [30])
);

FILL SFILL23880x82050 (
);

FILL FILL_1__9975_ (
);

FILL FILL_5__11853_ (
);

FILL FILL_1__9555_ (
);

FILL FILL_5__11433_ (
);

FILL FILL_1__9135_ (
);

FILL FILL_5__11013_ (
);

FILL FILL_4__7980_ (
);

FILL FILL_2__16325_ (
);

FILL FILL_4__7560_ (
);

FILL SFILL94360x69050 (
);

FILL SFILL94840x31050 (
);

FILL FILL_2__11880_ (
);

FILL FILL_4__10426_ (
);

FILL FILL_2__11460_ (
);

FILL FILL_4__10006_ (
);

FILL FILL_2__11040_ (
);

FILL FILL_1__15738_ (
);

FILL FILL_1__15318_ (
);

FILL FILL_1__10873_ (
);

FILL FILL_1__10453_ (
);

FILL FILL_1__10033_ (
);

FILL FILL_0__7880_ (
);

FILL FILL_2__7478_ (
);

FILL FILL_0__7460_ (
);

FILL FILL_0__7040_ (
);

FILL FILL_2__7058_ (
);

FILL SFILL23800x80050 (
);

FILL SFILL18760x5050 (
);

FILL FILL_5__12638_ (
);

FILL FILL_3__13672_ (
);

FILL FILL_5__12218_ (
);

FILL FILL_3__13252_ (
);

INVX1 _6938_ (
    .A(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_26_)
);

FILL FILL_4__8765_ (
);

FILL FILL_4__8345_ (
);

FILL FILL111800x53050 (
);

FILL FILL_2__12245_ (
);

FILL FILL_1__11658_ (
);

FILL FILL_1__11238_ (
);

FILL FILL_5__16051_ (
);

NAND3X1 _10936_ (
    .A(\control_1.op [0]),
    .B(_2063_),
    .C(_2069_),
    .Y(_2070_)
);

FILL FILL_0__8245_ (
);

FILL FILL_6__9632_ (
);

INVX1 _10516_ (
    .A(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_1842_)
);

FILL FILL_4__15884_ (
);

FILL FILL_4__15464_ (
);

FILL FILL_4__15044_ (
);

FILL FILL_3__14877_ (
);

FILL FILL_2__9624_ (
);

FILL FILL_3__14457_ (
);

FILL SFILL13880x80050 (
);

FILL SFILL29480x65050 (
);

FILL FILL_3__14037_ (
);

FILL FILL_1__15491_ (
);

FILL FILL_1__15071_ (
);

FILL FILL_0__14484_ (
);

FILL FILL_0__14064_ (
);

FILL SFILL53960x76050 (
);

FILL SFILL84360x67050 (
);

FILL FILL_1__7621_ (
);

FILL FILL_1__7201_ (
);

FILL FILL_2__14811_ (
);

FILL FILL_3__7967_ (
);

FILL FILL_3__7547_ (
);

FILL FILL_5__12391_ (
);

FILL FILL_1__13804_ (
);

FILL FILL_4__16249_ (
);

FILL FILL_4__11384_ (
);

FILL SFILL8760x41050 (
);

FILL FILL_1__16276_ (
);

FILL FILL_5__8834_ (
);

FILL FILL_3__10797_ (
);

FILL FILL_3__10377_ (
);

FILL FILL_0__15689_ (
);

OAI22X1 _15974_ (
    .A(_5480__bF$buf3),
    .B(_5042_),
    .C(_6430_),
    .D(_5569_),
    .Y(_6431_)
);

OAI22X1 _15554_ (
    .A(_5499__bF$buf1),
    .B(_6021_),
    .C(_5532__bF$buf0),
    .D(_6020_),
    .Y(_6022_)
);

FILL FILL_0__15269_ (
);

OAI22X1 _15134_ (
    .A(_4083_),
    .B(_5539__bF$buf2),
    .C(_5530__bF$buf0),
    .D(_5611_),
    .Y(_5612_)
);

FILL FILL_5__10704_ (
);

FILL FILL_1__8826_ (
);

FILL FILL_0__16210_ (
);

FILL FILL_5__13596_ (
);

FILL FILL_2__10311_ (
);

DFFSR _7896_ (
    .Q(\datapath_1.regfile_1.regOut[8] [2]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_458_[2])
);

OAI21X1 _7476_ (
    .A(_302_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .C(_303_),
    .Y(_263_[20])
);

OAI21X1 _7056_ (
    .A(_83_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .C(_84_),
    .Y(_68_[8])
);

FILL FILL_4__12589_ (
);

FILL FILL_4__12169_ (
);

FILL SFILL114520x48050 (
);

FILL FILL_5__9619_ (
);

FILL SFILL53880x38050 (
);

FILL FILL_1__12196_ (
);

FILL FILL_4__13950_ (
);

INVX1 _16339_ (
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_6780_)
);

FILL FILL_4__13530_ (
);

FILL FILL_4__13110_ (
);

NAND2X1 _11894_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[2]),
    .Y(_2971_)
);

FILL FILL_0__11189_ (
);

INVX1 _11474_ (
    .A(_2443_),
    .Y(_2589_)
);

FILL FILL_5__11909_ (
);

NOR2X1 _11054_ (
    .A(_2171_),
    .B(_2172_),
    .Y(_2173_)
);

FILL SFILL43960x74050 (
);

FILL FILL_6__15388_ (
);

FILL FILL_3__12523_ (
);

FILL FILL_3__12103_ (
);

FILL FILL_4__7616_ (
);

FILL FILL_2__11936_ (
);

FILL FILL_2__11516_ (
);

FILL FILL_0__12970_ (
);

FILL FILL_0__12130_ (
);

FILL FILL_1__10929_ (
);

FILL FILL_1__10509_ (
);

FILL FILL_5__15742_ (
);

FILL FILL_0__7936_ (
);

FILL FILL_5__15322_ (
);

FILL FILL_6__8903_ (
);

OAI21X1 _9622_ (
    .A(_1387_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .C(_1388_),
    .Y(_1368_[10])
);

DFFSR _9202_ (
    .Q(\datapath_1.regfile_1.regOut[18] [28]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_1108_[28])
);

FILL FILL_4__14735_ (
);

FILL FILL_4__14315_ (
);

DFFSR _12679_ (
    .Q(\datapath_1.Data [16]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3425_[16])
);

FILL FILL_3__8085_ (
);

NAND3X1 _12259_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3233_)
);

FILL SFILL3720x22050 (
);

FILL FILL_3__13728_ (
);

FILL FILL_3__13308_ (
);

FILL FILL_1__14762_ (
);

FILL FILL_1__14342_ (
);

FILL FILL_5__6900_ (
);

FILL FILL_0__13755_ (
);

FILL FILL_0__13335_ (
);

INVX8 _13620_ (
    .A(_3967__bF$buf2),
    .Y(_4129_)
);

DFFSR _13200_ (
    .Q(\datapath_1.mux_iord.din0 [25]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[25])
);

FILL FILL_5__9792_ (
);

FILL FILL_5__9372_ (
);

NOR2X1 _16092_ (
    .A(_6545_),
    .B(_5549__bF$buf3),
    .Y(_6546_)
);

FILL FILL_5__16107_ (
);

FILL SFILL3640x29050 (
);

FILL FILL_1__9784_ (
);

FILL FILL_5__11662_ (
);

FILL FILL_5__11242_ (
);

FILL FILL_1__9364_ (
);

FILL SFILL43880x36050 (
);

FILL FILL_2__16134_ (
);

FILL FILL_4__10655_ (
);

FILL FILL_4__10235_ (
);

FILL FILL_1__15967_ (
);

FILL FILL_1__15547_ (
);

FILL FILL_1__15127_ (
);

FILL FILL_1__10682_ (
);

FILL FILL_1__10262_ (
);

INVX1 _14825_ (
    .A(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_5309_)
);

INVX1 _14405_ (
    .A(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_4897_)
);

FILL FILL_2__7287_ (
);

FILL FILL_6__13874_ (
);

FILL FILL_6__13454_ (
);

FILL FILL_0__15901_ (
);

FILL FILL_5__12867_ (
);

FILL FILL_5__12447_ (
);

FILL FILL_5__12027_ (
);

FILL FILL_3__13481_ (
);

FILL FILL_4__8994_ (
);

FILL SFILL33880x79050 (
);

FILL FILL_4__8574_ (
);

FILL FILL_2__12894_ (
);

FILL FILL_2__12474_ (
);

FILL FILL_2__12054_ (
);

FILL FILL_1__11887_ (
);

FILL FILL_1__11467_ (
);

FILL FILL_1__11047_ (
);

FILL FILL_0__8894_ (
);

FILL FILL_3__6991_ (
);

FILL FILL_5__16280_ (
);

FILL FILL_0__8474_ (
);

FILL FILL_0__8054_ (
);

INVX1 _10745_ (
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_1954_)
);

OAI21X1 _10325_ (
    .A(_1754_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .C(_1755_),
    .Y(_1693_[31])
);

FILL FILL_4__15693_ (
);

FILL FILL_4__15273_ (
);

FILL FILL_2__9853_ (
);

FILL FILL_0__11821_ (
);

FILL FILL_3__14686_ (
);

FILL FILL_2__9013_ (
);

FILL FILL_3__14266_ (
);

FILL FILL_0__11401_ (
);

FILL FILL_4__9779_ (
);

FILL FILL_4__9359_ (
);

FILL FILL_2__13679_ (
);

FILL FILL_2__13259_ (
);

FILL FILL_0__14293_ (
);

FILL SFILL33880x34050 (
);

FILL FILL_1__7850_ (
);

FILL FILL_1__7430_ (
);

FILL FILL_2__14620_ (
);

FILL SFILL49000x48050 (
);

FILL FILL_0__9679_ (
);

FILL FILL_2__14200_ (
);

FILL FILL_3__7356_ (
);

FILL FILL_0__9259_ (
);

FILL FILL_1__13613_ (
);

FILL FILL_4__16058_ (
);

FILL FILL_6__10579_ (
);

FILL SFILL94440x57050 (
);

FILL FILL_4__11193_ (
);

FILL FILL_0__12606_ (
);

FILL FILL_1__16085_ (
);

FILL FILL_5__8643_ (
);

FILL FILL_3__10186_ (
);

FILL FILL_6_BUFX2_insert771 (
);

FILL FILL_5__8223_ (
);

FILL FILL_0__15498_ (
);

OAI22X1 _15783_ (
    .A(_6244_),
    .B(_5503__bF$buf1),
    .C(_5504__bF$buf4),
    .D(_6243_),
    .Y(_6245_)
);

OAI22X1 _15363_ (
    .A(_4325_),
    .B(_5518__bF$buf2),
    .C(_5478__bF$buf1),
    .D(_4324_),
    .Y(_5836_)
);

FILL FILL_0__15078_ (
);

FILL SFILL23880x77050 (
);

FILL FILL_6_BUFX2_insert776 (
);

FILL FILL_3__16412_ (
);

FILL FILL_5__10933_ (
);

FILL FILL_1__8635_ (
);

FILL FILL_5__10513_ (
);

FILL FILL_1__8215_ (
);

FILL FILL_2__15825_ (
);

FILL FILL_2__15405_ (
);

FILL FILL_2__10960_ (
);

FILL FILL_2__10540_ (
);

FILL FILL_2__10120_ (
);

FILL FILL_6__6986_ (
);

FILL FILL_1__14818_ (
);

DFFSR _7285_ (
    .Q(\datapath_1.regfile_1.regOut[3] [31]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_133_[31])
);

FILL FILL_4__12398_ (
);

FILL FILL_3__9922_ (
);

FILL FILL_3__9502_ (
);

FILL FILL_0__6960_ (
);

FILL FILL_2__6978_ (
);

FILL SFILL94440x12050 (
);

FILL FILL_5__9848_ (
);

FILL FILL_5__9428_ (
);

FILL FILL_5__9008_ (
);

FILL FILL_6__12305_ (
);

FILL SFILL23800x75050 (
);

NAND3X1 _16148_ (
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf1),
    .Y(_6601_)
);

NOR2X1 _11283_ (
    .A(_2401_),
    .B(_2212_),
    .Y(_2402_)
);

FILL FILL_5__11718_ (
);

FILL FILL_3__12752_ (
);

FILL FILL_3__12332_ (
);

FILL FILL_4__7845_ (
);

FILL FILL_4__7425_ (
);

FILL FILL111800x48050 (
);

FILL FILL_2__11745_ (
);

FILL FILL_2__11325_ (
);

FILL SFILL94360x19050 (
);

FILL FILL_1__10318_ (
);

FILL FILL_5__15971_ (
);

FILL FILL_5__15551_ (
);

FILL FILL_5__15131_ (
);

FILL FILL_0__7745_ (
);

FILL FILL_0__7325_ (
);

OAI21X1 _9851_ (
    .A(_1499_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .C(_1500_),
    .Y(_1498_[1])
);

DFFSR _9431_ (
    .Q(\datapath_1.regfile_1.regOut[20] [1]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_1238_[1])
);

NAND2X1 _9011_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1083_)
);

FILL FILL_4__14964_ (
);

FILL FILL_4__14544_ (
);

FILL FILL_4__14124_ (
);

NAND2X1 _12488_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [16]),
    .Y(_3392_)
);

NAND3X1 _12068_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [20]),
    .C(_3034__bF$buf4),
    .Y(_3097_)
);

FILL SFILL23800x30050 (
);

FILL FILL_2__8704_ (
);

FILL FILL_3__13957_ (
);

FILL FILL_1__14991_ (
);

FILL FILL_3__13537_ (
);

FILL FILL_1__14571_ (
);

FILL FILL_3__13117_ (
);

FILL FILL_1__14151_ (
);

FILL FILL_5_BUFX2_insert790 (
);

FILL FILL_5_BUFX2_insert791 (
);

FILL FILL_0__13984_ (
);

FILL FILL_5_BUFX2_insert792 (
);

FILL FILL_5_BUFX2_insert793 (
);

FILL FILL_0__13564_ (
);

FILL FILL_0__13144_ (
);

FILL FILL_5_BUFX2_insert794 (
);

FILL FILL_5_BUFX2_insert795 (
);

FILL FILL_5_BUFX2_insert796 (
);

FILL FILL_5_BUFX2_insert797 (
);

FILL FILL_5_BUFX2_insert798 (
);

FILL FILL_5_BUFX2_insert799 (
);

FILL FILL_5__16336_ (
);

FILL FILL_5__11891_ (
);

FILL FILL_1__9593_ (
);

FILL FILL_5__11471_ (
);

FILL FILL_1__9173_ (
);

FILL FILL_5__11051_ (
);

FILL FILL_4__15749_ (
);

FILL FILL_4__15329_ (
);

FILL FILL_2__16363_ (
);

FILL FILL_3__9099_ (
);

FILL FILL_4__10884_ (
);

FILL SFILL8760x36050 (
);

FILL FILL_2__9909_ (
);

FILL FILL_4__10044_ (
);

FILL SFILL13800x73050 (
);

FILL FILL_1__15776_ (
);

FILL FILL_1__15356_ (
);

FILL FILL_1__10491_ (
);

FILL FILL_0__14769_ (
);

INVX1 _14634_ (
    .A(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_5122_)
);

FILL FILL_0__14349_ (
);

AOI22X1 _14214_ (
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .B(_3885_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_4711_)
);

FILL FILL_2__7096_ (
);

FILL SFILL114600x36050 (
);

FILL FILL_0__15710_ (
);

FILL FILL_5__12256_ (
);

FILL FILL_3__13290_ (
);

OAI21X1 _6976_ (
    .A(_50_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_51_),
    .Y(_3_[24])
);

FILL FILL_4__8383_ (
);

FILL FILL_4__11669_ (
);

FILL FILL_4__11249_ (
);

FILL FILL_2__12283_ (
);

FILL FILL_1__11696_ (
);

FILL FILL_1__11276_ (
);

NOR2X1 _15839_ (
    .A(_6297_),
    .B(_6299_),
    .Y(_6300_)
);

FILL FILL_4__12610_ (
);

INVX1 _15419_ (
    .A(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_5890_)
);

OAI21X1 _10974_ (
    .A(_2099_),
    .B(vdd),
    .C(_2100_),
    .Y(_2098_[0])
);

FILL FILL_0__10689_ (
);

FILL FILL_6__9250_ (
);

OAI21X1 _10554_ (
    .A(_1866_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1867_),
    .Y(_1823_[22])
);

FILL FILL_0__10269_ (
);

OAI21X1 _10134_ (
    .A(_1647_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .C(_1648_),
    .Y(_1628_[10])
);

FILL SFILL43960x69050 (
);

FILL FILL_3__11603_ (
);

FILL FILL_4__15082_ (
);

FILL FILL_2__9662_ (
);

FILL FILL_3__14495_ (
);

FILL FILL_2__9242_ (
);

FILL FILL_0__11630_ (
);

FILL FILL_3__14075_ (
);

FILL FILL_0__11210_ (
);

FILL FILL_4__9168_ (
);

FILL FILL112360x73050 (
);

FILL FILL_2__13488_ (
);

FILL FILL_5__14822_ (
);

FILL FILL_5__14402_ (
);

OAI21X1 _8702_ (
    .A(_916_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .C(_917_),
    .Y(_913_[2])
);

FILL FILL_4__13815_ (
);

FILL FILL_0__9488_ (
);

FILL FILL_3__7585_ (
);

INVX1 _11759_ (
    .A(_2156_),
    .Y(_2854_)
);

FILL FILL_3__7165_ (
);

NAND2X1 _11339_ (
    .A(_2343_),
    .B(_2334_),
    .Y(_2458_)
);

FILL SFILL3720x17050 (
);

FILL FILL_1__13842_ (
);

FILL FILL_1__13422_ (
);

FILL FILL_4__16287_ (
);

FILL FILL_1__13002_ (
);

FILL SFILL43960x24050 (
);

FILL FILL_6__10388_ (
);

FILL SFILL74360x15050 (
);

FILL FILL_0__12835_ (
);

OAI21X1 _12700_ (
    .A(_3491_),
    .B(IRWrite_bF$buf2),
    .C(_3492_),
    .Y(_3490_[1])
);

FILL FILL_0__12415_ (
);

FILL FILL_5__8872_ (
);

FILL FILL_5__8452_ (
);

OAI22X1 _15592_ (
    .A(_5480__bF$buf1),
    .B(_6057_),
    .C(_6058_),
    .D(_5499__bF$buf0),
    .Y(_6059_)
);

INVX8 _15172_ (
    .A(_5530__bF$buf1),
    .Y(_5649_)
);

FILL FILL_5__15607_ (
);

FILL FILL_3__16221_ (
);

NAND2X1 _9907_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1538_)
);

FILL FILL_1__8864_ (
);

FILL FILL_5__10742_ (
);

FILL FILL_1__8444_ (
);

FILL FILL_5__10322_ (
);

FILL FILL_2__15634_ (
);

FILL FILL_2__15214_ (
);

FILL FILL_1__14627_ (
);

NAND2X1 _7094_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_110_)
);

FILL FILL_1__14207_ (
);

FILL FILL_3__9731_ (
);

OAI22X1 _13905_ (
    .A(_4406_),
    .B(_3936__bF$buf1),
    .C(_3935__bF$buf0),
    .D(_4407_),
    .Y(_4408_)
);

FILL FILL112280x35050 (
);

FILL FILL_5__9657_ (
);

FILL FILL_5__9237_ (
);

OAI21X1 _16377_ (
    .A(_6804_),
    .B(gnd),
    .C(_6805_),
    .Y(_6769_[18])
);

FILL FILL_5__11947_ (
);

NOR2X1 _11092_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(_2210_),
    .Y(_2211_)
);

FILL FILL_1__9649_ (
);

FILL FILL_3__12981_ (
);

FILL FILL_5__11527_ (
);

FILL FILL_1__9229_ (
);

FILL FILL_5__11107_ (
);

FILL FILL_3__12141_ (
);

FILL FILL_4__7234_ (
);

FILL FILL_2__11974_ (
);

FILL FILL_2__11554_ (
);

FILL FILL_2__11134_ (
);

FILL SFILL54040x80050 (
);

DFFSR _8299_ (
    .Q(\datapath_1.regfile_1.regOut[11] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_653_[21])
);

FILL FILL_1__10967_ (
);

FILL FILL_1__10547_ (
);

FILL FILL_1__10127_ (
);

FILL FILL_5__15780_ (
);

FILL FILL_0__7974_ (
);

FILL FILL_5__15360_ (
);

FILL FILL_0__7554_ (
);

NAND2X1 _9660_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1414_)
);

FILL FILL_6__8521_ (
);

NAND2X1 _9240_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1195_)
);

FILL FILL_4__14773_ (
);

FILL FILL_4__14353_ (
);

AOI22X1 _12297_ (
    .A(_2_[20]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3262_)
);

FILL FILL_0__10901_ (
);

FILL FILL_3__13766_ (
);

FILL FILL_2__8513_ (
);

FILL FILL_3__13346_ (
);

FILL FILL_1__14380_ (
);

FILL FILL_4__8859_ (
);

FILL FILL_4__8439_ (
);

FILL FILL_4__8019_ (
);

FILL FILL_2__12759_ (
);

FILL FILL_0__13793_ (
);

FILL FILL_2__12339_ (
);

FILL SFILL33880x29050 (
);

FILL FILL_0__13373_ (
);

FILL FILL_1__6930_ (
);

FILL FILL_4__9800_ (
);

FILL FILL_2__13700_ (
);

FILL FILL_0__8759_ (
);

FILL FILL_3__6856_ (
);

FILL FILL_5__16145_ (
);

FILL FILL_6__9726_ (
);

FILL FILL_0__8339_ (
);

FILL FILL_5__11280_ (
);

FILL FILL_4__15978_ (
);

FILL FILL_4__15558_ (
);

FILL FILL_4__15138_ (
);

FILL FILL_2__16172_ (
);

FILL FILL_4__10693_ (
);

FILL FILL_4__10273_ (
);

FILL FILL_2__9718_ (
);

FILL FILL_1__15585_ (
);

FILL FILL_1__15165_ (
);

FILL FILL_5__7723_ (
);

FILL FILL_5__7303_ (
);

FILL FILL_0__14998_ (
);

INVX1 _14863_ (
    .A(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_5346_)
);

FILL FILL_0__14578_ (
);

FILL FILL_0__14158_ (
);

INVX1 _14443_ (
    .A(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_4935_)
);

NOR2X1 _14023_ (
    .A(_4513_),
    .B(_4523_),
    .Y(_4524_)
);

FILL FILL_3__15912_ (
);

FILL FILL_1__7715_ (
);

FILL FILL_2__14905_ (
);

FILL FILL_5__12485_ (
);

FILL FILL_5__12065_ (
);

FILL FILL_4__8192_ (
);

FILL FILL_4__11898_ (
);

FILL FILL_4__11478_ (
);

FILL FILL_4__11058_ (
);

FILL FILL_2__12092_ (
);

FILL FILL_5__8508_ (
);

FILL FILL_1__11085_ (
);

FILL SFILL23080x44050 (
);

NOR2X1 _15648_ (
    .A(_6112_),
    .B(_6113_),
    .Y(_6114_)
);

NOR2X1 _15228_ (
    .A(_5703_),
    .B(_5702_),
    .Y(_5704_)
);

FILL FILL_0__8092_ (
);

FILL FILL_0__10498_ (
);

OAI21X1 _10783_ (
    .A(_1978_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .C(_1979_),
    .Y(_1953_[13])
);

OAI21X1 _10363_ (
    .A(_1759_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .C(_1760_),
    .Y(_1758_[1])
);

FILL SFILL23880x27050 (
);

FILL FILL_6__14697_ (
);

FILL FILL_3__11832_ (
);

FILL FILL_3__11412_ (
);

FILL SFILL8840x69050 (
);

FILL FILL_4__6925_ (
);

FILL FILL_0__16304_ (
);

FILL FILL_2__9891_ (
);

FILL FILL_2__10825_ (
);

FILL FILL_2__9471_ (
);

FILL FILL_2__10405_ (
);

FILL FILL112440x4050 (
);

FILL FILL_4__9397_ (
);

FILL FILL_2__13297_ (
);

FILL FILL_5__14631_ (
);

FILL FILL_5__14211_ (
);

DFFSR _8931_ (
    .Q(\datapath_1.regfile_1.regOut[16] [13]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_978_[13])
);

NAND2X1 _8511_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_831_)
);

FILL SFILL109320x72050 (
);

FILL FILL112040x3050 (
);

FILL FILL_4__13624_ (
);

AND2X2 _11988_ (
    .A(ALUOp_0_bF$buf0),
    .B(PCSource_1_bF$buf4),
    .Y(_3037_)
);

FILL FILL_0__9297_ (
);

NOR2X1 _11568_ (
    .A(_2518_),
    .B(_2507_),
    .Y(_2676_)
);

FILL SFILL23800x25050 (
);

NOR2X1 _11148_ (
    .A(\datapath_1.alu_1.ALUInB [16]),
    .B(_2254_),
    .Y(_2267_)
);

FILL FILL_3__12617_ (
);

FILL FILL_3_BUFX2_insert30 (
);

FILL FILL_1__13651_ (
);

FILL FILL_3_BUFX2_insert31 (
);

FILL FILL_1__13231_ (
);

FILL FILL_4__16096_ (
);

FILL FILL_3_BUFX2_insert32 (
);

FILL FILL_3_BUFX2_insert33 (
);

FILL FILL_3_BUFX2_insert34 (
);

FILL FILL_3_BUFX2_insert35 (
);

FILL FILL_3_BUFX2_insert36 (
);

FILL FILL_3_BUFX2_insert37 (
);

FILL FILL_0__12644_ (
);

FILL FILL_3_BUFX2_insert38 (
);

FILL FILL_0__12224_ (
);

FILL FILL_3_BUFX2_insert39 (
);

FILL FILL_3__15089_ (
);

FILL FILL_5__8261_ (
);

FILL SFILL74120x72050 (
);

FILL SFILL74200x6050 (
);

FILL FILL_5__15836_ (
);

FILL FILL_5__15416_ (
);

FILL FILL_3__16450_ (
);

FILL FILL_3__16030_ (
);

DFFSR _9716_ (
    .Q(\datapath_1.regfile_1.regOut[22] [30]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_1368_[30])
);

FILL FILL_5__10971_ (
);

FILL FILL_5__10551_ (
);

FILL FILL_1__8253_ (
);

FILL FILL_5__10131_ (
);

FILL FILL_4__14829_ (
);

FILL FILL_4__14409_ (
);

FILL FILL_2__15863_ (
);

FILL FILL_2__15443_ (
);

FILL FILL_2__15023_ (
);

FILL FILL_3__8599_ (
);

FILL FILL_1__14856_ (
);

FILL FILL_1__14436_ (
);

FILL FILL_1__14016_ (
);

FILL FILL_0__13849_ (
);

FILL FILL_3__9540_ (
);

FILL FILL_3__9120_ (
);

FILL FILL_0__13429_ (
);

NOR2X1 _13714_ (
    .A(_4220_),
    .B(_4205_),
    .Y(_4221_)
);

FILL FILL_0__13009_ (
);

FILL FILL_5__9886_ (
);

FILL FILL_5__9466_ (
);

FILL FILL_6__12763_ (
);

OAI21X1 _16186_ (
    .A(_5278_),
    .B(_5535__bF$buf0),
    .C(_6637_),
    .Y(_6638_)
);

FILL FILL_5__11756_ (
);

FILL FILL_1__9878_ (
);

FILL FILL_3__12790_ (
);

FILL FILL_5__11336_ (
);

FILL FILL_1__9038_ (
);

FILL FILL_3__12370_ (
);

FILL FILL_2__16228_ (
);

FILL FILL_4__7883_ (
);

FILL FILL_4__7463_ (
);

FILL FILL_4__7043_ (
);

FILL FILL_4__10749_ (
);

FILL FILL_2__11783_ (
);

FILL FILL_2__11363_ (
);

FILL SFILL13800x23050 (
);

FILL FILL_1__10776_ (
);

INVX1 _14919_ (
    .A(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_5401_)
);

FILL FILL_0__7363_ (
);

FILL FILL_6__8330_ (
);

FILL FILL_4__14582_ (
);

FILL FILL_4__14162_ (
);

FILL SFILL64120x70050 (
);

FILL FILL_2__8742_ (
);

FILL FILL_3__13995_ (
);

FILL FILL_2__8322_ (
);

FILL FILL_3__13575_ (
);

FILL FILL_3__13155_ (
);

FILL SFILL34680x28050 (
);

FILL FILL_4__8248_ (
);

FILL FILL112360x68050 (
);

FILL FILL_2__12988_ (
);

FILL FILL_2__12568_ (
);

FILL FILL_2__12148_ (
);

FILL FILL_5__13902_ (
);

FILL FILL_4_BUFX2_insert100 (
);

FILL FILL_4_BUFX2_insert101 (
);

FILL FILL_4_BUFX2_insert102 (
);

FILL SFILL64040x77050 (
);

FILL FILL_4_BUFX2_insert103 (
);

FILL FILL_0__8988_ (
);

FILL FILL_4_BUFX2_insert104 (
);

FILL FILL_5__16374_ (
);

FILL FILL_4_BUFX2_insert105 (
);

FILL FILL_0__8568_ (
);

FILL FILL_4_BUFX2_insert106 (
);

FILL FILL_0__8148_ (
);

DFFSR _10839_ (
    .Q(\datapath_1.regfile_1.regOut[31] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_1953_[1])
);

FILL FILL_4_BUFX2_insert107 (
);

NAND2X1 _10419_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1798_)
);

FILL FILL_4_BUFX2_insert108 (
);

FILL FILL_4_BUFX2_insert109 (
);

FILL FILL_4__15787_ (
);

FILL FILL_4__15367_ (
);

FILL FILL_1__12502_ (
);

FILL SFILL43960x19050 (
);

FILL FILL_2__9527_ (
);

FILL FILL_0__11915_ (
);

FILL FILL_2__9107_ (
);

FILL FILL_1__15394_ (
);

FILL FILL_5__7952_ (
);

FILL FILL_5__7112_ (
);

FILL FILL_0__14387_ (
);

AOI21X1 _14672_ (
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .B(_4038__bF$buf0),
    .C(_5158_),
    .Y(_5159_)
);

AOI22X1 _14252_ (
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .B(_3894_),
    .C(_3995__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_4748_)
);

FILL FILL112360x23050 (
);

FILL FILL_3__15721_ (
);

FILL FILL_3__15301_ (
);

FILL FILL_1__7944_ (
);

FILL FILL_1__7104_ (
);

FILL FILL_2__14714_ (
);

FILL SFILL64040x32050 (
);

FILL FILL_5__12294_ (
);

FILL FILL_1__13707_ (
);

FILL FILL_4__11287_ (
);

FILL SFILL89240x81050 (
);

FILL FILL_1__16179_ (
);

FILL FILL_5__8737_ (
);

FILL FILL_5__8317_ (
);

NAND2X1 _15877_ (
    .A(_6331_),
    .B(_6336_),
    .Y(_6337_)
);

NAND2X1 _15457_ (
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .B(_5693_),
    .Y(_5927_)
);

OAI21X1 _15037_ (
    .A(_5510_),
    .B(_5493_),
    .C(_5516_),
    .Y(_5517_)
);

DFFSR _10592_ (
    .Q(\datapath_1.regfile_1.regOut[29] [10]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1823_[10])
);

NAND2X1 _10172_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1674_)
);

FILL FILL_1__8729_ (
);

FILL FILL_3__11641_ (
);

FILL FILL_3__11221_ (
);

FILL FILL_2__15919_ (
);

FILL FILL_0__16113_ (
);

FILL FILL_2__10634_ (
);

FILL FILL_5__13499_ (
);

FILL SFILL54040x75050 (
);

FILL FILL_2__9280_ (
);

FILL FILL_5__13079_ (
);

NAND2X1 _7799_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .Y(_522_)
);

INVX1 _7379_ (
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_259_)
);

FILL FILL_5__14860_ (
);

FILL FILL_5__14440_ (
);

FILL FILL_5__14020_ (
);

NAND2X1 _8740_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_943_)
);

FILL FILL_6__7601_ (
);

NAND2X1 _8320_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_724_)
);

FILL FILL_1__12099_ (
);

FILL FILL_4__13853_ (
);

FILL FILL_4__13433_ (
);

FILL FILL_4__13013_ (
);

OAI21X1 _11797_ (
    .A(_2888_),
    .B(_2148_),
    .C(_2470__bF$buf1),
    .Y(_2890_)
);

AOI21X1 _11377_ (
    .A(_2492_),
    .B(_2489_),
    .C(_2493_),
    .Y(_2494_)
);

FILL FILL_3__12846_ (
);

FILL FILL_1__13880_ (
);

FILL FILL_3__12426_ (
);

FILL FILL_1__13460_ (
);

FILL FILL_3__12006_ (
);

FILL FILL_1__13040_ (
);

FILL FILL_4__7939_ (
);

FILL FILL_2__11839_ (
);

FILL FILL_0__12873_ (
);

FILL FILL_2__11419_ (
);

FILL FILL_0__12453_ (
);

FILL FILL_0__12033_ (
);

FILL FILL_6__16232_ (
);

FILL FILL_5__8490_ (
);

FILL SFILL54040x30050 (
);

FILL FILL_5__8070_ (
);

FILL FILL_5__15645_ (
);

FILL FILL_5__15225_ (
);

FILL FILL_0__7839_ (
);

DFFSR _9945_ (
    .Q(\datapath_1.regfile_1.regOut[24] [3]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_1498_[3])
);

FILL FILL_0__7419_ (
);

INVX1 _9525_ (
    .A(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_1344_)
);

FILL FILL_5__10780_ (
);

INVX1 _9105_ (
    .A(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_1125_)
);

FILL FILL_5__10360_ (
);

FILL FILL_1__8482_ (
);

FILL FILL_1__8062_ (
);

FILL FILL_4__14638_ (
);

FILL FILL_4__14218_ (
);

FILL FILL_2__15672_ (
);

FILL FILL_2__15252_ (
);

FILL FILL_1__14665_ (
);

FILL FILL_1__14245_ (
);

FILL FILL_0_BUFX2_insert250 (
);

FILL FILL_0_BUFX2_insert251 (
);

FILL FILL_0_BUFX2_insert252 (
);

FILL FILL_0_BUFX2_insert253 (
);

FILL FILL_0_BUFX2_insert254 (
);

FILL FILL_0__13658_ (
);

INVX1 _13943_ (
    .A(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_4445_)
);

FILL FILL_0__13238_ (
);

FILL FILL_0_BUFX2_insert255 (
);

INVX1 _13523_ (
    .A(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_4034_)
);

INVX1 _13103_ (
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_3700_)
);

FILL FILL_0_BUFX2_insert256 (
);

FILL FILL_0_BUFX2_insert257 (
);

FILL FILL_0_BUFX2_insert258 (
);

FILL FILL_5__9275_ (
);

FILL FILL_0_BUFX2_insert259 (
);

FILL SFILL44040x73050 (
);

FILL FILL_6__12152_ (
);

FILL FILL_5__11985_ (
);

FILL SFILL84120x69050 (
);

FILL FILL_5__11565_ (
);

FILL FILL_1__9267_ (
);

FILL FILL_5__11145_ (
);

FILL FILL_4__7692_ (
);

FILL FILL_2__16037_ (
);

FILL FILL_4__10978_ (
);

FILL FILL_4__10558_ (
);

FILL FILL_4__10138_ (
);

FILL FILL_2__11592_ (
);

FILL FILL_2__11172_ (
);

FILL FILL_6__7198_ (
);

FILL FILL_1__10165_ (
);

OAI22X1 _14728_ (
    .A(_5213_),
    .B(_3960_),
    .C(_3959_),
    .D(_5212_),
    .Y(_5214_)
);

NOR2X1 _14308_ (
    .A(_4802_),
    .B(_3944__bF$buf4),
    .Y(_4803_)
);

FILL FILL_0__7592_ (
);

BUFX2 BUFX2_insert990 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf0 )
);

BUFX2 BUFX2_insert991 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf4 )
);

FILL FILL_0__7172_ (
);

BUFX2 BUFX2_insert992 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf3 )
);

BUFX2 BUFX2_insert993 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf2 )
);

BUFX2 BUFX2_insert994 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf1 )
);

FILL FILL_3__10912_ (
);

FILL SFILL109400x60050 (
);

BUFX2 BUFX2_insert995 (
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf0 )
);

FILL FILL_6__13357_ (
);

BUFX2 BUFX2_insert996 (
    .A(_5478_),
    .Y(_5478__bF$buf3)
);

FILL FILL_4__14391_ (
);

BUFX2 BUFX2_insert997 (
    .A(_5478_),
    .Y(_5478__bF$buf2)
);

BUFX2 BUFX2_insert998 (
    .A(_5478_),
    .Y(_5478__bF$buf1)
);

FILL FILL_0__15804_ (
);

BUFX2 BUFX2_insert999 (
    .A(_5478_),
    .Y(_5478__bF$buf0)
);

FILL FILL_2__8971_ (
);

FILL FILL_3__13384_ (
);

FILL FILL_2__8131_ (
);

FILL FILL_4__8897_ (
);

FILL SFILL84120x24050 (
);

FILL FILL_4__8477_ (
);

FILL FILL_4__8057_ (
);

FILL FILL_2__12377_ (
);

FILL FILL_5__13711_ (
);

FILL FILL_4__12704_ (
);

FILL FILL_5__16183_ (
);

FILL FILL_3__6894_ (
);

FILL FILL_0__8377_ (
);

NAND2X1 _10648_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1910_)
);

DFFSR _10228_ (
    .Q(\datapath_1.regfile_1.regOut[26] [30]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_1628_[30])
);

FILL FILL_1__12731_ (
);

FILL FILL_4__15596_ (
);

FILL FILL_4__15176_ (
);

FILL FILL_1__12311_ (
);

FILL SFILL104440x2050 (
);

FILL FILL_2__9756_ (
);

FILL FILL_3__14589_ (
);

FILL FILL_2__9336_ (
);

FILL FILL_0__11724_ (
);

FILL FILL_3__14169_ (
);

FILL FILL_0__11304_ (
);

FILL SFILL104360x7050 (
);

FILL FILL_5__7761_ (
);

FILL SFILL74120x67050 (
);

FILL FILL_5__7341_ (
);

AOI22X1 _14481_ (
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .B(_3995__bF$buf1),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_4972_)
);

FILL FILL_0__14196_ (
);

OAI22X1 _14061_ (
    .A(_4559_),
    .B(_3955__bF$buf1),
    .C(_3983__bF$buf3),
    .D(_4560_),
    .Y(_4561_)
);

FILL FILL_5__14916_ (
);

FILL FILL_3__15950_ (
);

FILL FILL_3__15530_ (
);

FILL FILL_3__15110_ (
);

FILL FILL_1__7753_ (
);

FILL FILL_1__7333_ (
);

FILL FILL_4__13909_ (
);

FILL FILL_2__14943_ (
);

FILL FILL_2__14523_ (
);

FILL FILL_3__7679_ (
);

FILL FILL_2__14103_ (
);

FILL FILL_1__13936_ (
);

FILL FILL_1__13516_ (
);

FILL FILL_4__11096_ (
);

FILL FILL_3__8620_ (
);

FILL FILL_0__12509_ (
);

FILL FILL_3__8200_ (
);

FILL FILL_5__8966_ (
);

FILL FILL_5__8126_ (
);

OAI22X1 _15686_ (
    .A(_6150_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf1),
    .D(_4672_),
    .Y(_6151_)
);

NAND2X1 _15266_ (
    .A(\datapath_1.regfile_1.regOut[7] [5]),
    .B(_5490_),
    .Y(_5741_)
);

FILL SFILL74120x22050 (
);

FILL FILL_3__16315_ (
);

FILL FILL_5__10836_ (
);

FILL FILL_1__8958_ (
);

FILL FILL_3__11870_ (
);

FILL FILL_5__10416_ (
);

FILL FILL_1__8118_ (
);

FILL FILL_3__11450_ (
);

FILL FILL_3__11030_ (
);

FILL FILL_2__15728_ (
);

FILL FILL_2__15308_ (
);

FILL FILL_4__6963_ (
);

FILL SFILL99320x71050 (
);

FILL FILL_0__16342_ (
);

FILL FILL_2__10443_ (
);

FILL FILL_2__10023_ (
);

INVX1 _7188_ (
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_152_)
);

FILL SFILL13800x18050 (
);

FILL SFILL49800x9050 (
);

FILL FILL_3__9405_ (
);

FILL SFILL59160x82050 (
);

FILL FILL_0__6863_ (
);

FILL FILL_4__13662_ (
);

FILL FILL_6__12208_ (
);

FILL FILL_4__13242_ (
);

FILL SFILL64120x65050 (
);

NAND2X1 _11186_ (
    .A(\datapath_1.alu_1.ALUInA [24]),
    .B(_2299_),
    .Y(_2305_)
);

FILL FILL_2__7822_ (
);

FILL SFILL49400x8050 (
);

FILL FILL_3__12655_ (
);

FILL FILL_3__12235_ (
);

FILL FILL_4__7748_ (
);

FILL FILL_4__7328_ (
);

FILL FILL_2__11648_ (
);

FILL FILL_2__11228_ (
);

FILL FILL_0__12262_ (
);

FILL SFILL49000x7050 (
);

FILL SFILL23720x3050 (
);

FILL FILL_5__15874_ (
);

FILL FILL_5__15454_ (
);

FILL FILL_5__15034_ (
);

FILL FILL_0__7228_ (
);

INVX1 _9754_ (
    .A(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_1456_)
);

INVX1 _9334_ (
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_1301_)
);

FILL SFILL63880x6050 (
);

FILL FILL_4__14867_ (
);

FILL FILL_4__14447_ (
);

FILL FILL_4__14027_ (
);

FILL FILL_2__15481_ (
);

FILL FILL_2__15061_ (
);

FILL FILL_2__8607_ (
);

FILL SFILL64120x20050 (
);

FILL FILL_1__14894_ (
);

FILL FILL_1__14474_ (
);

FILL FILL_1__14054_ (
);

FILL FILL_0__13887_ (
);

AOI22X1 _13752_ (
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .B(_3894_),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_4258_)
);

FILL FILL_0__13467_ (
);

NAND2X1 _13332_ (
    .A(_3777_),
    .B(_3760_),
    .Y(_3857_)
);

FILL FILL112360x18050 (
);

FILL FILL_3__14801_ (
);

FILL FILL_5__9084_ (
);

FILL SFILL113800x74050 (
);

FILL FILL_5__16239_ (
);

FILL SFILL64040x27050 (
);

FILL FILL_5__11794_ (
);

FILL FILL_1__9496_ (
);

FILL FILL_5__11374_ (
);

FILL FILL_2__16266_ (
);

FILL FILL_4__10787_ (
);

FILL FILL_4__7081_ (
);

FILL FILL_4__10367_ (
);

FILL FILL_4_BUFX2_insert80 (
);

FILL SFILL89240x76050 (
);

FILL FILL_4_BUFX2_insert81 (
);

FILL FILL_1__15679_ (
);

FILL FILL_4_BUFX2_insert82 (
);

FILL FILL_1__15259_ (
);

FILL FILL_4_BUFX2_insert83 (
);

FILL FILL_4_BUFX2_insert84 (
);

FILL FILL_5__7817_ (
);

FILL FILL_4_BUFX2_insert85 (
);

FILL FILL_4_BUFX2_insert86 (
);

FILL FILL_4_BUFX2_insert87 (
);

FILL FILL_1__10394_ (
);

FILL SFILL9320x42050 (
);

FILL FILL_4_BUFX2_insert88 (
);

FILL FILL_4_BUFX2_insert89 (
);

INVX1 _14957_ (
    .A(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_5438_)
);

NAND3X1 _14537_ (
    .A(_5018_),
    .B(_5019_),
    .C(_5026_),
    .Y(_5027_)
);

INVX1 _14117_ (
    .A(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_4616_)
);

FILL FILL_1__16200_ (
);

FILL FILL_1__7809_ (
);

FILL FILL_3__10301_ (
);

FILL FILL_6__13166_ (
);

FILL FILL_0__15613_ (
);

FILL FILL_5__12999_ (
);

FILL FILL_5__12579_ (
);

FILL FILL_2__8780_ (
);

FILL FILL_2__8360_ (
);

FILL FILL_5__12159_ (
);

BUFX2 _6879_ (
    .A(_2_[9]),
    .Y(memoryWriteData[9])
);

FILL FILL_2__12186_ (
);

FILL FILL_5__13940_ (
);

FILL FILL_5__13520_ (
);

FILL FILL_5__13100_ (
);

NAND2X1 _7820_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_472_)
);

FILL SFILL89240x31050 (
);

DFFSR _7400_ (
    .Q(\datapath_1.regfile_1.regOut[4] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_198_[18])
);

FILL FILL_1__11599_ (
);

FILL FILL_1__11179_ (
);

FILL FILL_4__12513_ (
);

INVX1 _10877_ (
    .A(ALUOp_0_bF$buf5),
    .Y(_2025_)
);

FILL FILL_0__8186_ (
);

DFFSR _10457_ (
    .Q(\datapath_1.regfile_1.regOut[28] [3]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_1758_[3])
);

INVX1 _10037_ (
    .A(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_1604_)
);

FILL FILL_3__11926_ (
);

FILL FILL_1__12960_ (
);

FILL FILL_3__11506_ (
);

FILL SFILL18680x51050 (
);

FILL FILL_1__12120_ (
);

FILL FILL_2__9985_ (
);

FILL FILL_2__10919_ (
);

FILL FILL_0__11953_ (
);

FILL FILL_2__9145_ (
);

FILL FILL_3__14398_ (
);

FILL FILL_0__11533_ (
);

FILL FILL_0__11113_ (
);

FILL FILL_5__7990_ (
);

FILL SFILL54040x25050 (
);

FILL FILL_5__7570_ (
);

AOI22X1 _14290_ (
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .B(_4246_),
    .C(_4001__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_4785_)
);

FILL FILL_5__14725_ (
);

FILL FILL_5__14305_ (
);

FILL FILL_0__6919_ (
);

INVX1 _8605_ (
    .A(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_873_)
);

FILL SFILL79240x74050 (
);

FILL FILL_1__7982_ (
);

FILL FILL_1__7562_ (
);

FILL FILL_4__13718_ (
);

FILL FILL_2__14752_ (
);

FILL FILL_2__14332_ (
);

FILL FILL_3__7488_ (
);

FILL FILL_3__7068_ (
);

FILL FILL_1__13745_ (
);

FILL FILL_1__13325_ (
);

FILL SFILL59160x9050 (
);

FILL FILL_0__12738_ (
);

INVX1 _12603_ (
    .A(\datapath_1.Data [12]),
    .Y(_3448_)
);

FILL FILL_0__12318_ (
);

FILL FILL_5__8775_ (
);

FILL SFILL44040x68050 (
);

FILL FILL_5__8355_ (
);

NAND3X1 _15495_ (
    .A(_5957_),
    .B(_5964_),
    .C(_5952_),
    .Y(_5965_)
);

NAND2X1 _15075_ (
    .A(_5547_),
    .B(_5554_),
    .Y(_5555_)
);

FILL FILL_3__16124_ (
);

FILL FILL_1__8767_ (
);

FILL FILL_5__10645_ (
);

FILL FILL_1__8347_ (
);

FILL FILL_2__15957_ (
);

FILL FILL_2__15537_ (
);

FILL FILL_2__15117_ (
);

FILL FILL_0__16151_ (
);

FILL FILL_2__10672_ (
);

FILL FILL_2__10252_ (
);

FILL FILL111880x42050 (
);

FILL FILL_3__9634_ (
);

FILL FILL_3_BUFX2_insert500 (
);

FILL FILL_3_BUFX2_insert501 (
);

INVX1 _13808_ (
    .A(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_4313_)
);

FILL FILL_3__9214_ (
);

FILL FILL_3_BUFX2_insert502 (
);

FILL SFILL8520x38050 (
);

FILL FILL_3_BUFX2_insert503 (
);

FILL FILL_3_BUFX2_insert504 (
);

FILL FILL_3_BUFX2_insert505 (
);

FILL FILL_3_BUFX2_insert506 (
);

FILL SFILL109240x4050 (
);

FILL FILL_3_BUFX2_insert507 (
);

FILL SFILL109400x55050 (
);

FILL FILL_3_BUFX2_insert508 (
);

FILL FILL_6__12857_ (
);

FILL FILL_3_BUFX2_insert509 (
);

FILL FILL_4__13891_ (
);

FILL FILL_4__13471_ (
);

FILL SFILL44040x23050 (
);

FILL FILL_2__7631_ (
);

FILL FILL_3__12884_ (
);

FILL FILL_3__12464_ (
);

FILL FILL_2__7211_ (
);

FILL FILL_3__12044_ (
);

FILL FILL_4__7977_ (
);

FILL FILL_4__7557_ (
);

FILL FILL_2__11877_ (
);

FILL FILL_2__11457_ (
);

FILL FILL_0__12491_ (
);

FILL FILL_2__11037_ (
);

FILL FILL_0__12071_ (
);

FILL SFILL109800x24050 (
);

FILL FILL_5__15683_ (
);

FILL FILL_0__7877_ (
);

FILL FILL_5__15263_ (
);

INVX1 _9983_ (
    .A(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_1568_)
);

FILL FILL_0__7457_ (
);

FILL FILL_0__7037_ (
);

DFFSR _9563_ (
    .Q(\datapath_1.regfile_1.regOut[21] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1303_[5])
);

OAI21X1 _9143_ (
    .A(_1149_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1150_),
    .Y(_1108_[21])
);

FILL FILL_6__8004_ (
);

FILL FILL_1__11811_ (
);

FILL FILL_4__14676_ (
);

FILL FILL_4__14256_ (
);

FILL FILL_2__15290_ (
);

FILL SFILL109400x10050 (
);

FILL FILL_2__8836_ (
);

FILL FILL_3__13669_ (
);

FILL FILL_0__10804_ (
);

FILL FILL_3__13249_ (
);

FILL FILL_1__14283_ (
);

FILL FILL_5__6841_ (
);

FILL FILL_0_BUFX2_insert630 (
);

FILL FILL_0_BUFX2_insert631 (
);

FILL FILL_0_BUFX2_insert632 (
);

FILL FILL_0_BUFX2_insert633 (
);

FILL FILL_0_BUFX2_insert634 (
);

INVX1 _13981_ (
    .A(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_4482_)
);

FILL FILL_0__13696_ (
);

FILL FILL_0_BUFX2_insert635 (
);

FILL FILL_0__13276_ (
);

INVX1 _13561_ (
    .A(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_4071_)
);

FILL FILL_0_BUFX2_insert636 (
);

OAI21X1 _13141_ (
    .A(_3724_),
    .B(PCEn_bF$buf5),
    .C(_3725_),
    .Y(_3685_[20])
);

FILL FILL_0_BUFX2_insert637 (
);

FILL FILL_3__14610_ (
);

FILL FILL_0_BUFX2_insert638 (
);

FILL FILL_0_BUFX2_insert639 (
);

FILL FILL_2__13603_ (
);

FILL FILL_5__16048_ (
);

FILL FILL_6__9209_ (
);

FILL FILL_5__11183_ (
);

FILL FILL_2__16075_ (
);

FILL FILL_4__10176_ (
);

FILL SFILL69160x34050 (
);

FILL FILL_0__9603_ (
);

FILL FILL_3__7700_ (
);

FILL FILL_1__15488_ (
);

FILL FILL_1__15068_ (
);

FILL FILL_5__7626_ (
);

FILL FILL_5__7206_ (
);

FILL FILL_4__16402_ (
);

FILL SFILL93640x45050 (
);

INVX1 _14766_ (
    .A(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_5251_)
);

FILL SFILL74120x17050 (
);

INVX1 _14346_ (
    .A(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_4840_)
);

FILL FILL_3__15815_ (
);

FILL FILL_3__10950_ (
);

FILL FILL_1__7618_ (
);

FILL FILL_3__10530_ (
);

FILL FILL_3__10110_ (
);

FILL FILL_2__14808_ (
);

FILL SFILL99320x66050 (
);

FILL FILL_0__15842_ (
);

FILL FILL_0__15422_ (
);

FILL FILL_0__15002_ (
);

FILL FILL_5__12388_ (
);

FILL FILL_4__8095_ (
);

FILL SFILL8760x7050 (
);

FILL FILL_3__8905_ (
);

FILL FILL_4__12742_ (
);

FILL FILL_4__12322_ (
);

INVX1 _10686_ (
    .A(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_1935_)
);

INVX1 _10266_ (
    .A(\datapath_1.regfile_1.regOut[27] [12]),
    .Y(_1716_)
);

FILL FILL_2__6902_ (
);

FILL FILL_3__11735_ (
);

FILL FILL_3__11315_ (
);

FILL FILL_0__16207_ (
);

FILL SFILL59560x46050 (
);

FILL FILL_2__9794_ (
);

FILL FILL_2__10308_ (
);

FILL FILL_0__11762_ (
);

FILL FILL_2__9374_ (
);

FILL SFILL99320x21050 (
);

FILL FILL_0__11342_ (
);

FILL FILL_6__15961_ (
);

FILL FILL_6__15541_ (
);

FILL FILL_5__14954_ (
);

FILL FILL_5__14534_ (
);

FILL FILL_5__14114_ (
);

FILL SFILL28760x41050 (
);

INVX1 _8834_ (
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_985_)
);

FILL SFILL59160x32050 (
);

DFFSR _8414_ (
    .Q(\datapath_1.regfile_1.regOut[12] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_718_[8])
);

FILL FILL_1__7371_ (
);

FILL FILL_4__13947_ (
);

FILL FILL_4__13527_ (
);

FILL FILL_2__14981_ (
);

FILL FILL_2__14561_ (
);

FILL FILL_4__13107_ (
);

FILL FILL_2__14141_ (
);

FILL FILL_3__7297_ (
);

FILL SFILL64120x15050 (
);

FILL FILL_1__13974_ (
);

FILL FILL_1__13554_ (
);

FILL FILL_1__13134_ (
);

FILL FILL_0__12967_ (
);

INVX1 _12832_ (
    .A(\datapath_1.a [3]),
    .Y(_3560_)
);

FILL SFILL89320x64050 (
);

INVX1 _12412_ (
    .A(ALUOut[23]),
    .Y(_3340_)
);

FILL FILL_0__12127_ (
);

FILL FILL_5__8584_ (
);

FILL FILL_6__11881_ (
);

FILL FILL_6__11461_ (
);

FILL FILL_5__15739_ (
);

FILL FILL_5__15319_ (
);

FILL FILL_3__16353_ (
);

OAI21X1 _9619_ (
    .A(_1385_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .C(_1386_),
    .Y(_1368_[9])
);

FILL FILL_1__8996_ (
);

FILL FILL_5__10874_ (
);

FILL FILL_1__8576_ (
);

FILL FILL_5__10034_ (
);

FILL FILL_2__15766_ (
);

FILL FILL_2__15346_ (
);

FILL FILL_0__16380_ (
);

FILL SFILL54120x58050 (
);

FILL FILL_2__10061_ (
);

FILL FILL_1__14759_ (
);

FILL FILL_1__14339_ (
);

FILL FILL_3__9863_ (
);

OAI22X1 _13617_ (
    .A(_3890_),
    .B(_4125_),
    .C(_4124_),
    .D(_3931__bF$buf0),
    .Y(_4126_)
);

FILL FILL_3__9023_ (
);

FILL FILL_5__9789_ (
);

FILL FILL_1__15700_ (
);

FILL FILL_5__9369_ (
);

FILL FILL_4__13280_ (
);

NOR2X1 _16089_ (
    .A(_5205_),
    .B(_5534__bF$buf1),
    .Y(_6543_)
);

FILL FILL_2__7860_ (
);

FILL FILL_5__11659_ (
);

FILL FILL_2__7440_ (
);

FILL FILL_5__11239_ (
);

FILL FILL_3__12273_ (
);

FILL FILL_4__7366_ (
);

FILL FILL_2__11686_ (
);

FILL FILL_2__11266_ (
);

FILL FILL_5__12600_ (
);

BUFX2 _6900_ (
    .A(_2_[30]),
    .Y(memoryWriteData[30])
);

FILL SFILL54120x13050 (
);

FILL FILL_1__10679_ (
);

FILL FILL_1__10259_ (
);

FILL FILL_5__15492_ (
);

FILL FILL_5__15072_ (
);

FILL FILL_0__7686_ (
);

OAI21X1 _9792_ (
    .A(_1480_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .C(_1481_),
    .Y(_1433_[24])
);

OAI21X1 _9372_ (
    .A(_1261_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1262_),
    .Y(_1238_[12])
);

FILL SFILL79320x62050 (
);

FILL SFILL18680x46050 (
);

FILL FILL_4__14485_ (
);

FILL FILL_1__11620_ (
);

FILL FILL_4__14065_ (
);

FILL FILL_1__11200_ (
);

FILL FILL_2__8645_ (
);

FILL FILL_3__13898_ (
);

FILL FILL_2__8225_ (
);

FILL FILL_3__13478_ (
);

FILL FILL111960x75050 (
);

FILL FILL_1__14092_ (
);

INVX1 _13790_ (
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_4295_)
);

FILL FILL_0__13085_ (
);

INVX8 _13370_ (
    .A(_3881_),
    .Y(_3882_)
);

FILL FILL_5__13805_ (
);

FILL SFILL79240x69050 (
);

FILL FILL_4__9932_ (
);

FILL FILL_4__9512_ (
);

FILL FILL_2__13832_ (
);

FILL FILL_3__6988_ (
);

FILL FILL_2__13412_ (
);

FILL FILL_5__16277_ (
);

FILL FILL_1__12825_ (
);

FILL FILL_1__12405_ (
);

FILL FILL_0__9412_ (
);

FILL FILL_0__11818_ (
);

FILL FILL_1__15297_ (
);

FILL FILL_5__7855_ (
);

FILL FILL_5__7435_ (
);

FILL FILL_4__16211_ (
);

FILL FILL111960x30050 (
);

INVX2 _14995_ (
    .A(\datapath_1.PCJump [24]),
    .Y(_5475_)
);

OAI22X1 _14575_ (
    .A(_5062_),
    .B(_3955__bF$buf3),
    .C(_3954__bF$buf3),
    .D(_5063_),
    .Y(_5064_)
);

INVX1 _14155_ (
    .A(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_4653_)
);

FILL FILL_3__15624_ (
);

FILL FILL_3__15204_ (
);

FILL FILL_1__7847_ (
);

FILL FILL_1__7427_ (
);

FILL SFILL79240x24050 (
);

FILL FILL_2__14617_ (
);

FILL FILL_0__15651_ (
);

FILL FILL_0__15231_ (
);

FILL FILL_5__12197_ (
);

FILL FILL_3__8714_ (
);

FILL FILL_6__11937_ (
);

FILL FILL_4__12971_ (
);

FILL SFILL44040x18050 (
);

FILL FILL_4__12131_ (
);

FILL FILL_3__16409_ (
);

INVX1 _10495_ (
    .A(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_1828_)
);

DFFSR _10075_ (
    .Q(\datapath_1.regfile_1.regOut[25] [5]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_1563_[5])
);

FILL FILL_3__11964_ (
);

FILL FILL_3__11544_ (
);

FILL FILL_3__11124_ (
);

FILL SFILL69240x67050 (
);

FILL FILL_0__16016_ (
);

OAI22X1 _16301_ (
    .A(_5480__bF$buf1),
    .B(_5425_),
    .C(_6749_),
    .D(_5499__bF$buf3),
    .Y(_6750_)
);

FILL FILL_2__10957_ (
);

FILL FILL_0__11991_ (
);

FILL FILL_2__10537_ (
);

FILL FILL_0__11571_ (
);

FILL FILL_2__10117_ (
);

FILL FILL_0__11151_ (
);

FILL FILL_3__9919_ (
);

FILL FILL_5__14763_ (
);

FILL FILL_0__6957_ (
);

FILL FILL_5__14343_ (
);

OAI21X1 _8643_ (
    .A(_897_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_898_),
    .Y(_848_[25])
);

OAI21X1 _8223_ (
    .A(_678_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_679_),
    .Y(_653_[13])
);

FILL FILL_1__7180_ (
);

FILL FILL_4__13756_ (
);

FILL FILL_4__13336_ (
);

FILL FILL_2__14790_ (
);

FILL FILL_2__14370_ (
);

FILL FILL_3__12749_ (
);

FILL FILL_1__13783_ (
);

FILL FILL_3__12329_ (
);

FILL FILL_1__13363_ (
);

FILL FILL_0__12776_ (
);

OAI21X1 _12641_ (
    .A(_3472_),
    .B(vdd),
    .C(_3473_),
    .Y(_3425_[24])
);

FILL FILL_0__12356_ (
);

AOI22X1 _12221_ (
    .A(_2_[1]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf3),
    .D(gnd),
    .Y(_3205_)
);

FILL FILL_5__8393_ (
);

FILL FILL_6__16135_ (
);

FILL FILL_5__15968_ (
);

FILL FILL_5__15548_ (
);

FILL FILL_5__15128_ (
);

OAI21X1 _9848_ (
    .A(_1561_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .C(_1562_),
    .Y(_1498_[0])
);

FILL FILL_3__16162_ (
);

NAND2X1 _9428_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1300_)
);

FILL FILL_5__10683_ (
);

NAND2X1 _9008_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1081_)
);

FILL FILL_5__10263_ (
);

FILL FILL_1__8385_ (
);

FILL FILL_2__15995_ (
);

FILL FILL_2__15575_ (
);

FILL FILL_2__15155_ (
);

FILL SFILL99400x54050 (
);

FILL SFILL69160x29050 (
);

FILL FILL_2__10290_ (
);

FILL FILL_1__14988_ (
);

FILL FILL_1__14568_ (
);

FILL FILL_1__14148_ (
);

FILL FILL_4__15902_ (
);

FILL FILL_3__9672_ (
);

OAI22X1 _13846_ (
    .A(_3944__bF$buf2),
    .B(_4348_),
    .C(_4349_),
    .D(_3955__bF$buf3),
    .Y(_4350_)
);

FILL FILL_3__9252_ (
);

NOR2X1 _13426_ (
    .A(_3932_),
    .B(_3937_),
    .Y(_3938_)
);

NAND2X1 _13006_ (
    .A(vdd),
    .B(\datapath_1.rd2 [18]),
    .Y(_3656_)
);

FILL FILL_5__9598_ (
);

FILL FILL_6__12055_ (
);

FILL FILL_0__14922_ (
);

FILL FILL_0__14502_ (
);

FILL FILL_5__11888_ (
);

FILL FILL_5__11468_ (
);

FILL FILL_5__11048_ (
);

FILL FILL_3__12082_ (
);

FILL FILL_4__7595_ (
);

FILL FILL_4__7175_ (
);

FILL FILL_2__11495_ (
);

FILL FILL_2__11075_ (
);

FILL FILL_1__10488_ (
);

FILL FILL_1__10068_ (
);

FILL FILL_4__11822_ (
);

FILL FILL_4__11402_ (
);

FILL FILL_0__7495_ (
);

FILL FILL_0__7075_ (
);

DFFSR _9181_ (
    .Q(\datapath_1.regfile_1.regOut[18] [7]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1108_[7])
);

FILL FILL_3__10815_ (
);

FILL FILL_4__14294_ (
);

FILL FILL_0__15707_ (
);

FILL FILL_2__8874_ (
);

FILL SFILL99320x16050 (
);

FILL FILL_2__8454_ (
);

FILL FILL_0__10422_ (
);

FILL FILL_3__13287_ (
);

FILL FILL_0__10002_ (
);

FILL FILL_6__14201_ (
);

FILL SFILL49640x77050 (
);

FILL FILL_5__13614_ (
);

FILL SFILL59160x27050 (
);

DFFSR _7914_ (
    .Q(\datapath_1.regfile_1.regOut[8] [20]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_458_[20])
);

FILL FILL_1__6871_ (
);

FILL FILL_4__9741_ (
);

FILL FILL_4__12607_ (
);

FILL FILL_2__13641_ (
);

FILL FILL_2__13221_ (
);

FILL FILL_5__16086_ (
);

FILL FILL_1__12634_ (
);

FILL FILL_4__15499_ (
);

FILL FILL_1__12214_ (
);

FILL FILL_4__15079_ (
);

FILL FILL_2__9659_ (
);

FILL FILL_0__9641_ (
);

FILL SFILL89320x59050 (
);

NAND2X1 _11912_ (
    .A(IorD_bF$buf0),
    .B(ALUOut[8]),
    .Y(_2983_)
);

FILL FILL_2__9239_ (
);

FILL FILL_0__9221_ (
);

FILL FILL_0__11627_ (
);

FILL FILL_0__11207_ (
);

FILL FILL_5__7244_ (
);

FILL FILL_4__16020_ (
);

FILL FILL_6__10961_ (
);

INVX1 _14384_ (
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_4877_)
);

FILL FILL_0__14099_ (
);

FILL FILL_5__14819_ (
);

FILL FILL_3__15853_ (
);

FILL SFILL18760x79050 (
);

FILL FILL_3__15433_ (
);

FILL FILL_3__15013_ (
);

FILL FILL_1__7236_ (
);

FILL FILL_2__14846_ (
);

FILL FILL_2__14426_ (
);

FILL FILL_0__15880_ (
);

FILL FILL_2__14006_ (
);

FILL FILL_0__15460_ (
);

FILL FILL_0__15040_ (
);

FILL FILL_1__13839_ (
);

FILL FILL_1__13419_ (
);

FILL FILL_3__8523_ (
);

FILL SFILL79800x64050 (
);

FILL FILL_3__8103_ (
);

FILL SFILL33960x54050 (
);

FILL FILL_5__8869_ (
);

FILL FILL_5__8449_ (
);

FILL SFILL89320x14050 (
);

FILL FILL_4__12780_ (
);

OAI21X1 _15589_ (
    .A(_5524__bF$buf2),
    .B(_4578_),
    .C(_6055_),
    .Y(_6056_)
);

OAI22X1 _15169_ (
    .A(_5534__bF$buf2),
    .B(_4132_),
    .C(_5645_),
    .D(_5549__bF$buf2),
    .Y(_5646_)
);

FILL FILL_4__12360_ (
);

FILL FILL_3__16218_ (
);

FILL SFILL113800x19050 (
);

FILL FILL_2__6940_ (
);

FILL FILL_5__10319_ (
);

FILL FILL_3__11773_ (
);

FILL FILL_5__9810_ (
);

FILL FILL_3__11353_ (
);

FILL SFILL18760x34050 (
);

FILL FILL_4__6866_ (
);

FILL FILL_0__16245_ (
);

NOR2X1 _16110_ (
    .A(_6563_),
    .B(_6560_),
    .Y(_6564_)
);

FILL FILL_2__10766_ (
);

FILL FILL_0__11380_ (
);

FILL FILL_1__9802_ (
);

FILL FILL_3__9728_ (
);

FILL FILL_5__14992_ (
);

FILL FILL_5__14572_ (
);

FILL FILL_5__14152_ (
);

OAI21X1 _8872_ (
    .A(_1009_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .C(_1010_),
    .Y(_978_[16])
);

OAI21X1 _8452_ (
    .A(_790_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .C(_791_),
    .Y(_783_[4])
);

FILL SFILL79320x57050 (
);

DFFSR _8032_ (
    .Q(\datapath_1.regfile_1.regOut[9] [10]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_523_[10])
);

FILL FILL_4__13985_ (
);

FILL FILL_1__10700_ (
);

FILL FILL_4__13565_ (
);

FILL FILL_4__13145_ (
);

NOR2X1 _11089_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(_2183_),
    .Y(_2208_)
);

FILL FILL_2__7725_ (
);

FILL FILL_3__12978_ (
);

FILL FILL_2__7305_ (
);

FILL FILL_1__13592_ (
);

FILL FILL_3__12138_ (
);

FILL FILL_1__13172_ (
);

FILL FILL_0__12585_ (
);

OAI21X1 _12870_ (
    .A(_3584_),
    .B(vdd),
    .C(_3585_),
    .Y(_3555_[15])
);

OAI21X1 _12450_ (
    .A(_3365_),
    .B(vdd),
    .C(_3366_),
    .Y(_3360_[3])
);

FILL FILL_0__12165_ (
);

NAND3X1 _12030_ (
    .A(_3066_),
    .B(_3067_),
    .C(_3068_),
    .Y(\datapath_1.mux_pcsrc.dout [10])
);

FILL FILL_5_BUFX2_insert410 (
);

FILL FILL_2__12912_ (
);

FILL FILL_5_BUFX2_insert411 (
);

FILL FILL_5__15777_ (
);

FILL FILL_5__15357_ (
);

FILL FILL_5_BUFX2_insert412 (
);

FILL FILL_5_BUFX2_insert413 (
);

FILL FILL_3__16391_ (
);

NAND2X1 _9657_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1412_)
);

FILL FILL_5_BUFX2_insert414 (
);

FILL FILL_5_BUFX2_insert415 (
);

NAND2X1 _9237_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1193_)
);

FILL FILL_5_BUFX2_insert416 (
);

FILL FILL_5__10492_ (
);

FILL FILL_1__8194_ (
);

FILL FILL_5_BUFX2_insert417 (
);

FILL FILL_1__11905_ (
);

FILL FILL_5_BUFX2_insert418 (
);

FILL FILL_5_BUFX2_insert419 (
);

FILL FILL_2__15384_ (
);

FILL SFILL114440x82050 (
);

FILL SFILL79320x12050 (
);

FILL FILL_0__8912_ (
);

FILL FILL_1__14797_ (
);

FILL FILL_1__14377_ (
);

FILL FILL_5__6935_ (
);

FILL FILL_4__15711_ (
);

FILL FILL111960x25050 (
);

FILL FILL_3__9481_ (
);

NOR2X1 _13655_ (
    .A(_4159_),
    .B(_4162_),
    .Y(_4163_)
);

OAI21X1 _13235_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .C(_3777_),
    .Y(_3778_)
);

FILL FILL_3__14704_ (
);

FILL FILL_1__6927_ (
);

FILL SFILL63640x34050 (
);

FILL FILL_0__14731_ (
);

FILL FILL_0__14311_ (
);

FILL FILL_5__11697_ (
);

FILL FILL_1__9399_ (
);

FILL FILL_5__11277_ (
);

FILL FILL_2__16169_ (
);

FILL SFILL69320x55050 (
);

FILL FILL_2_BUFX2_insert540 (
);

FILL FILL_1__10297_ (
);

FILL FILL_2_BUFX2_insert541 (
);

FILL FILL_2_BUFX2_insert542 (
);

FILL FILL_2_BUFX2_insert543 (
);

FILL FILL_2_BUFX2_insert544 (
);

FILL FILL_4__11631_ (
);

FILL FILL_2_BUFX2_insert545 (
);

FILL FILL_4__11211_ (
);

FILL FILL_3__15909_ (
);

FILL FILL_2_BUFX2_insert546 (
);

FILL FILL_2_BUFX2_insert547 (
);

FILL FILL_2_BUFX2_insert548 (
);

FILL FILL_2_BUFX2_insert549 (
);

FILL FILL_1__16103_ (
);

FILL FILL_3__10624_ (
);

FILL FILL_0__15936_ (
);

FILL FILL_0__15516_ (
);

OAI22X1 _15801_ (
    .A(_5530__bF$buf0),
    .B(_4819_),
    .C(_5532__bF$buf1),
    .D(_4823_),
    .Y(_6263_)
);

FILL FILL_0__10651_ (
);

FILL FILL_2__8263_ (
);

FILL FILL_0__10231_ (
);

FILL FILL_3__13096_ (
);

FILL FILL_4__8189_ (
);

FILL FILL_2__12089_ (
);

FILL FILL_5__13843_ (
);

FILL FILL_5__13423_ (
);

FILL FILL_5__13003_ (
);

OAI21X1 _7723_ (
    .A(_426_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .C(_427_),
    .Y(_393_[17])
);

OAI21X1 _7303_ (
    .A(_207_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .C(_208_),
    .Y(_198_[5])
);

FILL FILL_4__9550_ (
);

FILL FILL_4__12836_ (
);

FILL FILL_4__9130_ (
);

FILL FILL_4__12416_ (
);

FILL FILL_2__13870_ (
);

FILL FILL_2__13450_ (
);

FILL FILL_6__9896_ (
);

FILL FILL_2__13030_ (
);

FILL FILL_0__8089_ (
);

FILL FILL_3__11829_ (
);

FILL FILL_1__12863_ (
);

FILL FILL_3__11409_ (
);

FILL FILL_1__12443_ (
);

FILL FILL_1__12023_ (
);

FILL FILL_0__9870_ (
);

FILL FILL_2__9888_ (
);

FILL SFILL69240x17050 (
);

FILL FILL_0__11856_ (
);

FILL FILL_2__9468_ (
);

FILL FILL_0__9030_ (
);

NAND3X1 _11721_ (
    .A(_2462__bF$buf3),
    .B(_2802_),
    .C(_2818_),
    .Y(_2819_)
);

FILL FILL_0__11436_ (
);

FILL FILL_0__11016_ (
);

NOR2X1 _11301_ (
    .A(_2257_),
    .B(_2419_),
    .Y(_2420_)
);

FILL FILL_5__7893_ (
);

FILL FILL_5__7473_ (
);

FILL FILL_5__7053_ (
);

FILL FILL_6__10770_ (
);

NOR2X1 _14193_ (
    .A(_4689_),
    .B(_4686_),
    .Y(_4690_)
);

FILL FILL_5__14628_ (
);

FILL FILL_3__15662_ (
);

FILL FILL_5__14208_ (
);

FILL FILL_3__15242_ (
);

DFFSR _8928_ (
    .Q(\datapath_1.regfile_1.regOut[16] [10]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_978_[10])
);

NAND2X1 _8508_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_829_)
);

FILL FILL_1__7885_ (
);

FILL FILL_1__7465_ (
);

FILL FILL_1__7045_ (
);

FILL FILL_2__14655_ (
);

FILL SFILL99400x49050 (
);

FILL FILL_2__14235_ (
);

FILL FILL_1__13648_ (
);

FILL FILL_1__13228_ (
);

FILL FILL_1_BUFX2_insert560 (
);

FILL FILL_3__8752_ (
);

FILL FILL_1_BUFX2_insert561 (
);

FILL FILL_3__8332_ (
);

DFFSR _12926_ (
    .Q(\datapath_1.a [7]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3555_[7])
);

FILL FILL_1_BUFX2_insert562 (
);

FILL FILL_1_BUFX2_insert563 (
);

NAND2X1 _12506_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [22]),
    .Y(_3404_)
);

FILL FILL_1_BUFX2_insert564 (
);

FILL FILL_1_BUFX2_insert565 (
);

FILL FILL_1_BUFX2_insert566 (
);

FILL FILL_1_BUFX2_insert567 (
);

FILL FILL_5__8258_ (
);

FILL FILL_1_BUFX2_insert568 (
);

FILL FILL_1_BUFX2_insert569 (
);

NAND3X1 _15398_ (
    .A(_5862_),
    .B(_5867_),
    .C(_5869_),
    .Y(_5870_)
);

FILL FILL_3__16027_ (
);

FILL FILL_5__10968_ (
);

FILL FILL_5__10548_ (
);

FILL FILL_5__10128_ (
);

FILL FILL_3__11582_ (
);

FILL FILL_3__11162_ (
);

FILL FILL_0__16054_ (
);

FILL FILL_2__10995_ (
);

FILL FILL_2__10575_ (
);

FILL FILL_2__10155_ (
);

FILL FILL_1__9611_ (
);

FILL FILL_3__9537_ (
);

FILL FILL_4__10902_ (
);

FILL FILL_3__9117_ (
);

FILL FILL_0__6995_ (
);

FILL FILL_5__14381_ (
);

DFFSR _8681_ (
    .Q(\datapath_1.regfile_1.regOut[14] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_848_[19])
);

FILL SFILL59240x15050 (
);

NAND2X1 _8261_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_705_)
);

FILL FILL_4__13794_ (
);

FILL FILL_4__13374_ (
);

FILL FILL_2__7954_ (
);

FILL FILL_3__12787_ (
);

BUFX2 BUFX2_insert230 (
    .A(_2347_),
    .Y(_2347__bF$buf3)
);

FILL FILL_2__7114_ (
);

FILL FILL_3__12367_ (
);

BUFX2 BUFX2_insert231 (
    .A(_2347_),
    .Y(_2347__bF$buf2)
);

BUFX2 BUFX2_insert232 (
    .A(_2347_),
    .Y(_2347__bF$buf1)
);

FILL SFILL89880x9050 (
);

BUFX2 BUFX2_insert233 (
    .A(_2347_),
    .Y(_2347__bF$buf0)
);

BUFX2 BUFX2_insert234 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf4 )
);

BUFX2 BUFX2_insert235 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf3 )
);

BUFX2 BUFX2_insert236 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf2 )
);

BUFX2 BUFX2_insert237 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf1 )
);

BUFX2 BUFX2_insert238 (
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf0 )
);

BUFX2 BUFX2_insert239 (
    .A(_5545_),
    .Y(_5545__bF$buf3)
);

FILL FILL_0__12394_ (
);

FILL FILL_4__8401_ (
);

FILL FILL_2__12721_ (
);

FILL FILL_5__15586_ (
);

FILL FILL_2__12301_ (
);

FILL FILL_5__15166_ (
);

NAND2X1 _9886_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1524_)
);

NAND2X1 _9466_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1305_)
);

DFFSR _9046_ (
    .Q(\datapath_1.regfile_1.regOut[17] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_1043_[0])
);

FILL FILL_4__14999_ (
);

FILL FILL_4__14579_ (
);

FILL FILL_1__11714_ (
);

FILL FILL_4__14159_ (
);

FILL FILL_2__15193_ (
);

FILL FILL_2__8739_ (
);

FILL FILL_0__8721_ (
);

FILL FILL_2__8319_ (
);

FILL FILL_0__10707_ (
);

FILL FILL_1__14186_ (
);

FILL FILL_4__15940_ (
);

FILL FILL_4__15520_ (
);

FILL FILL_4__15100_ (
);

FILL FILL_0__13599_ (
);

AOI22X1 _13884_ (
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .B(_4102_),
    .C(_3995__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_4388_)
);

FILL FILL_3__9290_ (
);

INVX1 _13464_ (
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_3976_)
);

INVX1 _13044_ (
    .A(_2_[31]),
    .Y(_3681_)
);

FILL FILL_3__14933_ (
);

FILL FILL_3__14513_ (
);

FILL FILL_4__9606_ (
);

FILL FILL_2__13926_ (
);

FILL FILL_0__14960_ (
);

FILL FILL_2__13506_ (
);

FILL FILL_0__14540_ (
);

FILL FILL_0__14120_ (
);

FILL FILL_5__11086_ (
);

FILL FILL_2__16398_ (
);

FILL SFILL33160x66050 (
);

FILL FILL_4__10499_ (
);

FILL FILL_0__9926_ (
);

FILL FILL_0__9506_ (
);

FILL FILL_3__7603_ (
);

FILL SFILL33960x49050 (
);

FILL FILL_5__7949_ (
);

FILL FILL_5__7109_ (
);

FILL FILL_4__16305_ (
);

FILL FILL_4__11860_ (
);

AOI22X1 _14669_ (
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .B(_4102_),
    .C(_4001__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_5156_)
);

OAI22X1 _14249_ (
    .A(_4743_),
    .B(_3905__bF$buf2),
    .C(_3909_),
    .D(_4744_),
    .Y(_4745_)
);

FILL FILL_4__11440_ (
);

FILL FILL_4__11020_ (
);

FILL FILL_3__15718_ (
);

FILL FILL_1__16332_ (
);

FILL SFILL18760x29050 (
);

FILL FILL_3__10433_ (
);

FILL FILL_3__10013_ (
);

FILL FILL_0__15745_ (
);

FILL FILL_0__15325_ (
);

AOI21X1 _15610_ (
    .A(_6053_),
    .B(_6076_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [13])
);

FILL FILL_0__10880_ (
);

FILL FILL_2__8492_ (
);

FILL FILL_2__8072_ (
);

FILL FILL_0__10040_ (
);

FILL FILL_5__13652_ (
);

FILL FILL_5__13232_ (
);

OAI21X1 _7952_ (
    .A(_538_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_539_),
    .Y(_523_[8])
);

DFFSR _7532_ (
    .Q(\datapath_1.regfile_1.regOut[5] [22]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_263_[22])
);

NAND2X1 _7112_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_122_)
);

FILL FILL_4__12645_ (
);

FILL FILL_4__12225_ (
);

DFFSR _10589_ (
    .Q(\datapath_1.regfile_1.regOut[29] [7]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1823_[7])
);

NAND2X1 _10169_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1672_)
);

FILL FILL_3__11638_ (
);

FILL FILL_3__11218_ (
);

FILL FILL_1__12252_ (
);

FILL SFILL84280x51050 (
);

FILL FILL_2__9277_ (
);

INVX1 _11950_ (
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3008_)
);

FILL FILL_0__11665_ (
);

FILL FILL_0__11245_ (
);

OAI21X1 _11530_ (
    .A(_2411_),
    .B(_2344__bF$buf2),
    .C(_2640_),
    .Y(_2641_)
);

NOR2X1 _11110_ (
    .A(_2227_),
    .B(_2228_),
    .Y(_2229_)
);

FILL FILL_6__15864_ (
);

FILL FILL_6__15444_ (
);

FILL FILL_5__14857_ (
);

FILL FILL_5__14437_ (
);

FILL FILL_3__15891_ (
);

FILL FILL_5__14017_ (
);

FILL FILL_3__15471_ (
);

NAND2X1 _8737_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_941_)
);

FILL FILL_3__15051_ (
);

NAND2X1 _8317_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_722_)
);

FILL FILL_1__7694_ (
);

FILL FILL_2__14884_ (
);

FILL FILL_2__14464_ (
);

FILL FILL_2__14044_ (
);

FILL FILL_1__13877_ (
);

FILL FILL_1__13457_ (
);

FILL FILL_1__13037_ (
);

FILL FILL_3__8981_ (
);

FILL FILL_3__8141_ (
);

NAND2X1 _12735_ (
    .A(IRWrite_bF$buf3),
    .B(memoryOutData[13]),
    .Y(_3516_)
);

NAND3X1 _12315_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3275_)
);

FILL FILL_5__8487_ (
);

FILL FILL_5__8067_ (
);

FILL FILL_6__11784_ (
);

FILL SFILL114840x46050 (
);

FILL FILL_6__11364_ (
);

FILL FILL_0__13811_ (
);

FILL FILL_3__16256_ (
);

FILL FILL_5__10777_ (
);

FILL FILL_1__8899_ (
);

FILL FILL_1__8479_ (
);

FILL FILL_3__11391_ (
);

FILL FILL_1__8059_ (
);

FILL FILL_2__15669_ (
);

FILL FILL_2__15249_ (
);

FILL FILL_0__16283_ (
);

FILL FILL_2__10384_ (
);

FILL SFILL114440x32050 (
);

FILL FILL_1__9420_ (
);

FILL FILL_1__9000_ (
);

FILL FILL_3__9766_ (
);

FILL FILL_3__9346_ (
);

FILL SFILL109560x2050 (
);

FILL FILL_5__14190_ (
);

NAND2X1 _8490_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_817_)
);

FILL FILL_1__15603_ (
);

NAND2X1 _8070_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_598_)
);

FILL FILL_2__7763_ (
);

FILL FILL_3__12596_ (
);

FILL FILL_2__7343_ (
);

FILL FILL_3__12176_ (
);

FILL FILL_6__13930_ (
);

FILL FILL_4__7689_ (
);

FILL FILL_6__13510_ (
);

FILL FILL_2__11589_ (
);

FILL FILL_2__11169_ (
);

FILL FILL_5__12503_ (
);

FILL FILL_4__8630_ (
);

FILL FILL_4__11916_ (
);

FILL FILL_4__8210_ (
);

FILL FILL_5__15395_ (
);

FILL FILL_2__12530_ (
);

FILL FILL_6__8976_ (
);

FILL FILL_0__7589_ (
);

FILL FILL_2__12110_ (
);

FILL FILL_0__7169_ (
);

DFFSR _9695_ (
    .Q(\datapath_1.regfile_1.regOut[22] [9]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_1368_[9])
);

FILL SFILL13560x31050 (
);

INVX1 _9275_ (
    .A(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_1218_)
);

FILL FILL_3__10909_ (
);

FILL FILL_1__11943_ (
);

FILL FILL_4__14388_ (
);

FILL FILL_1__11523_ (
);

FILL FILL_1__11103_ (
);

FILL FILL_0__8950_ (
);

FILL FILL_2__8968_ (
);

FILL FILL_0__10936_ (
);

FILL FILL_0__8530_ (
);

FILL FILL_2__8128_ (
);

FILL FILL_0__8110_ (
);

OAI21X1 _10801_ (
    .A(_1990_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1991_),
    .Y(_1953_[19])
);

FILL FILL_0__10516_ (
);

FILL FILL_5__6973_ (
);

OAI22X1 _13693_ (
    .A(_4198_),
    .B(_3916_),
    .C(_3959_),
    .D(_4199_),
    .Y(_4200_)
);

OAI21X1 _13273_ (
    .A(_3813_),
    .B(_3811_),
    .C(_3750_),
    .Y(_3814_)
);

FILL FILL_5__13708_ (
);

FILL FILL_3__14742_ (
);

FILL FILL_3__14322_ (
);

FILL FILL_1__6965_ (
);

FILL FILL_4__9415_ (
);

FILL FILL_2__13735_ (
);

FILL FILL_2__13315_ (
);

FILL FILL_1__12728_ (
);

FILL FILL_1__12308_ (
);

FILL FILL_3__7832_ (
);

FILL FILL_0__9735_ (
);

FILL SFILL64520x8050 (
);

FILL SFILL104360x37050 (
);

FILL FILL_5__7758_ (
);

FILL FILL_2_BUFX2_insert920 (
);

FILL FILL_5__7338_ (
);

FILL FILL_2_BUFX2_insert921 (
);

FILL FILL_4__16114_ (
);

FILL FILL_2_BUFX2_insert922 (
);

FILL FILL_2_BUFX2_insert923 (
);

NOR2X1 _14898_ (
    .A(_5379_),
    .B(_5376_),
    .Y(_5380_)
);

INVX1 _14478_ (
    .A(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_4969_)
);

FILL FILL_2_BUFX2_insert924 (
);

OAI22X1 _14058_ (
    .A(_4557_),
    .B(_3905__bF$buf1),
    .C(_3972__bF$buf2),
    .D(_4556_),
    .Y(_4558_)
);

FILL FILL_2_BUFX2_insert925 (
);

FILL FILL_3__15947_ (
);

FILL FILL_2_BUFX2_insert926 (
);

FILL FILL_3__15527_ (
);

FILL FILL_2_BUFX2_insert927 (
);

FILL SFILL64200x2050 (
);

FILL FILL_3__15107_ (
);

FILL FILL_2_BUFX2_insert928 (
);

FILL FILL_1__16141_ (
);

FILL FILL_2_BUFX2_insert929 (
);

FILL FILL_3__10662_ (
);

FILL FILL_3__10242_ (
);

FILL SFILL64120x7050 (
);

FILL FILL_0__15974_ (
);

FILL FILL_0__15554_ (
);

FILL FILL_0__15134_ (
);

FILL FILL_3__8617_ (
);

FILL FILL_5__13881_ (
);

FILL FILL_5__13461_ (
);

FILL FILL_5__13041_ (
);

FILL FILL112440x43050 (
);

NAND2X1 _7761_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_453_)
);

NAND2X1 _7341_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_234_)
);

FILL FILL_4__12874_ (
);

FILL FILL_4__12454_ (
);

FILL FILL_4__12034_ (
);

NAND2X1 _10398_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1784_)
);

FILL FILL_5__9904_ (
);

FILL FILL_3__11867_ (
);

FILL FILL_3__11447_ (
);

FILL FILL_1__12481_ (
);

FILL FILL_3__11027_ (
);

FILL FILL_1__12061_ (
);

FILL FILL_0__16339_ (
);

AOI22X1 _16204_ (
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .B(_5579_),
    .C(_5649_),
    .D(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_6655_)
);

FILL FILL_0__11894_ (
);

FILL FILL_2__9086_ (
);

FILL FILL_0__11474_ (
);

FILL FILL_0__11054_ (
);

FILL FILL_5__7091_ (
);

FILL FILL_2__11801_ (
);

FILL FILL_5__14666_ (
);

FILL FILL_5__14246_ (
);

FILL FILL_3__15280_ (
);

NAND2X1 _8966_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1053_)
);

DFFSR _8546_ (
    .Q(\datapath_1.regfile_1.regOut[13] [12]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_783_[12])
);

INVX1 _8126_ (
    .A(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_635_)
);

FILL FILL_1__7083_ (
);

FILL FILL_4__13659_ (
);

FILL FILL_4__13239_ (
);

FILL FILL_2__14693_ (
);

FILL FILL_2__14273_ (
);

FILL FILL_2__7819_ (
);

FILL FILL_0__7801_ (
);

FILL FILL_1__13686_ (
);

FILL FILL_1__13266_ (
);

FILL FILL_4__14600_ (
);

FILL FILL_1_BUFX2_insert940 (
);

FILL FILL_1_BUFX2_insert941 (
);

NAND2X1 _12964_ (
    .A(vdd),
    .B(\datapath_1.rd2 [4]),
    .Y(_3628_)
);

FILL FILL_1_BUFX2_insert942 (
);

FILL FILL_3__8370_ (
);

DFFSR _12544_ (
    .Q(ALUOut[9]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3360_[9])
);

FILL FILL_0__12259_ (
);

FILL FILL_1_BUFX2_insert943 (
);

INVX1 _12124_ (
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_3136_)
);

FILL FILL_1_BUFX2_insert944 (
);

FILL FILL_1_BUFX2_insert945 (
);

FILL FILL_1_BUFX2_insert946 (
);

FILL FILL_6__16038_ (
);

FILL FILL_1_BUFX2_insert947 (
);

FILL FILL_1_BUFX2_insert948 (
);

FILL FILL_1_BUFX2_insert949 (
);

FILL SFILL94280x48050 (
);

FILL FILL_0__13620_ (
);

FILL FILL_3__16065_ (
);

FILL FILL_5__10166_ (
);

FILL FILL_2__15898_ (
);

FILL FILL_2__15478_ (
);

FILL FILL_2__15058_ (
);

FILL FILL_0__16092_ (
);

FILL FILL_2__10193_ (
);

FILL FILL_4__15805_ (
);

FILL FILL_3__9995_ (
);

FILL FILL_4__10940_ (
);

NOR2X1 _13749_ (
    .A(_4251_),
    .B(_4254_),
    .Y(_4255_)
);

FILL FILL_3__9155_ (
);

NOR2X1 _13329_ (
    .A(_3798_),
    .B(_3855_),
    .Y(\datapath_1.regfile_1.regEn [17])
);

FILL FILL_4__10520_ (
);

FILL FILL_6__7580_ (
);

FILL FILL_1__15832_ (
);

FILL FILL_1__15412_ (
);

FILL FILL_0__14825_ (
);

FILL FILL_0__14405_ (
);

FILL FILL_2__7992_ (
);

BUFX2 BUFX2_insert610 (
    .A(_5515_),
    .Y(_5515__bF$buf1)
);

FILL FILL_2__7572_ (
);

BUFX2 BUFX2_insert611 (
    .A(_5515_),
    .Y(_5515__bF$buf0)
);

BUFX2 BUFX2_insert612 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf5)
);

BUFX2 BUFX2_insert613 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf4)
);

BUFX2 BUFX2_insert614 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf3)
);

FILL FILL_4__7498_ (
);

BUFX2 BUFX2_insert615 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf2)
);

FILL FILL_4__7078_ (
);

BUFX2 BUFX2_insert616 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf1)
);

BUFX2 BUFX2_insert617 (
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf0)
);

BUFX2 BUFX2_insert618 (
    .A(_3942_),
    .Y(_3942__bF$buf3)
);

FILL FILL_2__11398_ (
);

BUFX2 BUFX2_insert619 (
    .A(_3942_),
    .Y(_3942__bF$buf2)
);

FILL FILL_5__12732_ (
);

FILL SFILL33800x9050 (
);

FILL FILL_5__12312_ (
);

FILL SFILL74280x9050 (
);

FILL FILL_4__11725_ (
);

FILL FILL_4__11305_ (
);

INVX1 _9084_ (
    .A(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_1111_)
);

FILL FILL_1__11752_ (
);

FILL FILL_4__14197_ (
);

FILL FILL_1__11332_ (
);

FILL FILL_2__8777_ (
);

FILL FILL_2__8357_ (
);

FILL FILL_0__10745_ (
);

DFFSR _10610_ (
    .Q(\datapath_1.regfile_1.regOut[29] [28]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_1823_[28])
);

FILL FILL_0__10325_ (
);

FILL FILL_6__14104_ (
);

FILL SFILL23160x59050 (
);

INVX1 _13082_ (
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_3686_)
);

FILL FILL_5__13937_ (
);

FILL FILL_3__14971_ (
);

FILL FILL_5__13517_ (
);

FILL FILL_3__14551_ (
);

FILL SFILL8600x63050 (
);

FILL FILL_3__14131_ (
);

NAND2X1 _7817_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_470_)
);

FILL FILL_4_BUFX2_insert450 (
);

FILL FILL_4_BUFX2_insert451 (
);

FILL FILL_4__9644_ (
);

FILL FILL_4__9224_ (
);

FILL FILL_4_BUFX2_insert452 (
);

FILL FILL_4_BUFX2_insert453 (
);

FILL FILL_2__13964_ (
);

FILL SFILL8680x20050 (
);

FILL FILL_4_BUFX2_insert454 (
);

FILL FILL_2__13544_ (
);

FILL FILL_2__13124_ (
);

FILL FILL_4_BUFX2_insert455 (
);

FILL FILL_4_BUFX2_insert456 (
);

FILL FILL_4_BUFX2_insert457 (
);

FILL FILL_4_BUFX2_insert458 (
);

FILL FILL_4_BUFX2_insert459 (
);

FILL FILL_1__12957_ (
);

FILL FILL_1__12117_ (
);

FILL SFILL84200x44050 (
);

FILL FILL_0__9544_ (
);

FILL FILL_3__7221_ (
);

FILL FILL_0__9124_ (
);

NOR2X1 _11815_ (
    .A(_2905_),
    .B(_2904_),
    .Y(_2906_)
);

FILL SFILL114040x58050 (
);

FILL FILL_5__7987_ (
);

FILL FILL_5__7567_ (
);

FILL FILL_4__16343_ (
);

FILL FILL_6__10444_ (
);

NAND3X1 _14287_ (
    .A(_4778_),
    .B(_4781_),
    .C(_4777_),
    .Y(_4782_)
);

FILL FILL_3__15756_ (
);

FILL FILL_3__15336_ (
);

FILL FILL_1__16370_ (
);

FILL FILL_1__7979_ (
);

FILL FILL_3__10891_ (
);

FILL FILL_1__7559_ (
);

FILL FILL_3__10051_ (
);

FILL FILL_2__14749_ (
);

FILL FILL_0__15783_ (
);

FILL FILL_2__14329_ (
);

FILL FILL_0__15363_ (
);

FILL SFILL114440x27050 (
);

FILL SFILL23880x50 (
);

FILL FILL_1__8500_ (
);

FILL FILL_3__8846_ (
);

FILL FILL_3__8006_ (
);

FILL FILL_5__13690_ (
);

FILL FILL_5__13270_ (
);

FILL SFILL74280x44050 (
);

NAND2X1 _7990_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_565_)
);

NAND2X1 _7570_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_346_)
);

DFFSR _7150_ (
    .Q(\datapath_1.regfile_1.regOut[2] [24]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_68_[24])
);

FILL FILL_4__12263_ (
);

FILL FILL_2__6843_ (
);

FILL FILL_3__11676_ (
);

FILL FILL_3__11256_ (
);

FILL FILL_1__12290_ (
);

FILL SFILL74600x56050 (
);

DFFSR _16433_ (
    .Q(\datapath_1.regfile_1.regOut[0] [16]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_6769_[16])
);

FILL FILL_0__16148_ (
);

NAND2X1 _16013_ (
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .B(_5490_),
    .Y(_6469_)
);

FILL FILL_2__10669_ (
);

FILL FILL_2__10249_ (
);

FILL FILL_0__11283_ (
);

FILL FILL_3_BUFX2_insert470 (
);

FILL FILL_4__7710_ (
);

FILL FILL_3_BUFX2_insert471 (
);

FILL FILL_3_BUFX2_insert472 (
);

FILL FILL_5__14895_ (
);

FILL FILL_5__14475_ (
);

FILL FILL_3_BUFX2_insert473 (
);

FILL FILL_2__11610_ (
);

FILL SFILL74200x42050 (
);

FILL FILL_5__14055_ (
);

FILL FILL_3_BUFX2_insert474 (
);

FILL FILL_3_BUFX2_insert475 (
);

INVX1 _8775_ (
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_966_)
);

INVX1 _8355_ (
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_747_)
);

FILL FILL_3_BUFX2_insert476 (
);

FILL FILL_3_BUFX2_insert477 (
);

FILL FILL_3_BUFX2_insert478 (
);

FILL FILL_3_BUFX2_insert479 (
);

FILL FILL_4__13888_ (
);

FILL FILL_4__13468_ (
);

FILL FILL_2__14082_ (
);

FILL FILL_0__7610_ (
);

FILL FILL_2__7628_ (
);

FILL FILL_2__7208_ (
);

FILL FILL_1__13495_ (
);

INVX1 _12773_ (
    .A(\control_1.op [0]),
    .Y(_3541_)
);

FILL FILL_0__12488_ (
);

NAND2X1 _12353_ (
    .A(MemToReg_bF$buf2),
    .B(\datapath_1.Data [3]),
    .Y(_3301_)
);

FILL FILL_0__12068_ (
);

FILL FILL_3__13822_ (
);

FILL FILL_3__13402_ (
);

FILL FILL_4__8915_ (
);

FILL FILL_3__16294_ (
);

FILL FILL_5__10395_ (
);

FILL FILL112120x62050 (
);

FILL FILL_1__8097_ (
);

FILL FILL_1__11808_ (
);

FILL FILL_2__15287_ (
);

FILL FILL_3__6912_ (
);

FILL FILL_5__16201_ (
);

FILL FILL_5__6838_ (
);

FILL FILL_4__15614_ (
);

FILL FILL_3__9384_ (
);

NOR2X1 _13978_ (
    .A(_4478_),
    .B(_3935__bF$buf1),
    .Y(_4479_)
);

NOR2X1 _13558_ (
    .A(_4064_),
    .B(_4067_),
    .Y(_4068_)
);

OAI21X1 _13138_ (
    .A(_3722_),
    .B(PCEn_bF$buf5),
    .C(_3723_),
    .Y(_3685_[19])
);

FILL FILL_3__14607_ (
);

FILL FILL_1__15641_ (
);

FILL FILL112040x69050 (
);

FILL FILL_1__15221_ (
);

FILL FILL_0__14634_ (
);

FILL FILL_0__14214_ (
);

FILL FILL_2__7381_ (
);

FILL SFILL64200x40050 (
);

FILL FILL_5__12961_ (
);

FILL FILL112440x38050 (
);

FILL FILL_5__12121_ (
);

BUFX2 _6841_ (
    .A(_1_[3]),
    .Y(memoryAddress[3])
);

FILL FILL_4__11954_ (
);

FILL FILL_4__11534_ (
);

FILL FILL_4__11114_ (
);

FILL FILL_6__8594_ (
);

FILL FILL_1__16006_ (
);

FILL FILL_3__10947_ (
);

FILL FILL_1__11981_ (
);

FILL FILL_3__10527_ (
);

FILL FILL_1__11561_ (
);

FILL FILL_3__10107_ (
);

FILL FILL_1__11141_ (
);

FILL FILL_0__15839_ (
);

AOI22X1 _15704_ (
    .A(_5481_),
    .B(\datapath_1.regfile_1.regOut[30] [16]),
    .C(\datapath_1.regfile_1.regOut[29] [16]),
    .D(_5486_),
    .Y(_6168_)
);

FILL FILL_0__15419_ (
);

FILL FILL_0__10974_ (
);

FILL FILL_2__8586_ (
);

FILL FILL_0__10554_ (
);

FILL FILL_0__10134_ (
);

FILL FILL_6__14753_ (
);

FILL FILL_5__13746_ (
);

FILL FILL_5__13326_ (
);

FILL FILL_3__14780_ (
);

FILL FILL_3__14360_ (
);

INVX1 _7626_ (
    .A(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_383_)
);

INVX1 _7206_ (
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_164_)
);

FILL FILL_4__9873_ (
);

FILL FILL_4__12739_ (
);

FILL FILL_4__9033_ (
);

FILL FILL_2__13773_ (
);

FILL FILL_4__12319_ (
);

FILL FILL_2__13353_ (
);

FILL FILL_6__9379_ (
);

FILL FILL_1__12766_ (
);

FILL FILL_1__12346_ (
);

FILL FILL_3__7870_ (
);

FILL FILL_0__9773_ (
);

FILL FILL_0__9353_ (
);

FILL FILL_3__7450_ (
);

FILL FILL_0__11759_ (
);

FILL FILL_3__7030_ (
);

FILL FILL_0__11339_ (
);

OAI21X1 _11624_ (
    .A(_2254_),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .C(_2728_),
    .Y(_2729_)
);

NOR2X1 _11204_ (
    .A(_2322_),
    .B(_2321_),
    .Y(_2323_)
);

FILL FILL_5__7376_ (
);

FILL FILL_4__16152_ (
);

NOR2X1 _14096_ (
    .A(_4594_),
    .B(_4584_),
    .Y(_4595_)
);

FILL SFILL103560x80050 (
);

FILL FILL_3__15985_ (
);

FILL FILL_0__12700_ (
);

FILL FILL_3__15565_ (
);

FILL FILL_3__15145_ (
);

FILL FILL_1__7368_ (
);

FILL FILL_3__10280_ (
);

FILL FILL_2__14978_ (
);

FILL FILL_2__14558_ (
);

FILL FILL_2__14138_ (
);

FILL FILL_0__15592_ (
);

FILL FILL_0__15172_ (
);

FILL SFILL13640x4050 (
);

FILL FILL_3__8655_ (
);

FILL FILL_3__8235_ (
);

INVX1 _12829_ (
    .A(\datapath_1.a [2]),
    .Y(_3558_)
);

INVX1 _12409_ (
    .A(ALUOut[22]),
    .Y(_3338_)
);

FILL FILL_1__14912_ (
);

FILL FILL_4__12492_ (
);

FILL FILL_4__12072_ (
);

FILL FILL_0__13905_ (
);

FILL FILL_5__9522_ (
);

FILL FILL_3__11485_ (
);

FILL FILL_5__9102_ (
);

FILL FILL_3__11065_ (
);

FILL FILL_0__16377_ (
);

NAND2X1 _16242_ (
    .A(_6687_),
    .B(_6692_),
    .Y(_6693_)
);

FILL FILL_2__10898_ (
);

FILL FILL_2__10058_ (
);

FILL FILL_0__11092_ (
);

FILL FILL_1__9934_ (
);

FILL FILL_5__11812_ (
);

FILL FILL_1__9514_ (
);

FILL FILL_6__15291_ (
);

FILL FILL_4__10805_ (
);

FILL FILL_0__6898_ (
);

FILL FILL_5__14284_ (
);

INVX1 _8584_ (
    .A(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_859_)
);

DFFSR _8164_ (
    .Q(\datapath_1.regfile_1.regOut[10] [14]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_588_[14])
);

FILL FILL_1__10832_ (
);

FILL FILL_4__13697_ (
);

FILL FILL_4__13277_ (
);

FILL FILL_1__10412_ (
);

FILL FILL_2__7857_ (
);

FILL FILL_2__7437_ (
);

INVX1 _12582_ (
    .A(\datapath_1.Data [5]),
    .Y(_3434_)
);

FILL FILL_0__12297_ (
);

OAI21X1 _12162_ (
    .A(_3160_),
    .B(ALUSrcA_bF$buf7),
    .C(_3161_),
    .Y(\datapath_1.alu_1.ALUInA [15])
);

FILL SFILL8600x58050 (
);

FILL FILL_3__13631_ (
);

FILL FILL_3__13211_ (
);

FILL FILL_4__8724_ (
);

FILL SFILL8680x15050 (
);

FILL SFILL13720x52050 (
);

FILL FILL_2__12624_ (
);

FILL FILL_5__15489_ (
);

FILL FILL_2__12204_ (
);

FILL FILL_5__15069_ (
);

OAI21X1 _9789_ (
    .A(_1478_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .C(_1479_),
    .Y(_1433_[23])
);

OAI21X1 _9369_ (
    .A(_1259_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .C(_1260_),
    .Y(_1238_[11])
);

FILL SFILL109560x32050 (
);

FILL FILL_1__11617_ (
);

FILL SFILL53800x48050 (
);

FILL FILL_2__15096_ (
);

FILL SFILL84200x39050 (
);

FILL FILL_5__16010_ (
);

FILL FILL_0__8624_ (
);

FILL FILL_0__8204_ (
);

FILL FILL_1__14089_ (
);

FILL FILL_4__15843_ (
);

FILL FILL_4__15423_ (
);

FILL FILL_4__15003_ (
);

NAND2X1 _13787_ (
    .A(_4292_),
    .B(_4285_),
    .Y(_4293_)
);

AND2X2 _13367_ (
    .A(_3878_),
    .B(\datapath_1.PCJump [18]),
    .Y(_3879_)
);

FILL FILL_3__14836_ (
);

FILL SFILL109480x39050 (
);

FILL FILL_1__15870_ (
);

FILL FILL_3__14416_ (
);

FILL FILL_1__15450_ (
);

FILL FILL_1__15030_ (
);

FILL FILL_4__9929_ (
);

FILL FILL_4__9509_ (
);

FILL SFILL8600x13050 (
);

FILL FILL_2__13829_ (
);

FILL FILL_0__14863_ (
);

FILL FILL_2__13409_ (
);

FILL FILL_0__14443_ (
);

FILL FILL_0__14023_ (
);

FILL FILL_2__7190_ (
);

CLKBUF1 CLKBUF1_insert150 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf74)
);

CLKBUF1 CLKBUF1_insert151 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf73)
);

CLKBUF1 CLKBUF1_insert152 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf72)
);

FILL FILL_3__7926_ (
);

CLKBUF1 CLKBUF1_insert153 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf71)
);

FILL FILL_3__7506_ (
);

CLKBUF1 CLKBUF1_insert154 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf70)
);

FILL FILL_0__9409_ (
);

CLKBUF1 CLKBUF1_insert155 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert156 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf68)
);

FILL FILL_5__12770_ (
);

CLKBUF1 CLKBUF1_insert157 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf67)
);

FILL FILL_5__12350_ (
);

CLKBUF1 CLKBUF1_insert158 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert159 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf65)
);

FILL FILL_4__16208_ (
);

FILL FILL_4__11763_ (
);

FILL FILL_4__11343_ (
);

FILL SFILL13640x14050 (
);

FILL FILL_1__16235_ (
);

FILL FILL_3__10756_ (
);

FILL FILL_1__11790_ (
);

FILL FILL_1__11370_ (
);

FILL FILL_0__15648_ (
);

NOR2X1 _15933_ (
    .A(_6390_),
    .B(_6388_),
    .Y(_6391_)
);

FILL FILL_0__15228_ (
);

NAND3X1 _15513_ (
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf3),
    .Y(_5982_)
);

FILL SFILL38840x63050 (
);

FILL FILL_2__8395_ (
);

FILL FILL_0__10783_ (
);

FILL FILL_0__10363_ (
);

FILL SFILL43800x46050 (
);

FILL FILL_5__13975_ (
);

FILL SFILL74200x37050 (
);

FILL FILL_5__13555_ (
);

FILL FILL_5__13135_ (
);

INVX1 _7855_ (
    .A(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_495_)
);

INVX1 _7435_ (
    .A(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_276_)
);

FILL FILL_4_BUFX2_insert830 (
);

DFFSR _7015_ (
    .Q(\datapath_1.regfile_1.regOut[1] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_3_[17])
);

FILL FILL_4_BUFX2_insert831 (
);

FILL FILL_4__9682_ (
);

FILL FILL_4_BUFX2_insert832 (
);

FILL FILL_4__9262_ (
);

FILL FILL_4__12968_ (
);

FILL FILL_4_BUFX2_insert833 (
);

FILL FILL_4__12128_ (
);

FILL FILL_4_BUFX2_insert834 (
);

FILL FILL_2__13582_ (
);

FILL FILL_4_BUFX2_insert835 (
);

FILL FILL_2__13162_ (
);

FILL FILL_4_BUFX2_insert836 (
);

FILL FILL_4_BUFX2_insert837 (
);

FILL FILL_4_BUFX2_insert838 (
);

FILL FILL_4_BUFX2_insert839 (
);

FILL FILL_1__12995_ (
);

FILL SFILL43400x32050 (
);

FILL FILL112200x50050 (
);

FILL FILL_1__12575_ (
);

FILL FILL_1__12155_ (
);

FILL FILL_0__11988_ (
);

FILL FILL_0__9162_ (
);

NAND3X1 _11853_ (
    .A(_2849_),
    .B(_2892_),
    .C(_2939_),
    .Y(_2940_)
);

FILL FILL_0__11568_ (
);

FILL FILL_0__11148_ (
);

OAI21X1 _11433_ (
    .A(_2547_),
    .B(_2548_),
    .C(_2422_),
    .Y(_2549_)
);

NAND2X1 _11013_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2132_)
);

FILL FILL_3__12902_ (
);

FILL FILL_6__15347_ (
);

FILL FILL_5__7185_ (
);

FILL FILL_4__16381_ (
);

FILL FILL_6__10062_ (
);

FILL FILL_3__15794_ (
);

FILL FILL_3__15374_ (
);

FILL FILL112120x57050 (
);

FILL FILL_1__7597_ (
);

FILL FILL_1__7177_ (
);

FILL FILL_2__14787_ (
);

FILL FILL_2__14367_ (
);

FILL FILL_5__15701_ (
);

FILL FILL_3__8884_ (
);

FILL FILL_3__8464_ (
);

OAI21X1 _12638_ (
    .A(_3470_),
    .B(vdd),
    .C(_3471_),
    .Y(_3425_[23])
);

NAND3X1 _12218_ (
    .A(_3197_),
    .B(_3199_),
    .C(_3202_),
    .Y(\datapath_1.alu_1.ALUInB [0])
);

FILL FILL_1__14721_ (
);

FILL FILL_1__14301_ (
);

FILL FILL_6__11267_ (
);

FILL FILL_0__13714_ (
);

FILL FILL_3__16159_ (
);

FILL FILL_2__6881_ (
);

FILL FILL_5__9751_ (
);

FILL SFILL89880x55050 (
);

FILL FILL_3__11294_ (
);

FILL FILL112120x12050 (
);

FILL FILL_0__16186_ (
);

INVX1 _16051_ (
    .A(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_6506_)
);

FILL FILL_2__10287_ (
);

FILL FILL_1__9743_ (
);

FILL FILL_5__11621_ (
);

FILL FILL_5__11201_ (
);

FILL FILL_3__9669_ (
);

FILL FILL_3_BUFX2_insert850 (
);

FILL FILL_3__9249_ (
);

FILL FILL_3_BUFX2_insert851 (
);

FILL FILL_3_BUFX2_insert852 (
);

FILL FILL_4__10614_ (
);

FILL FILL_3_BUFX2_insert853 (
);

FILL FILL_3_BUFX2_insert854 (
);

FILL FILL_5__14093_ (
);

FILL FILL_1__15926_ (
);

FILL FILL_3_BUFX2_insert855 (
);

FILL FILL_6__7674_ (
);

FILL FILL_3_BUFX2_insert856 (
);

FILL FILL_1__15506_ (
);

OAI21X1 _8393_ (
    .A(_771_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_772_),
    .Y(_718_[27])
);

FILL FILL_3_BUFX2_insert857 (
);

FILL FILL_3_BUFX2_insert858 (
);

FILL FILL_3_BUFX2_insert859 (
);

FILL FILL_1__10641_ (
);

FILL FILL112040x19050 (
);

FILL FILL_4__13086_ (
);

FILL FILL_0__14919_ (
);

FILL FILL_2__7246_ (
);

FILL FILL_3__12499_ (
);

FILL FILL_3__12079_ (
);

FILL FILL_6__13833_ (
);

FILL FILL_6__13413_ (
);

FILL SFILL89880x10050 (
);

INVX1 _12391_ (
    .A(ALUOut[16]),
    .Y(_3326_)
);

FILL FILL_5__12826_ (
);

FILL FILL_5__12406_ (
);

FILL FILL_3__13860_ (
);

FILL FILL_3__13440_ (
);

FILL FILL_3__13020_ (
);

FILL FILL_4__8953_ (
);

FILL FILL_4__8533_ (
);

FILL FILL_4__8113_ (
);

FILL FILL_4__11819_ (
);

FILL FILL_2__12853_ (
);

FILL FILL_5__15298_ (
);

FILL FILL_2__12433_ (
);

FILL FILL_2__12013_ (
);

FILL FILL_6__8459_ (
);

OAI21X1 _9598_ (
    .A(_1371_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .C(_1372_),
    .Y(_1368_[2])
);

DFFSR _9178_ (
    .Q(\datapath_1.regfile_1.regOut[18] [4]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1108_[4])
);

FILL FILL_1__11846_ (
);

FILL FILL_1__11426_ (
);

FILL FILL_1__11006_ (
);

FILL FILL_3__6950_ (
);

FILL FILL_0__8853_ (
);

FILL SFILL79080x70050 (
);

FILL FILL_0__8013_ (
);

FILL FILL_6__9400_ (
);

FILL FILL_0__10419_ (
);

INVX1 _10704_ (
    .A(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_1947_)
);

FILL FILL_0_BUFX2_insert980 (
);

FILL FILL_5__6876_ (
);

FILL FILL_4__15652_ (
);

FILL FILL_0_BUFX2_insert981 (
);

FILL FILL_4__15232_ (
);

FILL FILL_0_BUFX2_insert982 (
);

FILL SFILL54200x33050 (
);

FILL FILL_0_BUFX2_insert983 (
);

FILL FILL_0_BUFX2_insert984 (
);

INVX1 _13596_ (
    .A(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_4105_)
);

FILL FILL_0_BUFX2_insert985 (
);

FILL FILL_0_BUFX2_insert986 (
);

DFFSR _13176_ (
    .Q(\datapath_1.mux_iord.din0 [1]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[1])
);

FILL FILL_2__9812_ (
);

FILL FILL_0_BUFX2_insert987 (
);

FILL FILL_0_BUFX2_insert988 (
);

FILL FILL_3__14645_ (
);

FILL FILL_3__14225_ (
);

FILL FILL_0_BUFX2_insert989 (
);

FILL FILL_1__6868_ (
);

FILL FILL_4__9738_ (
);

FILL FILL_2__13638_ (
);

FILL FILL_2__13218_ (
);

FILL FILL_0__14672_ (
);

FILL FILL_0__14252_ (
);

FILL SFILL23720x49050 (
);

FILL FILL_3__7735_ (
);

FILL FILL_0__9638_ (
);

FILL FILL_0__9218_ (
);

NAND2X1 _11909_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[7]),
    .Y(_2981_)
);

FILL FILL_3__7315_ (
);

FILL FILL_4__16017_ (
);

FILL SFILL44200x76050 (
);

FILL FILL_4__11992_ (
);

FILL FILL_6__10538_ (
);

FILL FILL_4__11572_ (
);

FILL FILL_4__11152_ (
);

FILL FILL_1__16044_ (
);

FILL FILL_5__8602_ (
);

FILL FILL_3__10565_ (
);

FILL FILL_3__10145_ (
);

FILL FILL_6_BUFX2_insert362 (
);

FILL FILL_0__15877_ (
);

AOI21X1 _15742_ (
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .B(_5494_),
    .C(_6204_),
    .Y(_6205_)
);

FILL FILL_0__15457_ (
);

OAI22X1 _15322_ (
    .A(_5472__bF$buf3),
    .B(_4287_),
    .C(_4286_),
    .D(_5552__bF$buf2),
    .Y(_5796_)
);

FILL FILL_0__15037_ (
);

FILL FILL_6_BUFX2_insert367 (
);

FILL FILL_0__10172_ (
);

FILL FILL_5__13784_ (
);

FILL FILL_5__13364_ (
);

FILL FILL_6__6945_ (
);

DFFSR _7664_ (
    .Q(\datapath_1.regfile_1.regOut[6] [26]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_328_[26])
);

OAI21X1 _7244_ (
    .A(_188_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .C(_189_),
    .Y(_133_[28])
);

FILL FILL_4__9491_ (
);

FILL FILL_4__12777_ (
);

FILL FILL_4__12357_ (
);

FILL FILL_2__13391_ (
);

FILL FILL_2__6937_ (
);

FILL FILL_5__9807_ (
);

FILL FILL_1__12384_ (
);

INVX1 _16107_ (
    .A(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_6561_)
);

FILL FILL_0__9391_ (
);

FILL FILL_0__11797_ (
);

FILL FILL_0__11377_ (
);

NOR2X1 _11662_ (
    .A(_2205_),
    .B(_2742_),
    .Y(_2764_)
);

OAI21X1 _11242_ (
    .A(_2355_),
    .B(_2132_),
    .C(_2122_),
    .Y(_2361_)
);

FILL FILL_3__12711_ (
);

FILL FILL_4__16190_ (
);

FILL FILL_4__7804_ (
);

FILL SFILL13720x47050 (
);

FILL FILL_5__14989_ (
);

FILL FILL_5__14569_ (
);

FILL FILL_2__11704_ (
);

FILL FILL_5__14149_ (
);

OAI21X1 _8869_ (
    .A(_1007_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1008_),
    .Y(_978_[15])
);

FILL FILL_3__15183_ (
);

FILL SFILL109560x27050 (
);

OAI21X1 _8449_ (
    .A(_788_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .C(_789_),
    .Y(_783_[3])
);

DFFSR _8029_ (
    .Q(\datapath_1.regfile_1.regOut[9] [7]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_523_[7])
);

FILL FILL_2__14596_ (
);

FILL FILL_2__14176_ (
);

FILL FILL_5__15930_ (
);

FILL FILL_5__15510_ (
);

FILL FILL_0__7704_ (
);

OAI21X1 _9810_ (
    .A(_1492_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .C(_1493_),
    .Y(_1433_[30])
);

FILL FILL_1__13589_ (
);

FILL FILL_1__13169_ (
);

FILL FILL_4__14923_ (
);

FILL FILL_4__14503_ (
);

OAI21X1 _12867_ (
    .A(_3582_),
    .B(vdd),
    .C(_3583_),
    .Y(_3555_[14])
);

FILL FILL_3__8273_ (
);

OAI21X1 _12447_ (
    .A(_3363_),
    .B(vdd),
    .C(_3364_),
    .Y(_3360_[2])
);

NAND3X1 _12027_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[10]),
    .C(_3032__bF$buf3),
    .Y(_3066_)
);

FILL FILL_3__13916_ (
);

FILL FILL_1__14950_ (
);

FILL FILL_1__14530_ (
);

FILL FILL_5__8199_ (
);

FILL FILL_1__14110_ (
);

FILL FILL_5_BUFX2_insert380 (
);

FILL FILL_5_BUFX2_insert381 (
);

FILL FILL_2__12909_ (
);

FILL FILL_5_BUFX2_insert382 (
);

FILL FILL_0__13943_ (
);

FILL FILL_3__16388_ (
);

FILL FILL_5_BUFX2_insert383 (
);

FILL FILL_0__13523_ (
);

FILL FILL_0__13103_ (
);

FILL FILL_5_BUFX2_insert384 (
);

FILL FILL_5_BUFX2_insert385 (
);

FILL FILL_5_BUFX2_insert386 (
);

FILL FILL_5__9980_ (
);

FILL FILL_5__10489_ (
);

FILL FILL_5__10069_ (
);

FILL FILL_5_BUFX2_insert387 (
);

FILL FILL_5_BUFX2_insert388 (
);

FILL FILL_5__9140_ (
);

FILL FILL_5_BUFX2_insert389 (
);

NOR2X1 _16280_ (
    .A(_6726_),
    .B(_6729_),
    .Y(_6730_)
);

FILL FILL_0__8909_ (
);

FILL FILL_5__11850_ (
);

FILL FILL_1__9552_ (
);

FILL FILL_5__11430_ (
);

FILL FILL_1__9132_ (
);

FILL FILL_5__11010_ (
);

FILL FILL_4__15708_ (
);

FILL FILL_2__16322_ (
);

FILL FILL_3__9898_ (
);

FILL FILL_3__9478_ (
);

FILL FILL_4__10423_ (
);

FILL FILL_4__10003_ (
);

FILL FILL_1__15735_ (
);

FILL FILL_1__15315_ (
);

FILL FILL_1__10870_ (
);

FILL FILL_1__10450_ (
);

FILL FILL_1__10030_ (
);

FILL FILL_0__14728_ (
);

FILL FILL_0__14308_ (
);

FILL SFILL38840x58050 (
);

FILL FILL_2__7475_ (
);

FILL FILL_2__7055_ (
);

FILL FILL_5__12635_ (
);

FILL FILL_5__12215_ (
);

INVX1 _6935_ (
    .A(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_24_)
);

FILL FILL_4__8762_ (
);

FILL FILL_4__8342_ (
);

FILL FILL_4__11628_ (
);

FILL FILL_2__12662_ (
);

FILL FILL_4__11208_ (
);

FILL FILL_2__12242_ (
);

FILL SFILL99480x38050 (
);

FILL FILL_1__11655_ (
);

FILL FILL_1__11235_ (
);

INVX1 _10933_ (
    .A(\control_1.op [3]),
    .Y(_2067_)
);

FILL FILL_0__10648_ (
);

FILL FILL_0__8242_ (
);

INVX1 _10513_ (
    .A(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_1840_)
);

FILL SFILL68600x76050 (
);

FILL FILL_4__15881_ (
);

FILL FILL_6__14007_ (
);

FILL FILL_4__15461_ (
);

FILL FILL_4__15041_ (
);

FILL FILL_3__14874_ (
);

FILL FILL_2__9621_ (
);

FILL FILL_3__14454_ (
);

FILL FILL_3__14034_ (
);

FILL FILL_4__9547_ (
);

FILL FILL_3_CLKBUF1_insert1074 (
);

FILL FILL_4__9127_ (
);

FILL FILL_3_CLKBUF1_insert1075 (
);

FILL FILL_2__13867_ (
);

FILL FILL_3_CLKBUF1_insert1076 (
);

FILL FILL_3_CLKBUF1_insert1077 (
);

FILL FILL_2__13447_ (
);

FILL FILL_3_CLKBUF1_insert1078 (
);

FILL FILL_0__14481_ (
);

FILL FILL_2__13027_ (
);

FILL FILL_0__14061_ (
);

FILL FILL_3_CLKBUF1_insert1079 (
);

FILL FILL_0__9867_ (
);

FILL FILL_3__7964_ (
);

FILL FILL_3__7544_ (
);

FILL FILL_3__7124_ (
);

INVX1 _11718_ (
    .A(_2816_),
    .Y(\datapath_1.ALUResult [11])
);

FILL FILL_0__9027_ (
);

FILL FILL_1__13801_ (
);

FILL SFILL3480x12050 (
);

FILL FILL_4__16246_ (
);

FILL FILL_4__11381_ (
);

FILL FILL_3__15659_ (
);

FILL FILL_3__15239_ (
);

FILL FILL_1__16273_ (
);

FILL FILL_5__8831_ (
);

FILL FILL_3__10794_ (
);

FILL FILL_3__10374_ (
);

INVX1 _15971_ (
    .A(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_6428_)
);

FILL FILL_0__15686_ (
);

OAI22X1 _15551_ (
    .A(_4541_),
    .B(_5501_),
    .C(_5524__bF$buf0),
    .D(_4526_),
    .Y(_6019_)
);

FILL FILL_0__15266_ (
);

INVX1 _15131_ (
    .A(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_5609_)
);

FILL FILL_5__10701_ (
);

FILL FILL_1__8823_ (
);

FILL FILL_1__8403_ (
);

FILL FILL_6__14180_ (
);

FILL FILL_3__8749_ (
);

FILL FILL_3__8329_ (
);

FILL FILL_5__13593_ (
);

FILL FILL_5__13173_ (
);

OAI21X1 _7893_ (
    .A(_519_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .C(_520_),
    .Y(_458_[31])
);

OAI21X1 _7473_ (
    .A(_300_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .C(_301_),
    .Y(_263_[19])
);

OAI21X1 _7053_ (
    .A(_81_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .C(_82_),
    .Y(_68_[7])
);

FILL FILL_4__12586_ (
);

FILL SFILL28840x11050 (
);

FILL FILL_4__12166_ (
);

FILL FILL_3__11999_ (
);

FILL FILL_5__9616_ (
);

FILL FILL_3__11579_ (
);

FILL FILL_3__11159_ (
);

FILL FILL_1__12193_ (
);

FILL FILL_6__12913_ (
);

INVX1 _16336_ (
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_6778_)
);

NAND2X1 _11891_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[1]),
    .Y(_2969_)
);

FILL FILL_0__11186_ (
);

AOI21X1 _11471_ (
    .A(_2554_),
    .B(_2549_),
    .C(_2443_),
    .Y(_2586_)
);

FILL FILL_5__11906_ (
);

NOR2X1 _11051_ (
    .A(_2168_),
    .B(_2169_),
    .Y(_2170_)
);

FILL FILL_1__9608_ (
);

FILL FILL_3__12520_ (
);

FILL FILL_3__12100_ (
);

FILL SFILL79480x79050 (
);

FILL FILL_4__7613_ (
);

FILL FILL_2__11933_ (
);

FILL FILL_5__14798_ (
);

FILL FILL_5__14378_ (
);

FILL FILL_2__11513_ (
);

DFFSR _8678_ (
    .Q(\datapath_1.regfile_1.regOut[14] [16]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_848_[16])
);

NAND2X1 _8258_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_703_)
);

FILL FILL_1__10926_ (
);

FILL FILL_1__10506_ (
);

FILL SFILL18840x54050 (
);

FILL FILL_0__7933_ (
);

FILL FILL_1__13398_ (
);

FILL FILL_4__14732_ (
);

FILL SFILL54200x28050 (
);

FILL FILL_4__14312_ (
);

DFFSR _12676_ (
    .Q(\datapath_1.Data [13]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3425_[13])
);

FILL FILL_3__8082_ (
);

NAND3X1 _12256_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [12]),
    .C(_3198__bF$buf3),
    .Y(_3231_)
);

FILL FILL_3__13725_ (
);

FILL FILL_3__13305_ (
);

FILL FILL_2__12718_ (
);

FILL FILL_0__13752_ (
);

FILL FILL_0__13332_ (
);

FILL FILL_3__16197_ (
);

FILL FILL_5__10298_ (
);

FILL FILL_0__8718_ (
);

FILL FILL_5__16104_ (
);

FILL FILL_1__9781_ (
);

FILL FILL_1__9361_ (
);

FILL FILL_4__15937_ (
);

FILL FILL_4__15517_ (
);

FILL FILL_2__16131_ (
);

FILL FILL_3__9287_ (
);

FILL FILL_4__10652_ (
);

FILL FILL_4__10232_ (
);

FILL FILL_1__15964_ (
);

FILL FILL_1__15544_ (
);

FILL FILL_1__15124_ (
);

FILL FILL_0__14957_ (
);

NAND3X1 _14822_ (
    .A(_5304_),
    .B(_5305_),
    .C(_5303_),
    .Y(_5306_)
);

FILL FILL_0__14537_ (
);

AOI21X1 _14402_ (
    .A(_4873_),
    .B(_4894_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [19])
);

FILL FILL_0__14117_ (
);

FILL FILL_5__12864_ (
);

FILL FILL_5__12444_ (
);

FILL FILL_5__12024_ (
);

FILL SFILL69080x63050 (
);

FILL FILL_4__8991_ (
);

FILL FILL_4__8571_ (
);

FILL FILL_4__11857_ (
);

FILL SFILL48920x48050 (
);

FILL FILL_2__12891_ (
);

FILL FILL_4__11437_ (
);

FILL FILL_2__12471_ (
);

FILL FILL_4__11017_ (
);

FILL FILL_2__12051_ (
);

FILL FILL_6__8077_ (
);

FILL FILL_1__16329_ (
);

FILL FILL_1__11884_ (
);

FILL FILL_1__11464_ (
);

FILL FILL_1__11044_ (
);

NOR2X1 _15607_ (
    .A(_6070_),
    .B(_6073_),
    .Y(_6074_)
);

FILL FILL_0__8891_ (
);

FILL FILL_0__8471_ (
);

FILL FILL_0__10877_ (
);

FILL FILL_2__8489_ (
);

INVX1 _10742_ (
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_2016_)
);

FILL FILL_2__8069_ (
);

FILL FILL_0__10037_ (
);

OAI21X1 _10322_ (
    .A(_1752_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .C(_1753_),
    .Y(_1693_[30])
);

FILL FILL_6__14656_ (
);

FILL FILL_4__15690_ (
);

FILL FILL_4__15270_ (
);

FILL FILL_5__13649_ (
);

FILL FILL_2__9850_ (
);

FILL FILL_5__13229_ (
);

FILL FILL_3__14683_ (
);

OAI21X1 _7949_ (
    .A(_536_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .C(_537_),
    .Y(_523_[7])
);

FILL FILL_3__14263_ (
);

FILL FILL_2__9010_ (
);

DFFSR _7529_ (
    .Q(\datapath_1.regfile_1.regOut[5] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_263_[19])
);

NAND2X1 _7109_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_120_)
);

FILL FILL_4__9776_ (
);

FILL FILL_4__9356_ (
);

FILL FILL_2__13676_ (
);

FILL FILL_2__13256_ (
);

FILL FILL_0__14290_ (
);

FILL FILL_1__12249_ (
);

FILL SFILL3640x83050 (
);

FILL FILL_0__9676_ (
);

FILL FILL_0__9256_ (
);

INVX1 _11947_ (
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3006_)
);

FILL FILL_3__7353_ (
);

OAI21X1 _11527_ (
    .A(_2637_),
    .B(_2280_),
    .C(_2411_),
    .Y(_2638_)
);

NOR2X1 _11107_ (
    .A(_2220_),
    .B(_2225_),
    .Y(_2226_)
);

FILL FILL_5__7699_ (
);

FILL FILL_1__13610_ (
);

FILL FILL_4__16055_ (
);

FILL FILL_6__10996_ (
);

FILL FILL_4__11190_ (
);

FILL FILL_3__15888_ (
);

FILL FILL_0__12603_ (
);

FILL FILL_3__15468_ (
);

FILL FILL_3__15048_ (
);

FILL FILL_1__16082_ (
);

FILL FILL_5__8640_ (
);

FILL FILL_5__8220_ (
);

FILL FILL_6_BUFX2_insert741 (
);

FILL FILL_3__10183_ (
);

OAI22X1 _15780_ (
    .A(_5569_),
    .B(_4843_),
    .C(_5483__bF$buf1),
    .D(_4840_),
    .Y(_6242_)
);

FILL FILL_0__15495_ (
);

AOI21X1 _15360_ (
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .B(_5570__bF$buf3),
    .C(_5832_),
    .Y(_5833_)
);

FILL FILL_0__15075_ (
);

FILL FILL_6_BUFX2_insert746 (
);

FILL SFILL38920x46050 (
);

FILL FILL_5__10930_ (
);

FILL FILL_5__10510_ (
);

FILL FILL_1__8632_ (
);

FILL FILL_1__8212_ (
);

FILL FILL_2__15822_ (
);

FILL FILL_2__15402_ (
);

FILL FILL_3__8978_ (
);

FILL FILL_3__8138_ (
);

FILL FILL_1__14815_ (
);

DFFSR _7282_ (
    .Q(\datapath_1.regfile_1.regOut[3] [28]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_133_[28])
);

FILL FILL_4__12395_ (
);

FILL FILL_0__13808_ (
);

FILL FILL_2__6975_ (
);

FILL FILL_5__9425_ (
);

FILL FILL_3__11388_ (
);

FILL FILL_5__9005_ (
);

FILL FILL_6__12722_ (
);

INVX1 _16145_ (
    .A(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_6598_)
);

FILL SFILL3560x45050 (
);

INVX1 _11280_ (
    .A(_2398_),
    .Y(_2399_)
);

FILL SFILL24200x67050 (
);

FILL FILL_5__11715_ (
);

FILL FILL_1__9417_ (
);

FILL FILL_4__7842_ (
);

FILL FILL_4__7422_ (
);

FILL FILL_4__10708_ (
);

FILL FILL_2__11742_ (
);

FILL FILL_5__14187_ (
);

FILL FILL_2__11322_ (
);

NAND2X1 _8487_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_815_)
);

FILL FILL_6__7348_ (
);

NAND2X1 _8067_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_596_)
);

FILL FILL_1__10315_ (
);

FILL FILL_0__7742_ (
);

FILL FILL_0__7322_ (
);

FILL FILL_4__14961_ (
);

FILL FILL_4__14541_ (
);

FILL FILL_4__14121_ (
);

FILL SFILL69240x7050 (
);

NAND2X1 _12485_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [15]),
    .Y(_3390_)
);

AOI22X1 _12065_ (
    .A(\datapath_1.ALUResult [19]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3095_)
);

FILL FILL_3__13954_ (
);

FILL FILL_2__8701_ (
);

FILL FILL_3__13534_ (
);

FILL FILL_3__13114_ (
);

FILL FILL_4__8627_ (
);

FILL FILL_4__8207_ (
);

FILL FILL_5_BUFX2_insert760 (
);

FILL FILL_5_BUFX2_insert761 (
);

FILL SFILL68600x4050 (
);

FILL FILL_2__12527_ (
);

FILL FILL_0__13981_ (
);

FILL FILL_5_BUFX2_insert762 (
);

FILL FILL_5_BUFX2_insert763 (
);

FILL FILL_2__12107_ (
);

FILL FILL_0__13561_ (
);

FILL FILL_5_BUFX2_insert764 (
);

FILL FILL_0__13141_ (
);

FILL FILL_5_BUFX2_insert765 (
);

FILL FILL_5_BUFX2_insert766 (
);

FILL FILL_5_BUFX2_insert767 (
);

FILL FILL_5_BUFX2_insert768 (
);

FILL FILL_5_BUFX2_insert769 (
);

FILL FILL_5__16333_ (
);

FILL FILL_0__8527_ (
);

FILL FILL_0__8107_ (
);

FILL FILL_1__9590_ (
);

FILL FILL_1__9170_ (
);

FILL FILL_4__15746_ (
);

FILL FILL_4__15326_ (
);

FILL FILL_2__16360_ (
);

FILL FILL_3__9096_ (
);

FILL FILL_4__10881_ (
);

FILL FILL_4__10041_ (
);

FILL FILL_2__9906_ (
);

FILL FILL_3__14739_ (
);

FILL FILL_3__14319_ (
);

FILL FILL_1__15773_ (
);

FILL FILL_1__15353_ (
);

FILL FILL_0__14766_ (
);

INVX1 _14631_ (
    .A(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_5119_)
);

FILL FILL_0__14346_ (
);

OAI22X1 _14211_ (
    .A(_3947__bF$buf3),
    .B(_4707_),
    .C(_3971__bF$buf4),
    .D(_4706_),
    .Y(_4708_)
);

FILL FILL_2__7093_ (
);

FILL FILL_6__13260_ (
);

FILL FILL_3__7829_ (
);

FILL SFILL113640x15050 (
);

FILL FILL_5__12253_ (
);

OAI21X1 _6973_ (
    .A(_48_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .C(_49_),
    .Y(_3_[23])
);

FILL FILL_2_BUFX2_insert890 (
);

FILL FILL_2_BUFX2_insert891 (
);

FILL FILL_2_BUFX2_insert892 (
);

FILL FILL_2_BUFX2_insert893 (
);

FILL FILL_4__8380_ (
);

FILL FILL_2_BUFX2_insert894 (
);

FILL FILL_4__11666_ (
);

FILL SFILL94360x73050 (
);

FILL FILL_2_BUFX2_insert895 (
);

FILL FILL_4__11246_ (
);

FILL FILL_2_BUFX2_insert896 (
);

FILL FILL_2__12280_ (
);

FILL FILL_2_BUFX2_insert897 (
);

FILL FILL_2_BUFX2_insert898 (
);

FILL FILL_2_BUFX2_insert899 (
);

FILL FILL_1__16138_ (
);

FILL FILL_3__10659_ (
);

FILL FILL_3__10239_ (
);

FILL FILL_1__11693_ (
);

FILL FILL_1__11273_ (
);

OAI21X1 _15836_ (
    .A(_6295_),
    .B(_5535__bF$buf3),
    .C(_6296_),
    .Y(_6297_)
);

NOR2X1 _15416_ (
    .A(_4392_),
    .B(_5534__bF$buf1),
    .Y(_5887_)
);

FILL FILL_0__10686_ (
);

NAND2X1 _10971_ (
    .A(_2096_),
    .B(_2045_),
    .Y(\control_1.next [3])
);

FILL SFILL79160x53050 (
);

OAI21X1 _10551_ (
    .A(_1864_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .C(_1865_),
    .Y(_1823_[21])
);

FILL FILL_0__10266_ (
);

OAI21X1 _10131_ (
    .A(_1645_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .C(_1646_),
    .Y(_1628_[9])
);

FILL FILL_3__11600_ (
);

FILL FILL_5__13878_ (
);

FILL FILL_5__13458_ (
);

FILL FILL_3__14492_ (
);

FILL FILL_5__13038_ (
);

NAND2X1 _7758_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_451_)
);

FILL FILL_3__14072_ (
);

NAND2X1 _7338_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_232_)
);

FILL FILL_4__9165_ (
);

FILL SFILL18840x49050 (
);

FILL FILL_2__13485_ (
);

FILL FILL_1__12898_ (
);

FILL FILL_1__12478_ (
);

FILL FILL_1__12058_ (
);

FILL FILL_4__13812_ (
);

FILL FILL_0__9485_ (
);

FILL FILL_3__7582_ (
);

OAI21X1 _11756_ (
    .A(_2850_),
    .B(_2145_),
    .C(_2153_),
    .Y(_2851_)
);

FILL FILL_3__7162_ (
);

OAI21X1 _11336_ (
    .A(_2317_),
    .B(_2318_),
    .C(_2454_),
    .Y(_2455_)
);

FILL FILL_4__16284_ (
);

FILL FILL_5__7088_ (
);

FILL FILL_3__15697_ (
);

FILL FILL_0__12832_ (
);

FILL FILL_0__12412_ (
);

FILL FILL_3__15277_ (
);

FILL SFILL79480x4050 (
);

FILL FILL_5__15604_ (
);

FILL SFILL53960x80050 (
);

NAND2X1 _9904_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1536_)
);

FILL FILL_1__8861_ (
);

FILL FILL_1__8441_ (
);

FILL SFILL79080x15050 (
);

FILL FILL_1__8021_ (
);

FILL FILL_2__15631_ (
);

FILL FILL_2__15211_ (
);

FILL FILL_3__8787_ (
);

FILL FILL_3__8367_ (
);

FILL FILL_1__14624_ (
);

FILL FILL_1__14204_ (
);

NAND2X1 _7091_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_108_)
);

FILL FILL_0__13617_ (
);

OAI22X1 _13902_ (
    .A(_4404_),
    .B(_3931__bF$buf1),
    .C(_3966__bF$buf1),
    .D(_4403_),
    .Y(_4405_)
);

FILL FILL_5__9654_ (
);

FILL FILL_3__11197_ (
);

FILL FILL_5__9234_ (
);

FILL FILL_6__12111_ (
);

FILL FILL_0__16089_ (
);

OAI21X1 _16374_ (
    .A(_6802_),
    .B(gnd),
    .C(_6803_),
    .Y(_6769_[17])
);

FILL FILL_5__11944_ (
);

FILL FILL_1__9646_ (
);

FILL FILL_5__11524_ (
);

FILL FILL_1__9226_ (
);

FILL FILL_5__11104_ (
);

FILL FILL_2__16416_ (
);

FILL FILL_4__10937_ (
);

FILL FILL_4__7231_ (
);

FILL FILL_2__11971_ (
);

FILL FILL_4__10517_ (
);

FILL FILL_2__11551_ (
);

FILL FILL_2__11131_ (
);

FILL FILL_1__15829_ (
);

FILL FILL_1__15409_ (
);

DFFSR _8296_ (
    .Q(\datapath_1.regfile_1.regOut[11] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_653_[18])
);

FILL FILL_1__10964_ (
);

FILL FILL_1__10544_ (
);

FILL FILL_1__10124_ (
);

FILL FILL_2__7989_ (
);

FILL FILL_0__7971_ (
);

FILL FILL_0__7551_ (
);

BUFX2 BUFX2_insert580 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf27)
);

FILL FILL_2__7569_ (
);

BUFX2 BUFX2_insert581 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf26)
);

FILL SFILL114520x52050 (
);

BUFX2 BUFX2_insert582 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf25)
);

BUFX2 BUFX2_insert583 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf24)
);

BUFX2 BUFX2_insert584 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf23)
);

FILL FILL_6__13316_ (
);

BUFX2 BUFX2_insert585 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf22)
);

FILL FILL_4__14770_ (
);

FILL FILL_4__14350_ (
);

BUFX2 BUFX2_insert586 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf21)
);

BUFX2 BUFX2_insert587 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf20)
);

BUFX2 BUFX2_insert588 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf19)
);

BUFX2 BUFX2_insert589 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf18)
);

NAND3X1 _12294_ (
    .A(_3257_),
    .B(_3258_),
    .C(_3259_),
    .Y(\datapath_1.alu_1.ALUInB [19])
);

FILL FILL_5__12729_ (
);

FILL FILL_2__8510_ (
);

FILL FILL_3__13763_ (
);

FILL FILL_5__12309_ (
);

FILL FILL_3__13343_ (
);

FILL FILL_4__8856_ (
);

FILL FILL_4__8016_ (
);

FILL FILL_2__12756_ (
);

FILL FILL_0__13790_ (
);

FILL FILL_2__12336_ (
);

FILL FILL_0__13370_ (
);

FILL FILL_1__11749_ (
);

FILL FILL_1__11329_ (
);

FILL SFILL93560x24050 (
);

FILL SFILL3640x78050 (
);

FILL FILL_3__6853_ (
);

FILL FILL_5__16142_ (
);

FILL FILL_0__8756_ (
);

FILL FILL_0__8336_ (
);

DFFSR _10607_ (
    .Q(\datapath_1.regfile_1.regOut[29] [25]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_1823_[25])
);

FILL SFILL69240x50 (
);

FILL FILL_4__15975_ (
);

FILL FILL_4__15555_ (
);

FILL FILL_4__15135_ (
);

INVX1 _13499_ (
    .A(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_4010_)
);

FILL FILL_4__10690_ (
);

INVX1 _13079_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3748_)
);

FILL FILL_4__10270_ (
);

FILL FILL_3__14968_ (
);

FILL FILL_3__14548_ (
);

FILL FILL_3__14128_ (
);

FILL FILL_1__15582_ (
);

FILL FILL_1__15162_ (
);

FILL FILL_5__7720_ (
);

FILL FILL_5__7300_ (
);

FILL SFILL59080x56050 (
);

FILL FILL_0__14995_ (
);

INVX1 _14860_ (
    .A(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_5343_)
);

FILL FILL_0__14575_ (
);

FILL FILL_0__14155_ (
);

INVX1 _14440_ (
    .A(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_4932_)
);

AOI22X1 _14020_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [11]),
    .C(\datapath_1.regfile_1.regOut[27] [11]),
    .D(_4129_),
    .Y(_4521_)
);

FILL FILL_1__7712_ (
);

FILL FILL_2__14902_ (
);

FILL FILL_3__7218_ (
);

FILL SFILL3640x33050 (
);

FILL FILL_5__12482_ (
);

FILL FILL_5__12062_ (
);

FILL SFILL104520x50050 (
);

FILL SFILL43880x40050 (
);

FILL FILL_4__11895_ (
);

FILL FILL_4__11475_ (
);

FILL FILL_4__11055_ (
);

FILL FILL_1__16367_ (
);

FILL FILL_3__10888_ (
);

FILL FILL_5__8505_ (
);

FILL FILL_3__10048_ (
);

FILL FILL_1__11082_ (
);

NOR2X1 _15645_ (
    .A(_6110_),
    .B(_6108_),
    .Y(_6111_)
);

AOI22X1 _15225_ (
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [4]),
    .C(\datapath_1.regfile_1.regOut[5] [4]),
    .D(_5700_),
    .Y(_5701_)
);

FILL SFILL59080x11050 (
);

FILL FILL_0__10495_ (
);

OAI21X1 _10780_ (
    .A(_1976_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1977_),
    .Y(_1953_[12])
);

OAI21X1 _10360_ (
    .A(_1821_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1822_),
    .Y(_1758_[0])
);

FILL FILL_1__8917_ (
);

FILL SFILL104440x57050 (
);

FILL FILL_4__6922_ (
);

FILL FILL_0__16301_ (
);

FILL FILL_2__10822_ (
);

FILL FILL_5__13687_ (
);

FILL FILL_5__13267_ (
);

FILL FILL_2__10402_ (
);

NAND2X1 _7987_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_563_)
);

NAND2X1 _7567_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_344_)
);

DFFSR _7147_ (
    .Q(\datapath_1.regfile_1.regOut[2] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_68_[21])
);

FILL FILL_4__9394_ (
);

FILL SFILL33880x83050 (
);

FILL SFILL49480x68050 (
);

FILL SFILL108760x65050 (
);

FILL FILL_2__13294_ (
);

FILL FILL_1__12287_ (
);

FILL FILL_4__13621_ (
);

FILL FILL_0__9294_ (
);

INVX8 _11985_ (
    .A(ALUOp_0_bF$buf2),
    .Y(_3034_)
);

FILL SFILL49080x54050 (
);

NOR2X1 _11565_ (
    .A(_2673_),
    .B(_2631_),
    .Y(_2674_)
);

NOR2X1 _11145_ (
    .A(_2246_),
    .B(_2244_),
    .Y(_2264_)
);

FILL FILL_6__15899_ (
);

FILL FILL_3__12614_ (
);

FILL SFILL28920x39050 (
);

FILL FILL_4__16093_ (
);

FILL FILL_4__7707_ (
);

FILL FILL_2__11607_ (
);

FILL FILL_0__12641_ (
);

FILL FILL_3__15086_ (
);

FILL FILL_0__12221_ (
);

FILL FILL_2__14499_ (
);

FILL FILL_2__14079_ (
);

FILL FILL_5__15833_ (
);

FILL FILL_5__15413_ (
);

FILL FILL_0__7607_ (
);

DFFSR _9713_ (
    .Q(\datapath_1.regfile_1.regOut[22] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_1368_[27])
);

FILL FILL_1__8250_ (
);

FILL FILL_4__14826_ (
);

FILL FILL_2__15860_ (
);

FILL FILL_4__14406_ (
);

FILL FILL_2__15440_ (
);

FILL FILL_2__15020_ (
);

FILL FILL_3__8596_ (
);

FILL SFILL49000x52050 (
);

FILL FILL_3__13819_ (
);

FILL FILL_1__14853_ (
);

FILL FILL_1__14433_ (
);

FILL FILL_1__14013_ (
);

FILL FILL_0__13846_ (
);

FILL FILL_0__13426_ (
);

OAI22X1 _13711_ (
    .A(_4217_),
    .B(_3960_),
    .C(_3983__bF$buf2),
    .D(_4216_),
    .Y(_4218_)
);

FILL FILL_0__13006_ (
);

FILL FILL_5__9883_ (
);

FILL FILL_5__9463_ (
);

FILL FILL_5__9043_ (
);

OAI22X1 _16183_ (
    .A(_5480__bF$buf0),
    .B(_5291_),
    .C(_6634_),
    .D(_5499__bF$buf2),
    .Y(_6635_)
);

FILL SFILL23880x81050 (
);

FILL FILL_3__6909_ (
);

FILL FILL_5__11753_ (
);

FILL FILL_1__9875_ (
);

FILL FILL_5__11333_ (
);

FILL FILL_1__9035_ (
);

FILL FILL_2__16225_ (
);

FILL FILL_4__7880_ (
);

FILL FILL_4__7460_ (
);

FILL FILL_4__7040_ (
);

FILL FILL_4__10746_ (
);

FILL FILL_2__11780_ (
);

FILL SFILL103720x46050 (
);

FILL FILL_2__11360_ (
);

FILL FILL_1__15638_ (
);

FILL FILL_1__15218_ (
);

FILL SFILL39080x52050 (
);

FILL FILL_1__10773_ (
);

NOR2X1 _14916_ (
    .A(_5397_),
    .B(_5394_),
    .Y(_5398_)
);

FILL FILL_2__7798_ (
);

FILL FILL_0__7360_ (
);

FILL FILL_2__7378_ (
);

FILL FILL_6__13125_ (
);

FILL FILL_5__12958_ (
);

FILL SFILL18760x4050 (
);

FILL FILL_3__13992_ (
);

FILL FILL_5__12118_ (
);

FILL FILL_3__13572_ (
);

BUFX2 _6838_ (
    .A(_1_[0]),
    .Y(memoryAddress[0])
);

FILL FILL_3__13152_ (
);

FILL FILL_4__8245_ (
);

FILL FILL_2__12985_ (
);

FILL FILL_2__12145_ (
);

FILL SFILL63960x32050 (
);

FILL SFILL39000x50050 (
);

FILL SFILL94360x23050 (
);

FILL FILL_1__11978_ (
);

FILL FILL_1__11558_ (
);

FILL FILL_1__11138_ (
);

FILL FILL_5__16371_ (
);

FILL FILL_0__8985_ (
);

NAND2X1 _10836_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_2015_)
);

FILL FILL_0__8145_ (
);

NAND2X1 _10416_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1796_)
);

FILL FILL_4__15784_ (
);

FILL FILL_4__15364_ (
);

FILL FILL_0__11912_ (
);

FILL FILL_2__9524_ (
);

FILL FILL_3__14777_ (
);

FILL FILL_2__9104_ (
);

FILL FILL_3__14357_ (
);

FILL FILL_1__15391_ (
);

FILL FILL_0__14384_ (
);

FILL SFILL53960x75050 (
);

FILL SFILL84360x66050 (
);

FILL FILL_1__7941_ (
);

FILL FILL_1__7101_ (
);

FILL FILL_2__14711_ (
);

FILL FILL_3__7867_ (
);

FILL FILL_3__7447_ (
);

FILL FILL_5__12291_ (
);

FILL SFILL88680x74050 (
);

FILL FILL_1__13704_ (
);

FILL FILL_4__16149_ (
);

FILL FILL_4__11284_ (
);

FILL SFILL8760x40050 (
);

FILL SFILL29400x62050 (
);

FILL SFILL84760x35050 (
);

FILL FILL_1__16176_ (
);

FILL FILL111720x14050 (
);

FILL FILL_3__10697_ (
);

FILL FILL_5__8734_ (
);

FILL FILL_3__10277_ (
);

FILL FILL_5__8314_ (
);

INVX1 _15874_ (
    .A(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_6334_)
);

FILL FILL_0__15589_ (
);

FILL FILL_0__15169_ (
);

NAND3X1 _15454_ (
    .A(_5917_),
    .B(_5924_),
    .C(_5912_),
    .Y(_5925_)
);

OAI21X1 _15034_ (
    .A(_5461_),
    .B(_5513_),
    .C(_5471__bF$buf5),
    .Y(_5514_)
);

FILL FILL_1__8726_ (
);

FILL SFILL53960x30050 (
);

FILL FILL_6__14083_ (
);

FILL FILL_2__15916_ (
);

FILL FILL_0__16110_ (
);

FILL FILL_5__13496_ (
);

FILL FILL_2__10631_ (
);

DFFSR _7796_ (
    .Q(\datapath_1.regfile_1.regOut[7] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_393_[30])
);

FILL FILL_1__14909_ (
);

INVX1 _7376_ (
    .A(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_257_)
);

FILL FILL_4__12489_ (
);

FILL FILL_4__12069_ (
);

FILL FILL_5__9939_ (
);

FILL FILL_5__9519_ (
);

FILL SFILL53880x37050 (
);

FILL FILL_1__12096_ (
);

FILL FILL_4__13850_ (
);

INVX1 _16239_ (
    .A(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_6690_)
);

FILL FILL_4__13430_ (
);

FILL SFILL3720x66050 (
);

FILL FILL_4__13010_ (
);

INVX1 _11794_ (
    .A(_2144_),
    .Y(_2887_)
);

AND2X2 _11374_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2491_)
);

FILL FILL_0__11089_ (
);

FILL FILL_5__11809_ (
);

FILL SFILL104600x83050 (
);

FILL FILL_3__12843_ (
);

FILL SFILL43960x73050 (
);

FILL FILL_3__12423_ (
);

FILL FILL_3__12003_ (
);

FILL FILL_4__7936_ (
);

FILL FILL_2__11836_ (
);

FILL FILL_0__12870_ (
);

FILL FILL_2__11416_ (
);

FILL FILL_0__12450_ (
);

FILL FILL_0__12030_ (
);

FILL FILL_1__10829_ (
);

FILL FILL_1__10409_ (
);

FILL FILL_5__15642_ (
);

FILL FILL_5__15222_ (
);

FILL FILL_0__7836_ (
);

FILL FILL_0__7416_ (
);

DFFSR _9942_ (
    .Q(\datapath_1.regfile_1.regOut[24] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_1498_[0])
);

INVX1 _9522_ (
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_1342_)
);

INVX1 _9102_ (
    .A(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_1123_)
);

FILL FILL_4__14635_ (
);

FILL FILL_4__14215_ (
);

INVX1 _12999_ (
    .A(_2_[16]),
    .Y(_3651_)
);

INVX1 _12579_ (
    .A(\datapath_1.Data [4]),
    .Y(_3432_)
);

OAI21X1 _12159_ (
    .A(_3158_),
    .B(ALUSrcA_bF$buf4),
    .C(_3159_),
    .Y(\datapath_1.alu_1.ALUInA [14])
);

FILL SFILL3720x21050 (
);

FILL FILL_3__13628_ (
);

FILL FILL_3__13208_ (
);

FILL FILL_1__14662_ (
);

FILL FILL_1__14242_ (
);

FILL FILL_0__13655_ (
);

OAI22X1 _13940_ (
    .A(_4440_),
    .B(_3931__bF$buf1),
    .C(_3977__bF$buf0),
    .D(_4441_),
    .Y(_4442_)
);

FILL FILL_0__13235_ (
);

FILL FILL_0_BUFX2_insert225 (
);

INVX1 _13520_ (
    .A(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_4031_)
);

FILL FILL_0_BUFX2_insert226 (
);

INVX1 _13100_ (
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_3698_)
);

FILL FILL_0_BUFX2_insert227 (
);

FILL FILL_0_BUFX2_insert228 (
);

FILL FILL_0_BUFX2_insert229 (
);

FILL FILL_5__9272_ (
);

FILL FILL_5__16007_ (
);

FILL FILL_5__11982_ (
);

FILL FILL_1__9684_ (
);

FILL FILL_5__11562_ (
);

FILL FILL_1__9264_ (
);

FILL FILL_5__11142_ (
);

FILL SFILL43880x35050 (
);

FILL FILL_2__16034_ (
);

FILL FILL_4__10975_ (
);

FILL FILL_4__10555_ (
);

FILL FILL_4__10135_ (
);

FILL FILL_1__15867_ (
);

FILL FILL_1__15447_ (
);

FILL FILL_1__15027_ (
);

FILL SFILL59000x49050 (
);

FILL FILL_1__10162_ (
);

OAI22X1 _14725_ (
    .A(_3902__bF$buf3),
    .B(_5210_),
    .C(_5209_),
    .D(_3955__bF$buf0),
    .Y(_5211_)
);

NOR2X1 _14305_ (
    .A(_4796_),
    .B(_4799_),
    .Y(_4800_)
);

BUFX2 BUFX2_insert960 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf5 )
);

BUFX2 BUFX2_insert961 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf4 )
);

FILL FILL_2__7187_ (
);

BUFX2 BUFX2_insert962 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf3 )
);

BUFX2 BUFX2_insert963 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf2 )
);

BUFX2 BUFX2_insert964 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf1 )
);

BUFX2 BUFX2_insert965 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf0 )
);

BUFX2 BUFX2_insert966 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf4 )
);

BUFX2 BUFX2_insert967 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf3 )
);

BUFX2 BUFX2_insert968 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf2 )
);

FILL FILL_0__15801_ (
);

BUFX2 BUFX2_insert969 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf1 )
);

FILL FILL_5__12767_ (
);

FILL FILL_5__12347_ (
);

FILL FILL_3__13381_ (
);

FILL FILL_4__8894_ (
);

FILL SFILL33880x78050 (
);

FILL FILL_4__8474_ (
);

FILL FILL_4__8054_ (
);

FILL FILL_2__12374_ (
);

FILL FILL_1__11787_ (
);

FILL FILL_1__11367_ (
);

FILL FILL_4__12701_ (
);

FILL FILL_3__6891_ (
);

FILL FILL_5__16180_ (
);

FILL FILL_0__8374_ (
);

NAND2X1 _10645_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1908_)
);

DFFSR _10225_ (
    .Q(\datapath_1.regfile_1.regOut[26] [27]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1628_[27])
);

FILL FILL_6__14979_ (
);

FILL FILL_6__14559_ (
);

FILL FILL_4__15593_ (
);

FILL FILL_4__15173_ (
);

FILL FILL_2__9753_ (
);

FILL FILL_3__14586_ (
);

FILL FILL_0__11721_ (
);

FILL FILL_3__14166_ (
);

FILL FILL_0__11301_ (
);

FILL FILL_6__15920_ (
);

FILL SFILL33080x50050 (
);

FILL FILL_4__9679_ (
);

FILL FILL_6__15500_ (
);

FILL FILL_4__9259_ (
);

FILL FILL_2__13999_ (
);

FILL FILL_2__13579_ (
);

FILL FILL_2__13159_ (
);

FILL FILL_0__14193_ (
);

FILL SFILL33880x33050 (
);

FILL FILL_5__14913_ (
);

FILL FILL_1__7750_ (
);

FILL FILL_1__7330_ (
);

FILL FILL_4__13906_ (
);

FILL FILL_2__14940_ (
);

FILL FILL_2__14520_ (
);

FILL FILL_0__9999_ (
);

FILL SFILL49000x47050 (
);

FILL FILL_2__14100_ (
);

FILL FILL_3__7676_ (
);

FILL FILL_0__9159_ (
);

FILL FILL_1__13933_ (
);

FILL FILL_4__16378_ (
);

FILL FILL_1__13513_ (
);

FILL SFILL94440x56050 (
);

FILL FILL_4__11093_ (
);

FILL FILL_0__12506_ (
);

FILL FILL_5__8963_ (
);

FILL FILL_5__8123_ (
);

FILL FILL_6__11840_ (
);

OAI22X1 _15683_ (
    .A(_6147_),
    .B(_5548__bF$buf0),
    .C(_5489__bF$buf1),
    .D(_4707_),
    .Y(_6148_)
);

FILL FILL_0__15398_ (
);

FILL FILL_6__11420_ (
);

OAI22X1 _15263_ (
    .A(_4239_),
    .B(_5539__bF$buf2),
    .C(_5530__bF$buf0),
    .D(_4198_),
    .Y(_5738_)
);

FILL SFILL23880x76050 (
);

FILL FILL_3__16312_ (
);

FILL FILL_5__10833_ (
);

FILL FILL_1__8955_ (
);

FILL FILL_5__10413_ (
);

FILL FILL_1__8115_ (
);

FILL FILL_2__15725_ (
);

FILL FILL_2__15305_ (
);

FILL FILL_4__6960_ (
);

FILL FILL_2__10440_ (
);

FILL FILL_2__10020_ (
);

FILL FILL_1__14718_ (
);

FILL SFILL23480x62050 (
);

INVX1 _7185_ (
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_150_)
);

FILL FILL_4__12298_ (
);

FILL FILL_3__9402_ (
);

FILL FILL_0__6860_ (
);

FILL FILL_2__6878_ (
);

FILL SFILL94440x11050 (
);

FILL FILL_5__9748_ (
);

FILL SFILL23800x74050 (
);

NOR2X1 _16048_ (
    .A(_5157_),
    .B(_5534__bF$buf1),
    .Y(_6503_)
);

OAI21X1 _11183_ (
    .A(_2300_),
    .B(_2301_),
    .C(_2297_),
    .Y(_2302_)
);

FILL FILL_5__11618_ (
);

FILL FILL_3__12652_ (
);

FILL FILL_3__12232_ (
);

FILL FILL_4__7745_ (
);

FILL FILL_4__7325_ (
);

FILL FILL_2__11645_ (
);

FILL FILL_2__11225_ (
);

FILL SFILL94360x18050 (
);

FILL FILL_1__10638_ (
);

FILL FILL_5__15871_ (
);

FILL FILL_5__15451_ (
);

FILL FILL_5__15031_ (
);

INVX1 _9751_ (
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_1454_)
);

FILL FILL_0__7225_ (
);

DFFSR _9331_ (
    .Q(\datapath_1.regfile_1.regOut[19] [29]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1173_[29])
);

FILL FILL_4__14864_ (
);

FILL FILL_4__14444_ (
);

FILL FILL_4__14024_ (
);

INVX1 _12388_ (
    .A(ALUOut[15]),
    .Y(_3324_)
);

FILL FILL_3__13857_ (
);

FILL FILL_2__8604_ (
);

FILL FILL_3__13437_ (
);

FILL FILL_1__14891_ (
);

FILL FILL_1__14471_ (
);

FILL FILL_3__13017_ (
);

FILL FILL_1__14051_ (
);

FILL FILL_0__13884_ (
);

FILL FILL_0__13464_ (
);

FILL FILL_0__13044_ (
);

FILL FILL_5__9081_ (
);

FILL FILL_5__16236_ (
);

FILL FILL_3__6947_ (
);

FILL FILL_5__11791_ (
);

FILL FILL_5__11371_ (
);

FILL FILL_1__9493_ (
);

FILL FILL_4__15649_ (
);

FILL FILL_4__15229_ (
);

FILL FILL_2__16263_ (
);

FILL FILL_4__10784_ (
);

FILL FILL_4__10364_ (
);

FILL SFILL8760x35050 (
);

FILL FILL_4_BUFX2_insert50 (
);

FILL FILL_2__9809_ (
);

FILL SFILL13800x72050 (
);

FILL FILL_4_BUFX2_insert51 (
);

FILL FILL_1__15676_ (
);

FILL FILL_4_BUFX2_insert52 (
);

FILL FILL_1__15256_ (
);

FILL FILL_4_BUFX2_insert53 (
);

FILL FILL_4_BUFX2_insert54 (
);

FILL FILL_4_BUFX2_insert55 (
);

FILL FILL_5__7814_ (
);

FILL SFILL74040x83050 (
);

FILL FILL_4_BUFX2_insert56 (
);

FILL FILL_4_BUFX2_insert57 (
);

FILL FILL_1__10391_ (
);

FILL FILL_4_BUFX2_insert58 (
);

FILL FILL_4_BUFX2_insert59 (
);

NOR2X1 _14954_ (
    .A(_5434_),
    .B(_3983__bF$buf3),
    .Y(_5435_)
);

FILL FILL_0__14669_ (
);

FILL FILL_0__14249_ (
);

INVX1 _14534_ (
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_5024_)
);

INVX1 _14114_ (
    .A(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_4613_)
);

FILL SFILL114600x35050 (
);

FILL SFILL53960x25050 (
);

FILL FILL_1__7806_ (
);

FILL SFILL84360x16050 (
);

FILL FILL_0__15610_ (
);

FILL FILL_5__12996_ (
);

FILL FILL_5__12576_ (
);

FILL FILL_5__12156_ (
);

BUFX2 _6876_ (
    .A(_2_[6]),
    .Y(memoryWriteData[6])
);

FILL SFILL74440x52050 (
);

FILL FILL_4__11989_ (
);

FILL FILL_4__11569_ (
);

FILL FILL_4__11149_ (
);

FILL FILL_2__12183_ (
);

FILL FILL_1__11596_ (
);

FILL FILL_1__11176_ (
);

AOI22X1 _15739_ (
    .A(_5567_),
    .B(\datapath_1.regfile_1.regOut[28] [17]),
    .C(\datapath_1.regfile_1.regOut[31] [17]),
    .D(_5571_),
    .Y(_6202_)
);

FILL FILL_4__12510_ (
);

INVX1 _15319_ (
    .A(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_5793_)
);

FILL FILL_0__8183_ (
);

NOR2X1 _10874_ (
    .A(_2019_),
    .B(_2021_),
    .Y(_2022_)
);

DFFSR _10454_ (
    .Q(\datapath_1.regfile_1.regOut[28] [0]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1758_[0])
);

FILL FILL_0__10169_ (
);

INVX1 _10034_ (
    .A(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_1602_)
);

FILL SFILL43960x68050 (
);

FILL FILL_3__11923_ (
);

FILL FILL_3__11503_ (
);

FILL FILL_2__10916_ (
);

FILL FILL_2__9982_ (
);

FILL FILL_0__11950_ (
);

FILL FILL_2__9142_ (
);

FILL FILL_3__14395_ (
);

FILL FILL_0__11530_ (
);

FILL FILL_0__11110_ (
);

FILL FILL_4__9488_ (
);

FILL FILL112360x72050 (
);

FILL FILL_2__13388_ (
);

FILL FILL_5__14722_ (
);

FILL FILL_0__6916_ (
);

FILL FILL_5__14302_ (
);

INVX1 _8602_ (
    .A(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_871_)
);

FILL FILL_4__13715_ (
);

FILL SFILL64040x81050 (
);

FILL FILL_3__7485_ (
);

FILL FILL_0__9388_ (
);

FILL FILL_3__7065_ (
);

OAI21X1 _11659_ (
    .A(_2759_),
    .B(_2178_),
    .C(_2161_),
    .Y(_2762_)
);

NAND2X1 _11239_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2358_)
);

FILL SFILL3720x16050 (
);

FILL FILL_3__12708_ (
);

FILL FILL_1__13742_ (
);

FILL FILL_1__13322_ (
);

FILL FILL_4__16187_ (
);

FILL SFILL43960x23050 (
);

FILL FILL_0__12735_ (
);

INVX1 _12600_ (
    .A(\datapath_1.Data [11]),
    .Y(_3446_)
);

FILL FILL_0__12315_ (
);

FILL FILL_5__8772_ (
);

FILL FILL_5__8352_ (
);

INVX1 _15492_ (
    .A(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_5962_)
);

FILL FILL_5__15927_ (
);

NAND3X1 _15072_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5471__bF$buf5),
    .C(_5476_),
    .Y(_5552_)
);

FILL FILL_5__15507_ (
);

OAI21X1 _9807_ (
    .A(_1490_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .C(_1491_),
    .Y(_1433_[29])
);

FILL FILL_3__16121_ (
);

FILL FILL_1__8764_ (
);

FILL FILL_5__10642_ (
);

FILL FILL_1__8344_ (
);

FILL FILL_2__15954_ (
);

FILL FILL_2__15534_ (
);

FILL FILL_2__15114_ (
);

FILL FILL_1__14947_ (
);

FILL FILL_1__14527_ (
);

FILL FILL_1__14107_ (
);

FILL FILL_3__9631_ (
);

NAND2X1 _13805_ (
    .A(_4309_),
    .B(_4301_),
    .Y(_4310_)
);

FILL FILL_3__9211_ (
);

FILL FILL112280x34050 (
);

FILL FILL_5__9977_ (
);

FILL FILL_5__9557_ (
);

FILL FILL_5__9137_ (
);

FILL FILL_6__12014_ (
);

INVX1 _16277_ (
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_6727_)
);

FILL FILL_5__11847_ (
);

FILL FILL_1__9549_ (
);

FILL FILL_3__12881_ (
);

FILL FILL_5__11427_ (
);

FILL FILL_3__12461_ (
);

FILL FILL_5__11007_ (
);

FILL FILL_1__9129_ (
);

FILL FILL_3__12041_ (
);

FILL FILL_4__7974_ (
);

FILL FILL_2__16319_ (
);

FILL FILL_4__7554_ (
);

FILL FILL_2__11874_ (
);

FILL FILL_2__11454_ (
);

FILL FILL_2__11034_ (
);

OAI21X1 _8199_ (
    .A(_662_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_663_),
    .Y(_653_[5])
);

FILL FILL_1__10447_ (
);

FILL FILL_1__10027_ (
);

FILL FILL_5__15680_ (
);

FILL FILL_5__15260_ (
);

FILL FILL_0__7874_ (
);

INVX1 _9980_ (
    .A(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_1566_)
);

FILL FILL_0__7454_ (
);

FILL FILL_0__7034_ (
);

DFFSR _9560_ (
    .Q(\datapath_1.regfile_1.regOut[21] [2]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1303_[2])
);

OAI21X1 _9140_ (
    .A(_1147_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1148_),
    .Y(_1108_[20])
);

FILL FILL_6__13219_ (
);

FILL FILL_4__14673_ (
);

FILL FILL_4__14253_ (
);

NAND2X1 _12197_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [27]),
    .Y(_3185_)
);

FILL FILL_2__8833_ (
);

FILL FILL_3__13666_ (
);

FILL FILL_0__10801_ (
);

FILL FILL_3__13246_ (
);

FILL FILL_1__14280_ (
);

FILL FILL_4__8759_ (
);

FILL FILL_0_BUFX2_insert600 (
);

FILL FILL_0_BUFX2_insert601 (
);

FILL FILL_4__8339_ (
);

FILL FILL_0_BUFX2_insert602 (
);

FILL FILL_0_BUFX2_insert603 (
);

FILL FILL_2__12659_ (
);

FILL FILL_0_BUFX2_insert604 (
);

FILL FILL_2__12239_ (
);

FILL FILL_0__13693_ (
);

FILL FILL_0_BUFX2_insert605 (
);

FILL FILL_0__13273_ (
);

FILL FILL_0_BUFX2_insert606 (
);

FILL FILL_0_BUFX2_insert607 (
);

FILL FILL_0_BUFX2_insert608 (
);

FILL FILL_0_BUFX2_insert609 (
);

FILL FILL_2__13600_ (
);

FILL FILL_5__16045_ (
);

FILL FILL_0__8659_ (
);

FILL FILL_0__8239_ (
);

FILL SFILL98840x52050 (
);

FILL FILL_5__11180_ (
);

FILL FILL_4__15878_ (
);

FILL FILL_4__15458_ (
);

FILL FILL_4__15038_ (
);

FILL FILL_2__16072_ (
);

FILL FILL_4__10173_ (
);

FILL FILL_0__9600_ (
);

FILL FILL_2__9618_ (
);

FILL FILL_1__15485_ (
);

FILL FILL_1__15065_ (
);

FILL FILL_5__7623_ (
);

FILL FILL_5__7203_ (
);

FILL FILL_6__10920_ (
);

FILL FILL_0__14898_ (
);

FILL FILL_0__14478_ (
);

AOI22X1 _14763_ (
    .A(_3882__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [27]),
    .C(\datapath_1.regfile_1.regOut[1] [27]),
    .D(_3997__bF$buf2),
    .Y(_5248_)
);

FILL FILL_0__14058_ (
);

AOI21X1 _14343_ (
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .B(_4115_),
    .C(_4836_),
    .Y(_4837_)
);

FILL FILL_3__15812_ (
);

FILL FILL_1__7615_ (
);

FILL FILL_2__14805_ (
);

FILL FILL_5__12385_ (
);

FILL FILL_4__8092_ (
);

FILL FILL_4__11798_ (
);

FILL FILL_4__11378_ (
);

FILL FILL_3__8902_ (
);

FILL FILL_5__8828_ (
);

AOI21X1 _15968_ (
    .A(_6401_),
    .B(_6425_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [22])
);

FILL SFILL23800x69050 (
);

NAND3X1 _15548_ (
    .A(_6014_),
    .B(_6015_),
    .C(_6013_),
    .Y(_6016_)
);

INVX4 _15128_ (
    .A(_5469__bF$buf2),
    .Y(_5606_)
);

INVX1 _10683_ (
    .A(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_1933_)
);

FILL FILL_0__10398_ (
);

INVX1 _10263_ (
    .A(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_1714_)
);

FILL FILL_3__11732_ (
);

FILL FILL_3__11312_ (
);

FILL FILL_0__16204_ (
);

FILL FILL_2__9791_ (
);

FILL FILL_2__9371_ (
);

FILL FILL_2__10305_ (
);

FILL FILL112440x3050 (
);

FILL FILL_4__9297_ (
);

FILL FILL_5__14951_ (
);

FILL FILL_5__14531_ (
);

FILL FILL_5__14111_ (
);

INVX1 _8831_ (
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_983_)
);

DFFSR _8411_ (
    .Q(\datapath_1.regfile_1.regOut[12] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_718_[5])
);

FILL FILL_4__13944_ (
);

FILL FILL_4__13524_ (
);

FILL FILL_4__13104_ (
);

NAND2X1 _11888_ (
    .A(ALUOut[0]),
    .B(IorD_bF$buf2),
    .Y(_3031_)
);

FILL FILL_3__7294_ (
);

OAI22X1 _11468_ (
    .A(_2290_),
    .B(_2346_),
    .C(_2480_),
    .D(_2582_),
    .Y(_2583_)
);

FILL SFILL23800x24050 (
);

NAND2X1 _11048_ (
    .A(_2163_),
    .B(_2166_),
    .Y(_2167_)
);

FILL FILL_3__12517_ (
);

FILL FILL_1__13971_ (
);

FILL FILL_1__13551_ (
);

FILL FILL_1__13131_ (
);

FILL FILL_0__12964_ (
);

FILL FILL_0__12124_ (
);

FILL FILL_5__8581_ (
);

FILL SFILL74200x5050 (
);

FILL FILL_5__15736_ (
);

FILL FILL_5__15316_ (
);

FILL FILL_3__16350_ (
);

OAI21X1 _9616_ (
    .A(_1383_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .C(_1384_),
    .Y(_1368_[8])
);

FILL FILL_1__8993_ (
);

FILL FILL_5__10871_ (
);

FILL FILL_5__10451_ (
);

FILL FILL_1__8573_ (
);

FILL FILL_5__10031_ (
);

FILL FILL_4__14729_ (
);

FILL FILL_2__15763_ (
);

FILL FILL_4__14309_ (
);

FILL FILL_2__15343_ (
);

FILL FILL_3__8499_ (
);

FILL FILL_3__8079_ (
);

FILL SFILL13800x67050 (
);

FILL FILL_1__14756_ (
);

FILL FILL_1__14336_ (
);

FILL SFILL13880x24050 (
);

FILL FILL_3__9860_ (
);

FILL FILL_0__13749_ (
);

FILL FILL_3__9020_ (
);

FILL FILL_0__13329_ (
);

OAI22X1 _13614_ (
    .A(_4122_),
    .B(_3910_),
    .C(_3982__bF$buf3),
    .D(_4121_),
    .Y(_4123_)
);

FILL FILL_5__9786_ (
);

FILL FILL_5__9366_ (
);

FILL SFILL29000x38050 (
);

NOR2X1 _16086_ (
    .A(_6530_),
    .B(_6540_),
    .Y(_6541_)
);

FILL FILL_1__9778_ (
);

FILL FILL_5__11656_ (
);

FILL FILL_1__9358_ (
);

FILL FILL_5__11236_ (
);

FILL FILL_3__12270_ (
);

FILL FILL_2__16128_ (
);

FILL FILL_4__7363_ (
);

FILL FILL_4__10649_ (
);

FILL FILL_2__11683_ (
);

FILL FILL_2__11263_ (
);

FILL SFILL13800x22050 (
);

FILL FILL_1__10676_ (
);

FILL FILL_1__10256_ (
);

NOR2X1 _14819_ (
    .A(_5299_),
    .B(_5302_),
    .Y(_5303_)
);

FILL FILL_0__7683_ (
);

FILL FILL_6__8650_ (
);

FILL FILL_6__13868_ (
);

FILL FILL_4__14482_ (
);

FILL FILL_4__14062_ (
);

FILL FILL_3__13895_ (
);

FILL FILL_2__8642_ (
);

FILL FILL_3__13475_ (
);

FILL FILL_2__8222_ (
);

FILL FILL_4__8988_ (
);

FILL FILL_4__8568_ (
);

FILL FILL_4__8148_ (
);

FILL FILL112360x67050 (
);

FILL FILL_2__12888_ (
);

FILL FILL_2__12468_ (
);

FILL FILL_2__12048_ (
);

FILL FILL_0__13082_ (
);

FILL FILL_5__13802_ (
);

FILL SFILL64040x76050 (
);

FILL FILL_0__8888_ (
);

FILL FILL_5__16274_ (
);

FILL FILL_3__6985_ (
);

FILL FILL_6__9855_ (
);

FILL FILL_0__8468_ (
);

DFFSR _10739_ (
    .Q(\datapath_1.regfile_1.regOut[30] [29]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_1888_[29])
);

OAI21X1 _10319_ (
    .A(_1750_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1751_),
    .Y(_1693_[29])
);

FILL FILL_4__15687_ (
);

FILL FILL_1__12402_ (
);

FILL FILL_4__15267_ (
);

FILL SFILL43960x18050 (
);

FILL FILL_2__9847_ (
);

FILL FILL_2__9427_ (
);

FILL FILL_0__11815_ (
);

FILL FILL_2__9007_ (
);

FILL FILL_1__15294_ (
);

FILL FILL_5__7852_ (
);

FILL FILL_5__7432_ (
);

NAND3X1 _14992_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5461_),
    .C(_5471__bF$buf5),
    .Y(_5472_)
);

AOI22X1 _14572_ (
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .B(_3942__bF$buf2),
    .C(_3995__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_5061_)
);

FILL FILL_0__14287_ (
);

OAI22X1 _14152_ (
    .A(_4648_),
    .B(_3890_),
    .C(_3960_),
    .D(_4649_),
    .Y(_4650_)
);

FILL FILL112360x22050 (
);

FILL FILL_3__15621_ (
);

FILL FILL_3__15201_ (
);

FILL FILL_1__7844_ (
);

FILL FILL_1__7424_ (
);

FILL FILL_2__14614_ (
);

FILL SFILL64040x31050 (
);

FILL FILL_5__12194_ (
);

FILL FILL_1__13607_ (
);

FILL FILL_4__11187_ (
);

FILL FILL_3__8711_ (
);

FILL SFILL89240x80050 (
);

FILL FILL112280x29050 (
);

FILL FILL_1__16079_ (
);

FILL FILL_5__8637_ (
);

FILL FILL_5__8217_ (
);

NAND3X1 _15777_ (
    .A(_6233_),
    .B(_6234_),
    .C(_6238_),
    .Y(_6239_)
);

AOI22X1 _15357_ (
    .A(\datapath_1.regfile_1.regOut[31] [7]),
    .B(_5571_),
    .C(_5481_),
    .D(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_5830_)
);

FILL FILL_3__16406_ (
);

INVX1 _10492_ (
    .A(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_1826_)
);

FILL FILL_5__10927_ (
);

DFFSR _10072_ (
    .Q(\datapath_1.regfile_1.regOut[25] [2]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_1563_[2])
);

FILL FILL_5__10507_ (
);

FILL FILL_1__8629_ (
);

FILL FILL_3__11961_ (
);

FILL FILL_3__11541_ (
);

FILL FILL_1__8209_ (
);

FILL FILL_3__11121_ (
);

FILL FILL_2__15819_ (
);

FILL FILL_0__16013_ (
);

FILL FILL_2__10954_ (
);

FILL FILL_2__10534_ (
);

FILL FILL_5__13399_ (
);

FILL FILL_2__10114_ (
);

OAI21X1 _7699_ (
    .A(_410_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_411_),
    .Y(_393_[9])
);

DFFSR _7279_ (
    .Q(\datapath_1.regfile_1.regOut[3] [25]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_133_[25])
);

FILL FILL_3__9916_ (
);

FILL FILL_5__14760_ (
);

FILL FILL_5__14340_ (
);

FILL FILL_0__6954_ (
);

OAI21X1 _8640_ (
    .A(_895_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_896_),
    .Y(_848_[24])
);

OAI21X1 _8220_ (
    .A(_676_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_677_),
    .Y(_653_[12])
);

FILL FILL_4__13753_ (
);

FILL FILL_4__13333_ (
);

OAI21X1 _11697_ (
    .A(_2165_),
    .B(_2757_),
    .C(_2796_),
    .Y(_2797_)
);

INVX1 _11277_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .Y(_2396_)
);

FILL FILL_3__12746_ (
);

FILL FILL_1__13780_ (
);

FILL FILL_3__12326_ (
);

FILL FILL_1__13360_ (
);

FILL FILL_4__7839_ (
);

FILL FILL_4__7419_ (
);

FILL FILL_2__11739_ (
);

FILL FILL_0__12773_ (
);

FILL FILL_2__11319_ (
);

FILL FILL_0__12353_ (
);

FILL FILL_5__8390_ (
);

FILL FILL_5__15965_ (
);

FILL FILL_5__15545_ (
);

FILL FILL_0__7739_ (
);

FILL FILL_5__15125_ (
);

FILL FILL_0__7319_ (
);

DFFSR _9845_ (
    .Q(\datapath_1.regfile_1.regOut[23] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_1433_[31])
);

NAND2X1 _9425_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1298_)
);

FILL FILL_5__10680_ (
);

NAND2X1 _9005_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1079_)
);

FILL FILL_1__8382_ (
);

FILL FILL_5__10260_ (
);

FILL FILL_4__14958_ (
);

FILL FILL_2__15992_ (
);

FILL FILL_4__14538_ (
);

FILL FILL_2__15572_ (
);

FILL FILL_4__14118_ (
);

FILL FILL_2__15152_ (
);

FILL FILL_1__14985_ (
);

FILL FILL_1__14565_ (
);

FILL FILL_1__14145_ (
);

FILL FILL_0__13978_ (
);

OAI22X1 _13843_ (
    .A(_4346_),
    .B(_3941_),
    .C(_3890_),
    .D(_4345_),
    .Y(_4347_)
);

FILL FILL_0__13558_ (
);

NAND3X1 _13423_ (
    .A(_3898_),
    .B(_3883_),
    .C(_3919_),
    .Y(_3935_)
);

FILL FILL_0__13138_ (
);

NAND2X1 _13003_ (
    .A(vdd),
    .B(\datapath_1.rd2 [17]),
    .Y(_3654_)
);

FILL FILL_5__9595_ (
);

FILL SFILL44040x72050 (
);

FILL FILL_6__12892_ (
);

FILL SFILL58280x44050 (
);

FILL FILL_5__11885_ (
);

FILL SFILL84120x68050 (
);

FILL FILL_5__11465_ (
);

FILL FILL_1__9167_ (
);

FILL FILL_5__11045_ (
);

FILL FILL_2__16357_ (
);

FILL FILL_4__7592_ (
);

FILL FILL_4__7172_ (
);

FILL FILL_4__10878_ (
);

FILL FILL_4__10038_ (
);

FILL FILL_2__11492_ (
);

FILL FILL_2__11072_ (
);

FILL FILL_1__10065_ (
);

NOR2X1 _14628_ (
    .A(_5115_),
    .B(_3955__bF$buf3),
    .Y(_5116_)
);

OAI22X1 _14208_ (
    .A(_4703_),
    .B(_3982__bF$buf0),
    .C(_3978_),
    .D(_4704_),
    .Y(_4705_)
);

FILL FILL_0__7492_ (
);

FILL FILL_0__7072_ (
);

FILL FILL_3__10812_ (
);

FILL FILL_4__14291_ (
);

FILL FILL_0__15704_ (
);

FILL FILL_2__8871_ (
);

FILL FILL_2__8451_ (
);

FILL FILL_3__13284_ (
);

FILL FILL_4__8377_ (
);

FILL FILL_2__12697_ (
);

FILL FILL_2__12277_ (
);

FILL FILL_5__13611_ (
);

DFFSR _7911_ (
    .Q(\datapath_1.regfile_1.regOut[8] [17]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_458_[17])
);

FILL SFILL105080x4050 (
);

FILL FILL_4__12604_ (
);

FILL FILL_5__16083_ (
);

FILL FILL_0__8697_ (
);

NAND2X1 _10968_ (
    .A(\control_1.op [1]),
    .B(_2042_),
    .Y(_2043_)
);

FILL FILL_0__8277_ (
);

OAI21X1 _10548_ (
    .A(_1862_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1863_),
    .Y(_1823_[20])
);

OAI21X1 _10128_ (
    .A(_1643_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1644_),
    .Y(_1628_[8])
);

FILL FILL_1__12631_ (
);

FILL FILL_4__15496_ (
);

FILL FILL_4__15076_ (
);

FILL FILL_1__12211_ (
);

FILL SFILL69160x83050 (
);

FILL FILL_2__9656_ (
);

FILL FILL_3__14489_ (
);

FILL FILL_2__9236_ (
);

FILL FILL_0__11624_ (
);

FILL FILL_3__14069_ (
);

FILL FILL_0__11204_ (
);

FILL FILL_6__15823_ (
);

FILL FILL_6__15403_ (
);

FILL SFILL74120x66050 (
);

FILL FILL_5__7241_ (
);

INVX1 _14381_ (
    .A(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_4874_)
);

FILL FILL_0__14096_ (
);

FILL FILL_5__14816_ (
);

FILL FILL_3__15850_ (
);

FILL FILL_3__15430_ (
);

FILL FILL_3__15010_ (
);

FILL FILL_1__7233_ (
);

FILL FILL_4__13809_ (
);

FILL FILL_2__14843_ (
);

FILL FILL_3__7999_ (
);

FILL FILL_2__14423_ (
);

FILL FILL_2__14003_ (
);

FILL FILL_3__7579_ (
);

FILL FILL_3__7159_ (
);

FILL FILL_1__13836_ (
);

FILL FILL_1__13416_ (
);

FILL FILL_3__8520_ (
);

FILL FILL_0__12829_ (
);

FILL FILL_3__8100_ (
);

FILL FILL_0__12409_ (
);

FILL FILL_5__8866_ (
);

FILL FILL_5__8446_ (
);

FILL FILL_6__11743_ (
);

NOR2X1 _15586_ (
    .A(_6052_),
    .B(_6047_),
    .Y(_6053_)
);

FILL FILL_6__11323_ (
);

NOR3X1 _15166_ (
    .A(_5634_),
    .B(_5623_),
    .C(_5643_),
    .Y(_5644_)
);

FILL SFILL74120x21050 (
);

FILL FILL_3__16215_ (
);

FILL FILL_1__8858_ (
);

FILL FILL_5__10316_ (
);

FILL FILL_1__8438_ (
);

FILL FILL_3__11770_ (
);

FILL FILL_3__11350_ (
);

FILL FILL_1__8018_ (
);

FILL FILL_2__15628_ (
);

FILL FILL_2__15208_ (
);

FILL FILL_4__6863_ (
);

FILL SFILL99320x70050 (
);

FILL FILL_0__16242_ (
);

FILL FILL_2__10763_ (
);

NAND2X1 _7088_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_106_)
);

FILL SFILL13800x17050 (
);

FILL FILL_3__9725_ (
);

FILL SFILL59160x81050 (
);

FILL FILL_6__7730_ (
);

FILL FILL_4__13982_ (
);

FILL FILL_4__13562_ (
);

FILL FILL_4__13142_ (
);

FILL SFILL64120x64050 (
);

OAI21X1 _11086_ (
    .A(_2200_),
    .B(_2193_),
    .C(_2204_),
    .Y(_2205_)
);

FILL FILL_3__12975_ (
);

FILL FILL_2__7722_ (
);

FILL FILL_2__7302_ (
);

FILL FILL_3__12135_ (
);

FILL FILL_4__7228_ (
);

FILL FILL_2__11968_ (
);

FILL FILL_2__11548_ (
);

FILL FILL_0__12582_ (
);

FILL FILL_2__11128_ (
);

FILL SFILL68440x72050 (
);

FILL FILL_0__12162_ (
);

FILL SFILL49000x6050 (
);

FILL SFILL23720x2050 (
);

FILL FILL_5__15774_ (
);

FILL FILL_5__15354_ (
);

FILL FILL_0__7968_ (
);

FILL FILL_0__7548_ (
);

NAND2X1 _9654_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1410_)
);

NAND2X1 _9234_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1191_)
);

FILL FILL_1__8191_ (
);

FILL FILL_1__11902_ (
);

FILL FILL_4__14767_ (
);

FILL FILL_4__14347_ (
);

FILL FILL_2__15381_ (
);

FILL FILL_2__8507_ (
);

FILL FILL_1__14794_ (
);

FILL FILL_1__14374_ (
);

FILL FILL_5__6932_ (
);

FILL FILL_0__13787_ (
);

INVX1 _13652_ (
    .A(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_4160_)
);

FILL FILL_0__13367_ (
);

OAI21X1 _13232_ (
    .A(_3773_),
    .B(_3770_),
    .C(_3774_),
    .Y(_3775_)
);

FILL FILL_3__14701_ (
);

FILL FILL_1__6924_ (
);

FILL FILL_5__16139_ (
);

FILL SFILL64040x26050 (
);

FILL FILL_5__11694_ (
);

FILL FILL_1__9396_ (
);

FILL FILL_5__11274_ (
);

FILL FILL_2__16166_ (
);

FILL SFILL64120x50 (
);

FILL FILL_4__10687_ (
);

FILL FILL_4__10267_ (
);

FILL FILL_1__15999_ (
);

FILL SFILL54120x62050 (
);

FILL FILL_1__15579_ (
);

FILL FILL_1__15159_ (
);

FILL FILL_5__7717_ (
);

FILL FILL_2_BUFX2_insert510 (
);

FILL FILL_1__10294_ (
);

FILL FILL_2_BUFX2_insert511 (
);

FILL FILL_2_BUFX2_insert512 (
);

NOR2X1 _14857_ (
    .A(_5339_),
    .B(_5336_),
    .Y(_5340_)
);

FILL FILL_2_BUFX2_insert513 (
);

NOR2X1 _14437_ (
    .A(_4928_),
    .B(_4925_),
    .Y(_4929_)
);

FILL FILL_2_BUFX2_insert514 (
);

FILL FILL_2_BUFX2_insert515 (
);

INVX1 _14017_ (
    .A(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_4518_)
);

FILL FILL_3__15906_ (
);

FILL FILL_2_BUFX2_insert516 (
);

FILL SFILL38920x50 (
);

FILL FILL_2_BUFX2_insert517 (
);

FILL FILL_2_BUFX2_insert518 (
);

FILL FILL_2_BUFX2_insert519 (
);

FILL FILL_1__16100_ (
);

FILL FILL_1__7709_ (
);

FILL FILL_3__10621_ (
);

FILL FILL_0_CLKBUF1_insert210 (
);

FILL FILL_0_CLKBUF1_insert211 (
);

FILL FILL_0_CLKBUF1_insert212 (
);

FILL FILL_0__15933_ (
);

FILL FILL_0_CLKBUF1_insert213 (
);

FILL FILL_0__15513_ (
);

FILL FILL_0_CLKBUF1_insert214 (
);

FILL FILL_0_CLKBUF1_insert215 (
);

FILL FILL_5__12899_ (
);

FILL SFILL54040x69050 (
);

FILL FILL_0_CLKBUF1_insert216 (
);

FILL FILL_5__12479_ (
);

FILL FILL_0_CLKBUF1_insert217 (
);

FILL FILL_5__12059_ (
);

FILL FILL_2__8260_ (
);

FILL FILL_0_CLKBUF1_insert218 (
);

FILL FILL_3__13093_ (
);

FILL FILL_0_CLKBUF1_insert219 (
);

FILL FILL_4__8186_ (
);

FILL FILL_2__12086_ (
);

FILL FILL_5__13840_ (
);

FILL FILL_5__13420_ (
);

FILL FILL_5__13000_ (
);

OAI21X1 _7720_ (
    .A(_424_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .C(_425_),
    .Y(_393_[16])
);

OAI21X1 _7300_ (
    .A(_205_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_206_),
    .Y(_198_[4])
);

FILL FILL_1__11499_ (
);

FILL FILL_1__11079_ (
);

FILL FILL_4__12833_ (
);

FILL FILL_4__12413_ (
);

OAI21X1 _10777_ (
    .A(_1974_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .C(_1975_),
    .Y(_1953_[11])
);

FILL FILL_0__8086_ (
);

DFFSR _10357_ (
    .Q(\datapath_1.regfile_1.regOut[27] [31]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_1693_[31])
);

FILL FILL_3__11826_ (
);

FILL FILL_1__12860_ (
);

FILL FILL_3__11406_ (
);

FILL SFILL18680x50050 (
);

FILL FILL_1__12440_ (
);

FILL FILL_1__12020_ (
);

FILL FILL_4__6919_ (
);

FILL FILL_2__9885_ (
);

FILL FILL_2__10819_ (
);

FILL FILL_0__11853_ (
);

FILL FILL_2__9465_ (
);

FILL FILL_3__14298_ (
);

FILL FILL_2__9045_ (
);

FILL FILL_0__11433_ (
);

FILL FILL_0__11013_ (
);

FILL FILL_5__7890_ (
);

FILL SFILL54040x24050 (
);

FILL FILL_5__7470_ (
);

FILL FILL_5__7050_ (
);

INVX1 _14190_ (
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_4687_)
);

FILL FILL_5__14625_ (
);

FILL FILL_5__14205_ (
);

DFFSR _8925_ (
    .Q(\datapath_1.regfile_1.regOut[16] [7]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_978_[7])
);

NAND2X1 _8505_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_827_)
);

FILL SFILL79240x73050 (
);

FILL FILL_1__7882_ (
);

FILL FILL_1__7462_ (
);

FILL FILL_1__7042_ (
);

FILL FILL_4__13618_ (
);

FILL FILL_2__14652_ (
);

FILL FILL_2__14232_ (
);

FILL FILL_1__13645_ (
);

FILL FILL_1__13225_ (
);

FILL FILL_1_BUFX2_insert530 (
);

FILL FILL_1_BUFX2_insert531 (
);

FILL FILL_0__12638_ (
);

FILL FILL_1_BUFX2_insert532 (
);

DFFSR _12923_ (
    .Q(\datapath_1.a [4]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_3555_[4])
);

NAND2X1 _12503_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [21]),
    .Y(_3402_)
);

FILL FILL_1_BUFX2_insert533 (
);

FILL FILL_0__12218_ (
);

FILL FILL_1_BUFX2_insert534 (
);

FILL FILL_1_BUFX2_insert535 (
);

FILL FILL_1_BUFX2_insert536 (
);

FILL SFILL44040x67050 (
);

FILL FILL_5__8255_ (
);

FILL FILL_1_BUFX2_insert537 (
);

FILL FILL_1_BUFX2_insert538 (
);

FILL FILL_1_BUFX2_insert539 (
);

NOR2X1 _15395_ (
    .A(_5864_),
    .B(_5866_),
    .Y(_5867_)
);

FILL FILL_3__16024_ (
);

FILL FILL_5__10965_ (
);

FILL FILL_5__10545_ (
);

FILL FILL_5__10125_ (
);

FILL FILL_1__8247_ (
);

FILL SFILL33480x3050 (
);

FILL FILL_2__15857_ (
);

FILL FILL_2__15437_ (
);

FILL FILL_2__15017_ (
);

FILL FILL_0__16051_ (
);

FILL FILL_2__10992_ (
);

FILL FILL_2__10572_ (
);

FILL SFILL109800x68050 (
);

FILL FILL_2__10152_ (
);

FILL FILL_3__9534_ (
);

FILL FILL_3__9114_ (
);

OAI22X1 _13708_ (
    .A(_4214_),
    .B(_3902__bF$buf2),
    .C(_3954__bF$buf2),
    .D(_4213_),
    .Y(_4215_)
);

FILL FILL_0__6992_ (
);

FILL FILL_4__13791_ (
);

FILL FILL_4__13371_ (
);

FILL SFILL44040x22050 (
);

FILL FILL_2__7951_ (
);

FILL FILL_3__12784_ (
);

FILL FILL_3__12364_ (
);

FILL FILL_2__7111_ (
);

FILL SFILL84120x18050 (
);

FILL FILL_4__7877_ (
);

FILL SFILL69240x71050 (
);

FILL FILL_4__7457_ (
);

FILL FILL_4__7037_ (
);

FILL FILL_2__11777_ (
);

FILL FILL_2__11357_ (
);

FILL FILL_0__12391_ (
);

FILL FILL_5__15583_ (
);

FILL FILL_5__15163_ (
);

FILL FILL_0__7357_ (
);

NAND2X1 _9883_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1522_)
);

NAND2X1 _9463_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .Y(_1367_)
);

INVX1 _9043_ (
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_1104_)
);

FILL FILL_4__14996_ (
);

FILL FILL_4__14576_ (
);

FILL FILL_1__11711_ (
);

FILL FILL_4__14156_ (
);

FILL FILL_2__15190_ (
);

FILL FILL_2__8736_ (
);

FILL FILL_3__13989_ (
);

FILL FILL_3__13569_ (
);

FILL FILL_0__10704_ (
);

FILL FILL_2__8316_ (
);

FILL FILL_3__13149_ (
);

FILL FILL_1__14183_ (
);

INVX1 _13881_ (
    .A(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_4385_)
);

FILL FILL_0__13596_ (
);

OAI22X1 _13461_ (
    .A(_3972__bF$buf2),
    .B(_3969_),
    .C(_3971__bF$buf3),
    .D(_3970_),
    .Y(_3973_)
);

INVX1 _13041_ (
    .A(_2_[30]),
    .Y(_3679_)
);

FILL FILL_3__14930_ (
);

FILL FILL_3__14510_ (
);

FILL FILL_4__9603_ (
);

FILL FILL_6__12090_ (
);

FILL FILL_2__13923_ (
);

FILL FILL_5__16368_ (
);

FILL FILL_2__13503_ (
);

FILL FILL_6__9529_ (
);

FILL FILL_5__11083_ (
);

FILL FILL_1__12916_ (
);

FILL FILL_2__16395_ (
);

FILL FILL_4__10496_ (
);

FILL FILL_0__9923_ (
);

FILL SFILL69160x33050 (
);

FILL FILL_0__11909_ (
);

FILL FILL_3__7600_ (
);

FILL FILL_0__9503_ (
);

FILL FILL_1__15388_ (
);

FILL FILL_5__7946_ (
);

FILL FILL_4__16302_ (
);

FILL FILL_5__7106_ (
);

FILL FILL_6__10403_ (
);

NOR2X1 _14666_ (
    .A(_5152_),
    .B(_5149_),
    .Y(_5153_)
);

FILL SFILL74120x16050 (
);

OAI22X1 _14246_ (
    .A(_3884__bF$buf0),
    .B(_4740_),
    .C(_3966__bF$buf3),
    .D(_4741_),
    .Y(_4742_)
);

FILL SFILL28920x5050 (
);

FILL FILL_3__15715_ (
);

FILL FILL_1__7938_ (
);

FILL FILL_6__13295_ (
);

FILL FILL_3__10430_ (
);

FILL FILL_3__10010_ (
);

FILL FILL_2__14708_ (
);

FILL SFILL99320x65050 (
);

FILL FILL_0__15742_ (
);

FILL FILL_0__15322_ (
);

FILL FILL_5__12288_ (
);

BUFX2 BUFX2_insert0 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf4 )
);

BUFX2 BUFX2_insert1 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf3 )
);

BUFX2 BUFX2_insert2 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf2 )
);

BUFX2 BUFX2_insert3 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf1 )
);

BUFX2 BUFX2_insert4 (
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf0 )
);

BUFX2 BUFX2_insert5 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf7 )
);

BUFX2 BUFX2_insert6 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf6 )
);

FILL SFILL8760x6050 (
);

BUFX2 BUFX2_insert7 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf5 )
);

BUFX2 BUFX2_insert8 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf4 )
);

FILL SFILL24040x63050 (
);

BUFX2 BUFX2_insert9 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf3 )
);

FILL FILL_4__12642_ (
);

FILL FILL_4__12222_ (
);

DFFSR _10586_ (
    .Q(\datapath_1.regfile_1.regOut[29] [4]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1823_[4])
);

NAND2X1 _10166_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1670_)
);

FILL FILL_3__11635_ (
);

FILL FILL_3__11215_ (
);

FILL FILL_0__16107_ (
);

FILL FILL_2__10628_ (
);

FILL FILL_2__9274_ (
);

FILL FILL_0__11662_ (
);

FILL SFILL99320x20050 (
);

FILL FILL_0__11242_ (
);

FILL FILL_5__14854_ (
);

FILL FILL_5__14434_ (
);

FILL FILL_5__14014_ (
);

FILL SFILL28760x40050 (
);

NAND2X1 _8734_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_939_)
);

FILL SFILL59160x31050 (
);

NAND2X1 _8314_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_720_)
);

FILL FILL_1__7691_ (
);

FILL FILL_4__13847_ (
);

FILL SFILL89720x77050 (
);

FILL FILL_2__14881_ (
);

FILL FILL_4__13427_ (
);

FILL FILL_2__14461_ (
);

FILL FILL_4__13007_ (
);

FILL FILL_2__14041_ (
);

FILL FILL_3__7197_ (
);

FILL SFILL64120x14050 (
);

FILL FILL_1__13874_ (
);

FILL FILL_1__13454_ (
);

FILL FILL_1__13034_ (
);

FILL FILL_0__12867_ (
);

NAND2X1 _12732_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[12]),
    .Y(_3514_)
);

FILL FILL_0__12447_ (
);

FILL SFILL89320x63050 (
);

FILL FILL_0__12027_ (
);

NAND3X1 _12312_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3198__bF$buf0),
    .Y(_3273_)
);

FILL FILL_5__8484_ (
);

FILL SFILL68440x22050 (
);

FILL FILL_5__8064_ (
);

FILL FILL_5__15639_ (
);

FILL FILL_5__15219_ (
);

INVX1 _9939_ (
    .A(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_1559_)
);

FILL FILL_3__16253_ (
);

FILL SFILL18760x83050 (
);

INVX1 _9519_ (
    .A(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_1340_)
);

FILL FILL_1__8896_ (
);

FILL FILL_5__10774_ (
);

FILL FILL_1__8476_ (
);

FILL FILL_1__8056_ (
);

FILL FILL_2__15666_ (
);

FILL FILL_2__15246_ (
);

FILL FILL_0__16280_ (
);

FILL FILL_2__10381_ (
);

FILL FILL_1__14659_ (
);

FILL FILL_1__14239_ (
);

FILL FILL_3__9763_ (
);

FILL FILL_3__9343_ (
);

OAI22X1 _13937_ (
    .A(_3947__bF$buf2),
    .B(_4438_),
    .C(_3954__bF$buf0),
    .D(_4437_),
    .Y(_4439_)
);

OAI22X1 _13517_ (
    .A(_4027_),
    .B(_3905__bF$buf3),
    .C(_3955__bF$buf2),
    .D(_4026_),
    .Y(_4028_)
);

FILL FILL_5__9269_ (
);

FILL FILL_1__15600_ (
);

FILL FILL_6__12986_ (
);

FILL FILL_5__11979_ (
);

FILL FILL_2__7760_ (
);

FILL FILL_5__11559_ (
);

FILL FILL_3__12593_ (
);

FILL FILL_2__7340_ (
);

FILL FILL_5__11139_ (
);

FILL FILL_3__12173_ (
);

FILL FILL_4__7686_ (
);

FILL FILL_2__11586_ (
);

FILL FILL_2__11166_ (
);

FILL FILL_5__12500_ (
);

FILL SFILL89240x25050 (
);

FILL FILL_1__10999_ (
);

FILL SFILL54120x12050 (
);

FILL FILL_1__10579_ (
);

FILL FILL_1__10159_ (
);

FILL FILL_4__11913_ (
);

FILL FILL_5__15392_ (
);

FILL FILL_0__7586_ (
);

DFFSR _9692_ (
    .Q(\datapath_1.regfile_1.regOut[22] [6]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_1368_[6])
);

FILL FILL_0__7166_ (
);

FILL SFILL38760x1050 (
);

INVX1 _9272_ (
    .A(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_1216_)
);

FILL FILL_6__8133_ (
);

FILL SFILL79320x61050 (
);

FILL FILL_3__10906_ (
);

FILL SFILL18680x45050 (
);

FILL FILL_1__11940_ (
);

FILL FILL_4__14385_ (
);

FILL FILL_1__11520_ (
);

FILL FILL_1__11100_ (
);

FILL FILL_2__8965_ (
);

FILL FILL_0__10933_ (
);

FILL FILL_3__13798_ (
);

FILL FILL_2__8125_ (
);

FILL FILL_3__13378_ (
);

FILL FILL_0__10513_ (
);

FILL SFILL54040x19050 (
);

FILL FILL_5__6970_ (
);

AOI21X1 _13690_ (
    .A(\datapath_1.regfile_1.regOut[6] [5]),
    .B(_4001__bF$buf1),
    .C(_4196_),
    .Y(_4197_)
);

INVX1 _13270_ (
    .A(_3800_),
    .Y(_3811_)
);

FILL FILL_5__13705_ (
);

FILL FILL_1__6962_ (
);

FILL FILL_4__9412_ (
);

FILL FILL_2__13732_ (
);

FILL FILL_2__13312_ (
);

FILL FILL_5__16177_ (
);

FILL FILL_3__6888_ (
);

FILL FILL_6__9338_ (
);

FILL FILL_1__12725_ (
);

FILL FILL_1__12305_ (
);

FILL FILL_0__9732_ (
);

FILL FILL_0__11718_ (
);

FILL FILL_1__15197_ (
);

FILL FILL_5__7755_ (
);

FILL FILL_5__7335_ (
);

FILL FILL_4__16111_ (
);

INVX1 _14895_ (
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_5377_)
);

INVX1 _14475_ (
    .A(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_4966_)
);

NOR2X1 _14055_ (
    .A(_4554_),
    .B(_4551_),
    .Y(_4555_)
);

FILL FILL_3__15944_ (
);

FILL FILL_3__15524_ (
);

FILL FILL_3__15104_ (
);

FILL FILL_1__7747_ (
);

FILL FILL_1__7327_ (
);

FILL FILL_2__14937_ (
);

FILL SFILL79240x23050 (
);

FILL FILL_0__15971_ (
);

FILL FILL_2__14517_ (
);

FILL FILL_0__15551_ (
);

FILL FILL_0__15131_ (
);

FILL FILL_5__12097_ (
);

FILL FILL_3__8614_ (
);

FILL SFILL109400x49050 (
);

FILL FILL_4__12871_ (
);

FILL SFILL44040x17050 (
);

FILL FILL_4__12451_ (
);

FILL FILL_4__12031_ (
);

FILL FILL_3__16309_ (
);

NAND2X1 _10395_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1782_)
);

FILL FILL_3__11864_ (
);

FILL FILL_5__9901_ (
);

FILL FILL_3__11444_ (
);

FILL FILL_3__11024_ (
);

FILL SFILL69240x66050 (
);

FILL FILL_4__6957_ (
);

FILL FILL_0__16336_ (
);

NAND2X1 _16201_ (
    .A(_6647_),
    .B(_6652_),
    .Y(_6653_)
);

FILL SFILL109000x35050 (
);

FILL FILL_2__10437_ (
);

FILL FILL_0__11891_ (
);

FILL FILL_2__10017_ (
);

FILL FILL_2__9083_ (
);

FILL FILL_0__11471_ (
);

FILL FILL_0__11051_ (
);

FILL FILL_6__15250_ (
);

FILL FILL_5__14663_ (
);

FILL FILL_5__14243_ (
);

FILL FILL_0__6857_ (
);

FILL FILL_6__7824_ (
);

NAND2X1 _8963_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1051_)
);

DFFSR _8543_ (
    .Q(\datapath_1.regfile_1.regOut[13] [9]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_783_[9])
);

INVX1 _8123_ (
    .A(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_633_)
);

FILL FILL_1__7080_ (
);

FILL FILL_4__13656_ (
);

FILL FILL_4__13236_ (
);

FILL FILL_2__14690_ (
);

FILL FILL_2__14270_ (
);

FILL SFILL114280x55050 (
);

FILL FILL_2__7816_ (
);

FILL FILL_3__12649_ (
);

FILL FILL_1__13683_ (
);

FILL FILL_3__12229_ (
);

FILL FILL_1__13263_ (
);

FILL FILL_1_BUFX2_insert910 (
);

FILL FILL_1_BUFX2_insert911 (
);

NAND2X1 _12961_ (
    .A(vdd),
    .B(\datapath_1.rd2 [3]),
    .Y(_3626_)
);

FILL FILL_1_BUFX2_insert912 (
);

DFFSR _12541_ (
    .Q(ALUOut[6]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3360_[6])
);

FILL FILL_0__12256_ (
);

FILL FILL_1_BUFX2_insert913 (
);

INVX1 _12121_ (
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_3134_)
);

FILL FILL_1_BUFX2_insert914 (
);

FILL FILL_1_BUFX2_insert915 (
);

FILL FILL_1_BUFX2_insert916 (
);

FILL FILL_1_BUFX2_insert917 (
);

FILL FILL_1_BUFX2_insert918 (
);

FILL FILL_1_BUFX2_insert919 (
);

FILL FILL_6__11170_ (
);

FILL FILL_5__15868_ (
);

FILL FILL_5__15448_ (
);

FILL FILL_5__15028_ (
);

FILL FILL_6__8609_ (
);

FILL FILL_3__16062_ (
);

INVX1 _9748_ (
    .A(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_1452_)
);

DFFSR _9328_ (
    .Q(\datapath_1.regfile_1.regOut[19] [26]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_1173_[26])
);

FILL FILL_5__10163_ (
);

FILL FILL_2__15895_ (
);

FILL FILL_2__15475_ (
);

FILL FILL_2__15055_ (
);

FILL SFILL99400x53050 (
);

FILL SFILL69160x28050 (
);

FILL FILL_2__10190_ (
);

FILL FILL_1__14888_ (
);

FILL FILL_1__14468_ (
);

FILL FILL_1__14048_ (
);

FILL SFILL3400x72050 (
);

FILL FILL_4__15802_ (
);

FILL FILL_3__9992_ (
);

FILL FILL_3__9152_ (
);

INVX1 _13746_ (
    .A(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_4252_)
);

NOR2X1 _13326_ (
    .A(_3797_),
    .B(_3854_),
    .Y(\datapath_1.regfile_1.regEn [15])
);

FILL FILL_5__9498_ (
);

FILL FILL_5__9078_ (
);

FILL FILL_0__14822_ (
);

FILL FILL_0__14402_ (
);

FILL FILL_5__11788_ (
);

FILL FILL_5__11368_ (
);

FILL FILL_4__7495_ (
);

FILL FILL_4__7075_ (
);

FILL FILL_2__11395_ (
);

FILL FILL_1__10388_ (
);

FILL FILL_4__11722_ (
);

FILL FILL_4__11302_ (
);

INVX1 _9081_ (
    .A(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_1109_)
);

FILL FILL_4__14194_ (
);

FILL FILL_0__15607_ (
);

FILL FILL_2__8774_ (
);

FILL FILL_2__8354_ (
);

FILL FILL_0__10742_ (
);

FILL FILL_0__10322_ (
);

FILL FILL_5__13934_ (
);

FILL SFILL89400x51050 (
);

FILL FILL_5__13514_ (
);

FILL SFILL28760x35050 (
);

FILL SFILL59160x26050 (
);

NAND2X1 _7814_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_468_)
);

FILL FILL_4_BUFX2_insert420 (
);

FILL FILL_4_BUFX2_insert421 (
);

FILL FILL_4__9641_ (
);

FILL FILL_4_BUFX2_insert422 (
);

FILL FILL_4__9221_ (
);

FILL FILL_4__12507_ (
);

FILL FILL_4_BUFX2_insert423 (
);

FILL FILL_2__13961_ (
);

FILL FILL_4_BUFX2_insert424 (
);

FILL FILL_2__13541_ (
);

FILL FILL_4_BUFX2_insert425 (
);

FILL FILL_2__13121_ (
);

FILL FILL_4_BUFX2_insert426 (
);

FILL FILL_4_BUFX2_insert427 (
);

FILL FILL_4_BUFX2_insert428 (
);

FILL FILL_4_BUFX2_insert429 (
);

FILL FILL_1__12954_ (
);

FILL FILL_4__15399_ (
);

FILL FILL_1__12534_ (
);

FILL FILL_1__12114_ (
);

FILL FILL_2__9979_ (
);

FILL FILL_0__11947_ (
);

FILL FILL_0__9541_ (
);

FILL SFILL89320x58050 (
);

FILL FILL_0__9121_ (
);

FILL FILL_2__9139_ (
);

OAI21X1 _11812_ (
    .A(_2901_),
    .B(_2124_),
    .C(_2462__bF$buf0),
    .Y(_2903_)
);

FILL FILL_0__11527_ (
);

FILL FILL_0__11107_ (
);

FILL FILL_5__7984_ (
);

FILL FILL_5__7564_ (
);

FILL FILL_6__15306_ (
);

FILL FILL_4__16340_ (
);

FILL FILL_6__10021_ (
);

INVX1 _14284_ (
    .A(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_4779_)
);

FILL FILL_5__14719_ (
);

FILL FILL_3__15753_ (
);

FILL FILL_3__15333_ (
);

FILL FILL_1__7976_ (
);

FILL FILL_1__7556_ (
);

FILL FILL_2__14746_ (
);

FILL FILL_0__15780_ (
);

FILL FILL_2__14326_ (
);

FILL FILL_0__15360_ (
);

FILL FILL_1__13739_ (
);

FILL FILL_1__13319_ (
);

FILL FILL_3__8843_ (
);

FILL FILL_3__8003_ (
);

FILL SFILL33960x53050 (
);

FILL FILL_5__8769_ (
);

FILL FILL_5__8349_ (
);

FILL SFILL89320x13050 (
);

FILL FILL_6__11226_ (
);

INVX1 _15489_ (
    .A(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_5959_)
);

NAND3X1 _15069_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5477_),
    .C(_5476_),
    .Y(_5549_)
);

FILL FILL_4__12260_ (
);

FILL FILL_3__16118_ (
);

FILL SFILL113800x18050 (
);

FILL FILL_5__10639_ (
);

FILL FILL_2__6840_ (
);

FILL FILL_3__11673_ (
);

FILL FILL_3__11253_ (
);

FILL SFILL18760x33050 (
);

FILL FILL_0__16145_ (
);

DFFSR _16430_ (
    .Q(\datapath_1.regfile_1.regOut[0] [13]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_6769_[13])
);

AOI22X1 _16010_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [24]),
    .C(\datapath_1.regfile_1.regOut[22] [24]),
    .D(_5650_),
    .Y(_6466_)
);

FILL FILL_2__10666_ (
);

FILL FILL_2__10246_ (
);

FILL FILL_0__11280_ (
);

FILL FILL_3__9628_ (
);

FILL FILL_3_BUFX2_insert440 (
);

FILL FILL_3__9208_ (
);

FILL FILL_3_BUFX2_insert441 (
);

FILL FILL_3_BUFX2_insert442 (
);

FILL FILL_5__14892_ (
);

FILL FILL_5__14472_ (
);

FILL FILL_3_BUFX2_insert443 (
);

FILL FILL_3_BUFX2_insert444 (
);

FILL FILL_5__14052_ (
);

FILL FILL_3_BUFX2_insert445 (
);

INVX1 _8772_ (
    .A(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_964_)
);

INVX1 _8352_ (
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_745_)
);

FILL FILL_3_BUFX2_insert446 (
);

FILL FILL_6__7213_ (
);

FILL SFILL79320x56050 (
);

FILL FILL_3_BUFX2_insert447 (
);

FILL FILL_3_BUFX2_insert448 (
);

FILL FILL_4__13885_ (
);

FILL FILL_3_BUFX2_insert449 (
);

FILL FILL_4__13465_ (
);

FILL FILL_4__13045_ (
);

FILL FILL_3__12878_ (
);

FILL FILL_2__7625_ (
);

FILL FILL111960x69050 (
);

FILL FILL_2__7205_ (
);

FILL FILL_3__12458_ (
);

FILL FILL_3__12038_ (
);

FILL FILL_1__13492_ (
);

FILL SFILL39160x67050 (
);

INVX1 _12770_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_3539_)
);

FILL FILL_0__12485_ (
);

NAND2X1 _12350_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [2]),
    .Y(_3299_)
);

FILL FILL_0__12065_ (
);

FILL FILL_4__8912_ (
);

FILL FILL_5__15677_ (
);

FILL FILL_5__15257_ (
);

FILL FILL_3__16291_ (
);

INVX1 _9977_ (
    .A(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_1564_)
);

OAI21X1 _9557_ (
    .A(_1364_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .C(_1365_),
    .Y(_1303_[31])
);

OAI21X1 _9137_ (
    .A(_1145_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1146_),
    .Y(_1108_[19])
);

FILL FILL_5__10392_ (
);

FILL FILL_1__8094_ (
);

FILL FILL_1__11805_ (
);

FILL FILL_2__15284_ (
);

FILL SFILL114440x81050 (
);

FILL SFILL79320x11050 (
);

FILL FILL_1__14697_ (
);

FILL FILL_1__14277_ (
);

FILL FILL_0_BUFX2_insert570 (
);

FILL FILL_4__15611_ (
);

FILL FILL_0_BUFX2_insert571 (
);

FILL FILL_0_BUFX2_insert572 (
);

FILL FILL_0_BUFX2_insert573 (
);

FILL FILL_3__9381_ (
);

AOI21X1 _13975_ (
    .A(_4476_),
    .B(_4455_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [10])
);

FILL FILL_0_BUFX2_insert574 (
);

FILL FILL_0_BUFX2_insert575 (
);

INVX1 _13555_ (
    .A(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_4065_)
);

OAI21X1 _13135_ (
    .A(_3720_),
    .B(PCEn_bF$buf5),
    .C(_3721_),
    .Y(_3685_[18])
);

FILL FILL_0_BUFX2_insert576 (
);

FILL FILL_0_BUFX2_insert577 (
);

FILL FILL_0_BUFX2_insert578 (
);

FILL FILL_3__14604_ (
);

FILL FILL_0_BUFX2_insert579 (
);

FILL SFILL79240x18050 (
);

FILL FILL_0__14631_ (
);

FILL FILL_0__14211_ (
);

FILL FILL_5__11597_ (
);

FILL FILL_1__9299_ (
);

FILL FILL_5__11177_ (
);

FILL FILL_2__16069_ (
);

FILL FILL_1__10197_ (
);

FILL FILL_4__11951_ (
);

FILL FILL_4__11531_ (
);

FILL FILL_4__11111_ (
);

FILL FILL_3__15809_ (
);

FILL FILL_1__16003_ (
);

FILL FILL_3__10944_ (
);

FILL FILL_3__10524_ (
);

FILL FILL_3__10104_ (
);

FILL FILL_0__15836_ (
);

NOR3X1 _15701_ (
    .A(_4735_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6165_)
);

FILL FILL_0__15416_ (
);

FILL FILL_0__10971_ (
);

FILL FILL_2__8583_ (
);

FILL FILL_0__10551_ (
);

FILL FILL_0__10131_ (
);

FILL FILL_4__8089_ (
);

FILL FILL_5__13743_ (
);

FILL FILL_5__13323_ (
);

FILL FILL_6__6904_ (
);

INVX1 _7623_ (
    .A(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_381_)
);

INVX1 _7203_ (
    .A(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_162_)
);

FILL FILL_4__9870_ (
);

FILL FILL_4__12736_ (
);

FILL FILL_4__9030_ (
);

FILL FILL_2__13770_ (
);

FILL FILL_4__12316_ (
);

FILL FILL_2__13350_ (
);

FILL FILL_3__11729_ (
);

FILL FILL_1__12763_ (
);

FILL FILL_3__11309_ (
);

FILL FILL_1__12343_ (
);

FILL FILL_0__9770_ (
);

FILL FILL_2__9788_ (
);

FILL SFILL53640x31050 (
);

FILL SFILL69240x16050 (
);

FILL FILL_2__9368_ (
);

FILL FILL_0__11756_ (
);

FILL FILL_0__9350_ (
);

FILL FILL_0__11336_ (
);

OAI22X1 _11621_ (
    .A(_2250_),
    .B(_2346_),
    .C(_2347__bF$buf1),
    .D(_2252_),
    .Y(_2726_)
);

NOR2X1 _11201_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .Y(_2320_)
);

FILL FILL_5__7373_ (
);

FILL FILL_5__14948_ (
);

AOI22X1 _14093_ (
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .B(_4135_),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_4592_)
);

FILL FILL_3__15982_ (
);

FILL FILL_5__14528_ (
);

FILL FILL_3__15562_ (
);

FILL FILL_5__14108_ (
);

FILL FILL_3__15142_ (
);

INVX1 _8828_ (
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_981_)
);

DFFSR _8408_ (
    .Q(\datapath_1.regfile_1.regOut[12] [2]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_718_[2])
);

FILL FILL_1__7365_ (
);

FILL FILL_2__14975_ (
);

FILL FILL_2__14555_ (
);

FILL SFILL99400x48050 (
);

FILL FILL_2__14135_ (
);

FILL FILL_1__13968_ (
);

FILL FILL_1__13548_ (
);

FILL SFILL3400x67050 (
);

FILL FILL_1__13128_ (
);

FILL FILL_1_CLKBUF1_insert1080 (
);

FILL FILL_1_CLKBUF1_insert1081 (
);

FILL FILL_1_CLKBUF1_insert1082 (
);

FILL FILL_1_CLKBUF1_insert1083 (
);

FILL FILL_3__8652_ (
);

FILL FILL_3__8232_ (
);

INVX1 _12826_ (
    .A(\datapath_1.a [1]),
    .Y(_3556_)
);

INVX1 _12406_ (
    .A(ALUOut[21]),
    .Y(_3336_)
);

FILL FILL_5__8998_ (
);

FILL FILL_5__8578_ (
);

FILL SFILL104360x41050 (
);

AOI22X1 _15298_ (
    .A(\datapath_1.regfile_1.regOut[31] [6]),
    .B(_5571_),
    .C(_5486_),
    .D(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_5772_)
);

FILL FILL_0__13902_ (
);

FILL FILL_3__16347_ (
);

FILL FILL_5__10448_ (
);

FILL FILL_5__10028_ (
);

FILL FILL_3__11482_ (
);

FILL FILL_3__11062_ (
);

FILL FILL_4__6995_ (
);

FILL FILL_0__16374_ (
);

FILL FILL_2__10895_ (
);

FILL FILL_2__10055_ (
);

FILL FILL_1__9931_ (
);

FILL FILL_1__9511_ (
);

FILL FILL_3__9857_ (
);

FILL SFILL49720x64050 (
);

FILL FILL_3__9017_ (
);

FILL FILL_4__10802_ (
);

FILL FILL_5__14281_ (
);

FILL FILL_0__6895_ (
);

INVX1 _8581_ (
    .A(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_857_)
);

DFFSR _8161_ (
    .Q(\datapath_1.regfile_1.regOut[10] [11]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_588_[11])
);

FILL SFILL85000x9050 (
);

FILL FILL_4__13694_ (
);

FILL FILL_4__13274_ (
);

FILL FILL_2__7854_ (
);

FILL FILL_2__7434_ (
);

FILL SFILL104680x17050 (
);

FILL FILL_3__12267_ (
);

FILL FILL_0__12294_ (
);

FILL SFILL89400x46050 (
);

FILL FILL_6__16073_ (
);

FILL FILL_4__8721_ (
);

FILL FILL_2__12621_ (
);

FILL FILL_5__15486_ (
);

FILL FILL_5__15066_ (
);

FILL FILL_2__12201_ (
);

OAI21X1 _9786_ (
    .A(_1476_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .C(_1477_),
    .Y(_1433_[22])
);

OAI21X1 _9366_ (
    .A(_1257_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .C(_1258_),
    .Y(_1238_[10])
);

FILL FILL_4__14899_ (
);

FILL FILL_4__14479_ (
);

FILL FILL_1__11614_ (
);

FILL SFILL28360x16050 (
);

FILL FILL_4__14059_ (
);

FILL FILL_2__15093_ (
);

FILL FILL_2__8639_ (
);

FILL FILL_0__8621_ (
);

FILL FILL_0__8201_ (
);

FILL FILL_2__8219_ (
);

FILL FILL_1__14086_ (
);

FILL FILL_4__15840_ (
);

FILL FILL_4__15420_ (
);

FILL FILL_4__15000_ (
);

INVX1 _13784_ (
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_4290_)
);

FILL FILL_0__13499_ (
);

NOR2X1 _13364_ (
    .A(_3874_),
    .B(_3877_),
    .Y(\datapath_1.regfile_1.regEn [30])
);

FILL FILL_0__13079_ (
);

FILL FILL_3__14833_ (
);

FILL FILL_3__14413_ (
);

FILL FILL_4__9926_ (
);

FILL FILL_4__9506_ (
);

FILL SFILL94280x52050 (
);

FILL FILL_2__13826_ (
);

FILL FILL_0__14860_ (
);

FILL FILL_2__13406_ (
);

FILL FILL_0__14440_ (
);

FILL FILL_0__14020_ (
);

FILL FILL_2__16298_ (
);

CLKBUF1 CLKBUF1_insert120 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf104)
);

CLKBUF1 CLKBUF1_insert121 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf103)
);

CLKBUF1 CLKBUF1_insert122 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf102)
);

FILL FILL_4__10399_ (
);

CLKBUF1 CLKBUF1_insert123 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf101)
);

FILL FILL_3__7503_ (
);

FILL FILL_0__9406_ (
);

CLKBUF1 CLKBUF1_insert124 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf100)
);

CLKBUF1 CLKBUF1_insert125 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf99)
);

CLKBUF1 CLKBUF1_insert126 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf98)
);

CLKBUF1 CLKBUF1_insert127 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf97)
);

CLKBUF1 CLKBUF1_insert128 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf96)
);

FILL FILL_5__7849_ (
);

CLKBUF1 CLKBUF1_insert129 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf95)
);

FILL FILL_5__7429_ (
);

FILL FILL_4__16205_ (
);

NAND3X1 _14989_ (
    .A(_5459__bF$buf1),
    .B(_5462_),
    .C(_5468_),
    .Y(_5469_)
);

NAND3X1 _14569_ (
    .A(_5049_),
    .B(_5050_),
    .C(_5057_),
    .Y(_5058_)
);

FILL FILL_4__11760_ (
);

OAI22X1 _14149_ (
    .A(_4645_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf3),
    .D(_4646_),
    .Y(_4647_)
);

FILL FILL_4__11340_ (
);

FILL FILL_3__15618_ (
);

FILL FILL_1__16232_ (
);

FILL FILL_3__10753_ (
);

FILL SFILL18760x28050 (
);

FILL FILL_0__15645_ (
);

OAI22X1 _15930_ (
    .A(_5504__bF$buf3),
    .B(_5030_),
    .C(_5527__bF$buf1),
    .D(_5010_),
    .Y(_6388_)
);

FILL FILL_0__15225_ (
);

NAND3X1 _15510_ (
    .A(_5977_),
    .B(_5978_),
    .C(_5976_),
    .Y(_5979_)
);

FILL FILL_0__10780_ (
);

FILL FILL_2__8392_ (
);

FILL FILL_0__10360_ (
);

FILL FILL_3__8708_ (
);

FILL FILL_5__13972_ (
);

FILL FILL_5__13552_ (
);

FILL FILL_5__13132_ (
);

INVX1 _7852_ (
    .A(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_493_)
);

INVX1 _7432_ (
    .A(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_274_)
);

FILL FILL_4_BUFX2_insert800 (
);

DFFSR _7012_ (
    .Q(\datapath_1.regfile_1.regOut[1] [14]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_3_[14])
);

FILL FILL_4_BUFX2_insert801 (
);

FILL FILL_4__12965_ (
);

FILL FILL_4_BUFX2_insert802 (
);

FILL FILL_4_BUFX2_insert803 (
);

FILL FILL_4__12125_ (
);

FILL FILL_4_BUFX2_insert804 (
);

FILL FILL_4_BUFX2_insert805 (
);

FILL FILL_4_BUFX2_insert806 (
);

FILL FILL_4_BUFX2_insert807 (
);

INVX1 _10489_ (
    .A(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_1824_)
);

FILL FILL_4_BUFX2_insert808 (
);

OAI21X1 _10069_ (
    .A(_1624_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .C(_1625_),
    .Y(_1563_[31])
);

FILL FILL_4_BUFX2_insert809 (
);

FILL FILL_3__11958_ (
);

FILL FILL_1__12992_ (
);

FILL FILL_3__11538_ (
);

FILL FILL_1__12572_ (
);

FILL FILL_3__11118_ (
);

FILL FILL_1__12152_ (
);

FILL FILL_0__11985_ (
);

FILL FILL_2__9597_ (
);

NOR3X1 _11850_ (
    .A(_2923_),
    .B(\datapath_1.ALUResult [0]),
    .C(_2929_),
    .Y(_2937_)
);

FILL FILL_0__11565_ (
);

INVX1 _11430_ (
    .A(_2375_),
    .Y(_2546_)
);

FILL FILL_0__11145_ (
);

NAND2X1 _11010_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2129_)
);

FILL FILL_5__7182_ (
);

FILL FILL_5__14757_ (
);

FILL FILL_3__15791_ (
);

FILL FILL_5__14337_ (
);

FILL FILL_3__15371_ (
);

OAI21X1 _8637_ (
    .A(_893_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .C(_894_),
    .Y(_848_[23])
);

OAI21X1 _8217_ (
    .A(_674_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .C(_675_),
    .Y(_653_[11])
);

FILL FILL_1__7594_ (
);

FILL FILL_1__7174_ (
);

FILL FILL_2__14784_ (
);

FILL FILL_2__14364_ (
);

FILL FILL_1__13777_ (
);

FILL FILL_1__13357_ (
);

FILL SFILL94200x2050 (
);

FILL FILL111960x19050 (
);

FILL FILL_3__8881_ (
);

FILL FILL_3__8461_ (
);

OAI21X1 _12635_ (
    .A(_3468_),
    .B(vdd),
    .C(_3469_),
    .Y(_3425_[22])
);

NOR2X1 _12215_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(ALUSrcB_1_bF$buf0),
    .Y(_3200_)
);

FILL FILL_5__8387_ (
);

FILL FILL_0__13711_ (
);

FILL FILL_3__16156_ (
);

FILL FILL_5__10677_ (
);

FILL FILL_1__8379_ (
);

FILL FILL_5__10257_ (
);

FILL FILL_3__11291_ (
);

FILL FILL_2__15989_ (
);

FILL FILL_2__15569_ (
);

FILL SFILL69320x49050 (
);

FILL FILL_2__15149_ (
);

FILL FILL_0__16183_ (
);

FILL FILL_2__10284_ (
);

FILL SFILL114440x31050 (
);

FILL FILL_1__9740_ (
);

FILL FILL_3_BUFX2_insert820 (
);

FILL FILL_3__9666_ (
);

FILL FILL_3_BUFX2_insert821 (
);

FILL FILL_3__9246_ (
);

FILL FILL_3_BUFX2_insert822 (
);

FILL SFILL109560x1050 (
);

FILL FILL_3_BUFX2_insert823 (
);

FILL FILL_3_BUFX2_insert824 (
);

FILL FILL_5__14090_ (
);

FILL FILL_3_BUFX2_insert825 (
);

FILL FILL_1__15923_ (
);

FILL FILL_1__15503_ (
);

OAI21X1 _8390_ (
    .A(_769_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .C(_770_),
    .Y(_718_[26])
);

FILL FILL_3_BUFX2_insert826 (
);

FILL FILL_3_BUFX2_insert827 (
);

FILL FILL_3_BUFX2_insert828 (
);

FILL FILL_3_BUFX2_insert829 (
);

FILL FILL_6__12469_ (
);

FILL FILL_4__13083_ (
);

FILL FILL_0__14916_ (
);

FILL FILL_2__7243_ (
);

FILL FILL_3__12496_ (
);

FILL FILL_3__12076_ (
);

FILL SFILL59800x54050 (
);

FILL FILL_4__7589_ (
);

FILL FILL_4__7169_ (
);

FILL FILL_2__11489_ (
);

FILL FILL_2__11069_ (
);

FILL FILL_5__12823_ (
);

FILL FILL_5__12403_ (
);

FILL FILL_4__8950_ (
);

FILL FILL_4__8530_ (
);

FILL FILL_4__8110_ (
);

FILL FILL_4__11816_ (
);

FILL FILL_2__12850_ (
);

FILL FILL_2__12430_ (
);

FILL FILL_5__15295_ (
);

FILL FILL_2__12010_ (
);

FILL FILL_0__7489_ (
);

OAI21X1 _9595_ (
    .A(_1369_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .C(_1370_),
    .Y(_1368_[1])
);

FILL FILL_0__7069_ (
);

DFFSR _9175_ (
    .Q(\datapath_1.regfile_1.regOut[18] [1]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_1108_[1])
);

FILL FILL_3__10809_ (
);

FILL FILL_1__11843_ (
);

FILL FILL_4__14288_ (
);

FILL FILL_1__11423_ (
);

FILL FILL_1__11003_ (
);

FILL FILL_2__8868_ (
);

FILL FILL_0__8850_ (
);

FILL FILL_2__8448_ (
);

FILL FILL_0__10836_ (
);

INVX1 _10701_ (
    .A(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_1945_)
);

FILL FILL_0__8010_ (
);

FILL FILL_0__10416_ (
);

FILL FILL_5__6873_ (
);

FILL FILL_6__14615_ (
);

FILL FILL_0_BUFX2_insert950 (
);

FILL FILL_0_BUFX2_insert951 (
);

FILL FILL_0_BUFX2_insert952 (
);

FILL FILL_0_BUFX2_insert953 (
);

FILL FILL_0_BUFX2_insert954 (
);

FILL FILL_0_BUFX2_insert955 (
);

AND2X2 _13593_ (
    .A(_3889_),
    .B(_3904_),
    .Y(_4102_)
);

FILL FILL_0_BUFX2_insert956 (
);

NAND2X1 _13173_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_pcsrc.dout [31]),
    .Y(_3747_)
);

FILL FILL_5__13608_ (
);

FILL FILL_0_BUFX2_insert957 (
);

FILL SFILL64680x60050 (
);

FILL FILL_3__14642_ (
);

FILL FILL_0_BUFX2_insert958 (
);

FILL FILL_3__14222_ (
);

DFFSR _7908_ (
    .Q(\datapath_1.regfile_1.regOut[8] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_458_[14])
);

FILL FILL_0_BUFX2_insert959 (
);

FILL FILL_1__6865_ (
);

FILL FILL_4__9735_ (
);

FILL FILL_2__13635_ (
);

FILL FILL_2__13215_ (
);

FILL FILL_1__12628_ (
);

FILL FILL_1__12208_ (
);

FILL FILL_0__9635_ (
);

FILL FILL_3__7732_ (
);

FILL FILL_0__9215_ (
);

FILL FILL_3__7312_ (
);

NAND2X1 _11906_ (
    .A(IorD_bF$buf0),
    .B(ALUOut[6]),
    .Y(_2979_)
);

FILL SFILL104360x36050 (
);

FILL FILL_5__7238_ (
);

FILL FILL_4__16014_ (
);

INVX1 _14798_ (
    .A(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_5282_)
);

AOI21X1 _14378_ (
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .B(_4225_),
    .C(_4870_),
    .Y(_4871_)
);

FILL FILL_3__15847_ (
);

FILL FILL_3__15427_ (
);

FILL SFILL64200x1050 (
);

FILL FILL_3__15007_ (
);

FILL FILL_1__16041_ (
);

FILL FILL112040x73050 (
);

FILL FILL_3__10982_ (
);

FILL FILL_3__10562_ (
);

FILL FILL_6_BUFX2_insert331 (
);

FILL FILL_3__10142_ (
);

FILL FILL_0__15874_ (
);

FILL FILL_0__15454_ (
);

FILL FILL_0__15034_ (
);

FILL FILL_6_BUFX2_insert336 (
);

FILL FILL_3__8517_ (
);

FILL FILL_5__13781_ (
);

FILL FILL_5__13361_ (
);

FILL FILL112440x42050 (
);

DFFSR _7661_ (
    .Q(\datapath_1.regfile_1.regOut[6] [23]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_328_[23])
);

OAI21X1 _7241_ (
    .A(_186_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .C(_187_),
    .Y(_133_[27])
);

FILL FILL_4__12774_ (
);

FILL FILL_4__12354_ (
);

OAI21X1 _10298_ (
    .A(_1736_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1737_),
    .Y(_1693_[22])
);

FILL FILL_2__6934_ (
);

FILL SFILL49320x45050 (
);

FILL FILL_5__9804_ (
);

FILL FILL_3__11767_ (
);

FILL FILL_3__11347_ (
);

FILL FILL_1__12381_ (
);

FILL FILL_0__16239_ (
);

OAI22X1 _16104_ (
    .A(_5466__bF$buf4),
    .B(_5220_),
    .C(_5218_),
    .D(_5483__bF$buf2),
    .Y(_6558_)
);

FILL FILL_0__11794_ (
);

FILL FILL_0__11374_ (
);

FILL FILL_6__15153_ (
);

FILL FILL_4__7801_ (
);

FILL FILL_5__14986_ (
);

FILL FILL_5__14566_ (
);

FILL FILL_2__11701_ (
);

FILL FILL_5__14146_ (
);

FILL FILL_3__15180_ (
);

OAI21X1 _8866_ (
    .A(_1005_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1006_),
    .Y(_978_[14])
);

FILL SFILL33640x67050 (
);

FILL FILL_6__7307_ (
);

OAI21X1 _8446_ (
    .A(_786_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_787_),
    .Y(_783_[2])
);

DFFSR _8026_ (
    .Q(\datapath_1.regfile_1.regOut[9] [4]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_523_[4])
);

FILL FILL_4__13979_ (
);

FILL FILL_4__13559_ (
);

FILL FILL_2__14593_ (
);

FILL FILL_4__13139_ (
);

FILL FILL_2__14173_ (
);

FILL FILL_2__7719_ (
);

FILL FILL_0__7701_ (
);

FILL FILL_1__13586_ (
);

FILL FILL_1__13166_ (
);

FILL FILL_4__14920_ (
);

FILL FILL_4__14500_ (
);

FILL FILL_0__12999_ (
);

FILL FILL_3__8270_ (
);

FILL FILL_0__12579_ (
);

OAI21X1 _12864_ (
    .A(_3580_),
    .B(vdd),
    .C(_3581_),
    .Y(_3555_[13])
);

FILL FILL_0__12159_ (
);

OAI21X1 _12444_ (
    .A(_3361_),
    .B(vdd),
    .C(_3362_),
    .Y(_3360_[1])
);

NAND3X1 _12024_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [9]),
    .C(_3034__bF$buf3),
    .Y(_3064_)
);

FILL FILL_3__13913_ (
);

FILL FILL_5__8196_ (
);

FILL FILL_5_BUFX2_insert350 (
);

FILL FILL_2__12906_ (
);

FILL FILL_5_BUFX2_insert351 (
);

FILL FILL_5_BUFX2_insert352 (
);

FILL FILL_0__13940_ (
);

FILL FILL_5_BUFX2_insert353 (
);

FILL FILL_3__16385_ (
);

FILL FILL_0__13520_ (
);

FILL FILL_5_BUFX2_insert354 (
);

FILL FILL_0__13100_ (
);

FILL FILL_5_BUFX2_insert355 (
);

FILL FILL_5_BUFX2_insert356 (
);

FILL FILL_5__10486_ (
);

FILL FILL_5_BUFX2_insert357 (
);

FILL FILL_5__10066_ (
);

FILL FILL_1__8188_ (
);

FILL FILL_5_BUFX2_insert358 (
);

FILL FILL_2__15798_ (
);

FILL FILL_5_BUFX2_insert359 (
);

FILL SFILL33640x22050 (
);

FILL FILL_2__15378_ (
);

FILL FILL_0__8906_ (
);

FILL SFILL94600x59050 (
);

FILL FILL_5__6929_ (
);

FILL FILL_4__15705_ (
);

FILL SFILL39320x43050 (
);

FILL FILL_3__9895_ (
);

FILL FILL_3__9475_ (
);

INVX1 _13649_ (
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_4157_)
);

NOR2X1 _13229_ (
    .A(\datapath_1.a3 [3]),
    .B(_3771_),
    .Y(_3772_)
);

FILL FILL_4__10420_ (
);

FILL FILL_4__10000_ (
);

FILL FILL_1__15732_ (
);

FILL FILL_1__15312_ (
);

FILL FILL_0__14725_ (
);

FILL FILL_0__14305_ (
);

FILL FILL_2__7892_ (
);

FILL FILL_2__7472_ (
);

FILL FILL_2__7052_ (
);

FILL SFILL103880x60050 (
);

FILL FILL_2__11298_ (
);

FILL FILL_5__12632_ (
);

FILL SFILL33800x8050 (
);

FILL FILL_5__12212_ (
);

INVX1 _6932_ (
    .A(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_22_)
);

FILL SFILL8680x64050 (
);

FILL FILL_2_BUFX2_insert480 (
);

FILL FILL_2_BUFX2_insert481 (
);

FILL FILL_2_BUFX2_insert482 (
);

FILL FILL_2_BUFX2_insert483 (
);

FILL SFILL74280x8050 (
);

FILL FILL_4__11625_ (
);

FILL FILL_2_BUFX2_insert484 (
);

FILL FILL_2_BUFX2_insert485 (
);

FILL FILL_4__11205_ (
);

FILL FILL_2_BUFX2_insert486 (
);

FILL FILL_0__7298_ (
);

FILL FILL_2_BUFX2_insert487 (
);

FILL FILL_2_BUFX2_insert488 (
);

FILL FILL_2_BUFX2_insert489 (
);

FILL FILL_3__10618_ (
);

FILL FILL_0_CLKBUF1_insert180 (
);

FILL FILL_1__11652_ (
);

FILL SFILL33800x50 (
);

FILL FILL_0_CLKBUF1_insert181 (
);

FILL FILL_1__11232_ (
);

FILL FILL_4__14097_ (
);

FILL FILL_0_CLKBUF1_insert182 (
);

FILL FILL_0_CLKBUF1_insert183 (
);

FILL FILL_0_CLKBUF1_insert184 (
);

FILL SFILL84280x45050 (
);

FILL FILL_0_CLKBUF1_insert185 (
);

FILL FILL_0_CLKBUF1_insert186 (
);

NOR2X1 _10930_ (
    .A(\control_1.op [4]),
    .B(\control_1.op [5]),
    .Y(_2064_)
);

FILL FILL_0_CLKBUF1_insert187 (
);

FILL FILL_0__10645_ (
);

FILL FILL_2__8257_ (
);

INVX1 _10510_ (
    .A(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_1838_)
);

FILL FILL_0_CLKBUF1_insert188 (
);

FILL FILL_0_CLKBUF1_insert189 (
);

FILL FILL_5__13837_ (
);

FILL FILL_3__14871_ (
);

FILL FILL_5__13417_ (
);

FILL FILL_3__14451_ (
);

FILL SFILL8600x62050 (
);

OAI21X1 _7717_ (
    .A(_422_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .C(_423_),
    .Y(_393_[15])
);

FILL FILL_3__14031_ (
);

FILL FILL_4__9544_ (
);

FILL FILL_4__9124_ (
);

FILL FILL_2__13864_ (
);

FILL FILL_2__13444_ (
);

FILL FILL_2__13024_ (
);

FILL FILL_1__12857_ (
);

FILL FILL_1__12437_ (
);

FILL FILL_1__12017_ (
);

FILL SFILL84200x43050 (
);

FILL FILL_0__9864_ (
);

FILL FILL_3__7961_ (
);

FILL FILL_3__7121_ (
);

OAI21X1 _11715_ (
    .A(_2812_),
    .B(_2188_),
    .C(_2470__bF$buf1),
    .Y(_2814_)
);

FILL FILL_0__9024_ (
);

FILL FILL_5__7887_ (
);

FILL FILL_6__15209_ (
);

FILL FILL_5__7467_ (
);

FILL FILL_4__16243_ (
);

FILL FILL_5__7047_ (
);

FILL SFILL13640x63050 (
);

INVX1 _14187_ (
    .A(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_4684_)
);

FILL FILL_3__15656_ (
);

FILL FILL_3__15236_ (
);

FILL SFILL109480x43050 (
);

FILL FILL_1__16270_ (
);

FILL FILL_1__7879_ (
);

FILL FILL_1__7459_ (
);

FILL FILL_3__10791_ (
);

FILL FILL_1__7039_ (
);

FILL FILL_3__10371_ (
);

FILL FILL_2__14649_ (
);

FILL FILL_2__14229_ (
);

FILL FILL_0__15683_ (
);

FILL FILL_0__15263_ (
);

FILL SFILL114440x26050 (
);

FILL FILL_1__8400_ (
);

FILL FILL_3__8746_ (
);

FILL FILL_3__8326_ (
);

FILL SFILL88920x20050 (
);

FILL FILL_5__13590_ (
);

FILL FILL_5__13170_ (
);

OAI21X1 _7890_ (
    .A(_517_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_518_),
    .Y(_458_[30])
);

OAI21X1 _7470_ (
    .A(_298_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .C(_299_),
    .Y(_263_[18])
);

OAI21X1 _7050_ (
    .A(_79_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_80_),
    .Y(_68_[6])
);

FILL FILL_4__12583_ (
);

FILL FILL_6__11129_ (
);

FILL FILL_4__12163_ (
);

FILL FILL_3__11996_ (
);

FILL FILL_5__9613_ (
);

FILL FILL_3__11576_ (
);

FILL FILL_3__11156_ (
);

FILL FILL_1__12190_ (
);

INVX1 _16333_ (
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .Y(_6776_)
);

FILL FILL_0__16048_ (
);

FILL FILL_2__10989_ (
);

FILL FILL_2__10569_ (
);

FILL FILL_2__10149_ (
);

FILL FILL_0__11183_ (
);

FILL FILL_5__11903_ (
);

FILL FILL_1__9605_ (
);

FILL FILL_4__7610_ (
);

FILL FILL_5__14795_ (
);

FILL FILL_2__11930_ (
);

FILL FILL_0__6989_ (
);

FILL FILL_5__14375_ (
);

FILL FILL_2__11510_ (
);

DFFSR _8675_ (
    .Q(\datapath_1.regfile_1.regOut[14] [13]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_848_[13])
);

NAND2X1 _8255_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_701_)
);

FILL FILL_1__10923_ (
);

FILL FILL_4__13788_ (
);

FILL FILL_4__13368_ (
);

FILL FILL_1__10503_ (
);

FILL FILL_2__7948_ (
);

FILL FILL_0__7930_ (
);

FILL FILL_2__7108_ (
);

FILL FILL_1__13395_ (
);

FILL SFILL69000x3050 (
);

FILL SFILL43720x57050 (
);

FILL FILL_0__12388_ (
);

DFFSR _12673_ (
    .Q(\datapath_1.Data [10]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3425_[10])
);

AOI22X1 _12253_ (
    .A(_2_[9]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump [9]),
    .Y(_3229_)
);

FILL FILL_3__13722_ (
);

FILL FILL_3__13302_ (
);

FILL FILL_2__12715_ (
);

FILL FILL_3__16194_ (
);

FILL FILL_5__10295_ (
);

FILL FILL112120x61050 (
);

FILL FILL_1__11708_ (
);

FILL FILL_2__15187_ (
);

FILL FILL_0__8715_ (
);

FILL FILL_5__16101_ (
);

FILL FILL_4__15934_ (
);

FILL FILL_4__15514_ (
);

INVX1 _13878_ (
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_4382_)
);

FILL FILL_3__9284_ (
);

INVX1 _13458_ (
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_3970_)
);

FILL SFILL18760x50 (
);

INVX1 _13038_ (
    .A(_2_[29]),
    .Y(_3677_)
);

FILL FILL_3__14927_ (
);

FILL FILL_3__14507_ (
);

FILL FILL_1__15961_ (
);

FILL FILL_1__15541_ (
);

FILL FILL112040x68050 (
);

FILL FILL_1__15121_ (
);

FILL FILL_0__14954_ (
);

FILL FILL_0__14534_ (
);

FILL FILL_0__14114_ (
);

FILL FILL_5__12861_ (
);

FILL FILL_5__12441_ (
);

FILL FILL112440x37050 (
);

FILL FILL_5__12021_ (
);

FILL FILL_4__11854_ (
);

FILL FILL_4__11434_ (
);

FILL FILL_4__11014_ (
);

FILL FILL_1__16326_ (
);

FILL SFILL33720x55050 (
);

FILL FILL_3__10427_ (
);

FILL FILL_1__11881_ (
);

FILL FILL_3__10007_ (
);

FILL FILL_1__11461_ (
);

FILL FILL_1__11041_ (
);

FILL FILL_0__15739_ (
);

FILL FILL_0__15319_ (
);

INVX1 _15604_ (
    .A(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_6071_)
);

FILL FILL_2__8486_ (
);

FILL FILL_0__10874_ (
);

FILL FILL_2__8066_ (
);

FILL FILL_0__10034_ (
);

FILL FILL_5__13646_ (
);

FILL FILL_5__13226_ (
);

FILL FILL_3__14680_ (
);

OAI21X1 _7946_ (
    .A(_534_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_535_),
    .Y(_523_[6])
);

FILL FILL_3__14260_ (
);

DFFSR _7526_ (
    .Q(\datapath_1.regfile_1.regOut[5] [16]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_263_[16])
);

NAND2X1 _7106_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_118_)
);

FILL FILL_4__9773_ (
);

FILL FILL_4__9353_ (
);

FILL FILL_4__12639_ (
);

FILL FILL_2__13673_ (
);

FILL FILL_4__12219_ (
);

FILL FILL_2__13253_ (
);

FILL FILL_1__12246_ (
);

FILL FILL_0__9673_ (
);

FILL FILL_3__7350_ (
);

FILL FILL_0__9253_ (
);

INVX1 _11944_ (
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3004_)
);

FILL FILL_0__11659_ (
);

FILL FILL_0__11239_ (
);

AOI21X1 _11524_ (
    .A(_2216_),
    .B(_2176_),
    .C(_2520_),
    .Y(_2635_)
);

NOR2X1 _11104_ (
    .A(_2221_),
    .B(_2222_),
    .Y(_2223_)
);

FILL FILL_5__7696_ (
);

FILL FILL_4__16052_ (
);

FILL FILL_6__10573_ (
);

FILL FILL_3__15885_ (
);

FILL FILL_0__12600_ (
);

FILL FILL_3__15465_ (
);

FILL FILL_3__15045_ (
);

FILL SFILL39000x2050 (
);

FILL FILL_1__7688_ (
);

FILL FILL_6_BUFX2_insert710 (
);

FILL FILL_3__10180_ (
);

FILL FILL_2__14878_ (
);

FILL FILL_2__14458_ (
);

FILL FILL_2__14038_ (
);

FILL FILL_0__15492_ (
);

FILL FILL_6_BUFX2_insert715 (
);

FILL FILL_0__15072_ (
);

FILL SFILL13640x3050 (
);

FILL SFILL23720x53050 (
);

FILL FILL_3__8975_ (
);

NAND2X1 _12729_ (
    .A(IRWrite_bF$buf5),
    .B(memoryOutData[11]),
    .Y(_3512_)
);

FILL FILL_3__8135_ (
);

AOI22X1 _12309_ (
    .A(_2_[23]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3271_)
);

FILL FILL_1__14812_ (
);

FILL FILL_6__11778_ (
);

FILL FILL_4__12392_ (
);

FILL FILL_0__13805_ (
);

FILL FILL_2__6972_ (
);

FILL FILL_5__9422_ (
);

FILL FILL_3__11385_ (
);

FILL FILL_5__9002_ (
);

FILL FILL_4__6898_ (
);

FILL FILL_0__16277_ (
);

NAND3X1 _16142_ (
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf4),
    .Y(_6595_)
);

FILL FILL_2__10798_ (
);

FILL FILL_2__10378_ (
);

FILL FILL_5__11712_ (
);

FILL FILL_1__9414_ (
);

FILL SFILL8680x59050 (
);

FILL SFILL109560x76050 (
);

FILL FILL_4__10705_ (
);

FILL FILL_5__14184_ (
);

NAND2X1 _8484_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_813_)
);

NAND2X1 _8064_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_594_)
);

FILL FILL_4__13597_ (
);

FILL FILL_1__10312_ (
);

FILL FILL_2__7757_ (
);

FILL FILL_2__7337_ (
);

NAND2X1 _12482_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [14]),
    .Y(_3388_)
);

FILL FILL_0__12197_ (
);

NAND3X1 _12062_ (
    .A(_3090_),
    .B(_3091_),
    .C(_3092_),
    .Y(\datapath_1.mux_pcsrc.dout [18])
);

FILL FILL_5__12917_ (
);

FILL FILL_3__13951_ (
);

FILL FILL_3__13531_ (
);

FILL FILL_6__16396_ (
);

FILL FILL_3__13111_ (
);

FILL FILL_4__8624_ (
);

FILL FILL_4__8204_ (
);

FILL FILL_5_BUFX2_insert730 (
);

FILL FILL_5_BUFX2_insert731 (
);

FILL SFILL13720x51050 (
);

FILL FILL_5__15389_ (
);

FILL FILL_2__12524_ (
);

FILL FILL_5_BUFX2_insert732 (
);

FILL FILL_2__12104_ (
);

FILL FILL_5_BUFX2_insert733 (
);

DFFSR _9689_ (
    .Q(\datapath_1.regfile_1.regOut[22] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1368_[3])
);

FILL FILL_5_BUFX2_insert734 (
);

INVX1 _9269_ (
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_1214_)
);

FILL FILL_5_BUFX2_insert735 (
);

FILL FILL_5_BUFX2_insert736 (
);

FILL FILL_5_BUFX2_insert737 (
);

FILL FILL_1__11937_ (
);

FILL FILL_5_BUFX2_insert738 (
);

FILL FILL_5_BUFX2_insert739 (
);

FILL FILL_1__11517_ (
);

FILL SFILL53800x47050 (
);

FILL FILL_5__16330_ (
);

FILL FILL_6__9911_ (
);

FILL FILL_0__8524_ (
);

FILL FILL_0__8104_ (
);

FILL FILL_5__6967_ (
);

FILL FILL_4__15743_ (
);

FILL FILL_4__15323_ (
);

FILL SFILL13640x58050 (
);

AOI22X1 _13687_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [5]),
    .C(\datapath_1.regfile_1.regOut[31] [5]),
    .D(_3995__bF$buf0),
    .Y(_4194_)
);

FILL FILL_3__9093_ (
);

NAND2X1 _13267_ (
    .A(_3802_),
    .B(_3808_),
    .Y(_3809_)
);

FILL FILL_2__9903_ (
);

FILL FILL_3__14736_ (
);

FILL FILL_3__14316_ (
);

FILL FILL_1__15770_ (
);

FILL FILL_1__15350_ (
);

FILL FILL_1__6959_ (
);

FILL FILL_4__9409_ (
);

FILL SFILL8600x12050 (
);

FILL FILL_2__13729_ (
);

FILL FILL_2__13309_ (
);

FILL FILL_0__14763_ (
);

FILL FILL_0__14343_ (
);

FILL SFILL99560x80050 (
);

FILL FILL_2__7090_ (
);

FILL FILL_0__9729_ (
);

FILL FILL_3__7826_ (
);

FILL SFILL74280x38050 (
);

FILL FILL_5__12250_ (
);

OAI21X1 _6970_ (
    .A(_46_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_47_),
    .Y(_3_[22])
);

FILL FILL_2_BUFX2_insert860 (
);

FILL FILL_4__16108_ (
);

FILL FILL_2_BUFX2_insert861 (
);

FILL FILL_2_BUFX2_insert862 (
);

FILL FILL_2_BUFX2_insert863 (
);

FILL FILL_2_BUFX2_insert864 (
);

FILL FILL_4__11663_ (
);

FILL FILL_2_BUFX2_insert865 (
);

FILL FILL_4__11243_ (
);

FILL FILL_2_BUFX2_insert866 (
);

FILL FILL_2_BUFX2_insert867 (
);

FILL FILL_2_BUFX2_insert868 (
);

FILL SFILL13640x13050 (
);

FILL FILL_2_BUFX2_insert869 (
);

FILL FILL_1__16135_ (
);

FILL FILL_3__10656_ (
);

FILL FILL_1__11690_ (
);

FILL FILL_3__10236_ (
);

FILL FILL_1__11270_ (
);

FILL FILL_0__15968_ (
);

FILL FILL_0__15548_ (
);

NOR2X1 _15833_ (
    .A(_6290_),
    .B(_6293_),
    .Y(_6294_)
);

NOR2X1 _15413_ (
    .A(_5870_),
    .B(_5884_),
    .Y(_5885_)
);

FILL FILL_0__15128_ (
);

FILL FILL_0__10683_ (
);

FILL FILL_0__10263_ (
);

FILL FILL_6__14462_ (
);

FILL FILL_6__14042_ (
);

FILL FILL_5__13875_ (
);

FILL FILL_5__13455_ (
);

FILL FILL_5__13035_ (
);

NAND2X1 _7755_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_449_)
);

NAND2X1 _7335_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_230_)
);

FILL FILL_4__9162_ (
);

FILL FILL_4__12868_ (
);

FILL FILL_4__12448_ (
);

FILL FILL_4__12028_ (
);

FILL FILL_2__13482_ (
);

FILL FILL_1__12895_ (
);

FILL FILL_1__12475_ (
);

FILL SFILL99480x42050 (
);

FILL FILL_1__12055_ (
);

FILL FILL_0__11888_ (
);

FILL FILL_0__9482_ (
);

FILL FILL_0__11468_ (
);

NOR2X1 _11753_ (
    .A(_2848_),
    .B(_2840_),
    .Y(_2849_)
);

FILL SFILL3480x61050 (
);

INVX2 _11333_ (
    .A(_2451_),
    .Y(_2452_)
);

FILL FILL_0__11048_ (
);

FILL FILL_5__7085_ (
);

FILL FILL_4__16281_ (
);

FILL SFILL64200x79050 (
);

FILL FILL_3__15694_ (
);

FILL FILL_3__15274_ (
);

FILL FILL112120x56050 (
);

FILL FILL_1__7497_ (
);

FILL FILL_1__7077_ (
);

FILL FILL_2__14687_ (
);

FILL FILL_2__14267_ (
);

FILL FILL_5__15601_ (
);

NAND2X1 _9901_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1534_)
);

FILL FILL_1_BUFX2_insert880 (
);

FILL FILL_1_BUFX2_insert881 (
);

FILL FILL_3__8784_ (
);

FILL FILL_3__8364_ (
);

FILL FILL_1_BUFX2_insert882 (
);

NAND2X1 _12958_ (
    .A(vdd),
    .B(\datapath_1.rd2 [2]),
    .Y(_3624_)
);

DFFSR _12538_ (
    .Q(ALUOut[3]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3360_[3])
);

FILL FILL_1_BUFX2_insert883 (
);

INVX1 _12118_ (
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_3132_)
);

FILL FILL_1_BUFX2_insert884 (
);

FILL FILL_1_BUFX2_insert885 (
);

FILL FILL_1_BUFX2_insert886 (
);

FILL FILL_1__14621_ (
);

FILL FILL_1_BUFX2_insert887 (
);

FILL SFILL28840x60050 (
);

FILL FILL_1__14201_ (
);

FILL FILL_1_BUFX2_insert888 (
);

FILL FILL_1_BUFX2_insert889 (
);

FILL FILL_0__13614_ (
);

FILL FILL_3__16059_ (
);

FILL SFILL33800x43050 (
);

FILL FILL_5__9651_ (
);

FILL FILL_5__9231_ (
);

FILL FILL_3__11194_ (
);

FILL FILL112120x11050 (
);

OAI21X1 _16371_ (
    .A(_6800_),
    .B(gnd),
    .C(_6801_),
    .Y(_6769_[16])
);

FILL FILL_0__16086_ (
);

FILL FILL_2__10187_ (
);

FILL FILL_5__11941_ (
);

FILL FILL_1__9643_ (
);

FILL FILL_5__11521_ (
);

FILL FILL_1__9223_ (
);

FILL FILL_5__11101_ (
);

FILL FILL_3__9989_ (
);

FILL FILL_2__16413_ (
);

FILL FILL_3__9149_ (
);

FILL FILL_4__10934_ (
);

FILL FILL_4__10514_ (
);

FILL FILL_6__7994_ (
);

FILL FILL_1__15826_ (
);

DFFSR _8293_ (
    .Q(\datapath_1.regfile_1.regOut[11] [15]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_653_[15])
);

FILL FILL_1__15406_ (
);

FILL FILL_1__10961_ (
);

FILL FILL_1__10541_ (
);

FILL FILL112040x18050 (
);

FILL FILL_1__10121_ (
);

FILL FILL_0__14819_ (
);

FILL FILL_2__7986_ (
);

FILL FILL_2__7566_ (
);

BUFX2 BUFX2_insert550 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf57)
);

FILL FILL_3__12399_ (
);

BUFX2 BUFX2_insert551 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf56)
);

BUFX2 BUFX2_insert552 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf55)
);

BUFX2 BUFX2_insert553 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf54)
);

BUFX2 BUFX2_insert554 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf53)
);

BUFX2 BUFX2_insert555 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf52)
);

BUFX2 BUFX2_insert556 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf51)
);

BUFX2 BUFX2_insert557 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf50)
);

BUFX2 BUFX2_insert558 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf49)
);

BUFX2 BUFX2_insert559 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf48)
);

NAND3X1 _12291_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3257_)
);

FILL FILL_5__12726_ (
);

FILL FILL_3__13760_ (
);

FILL FILL_5__12306_ (
);

FILL FILL_3__13340_ (
);

FILL FILL_4__8853_ (
);

FILL SFILL79480x83050 (
);

FILL FILL_4__8013_ (
);

FILL FILL_4__11719_ (
);

FILL FILL_2__12753_ (
);

FILL FILL_5__15198_ (
);

FILL FILL_2__12333_ (
);

FILL FILL_6__8779_ (
);

INVX1 _9498_ (
    .A(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_1326_)
);

INVX1 _9078_ (
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_1171_)
);

FILL FILL_1__11746_ (
);

FILL FILL_1__11326_ (
);

FILL FILL_3__6850_ (
);

FILL FILL_0__8753_ (
);

FILL FILL_0__8333_ (
);

FILL FILL_0__10319_ (
);

DFFSR _10604_ (
    .Q(\datapath_1.regfile_1.regOut[29] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_1823_[22])
);

FILL FILL_0_BUFX2_insert70 (
);

FILL FILL_0_BUFX2_insert71 (
);

FILL FILL_6__14938_ (
);

FILL FILL_0_BUFX2_insert72 (
);

FILL FILL_4__15972_ (
);

FILL FILL_6__14518_ (
);

FILL FILL_0_BUFX2_insert73 (
);

FILL FILL_4__15552_ (
);

FILL FILL_0_BUFX2_insert74 (
);

FILL FILL_4__15132_ (
);

FILL FILL_0_BUFX2_insert75 (
);

FILL FILL_0_BUFX2_insert76 (
);

FILL FILL_0_BUFX2_insert77 (
);

INVX1 _13496_ (
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_4007_)
);

FILL SFILL103560x74050 (
);

FILL FILL_0_BUFX2_insert78 (
);

DFFSR _13076_ (
    .Q(_2_[29]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3620_[29])
);

FILL FILL_0_BUFX2_insert79 (
);

FILL FILL_3__14965_ (
);

FILL FILL_3__14545_ (
);

FILL FILL_3__14125_ (
);

FILL FILL_4_BUFX2_insert390 (
);

FILL FILL_4__9638_ (
);

FILL FILL_4_BUFX2_insert391 (
);

FILL FILL_4__9218_ (
);

FILL FILL_4_BUFX2_insert392 (
);

FILL FILL_4_BUFX2_insert393 (
);

FILL FILL_2__13958_ (
);

FILL FILL_0__14992_ (
);

FILL FILL_2__13538_ (
);

FILL FILL_4_BUFX2_insert394 (
);

FILL FILL_0__14572_ (
);

FILL FILL_2__13118_ (
);

FILL FILL_4_BUFX2_insert395 (
);

FILL FILL_4_BUFX2_insert396 (
);

FILL FILL_0__14152_ (
);

FILL FILL_4_BUFX2_insert397 (
);

FILL FILL_4_BUFX2_insert398 (
);

FILL FILL_4_BUFX2_insert399 (
);

FILL FILL_3__7635_ (
);

FILL FILL_0__9538_ (
);

FILL FILL_3__7215_ (
);

OAI21X1 _11809_ (
    .A(_2131_),
    .B(_2127_),
    .C(_2541_),
    .Y(_2900_)
);

FILL FILL_0__9118_ (
);

FILL FILL_4__16337_ (
);

FILL FILL_4__11892_ (
);

FILL FILL_4__11472_ (
);

FILL FILL_4__11052_ (
);

FILL FILL_1__16364_ (
);

FILL FILL_3__10885_ (
);

FILL FILL_5__8502_ (
);

FILL FILL_3__10045_ (
);

FILL FILL_0__15777_ (
);

FILL FILL_0__15357_ (
);

OAI22X1 _15642_ (
    .A(_4634_),
    .B(_5548__bF$buf3),
    .C(_5526__bF$buf0),
    .D(_4657_),
    .Y(_6108_)
);

INVX4 _15222_ (
    .A(_5501_),
    .Y(_5698_)
);

FILL FILL_0__10492_ (
);

FILL FILL_1__8914_ (
);

FILL FILL_5__13684_ (
);

FILL FILL_5__13264_ (
);

NAND2X1 _7984_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_561_)
);

NAND2X1 _7564_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_342_)
);

DFFSR _7144_ (
    .Q(\datapath_1.regfile_1.regOut[2] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_68_[18])
);

FILL FILL_4__9391_ (
);

FILL FILL_4__12257_ (
);

FILL SFILL48920x52050 (
);

FILL FILL_2__13291_ (
);

FILL FILL_2__6837_ (
);

FILL FILL_1__12284_ (
);

DFFSR _16427_ (
    .Q(\datapath_1.regfile_1.regOut[0] [10]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_6769_[10])
);

OAI22X1 _16007_ (
    .A(_5102_),
    .B(_5469__bF$buf1),
    .C(_5463__bF$buf3),
    .D(_5126_),
    .Y(_6463_)
);

OAI21X1 _11982_ (
    .A(_3028_),
    .B(IorD_bF$buf6),
    .C(_3029_),
    .Y(_1_[31])
);

FILL FILL_0__9291_ (
);

FILL FILL_0__11697_ (
);

FILL FILL_0__11277_ (
);

OAI21X1 _11562_ (
    .A(_2635_),
    .B(_2524_),
    .C(_2670_),
    .Y(_2671_)
);

AOI21X1 _11142_ (
    .A(_2216_),
    .B(_2176_),
    .C(_2260_),
    .Y(_2261_)
);

FILL FILL_3__12611_ (
);

FILL FILL_4__16090_ (
);

FILL FILL_4__7704_ (
);

FILL SFILL94920x1050 (
);

FILL FILL_6__10191_ (
);

FILL SFILL13720x46050 (
);

FILL FILL_5__14889_ (
);

FILL SFILL44120x37050 (
);

FILL FILL_5__14469_ (
);

FILL FILL_2__11604_ (
);

FILL FILL_5__14049_ (
);

FILL FILL_3__15083_ (
);

INVX1 _8769_ (
    .A(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_962_)
);

INVX1 _8349_ (
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_743_)
);

FILL FILL_2__14496_ (
);

FILL FILL_2__14076_ (
);

FILL FILL_5__15830_ (
);

FILL FILL_5__15410_ (
);

FILL FILL_0__7604_ (
);

DFFSR _9710_ (
    .Q(\datapath_1.regfile_1.regOut[22] [24]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1368_[24])
);

FILL FILL_1__13489_ (
);

FILL FILL_4__14823_ (
);

FILL FILL_4__14403_ (
);

FILL FILL_3__8593_ (
);

INVX1 _12767_ (
    .A(\datapath_1.PCJump [26]),
    .Y(_3537_)
);

NAND2X1 _12347_ (
    .A(MemToReg_bF$buf6),
    .B(\datapath_1.Data [1]),
    .Y(_3297_)
);

FILL FILL_3__13816_ (
);

FILL FILL_1__14850_ (
);

FILL FILL_5__8099_ (
);

FILL FILL_1__14430_ (
);

FILL FILL_1__14010_ (
);

FILL FILL_4__8909_ (
);

FILL FILL_0__13843_ (
);

FILL FILL_0__13423_ (
);

FILL FILL_3__16288_ (
);

FILL FILL_0__13003_ (
);

FILL FILL_5__9880_ (
);

FILL FILL_5__10389_ (
);

FILL FILL_5__9040_ (
);

NOR3X1 _16180_ (
    .A(_5515__bF$buf3),
    .B(_5300_),
    .C(_5521__bF$buf3),
    .Y(_6632_)
);

FILL FILL_3__6906_ (
);

FILL SFILL38920x50050 (
);

FILL FILL_1__9872_ (
);

FILL FILL_5__11750_ (
);

FILL FILL_5__11330_ (
);

FILL FILL_1__9032_ (
);

FILL FILL_4__15608_ (
);

FILL SFILL99160x61050 (
);

FILL FILL_2__16222_ (
);

FILL FILL_3__9798_ (
);

FILL FILL_3__9378_ (
);

FILL FILL_4__10743_ (
);

FILL FILL_4__10323_ (
);

FILL FILL_1__15635_ (
);

FILL FILL_1__15215_ (
);

FILL FILL_1__10770_ (
);

FILL FILL_0__14628_ (
);

INVX1 _14913_ (
    .A(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_5395_)
);

FILL FILL_0__14208_ (
);

FILL FILL_2__7375_ (
);

FILL FILL_5__12955_ (
);

FILL SFILL24200x71050 (
);

FILL FILL_5__12115_ (
);

FILL FILL_4__11948_ (
);

FILL FILL_4__8242_ (
);

FILL FILL_2__12982_ (
);

FILL FILL_4__11528_ (
);

FILL FILL_4__11108_ (
);

FILL FILL_2__12142_ (
);

FILL FILL112200x44050 (
);

FILL FILL_1__11975_ (
);

FILL SFILL99480x37050 (
);

FILL FILL_1__11555_ (
);

FILL FILL_1__11135_ (
);

FILL FILL_0__8982_ (
);

FILL FILL_0__10968_ (
);

FILL FILL_0__8142_ (
);

FILL FILL_0__10548_ (
);

NAND2X1 _10833_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_2013_)
);

FILL FILL_0__10128_ (
);

NAND2X1 _10413_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1794_)
);

FILL SFILL38840x12050 (
);

FILL FILL_4__15781_ (
);

FILL FILL_4__15361_ (
);

FILL FILL_2__9941_ (
);

FILL FILL_2__9521_ (
);

FILL FILL_3__14774_ (
);

FILL FILL_2__9101_ (
);

FILL FILL_3__14354_ (
);

FILL FILL_1__6997_ (
);

FILL FILL_4__9867_ (
);

FILL FILL_4__9027_ (
);

FILL FILL_2__13767_ (
);

FILL FILL_2__13347_ (
);

FILL FILL_0__14381_ (
);

FILL FILL_0__9767_ (
);

FILL FILL_3__7864_ (
);

FILL FILL_0__9347_ (
);

FILL FILL_3__7444_ (
);

OR2X2 _11618_ (
    .A(_2722_),
    .B(_2719_),
    .Y(_2723_)
);

FILL SFILL28840x55050 (
);

FILL FILL_1__13701_ (
);

FILL FILL_4__16146_ (
);

FILL FILL_6__10667_ (
);

FILL FILL_4__11281_ (
);

FILL FILL_3__15979_ (
);

FILL FILL_3__15559_ (
);

FILL FILL_3__15139_ (
);

FILL FILL_1__16173_ (
);

FILL SFILL33800x38050 (
);

FILL FILL_3__10694_ (
);

FILL FILL_5__8731_ (
);

FILL FILL_3__10274_ (
);

FILL FILL_5__8311_ (
);

NOR2X1 _15871_ (
    .A(_6329_),
    .B(_6330_),
    .Y(_6331_)
);

FILL FILL_0__15586_ (
);

INVX1 _15451_ (
    .A(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_5922_)
);

FILL FILL_0__15166_ (
);

AOI21X1 _15031_ (
    .A(_5492_),
    .B(_5510_),
    .C(_5509_),
    .Y(_5511_)
);

FILL FILL_1__8723_ (
);

FILL FILL_2__15913_ (
);

FILL FILL_3__8649_ (
);

FILL FILL_3__8229_ (
);

FILL FILL_5__13493_ (
);

FILL FILL_1__14906_ (
);

DFFSR _7793_ (
    .Q(\datapath_1.regfile_1.regOut[7] [27]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_393_[27])
);

INVX1 _7373_ (
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_255_)
);

FILL FILL_4__12486_ (
);

FILL SFILL28840x10050 (
);

FILL FILL_4__12066_ (
);

FILL FILL_3__11899_ (
);

FILL FILL_5__9936_ (
);

FILL FILL_5__9516_ (
);

FILL FILL_3__11479_ (
);

FILL FILL_3__11059_ (
);

FILL FILL_1__12093_ (
);

NOR2X1 _16236_ (
    .A(_6684_),
    .B(_6686_),
    .Y(_6687_)
);

AOI22X1 _11791_ (
    .A(_2141_),
    .B(_2481__bF$buf0),
    .C(_2341__bF$buf3),
    .D(_2142_),
    .Y(_2884_)
);

OAI21X1 _11371_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2118_),
    .C(_2487_),
    .Y(_2488_)
);

FILL FILL_0__11086_ (
);

FILL FILL_1__9928_ (
);

FILL FILL_5__11806_ (
);

FILL FILL_1__9508_ (
);

FILL FILL_3__12840_ (
);

FILL FILL_3__12420_ (
);

FILL FILL_3__12000_ (
);

FILL FILL_4__7933_ (
);

FILL FILL_5__14698_ (
);

FILL FILL_2__11833_ (
);

FILL FILL_5__14278_ (
);

FILL FILL_2__11413_ (
);

INVX1 _8998_ (
    .A(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_1074_)
);

FILL FILL_6__7859_ (
);

INVX1 _8578_ (
    .A(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_855_)
);

DFFSR _8158_ (
    .Q(\datapath_1.regfile_1.regOut[10] [8]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_588_[8])
);

FILL FILL_1__10826_ (
);

FILL FILL_1__10406_ (
);

FILL SFILL18840x53050 (
);

FILL FILL_0__7833_ (
);

FILL FILL_1__13298_ (
);

FILL SFILL58920x49050 (
);

FILL FILL_4__14632_ (
);

FILL FILL_4__14212_ (
);

INVX1 _12996_ (
    .A(_2_[15]),
    .Y(_3649_)
);

INVX1 _12576_ (
    .A(\datapath_1.Data [3]),
    .Y(_3430_)
);

OAI21X1 _12156_ (
    .A(_3156_),
    .B(ALUSrcA_bF$buf3),
    .C(_3157_),
    .Y(\datapath_1.alu_1.ALUInA [13])
);

FILL FILL_3__13625_ (
);

FILL FILL_4__8718_ (
);

FILL FILL_2__12618_ (
);

FILL FILL_0__13652_ (
);

FILL FILL_0__13232_ (
);

FILL FILL_3__16097_ (
);

FILL SFILL48600x71050 (
);

FILL FILL_5__16004_ (
);

FILL FILL_0__8618_ (
);

FILL FILL_1__9681_ (
);

FILL FILL_1__9261_ (
);

FILL FILL_4__15837_ (
);

FILL FILL_4__15417_ (
);

FILL FILL_2__16451_ (
);

FILL FILL_2__16031_ (
);

FILL FILL_4__10972_ (
);

FILL SFILL109640x59050 (
);

FILL FILL_4__10552_ (
);

FILL FILL_4__10132_ (
);

FILL FILL_1__15864_ (
);

FILL FILL_1__15444_ (
);

FILL FILL_1__15024_ (
);

FILL FILL_0__14857_ (
);

NOR2X1 _14722_ (
    .A(_5207_),
    .B(_5204_),
    .Y(_5208_)
);

FILL FILL_0__14437_ (
);

FILL FILL_0__14017_ (
);

INVX1 _14302_ (
    .A(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_4797_)
);

BUFX2 BUFX2_insert930 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf4 )
);

FILL FILL_2__7184_ (
);

BUFX2 BUFX2_insert931 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf3 )
);

BUFX2 BUFX2_insert932 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf2 )
);

BUFX2 BUFX2_insert933 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf1 )
);

FILL FILL_6__13771_ (
);

BUFX2 BUFX2_insert934 (
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf0 )
);

BUFX2 BUFX2_insert935 (
    .A(_3935_),
    .Y(_3935__bF$buf4)
);

BUFX2 BUFX2_insert936 (
    .A(_3935_),
    .Y(_3935__bF$buf3)
);

BUFX2 BUFX2_insert937 (
    .A(_3935_),
    .Y(_3935__bF$buf2)
);

BUFX2 BUFX2_insert938 (
    .A(_3935_),
    .Y(_3935__bF$buf1)
);

BUFX2 BUFX2_insert939 (
    .A(_3935_),
    .Y(_3935__bF$buf0)
);

FILL FILL_5__12764_ (
);

FILL FILL_5__12344_ (
);

FILL SFILL69080x62050 (
);

FILL FILL_4__8891_ (
);

FILL FILL_4__8471_ (
);

FILL FILL_4__11757_ (
);

FILL SFILL48920x47050 (
);

FILL FILL_4__11337_ (
);

FILL FILL_2__12371_ (
);

FILL FILL_6__8397_ (
);

FILL FILL_1__16229_ (
);

FILL FILL_1__11784_ (
);

FILL FILL_1__11364_ (
);

NAND3X1 _15927_ (
    .A(_6382_),
    .B(_6385_),
    .C(_6377_),
    .Y(_6386_)
);

AOI21X1 _15507_ (
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .B(_5649_),
    .C(_5975_),
    .Y(_5976_)
);

FILL FILL_0__10777_ (
);

FILL FILL_2__8389_ (
);

FILL FILL_0__8371_ (
);

NAND2X1 _10642_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1906_)
);

DFFSR _10222_ (
    .Q(\datapath_1.regfile_1.regOut[26] [24]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_1628_[24])
);

FILL FILL_4__15590_ (
);

FILL FILL_4__15170_ (
);

FILL FILL_5__13969_ (
);

FILL FILL_2__9750_ (
);

FILL FILL_5__13549_ (
);

FILL FILL_3__14583_ (
);

FILL FILL_5__13129_ (
);

FILL FILL_3__14163_ (
);

INVX1 _7849_ (
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_491_)
);

FILL SFILL69000x60050 (
);

INVX1 _7429_ (
    .A(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_272_)
);

DFFSR _7009_ (
    .Q(\datapath_1.regfile_1.regOut[1] [11]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_3_[11])
);

FILL FILL_4_BUFX2_insert770 (
);

FILL FILL_4__9676_ (
);

FILL FILL_4_BUFX2_insert771 (
);

FILL FILL_4__9256_ (
);

FILL FILL_4_BUFX2_insert772 (
);

FILL FILL_4_BUFX2_insert773 (
);

FILL FILL_2__13996_ (
);

FILL FILL_4_BUFX2_insert774 (
);

FILL FILL_2__13576_ (
);

FILL FILL_2__13156_ (
);

FILL FILL_4_BUFX2_insert775 (
);

FILL FILL_0__14190_ (
);

FILL FILL_4_BUFX2_insert776 (
);

FILL FILL_4_BUFX2_insert777 (
);

FILL FILL_5__14910_ (
);

FILL FILL_4_BUFX2_insert778 (
);

FILL FILL_4_BUFX2_insert779 (
);

FILL FILL_1__12989_ (
);

FILL FILL_1__12569_ (
);

FILL FILL_1__12149_ (
);

FILL FILL_4__13903_ (
);

FILL FILL_0__9996_ (
);

FILL FILL_3__7673_ (
);

FILL FILL_0__9156_ (
);

FILL FILL_3__7253_ (
);

NOR2X1 _11847_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2935_)
);

AOI21X1 _11427_ (
    .A(_2542_),
    .B(_2130_),
    .C(_2491_),
    .Y(_2543_)
);

INVX1 _11007_ (
    .A(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2126_)
);

FILL FILL_5__7599_ (
);

FILL FILL_1__13930_ (
);

FILL FILL_5__7179_ (
);

FILL FILL_4__16375_ (
);

FILL FILL_1__13510_ (
);

FILL FILL_4__11090_ (
);

FILL FILL_3__15788_ (
);

FILL FILL_3__15368_ (
);

FILL FILL_0__12503_ (
);

FILL FILL_5__8960_ (
);

FILL FILL_5__8120_ (
);

FILL SFILL38120x62050 (
);

FILL SFILL59080x60050 (
);

FILL FILL_0__15395_ (
);

NAND3X1 _15680_ (
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6145_)
);

AOI22X1 _15260_ (
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_5735_)
);

FILL FILL_5__10830_ (
);

FILL FILL_1__8952_ (
);

FILL FILL_1__8532_ (
);

FILL FILL_5__10410_ (
);

FILL FILL_1__8112_ (
);

FILL FILL_2__15722_ (
);

FILL FILL_2__15302_ (
);

FILL FILL_3__8878_ (
);

FILL FILL_3__8458_ (
);

FILL SFILL59400x72050 (
);

FILL FILL_6__6883_ (
);

FILL FILL_1__14715_ (
);

INVX1 _7182_ (
    .A(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_148_)
);

FILL FILL_4__12295_ (
);

FILL FILL_0__13708_ (
);

FILL FILL_2__6875_ (
);

FILL FILL_5__9745_ (
);

FILL FILL_3__11288_ (
);

FILL SFILL99560x25050 (
);

NOR3X1 _16045_ (
    .A(_6500_),
    .B(_6478_),
    .C(_6489_),
    .Y(_6501_)
);

INVX1 _11180_ (
    .A(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2299_)
);

FILL FILL_1__9737_ (
);

FILL FILL_5__11615_ (
);

FILL FILL_4__7742_ (
);

FILL FILL_3_BUFX2_insert790 (
);

FILL FILL_4__7322_ (
);

FILL FILL_3_BUFX2_insert791 (
);

FILL FILL_3_BUFX2_insert792 (
);

FILL FILL_3_BUFX2_insert793 (
);

FILL FILL_2__11642_ (
);

FILL FILL_3_BUFX2_insert794 (
);

FILL FILL_2__11222_ (
);

FILL FILL_5__14087_ (
);

FILL FILL_3_BUFX2_insert795 (
);

FILL FILL_3_BUFX2_insert796 (
);

OAI21X1 _8387_ (
    .A(_767_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_768_),
    .Y(_718_[25])
);

FILL FILL_3_BUFX2_insert797 (
);

FILL FILL_3_BUFX2_insert798 (
);

FILL FILL_3_BUFX2_insert799 (
);

FILL FILL_1__10635_ (
);

FILL FILL_0__7222_ (
);

FILL SFILL73960x83050 (
);

FILL FILL_6__13827_ (
);

FILL FILL_4__14861_ (
);

FILL FILL_4__14441_ (
);

FILL FILL_4__14021_ (
);

FILL SFILL43960x2050 (
);

INVX1 _12385_ (
    .A(ALUOut[14]),
    .Y(_3322_)
);

FILL FILL_3__13854_ (
);

FILL FILL_2__8601_ (
);

FILL FILL_3__13434_ (
);

FILL FILL_3__13014_ (
);

FILL FILL_4__8527_ (
);

FILL FILL_4__8107_ (
);

FILL FILL_2__12847_ (
);

FILL SFILL89160x54050 (
);

FILL FILL_0__13881_ (
);

FILL FILL_2__12427_ (
);

FILL FILL_0__13461_ (
);

FILL FILL_2__12007_ (
);

FILL FILL_0__13041_ (
);

FILL FILL_0__8847_ (
);

FILL FILL_5__16233_ (
);

FILL FILL_3__6944_ (
);

FILL FILL_0__8007_ (
);

FILL FILL_1__9490_ (
);

FILL FILL_4__15646_ (
);

FILL FILL_4__15226_ (
);

FILL FILL_2__16260_ (
);

FILL SFILL73480x76050 (
);

FILL FILL_4__10781_ (
);

FILL FILL_4__10361_ (
);

FILL FILL_2__9806_ (
);

FILL FILL_4_BUFX2_insert20 (
);

FILL FILL_3__14639_ (
);

FILL FILL_4_BUFX2_insert21 (
);

FILL FILL_1__15673_ (
);

FILL FILL_3__14219_ (
);

FILL FILL_4_BUFX2_insert22 (
);

FILL FILL_1__15253_ (
);

FILL FILL_4_BUFX2_insert23 (
);

FILL FILL_4_BUFX2_insert24 (
);

FILL FILL_5__7811_ (
);

FILL FILL_4_BUFX2_insert25 (
);

FILL FILL_4_BUFX2_insert26 (
);

FILL FILL_4_BUFX2_insert27 (
);

FILL FILL_4_BUFX2_insert28 (
);

FILL FILL_4_BUFX2_insert29 (
);

NAND3X1 _14951_ (
    .A(_5423_),
    .B(_5424_),
    .C(_5431_),
    .Y(_5432_)
);

FILL FILL_0__14666_ (
);

FILL FILL_0__14246_ (
);

INVX1 _14531_ (
    .A(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_5021_)
);

NOR2X1 _14111_ (
    .A(_4609_),
    .B(_3935__bF$buf0),
    .Y(_4610_)
);

FILL FILL_1__7803_ (
);

FILL FILL_3__7729_ (
);

FILL FILL_3__7309_ (
);

FILL FILL_5__12993_ (
);

FILL FILL_5__12573_ (
);

FILL FILL_5__12153_ (
);

BUFX2 _6873_ (
    .A(_2_[3]),
    .Y(memoryWriteData[3])
);

FILL FILL_4__11986_ (
);

FILL FILL_4__11566_ (
);

FILL SFILL94360x72050 (
);

FILL FILL_4__11146_ (
);

FILL FILL_2__12180_ (
);

FILL FILL_1__16038_ (
);

FILL FILL_3__10979_ (
);

FILL FILL_3__10559_ (
);

FILL FILL_1__11593_ (
);

FILL FILL_3__10139_ (
);

FILL FILL_1__11173_ (
);

NAND3X1 _15736_ (
    .A(_6197_),
    .B(_6198_),
    .C(_6196_),
    .Y(_6199_)
);

INVX1 _15316_ (
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_5790_)
);

NAND2X1 _10871_ (
    .A(\aluControl_1.inst [5]),
    .B(_2018_),
    .Y(_2019_)
);

FILL FILL_2__8198_ (
);

FILL SFILL79160x52050 (
);

FILL FILL_0__10166_ (
);

INVX1 _10451_ (
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_1819_)
);

INVX1 _10031_ (
    .A(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_1600_)
);

FILL FILL_3__11920_ (
);

BUFX2 BUFX2_insert80 (
    .A(_5495_),
    .Y(_5495__bF$buf0)
);

BUFX2 BUFX2_insert81 (
    .A(_3884_),
    .Y(_3884__bF$buf3)
);

FILL FILL_6__14365_ (
);

FILL FILL_3__11500_ (
);

BUFX2 BUFX2_insert82 (
    .A(_3884_),
    .Y(_3884__bF$buf2)
);

BUFX2 BUFX2_insert83 (
    .A(_3884_),
    .Y(_3884__bF$buf1)
);

BUFX2 BUFX2_insert84 (
    .A(_3884_),
    .Y(_3884__bF$buf0)
);

BUFX2 BUFX2_insert85 (
    .A(_3902_),
    .Y(_3902__bF$buf3)
);

BUFX2 BUFX2_insert86 (
    .A(_3902_),
    .Y(_3902__bF$buf2)
);

FILL FILL_2__10913_ (
);

FILL FILL_5__13778_ (
);

BUFX2 BUFX2_insert87 (
    .A(_3902_),
    .Y(_3902__bF$buf1)
);

FILL FILL_5__13358_ (
);

BUFX2 BUFX2_insert88 (
    .A(_3902_),
    .Y(_3902__bF$buf0)
);

BUFX2 BUFX2_insert89 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf4 )
);

FILL FILL_3__14392_ (
);

DFFSR _7658_ (
    .Q(\datapath_1.regfile_1.regOut[6] [20]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_328_[20])
);

OAI21X1 _7238_ (
    .A(_184_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_185_),
    .Y(_133_[26])
);

FILL FILL_4__9485_ (
);

FILL FILL_2__13385_ (
);

FILL FILL_0__6913_ (
);

FILL FILL_1__12378_ (
);

FILL FILL_4__13712_ (
);

FILL FILL_3__7482_ (
);

FILL FILL_0__9385_ (
);

FILL FILL_3__7062_ (
);

NOR2X1 _11656_ (
    .A(_2752_),
    .B(_2758_),
    .Y(_2759_)
);

NOR2X1 _11236_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2355_)
);

FILL FILL_3__12705_ (
);

FILL FILL_4__16184_ (
);

FILL FILL_0__12732_ (
);

FILL FILL_3__15597_ (
);

FILL FILL_3__15177_ (
);

FILL FILL_0__12312_ (
);

FILL SFILL38920x8050 (
);

FILL FILL_5__15924_ (
);

FILL FILL_5__15504_ (
);

FILL SFILL84360x70050 (
);

OAI21X1 _9804_ (
    .A(_1488_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1489_),
    .Y(_1433_[28])
);

FILL FILL_1__8761_ (
);

FILL FILL_1__8341_ (
);

FILL FILL_4__14917_ (
);

FILL FILL_2__15951_ (
);

FILL FILL_2__15531_ (
);

FILL FILL_2__15111_ (
);

FILL FILL_3__8267_ (
);

FILL FILL_1__14944_ (
);

FILL FILL_1__14524_ (
);

FILL FILL_1__14104_ (
);

FILL FILL_0__13937_ (
);

INVX1 _13802_ (
    .A(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_4307_)
);

FILL FILL_0__13517_ (
);

FILL FILL_5__9974_ (
);

FILL FILL_5__9554_ (
);

FILL FILL_5__9134_ (
);

FILL FILL_3__11097_ (
);

INVX1 _16274_ (
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_6724_)
);

FILL FILL_5__11844_ (
);

FILL FILL_1__9546_ (
);

FILL FILL_5__11424_ (
);

FILL FILL_1__9126_ (
);

FILL FILL_5__11004_ (
);

FILL SFILL69080x57050 (
);

FILL FILL_4__7971_ (
);

FILL FILL_2__16316_ (
);

FILL FILL_4__7551_ (
);

FILL FILL_4__10837_ (
);

FILL FILL_2__11871_ (
);

FILL FILL_4__10417_ (
);

FILL FILL_2__11451_ (
);

FILL FILL_2__11031_ (
);

FILL FILL_6__7477_ (
);

FILL FILL_1__15729_ (
);

OAI21X1 _8196_ (
    .A(_660_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .C(_661_),
    .Y(_653_[4])
);

FILL FILL_1__15309_ (
);

FILL FILL_1__10444_ (
);

FILL FILL_1__10024_ (
);

FILL FILL_0__7871_ (
);

FILL FILL_2__7889_ (
);

FILL FILL_0__7451_ (
);

FILL FILL_2__7469_ (
);

FILL FILL_2__7049_ (
);

FILL FILL_0__7031_ (
);

FILL SFILL114520x51050 (
);

FILL FILL_4__14670_ (
);

FILL FILL_4__14250_ (
);

FILL SFILL3720x70050 (
);

NAND2X1 _12194_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.a [26]),
    .Y(_3183_)
);

FILL FILL_5__12629_ (
);

FILL FILL_2__8830_ (
);

FILL FILL_3__13663_ (
);

FILL FILL_5__12209_ (
);

FILL FILL_3__13243_ (
);

INVX1 _6929_ (
    .A(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_20_)
);

FILL FILL_4__8756_ (
);

FILL FILL_4__8336_ (
);

FILL FILL_2__12656_ (
);

FILL FILL_2__12236_ (
);

FILL FILL_0__13690_ (
);

FILL FILL_0__13270_ (
);

FILL FILL_1__11649_ (
);

FILL FILL_1__11229_ (
);

FILL SFILL3640x77050 (
);

FILL FILL_5__16042_ (
);

FILL FILL_0__8656_ (
);

NOR2X1 _10927_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2057_),
    .Y(ALUSrcB[0])
);

FILL FILL_0__8236_ (
);

INVX1 _10507_ (
    .A(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_1836_)
);

FILL FILL_4__15875_ (
);

FILL FILL_4__15455_ (
);

FILL FILL_4__15035_ (
);

OAI22X1 _13399_ (
    .A(_3907_),
    .B(_3910_),
    .C(_3909_),
    .D(_3908_),
    .Y(_3911_)
);

FILL FILL_4__10170_ (
);

FILL FILL_2__9615_ (
);

FILL FILL_3__14868_ (
);

FILL FILL_3__14448_ (
);

FILL FILL_3__14028_ (
);

FILL FILL_1__15482_ (
);

FILL FILL_1__15062_ (
);

FILL FILL_5__7620_ (
);

FILL FILL_5__7200_ (
);

FILL SFILL59080x55050 (
);

FILL FILL_0__14895_ (
);

FILL FILL_0__14475_ (
);

OAI22X1 _14760_ (
    .A(_5244_),
    .B(_3972__bF$buf3),
    .C(_3920_),
    .D(_5243_),
    .Y(_5245_)
);

FILL FILL_0__14055_ (
);

NOR2X1 _14340_ (
    .A(_4833_),
    .B(_4830_),
    .Y(_4834_)
);

FILL SFILL59880x38050 (
);

FILL FILL_1__7612_ (
);

FILL FILL_2__14802_ (
);

FILL FILL_3__7958_ (
);

FILL FILL_3__7118_ (
);

FILL SFILL3640x32050 (
);

FILL FILL_5__12382_ (
);

FILL FILL_4__11795_ (
);

FILL FILL_4__11375_ (
);

FILL FILL_1__16267_ (
);

FILL FILL_3__10788_ (
);

FILL FILL_5__8825_ (
);

FILL FILL_3__10368_ (
);

FILL FILL_5__8405_ (
);

FILL SFILL49080x1050 (
);

FILL SFILL59000x53050 (
);

NOR2X1 _15965_ (
    .A(_6422_),
    .B(_6419_),
    .Y(_6423_)
);

FILL FILL_6__11702_ (
);

AOI21X1 _15545_ (
    .A(\datapath_1.regfile_1.regOut[29] [12]),
    .B(_5486_),
    .C(_6012_),
    .Y(_6013_)
);

NAND2X1 _15125_ (
    .A(_5598_),
    .B(_5603_),
    .Y(_5604_)
);

FILL SFILL59080x10050 (
);

FILL FILL_0__10395_ (
);

INVX1 _10680_ (
    .A(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_1931_)
);

INVX1 _10260_ (
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_1712_)
);

FILL SFILL104440x56050 (
);

FILL FILL_0__16201_ (
);

FILL FILL_5__13587_ (
);

FILL FILL_2__10302_ (
);

FILL FILL_5__13167_ (
);

OAI21X1 _7887_ (
    .A(_515_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_516_),
    .Y(_458_[29])
);

OAI21X1 _7467_ (
    .A(_296_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .C(_297_),
    .Y(_263_[17])
);

OAI21X1 _7047_ (
    .A(_77_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_78_),
    .Y(_68_[5])
);

FILL FILL_4__9294_ (
);

FILL SFILL33880x82050 (
);

FILL FILL_1__12187_ (
);

FILL FILL_4__13941_ (
);

FILL FILL_4__13521_ (
);

FILL FILL_4__13101_ (
);

NAND2X1 _11885_ (
    .A(RegDst),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_2967_)
);

FILL FILL_3__7291_ (
);

FILL SFILL49080x53050 (
);

OAI21X1 _11465_ (
    .A(_2579_),
    .B(_2313_),
    .C(_2439_),
    .Y(_2580_)
);

XOR2X1 _11045_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2164_)
);

FILL FILL_3__12514_ (
);

FILL FILL_4__7607_ (
);

FILL FILL_2__11927_ (
);

FILL FILL_0__12961_ (
);

FILL FILL_2__11507_ (
);

FILL FILL_0__12121_ (
);

FILL FILL_2__14399_ (
);

FILL SFILL28520x24050 (
);

FILL FILL_5__15733_ (
);

FILL FILL_5__15313_ (
);

FILL FILL_0__7927_ (
);

FILL FILL_0__7507_ (
);

OAI21X1 _9613_ (
    .A(_1381_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1382_),
    .Y(_1368_[7])
);

FILL FILL_1__8990_ (
);

FILL FILL_1__8570_ (
);

FILL FILL_4__14726_ (
);

FILL FILL_2__15760_ (
);

FILL FILL_4__14306_ (
);

FILL FILL_2__15340_ (
);

FILL FILL_3__8496_ (
);

FILL FILL_3__8076_ (
);

FILL FILL_3__13719_ (
);

FILL FILL_1__14753_ (
);

FILL FILL_1__14333_ (
);

FILL SFILL14200x59050 (
);

FILL SFILL94440x60050 (
);

FILL FILL_0__13746_ (
);

FILL FILL_0__13326_ (
);

NOR2X1 _13611_ (
    .A(_4104_),
    .B(_4119_),
    .Y(_4120_)
);

FILL FILL_5__9783_ (
);

FILL FILL_5__9363_ (
);

FILL FILL_6__12660_ (
);

OAI22X1 _16083_ (
    .A(_5463__bF$buf2),
    .B(_5168_),
    .C(_5171_),
    .D(_5504__bF$buf2),
    .Y(_6538_)
);

FILL FILL_1__9775_ (
);

FILL FILL_5__11653_ (
);

FILL FILL_1__9355_ (
);

FILL FILL_5__11233_ (
);

FILL FILL_2__16125_ (
);

FILL FILL_4__7360_ (
);

FILL SFILL94360x67050 (
);

FILL FILL_4__10646_ (
);

FILL FILL_2__11680_ (
);

FILL FILL_2__11260_ (
);

FILL FILL_1__15958_ (
);

FILL FILL_6__7286_ (
);

FILL FILL_1__15538_ (
);

FILL FILL_1__15118_ (
);

FILL FILL_2_BUFX2_insert100 (
);

FILL FILL_1__10673_ (
);

FILL FILL_1__10253_ (
);

FILL FILL_2_BUFX2_insert101 (
);

FILL FILL_2_BUFX2_insert102 (
);

INVX1 _14816_ (
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_5300_)
);

FILL FILL_2_BUFX2_insert103 (
);

FILL FILL_2_BUFX2_insert104 (
);

FILL FILL_2_BUFX2_insert105 (
);

FILL FILL_0__7680_ (
);

FILL FILL_2_BUFX2_insert106 (
);

FILL FILL_2__7698_ (
);

FILL FILL_2_BUFX2_insert107 (
);

FILL FILL_2_BUFX2_insert108 (
);

FILL FILL_2_BUFX2_insert109 (
);

FILL FILL_5__12858_ (
);

FILL SFILL18760x3050 (
);

FILL FILL_5__12438_ (
);

FILL FILL_3__13892_ (
);

FILL FILL_5__12018_ (
);

FILL FILL_3__13472_ (
);

FILL FILL_4__8985_ (
);

FILL SFILL18680x8050 (
);

FILL FILL_4__8145_ (
);

FILL FILL_2__12885_ (
);

FILL FILL_2__12465_ (
);

FILL SFILL80120x50050 (
);

FILL FILL111800x51050 (
);

FILL FILL_2__12045_ (
);

FILL SFILL94360x22050 (
);

FILL FILL_1__11878_ (
);

FILL FILL_1__11458_ (
);

FILL FILL_1__11038_ (
);

FILL FILL_0__8885_ (
);

FILL FILL_3__6982_ (
);

FILL FILL_5__16271_ (
);

FILL FILL_0__8465_ (
);

DFFSR _10736_ (
    .Q(\datapath_1.regfile_1.regOut[30] [26]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_1888_[26])
);

OAI21X1 _10316_ (
    .A(_1748_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1749_),
    .Y(_1693_[28])
);

FILL FILL_6__9012_ (
);

FILL FILL_4__15684_ (
);

FILL FILL_4__15264_ (
);

FILL SFILL4040x62050 (
);

FILL FILL_2__9424_ (
);

FILL FILL_0__11812_ (
);

FILL FILL_3__14677_ (
);

FILL FILL_3__14257_ (
);

FILL FILL_2__9004_ (
);

FILL FILL_1__15291_ (
);

FILL FILL_0__14284_ (
);

FILL SFILL84360x65050 (
);

FILL FILL_1__7841_ (
);

FILL FILL_1__7421_ (
);

FILL FILL_2__14611_ (
);

FILL FILL_3__7347_ (
);

FILL FILL_5__12191_ (
);

FILL FILL_1__13604_ (
);

FILL FILL_4__16049_ (
);

FILL FILL_4__11184_ (
);

FILL SFILL29400x61050 (
);

FILL FILL_1__16076_ (
);

FILL FILL_5__8634_ (
);

FILL FILL_3__10177_ (
);

FILL FILL_5__8214_ (
);

FILL FILL_6_BUFX2_insert684 (
);

OAI22X1 _15774_ (
    .A(_5478__bF$buf2),
    .B(_6235_),
    .C(_5527__bF$buf3),
    .D(_4812_),
    .Y(_6236_)
);

FILL FILL_0__15489_ (
);

NAND3X1 _15354_ (
    .A(_5822_),
    .B(_5823_),
    .C(_5826_),
    .Y(_5827_)
);

FILL FILL_0__15069_ (
);

FILL FILL_3__16403_ (
);

FILL FILL_6_BUFX2_insert689 (
);

FILL FILL_5__10924_ (
);

FILL FILL_5__10504_ (
);

FILL FILL_1__8626_ (
);

FILL FILL_1__8206_ (
);

FILL SFILL84360x20050 (
);

FILL FILL_2__15816_ (
);

FILL FILL_0__16010_ (
);

FILL FILL_2__10951_ (
);

FILL FILL_2__10531_ (
);

FILL FILL_5__13396_ (
);

FILL FILL_2__10111_ (
);

OAI21X1 _7696_ (
    .A(_408_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .C(_409_),
    .Y(_393_[8])
);

FILL FILL_1__14809_ (
);

DFFSR _7276_ (
    .Q(\datapath_1.regfile_1.regOut[3] [22]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_133_[22])
);

FILL FILL_4__12389_ (
);

FILL FILL_3__9913_ (
);

FILL FILL_0__6951_ (
);

FILL FILL_2__6969_ (
);

FILL FILL_5__9419_ (
);

FILL FILL_4__13750_ (
);

FILL FILL_4__13330_ (
);

NAND3X1 _16139_ (
    .A(_6585_),
    .B(_6586_),
    .C(_6591_),
    .Y(_6592_)
);

FILL SFILL3720x65050 (
);

OAI21X1 _11694_ (
    .A(_2185_),
    .B(_2620_),
    .C(_2793_),
    .Y(_2794_)
);

NAND2X1 _11274_ (
    .A(_2391_),
    .B(_2202_),
    .Y(_2393_)
);

FILL FILL_5__11709_ (
);

FILL FILL_3__12743_ (
);

FILL SFILL43960x72050 (
);

FILL FILL_6__15188_ (
);

FILL FILL_3__12323_ (
);

FILL FILL_4__7836_ (
);

FILL FILL_4__7416_ (
);

FILL FILL_2__11736_ (
);

FILL FILL_0__12770_ (
);

FILL FILL_2__11316_ (
);

FILL FILL_0__12350_ (
);

FILL FILL_1__10309_ (
);

FILL FILL_5__15962_ (
);

FILL FILL_5__15542_ (
);

FILL FILL_0__7736_ (
);

FILL FILL_5__15122_ (
);

DFFSR _9842_ (
    .Q(\datapath_1.regfile_1.regOut[23] [28]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1433_[28])
);

FILL FILL_0__7316_ (
);

NAND2X1 _9422_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1296_)
);

FILL SFILL43880x79050 (
);

NAND2X1 _9002_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1077_)
);

FILL FILL_4__14955_ (
);

FILL FILL_4__14535_ (
);

FILL FILL_4__14115_ (
);

NAND2X1 _12899_ (
    .A(vdd),
    .B(\datapath_1.rd1 [25]),
    .Y(_3605_)
);

NAND2X1 _12479_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [13]),
    .Y(_3386_)
);

NAND3X1 _12059_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[18]),
    .C(_3032__bF$buf2),
    .Y(_3090_)
);

FILL FILL_3__13948_ (
);

FILL SFILL3720x20050 (
);

FILL FILL_1__14982_ (
);

FILL FILL_3__13528_ (
);

FILL FILL_1__14562_ (
);

FILL FILL_3__13108_ (
);

FILL FILL_1__14142_ (
);

FILL FILL112280x83050 (
);

FILL FILL_0__13975_ (
);

AOI21X1 _13840_ (
    .A(_4321_),
    .B(_4344_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [7])
);

FILL FILL_0__13555_ (
);

OAI22X1 _13420_ (
    .A(_3928_),
    .B(_3930__bF$buf0),
    .C(_3931__bF$buf3),
    .D(_3929_),
    .Y(_3932_)
);

FILL FILL_0__13135_ (
);

NAND2X1 _13000_ (
    .A(vdd),
    .B(\datapath_1.rd2 [16]),
    .Y(_3652_)
);

FILL FILL_5__9592_ (
);

FILL FILL_5__9172_ (
);

FILL FILL_5__16327_ (
);

FILL SFILL3640x27050 (
);

FILL FILL_5__11882_ (
);

FILL FILL_5__11462_ (
);

FILL FILL_1__9164_ (
);

FILL FILL_5__11042_ (
);

FILL SFILL104520x44050 (
);

FILL FILL_2__16354_ (
);

FILL SFILL43880x34050 (
);

FILL FILL_4__10875_ (
);

FILL FILL_4__10035_ (
);

FILL FILL_1__15767_ (
);

FILL FILL_1__15347_ (
);

FILL SFILL59000x48050 (
);

FILL FILL_1__10062_ (
);

FILL SFILL108840x52050 (
);

NOR2X1 _14625_ (
    .A(_5109_),
    .B(_5112_),
    .Y(_5113_)
);

NAND3X1 _14205_ (
    .A(_4693_),
    .B(_4694_),
    .C(_4701_),
    .Y(_4702_)
);

FILL FILL_2__7087_ (
);

FILL FILL_6__13674_ (
);

FILL FILL_0__15701_ (
);

FILL FILL_5__12247_ (
);

FILL FILL_3__13281_ (
);

OAI21X1 _6967_ (
    .A(_44_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .C(_45_),
    .Y(_3_[21])
);

FILL SFILL33880x77050 (
);

FILL FILL_4__8374_ (
);

FILL FILL_2__12274_ (
);

FILL FILL_1__11687_ (
);

FILL FILL_1__11267_ (
);

FILL FILL_4__12601_ (
);

FILL FILL_0__8694_ (
);

FILL FILL_5__16080_ (
);

FILL SFILL33480x63050 (
);

FILL SFILL49080x48050 (
);

OR2X2 _10965_ (
    .A(_2047_),
    .B(_2054_),
    .Y(_2096_)
);

FILL FILL_0__8274_ (
);

OAI21X1 _10545_ (
    .A(_1860_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .C(_1861_),
    .Y(_1823_[19])
);

OAI21X1 _10125_ (
    .A(_1641_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .C(_1642_),
    .Y(_1628_[7])
);

FILL FILL_4__15493_ (
);

FILL FILL_4__15073_ (
);

FILL FILL_2__9653_ (
);

FILL FILL_3__14486_ (
);

FILL FILL_0__11621_ (
);

FILL FILL_2__9233_ (
);

FILL FILL_3__14066_ (
);

FILL FILL_0__11201_ (
);

FILL FILL_4__9999_ (
);

FILL FILL_4__9159_ (
);

FILL FILL_2__13899_ (
);

FILL FILL_2__13479_ (
);

FILL FILL_0__14093_ (
);

FILL SFILL33880x32050 (
);

FILL FILL_5__14813_ (
);

FILL FILL_1__7230_ (
);

FILL FILL_4__13806_ (
);

FILL FILL_2__14840_ (
);

FILL FILL_3__7996_ (
);

FILL FILL_2__14420_ (
);

FILL FILL_0__9899_ (
);

FILL SFILL49000x46050 (
);

FILL FILL_2__14000_ (
);

FILL FILL_3__7576_ (
);

FILL FILL_0__9479_ (
);

FILL FILL_1__13833_ (
);

FILL FILL_1__13413_ (
);

FILL FILL_4__16278_ (
);

FILL SFILL94440x55050 (
);

FILL FILL_0__12826_ (
);

FILL FILL_0__12406_ (
);

FILL FILL_5__8863_ (
);

FILL FILL_5__8443_ (
);

FILL FILL_0__15298_ (
);

AOI22X1 _15583_ (
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .B(_5571_),
    .C(_5570__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_6050_)
);

OAI22X1 _15163_ (
    .A(_5485__bF$buf2),
    .B(_4062_),
    .C(_4072_),
    .D(_5549__bF$buf1),
    .Y(_5641_)
);

FILL FILL_3__16212_ (
);

FILL FILL_1__8855_ (
);

FILL FILL_5__10313_ (
);

FILL FILL_1__8015_ (
);

FILL FILL_2__15625_ (
);

FILL SFILL2760x82050 (
);

FILL FILL_2__15205_ (
);

FILL FILL_4__6860_ (
);

FILL FILL_2__10760_ (
);

FILL FILL_1__14618_ (
);

NAND2X1 _7085_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_104_)
);

FILL FILL_4__12198_ (
);

FILL FILL_3__9722_ (
);

FILL SFILL94440x10050 (
);

FILL FILL_5__9648_ (
);

FILL FILL_5__9228_ (
);

FILL FILL_6__12525_ (
);

OAI21X1 _16368_ (
    .A(_6798_),
    .B(gnd),
    .C(_6799_),
    .Y(_6769_[15])
);

FILL SFILL23800x73050 (
);

FILL FILL_5__11938_ (
);

INVX2 _11083_ (
    .A(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2202_)
);

FILL FILL_3__12972_ (
);

FILL FILL_5__11518_ (
);

FILL FILL_3__12132_ (
);

FILL FILL_4__7225_ (
);

FILL FILL_2__11965_ (
);

FILL FILL111800x46050 (
);

FILL FILL_2__11545_ (
);

FILL FILL_2__11125_ (
);

FILL SFILL39000x44050 (
);

FILL SFILL94360x17050 (
);

FILL FILL_1__10958_ (
);

FILL FILL_1__10538_ (
);

FILL FILL_1__10118_ (
);

FILL SFILL109400x50 (
);

FILL FILL_5__15771_ (
);

FILL FILL_5__15351_ (
);

FILL FILL_0__7965_ (
);

FILL FILL_0__7545_ (
);

FILL FILL_0__7125_ (
);

NAND2X1 _9651_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1408_)
);

NAND2X1 _9231_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1189_)
);

FILL FILL_4__14764_ (
);

FILL SFILL8760x79050 (
);

FILL FILL_4__14344_ (
);

NAND3X1 _12288_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf4),
    .Y(_3255_)
);

FILL SFILL39400x13050 (
);

FILL FILL_2__8504_ (
);

FILL FILL_3__13757_ (
);

FILL FILL_3__13337_ (
);

FILL FILL_1__14791_ (
);

FILL FILL_1__14371_ (
);

FILL FILL_0__13784_ (
);

FILL SFILL114600x79050 (
);

FILL FILL_0__13364_ (
);

FILL SFILL53960x69050 (
);

FILL FILL_1__6921_ (
);

FILL FILL_3__6847_ (
);

FILL FILL_5__16136_ (
);

FILL FILL_5__11691_ (
);

FILL FILL_1__9393_ (
);

FILL FILL_5__11271_ (
);

FILL FILL_4__15969_ (
);

FILL FILL_4__15549_ (
);

FILL FILL_4__15129_ (
);

FILL FILL_2__16163_ (
);

FILL FILL_4__10684_ (
);

FILL FILL_4__10264_ (
);

FILL SFILL8760x34050 (
);

FILL SFILL13800x71050 (
);

FILL FILL_1__15996_ (
);

FILL FILL_1__15576_ (
);

FILL FILL_1__15156_ (
);

FILL FILL_5__7714_ (
);

FILL SFILL74040x82050 (
);

FILL FILL_1__10291_ (
);

FILL FILL_0__14989_ (
);

FILL FILL_0__14569_ (
);

INVX1 _14854_ (
    .A(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_5337_)
);

FILL FILL_0__14149_ (
);

INVX1 _14434_ (
    .A(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_4926_)
);

INVX1 _14014_ (
    .A(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_4515_)
);

FILL FILL_3__15903_ (
);

FILL SFILL53960x24050 (
);

FILL FILL_1__7706_ (
);

FILL SFILL84360x15050 (
);

FILL FILL_0__15930_ (
);

FILL FILL_0__15510_ (
);

FILL FILL_5__12896_ (
);

FILL FILL_5__12476_ (
);

FILL FILL_5__12056_ (
);

FILL FILL_3__13090_ (
);

FILL FILL_4__11889_ (
);

FILL FILL_4__8183_ (
);

FILL SFILL88680x23050 (
);

FILL FILL_4__11469_ (
);

FILL FILL_4__11049_ (
);

FILL FILL_2__12083_ (
);

FILL FILL_1__11496_ (
);

FILL FILL_1__11076_ (
);

OAI22X1 _15639_ (
    .A(_5485__bF$buf3),
    .B(_6104_),
    .C(_5483__bF$buf4),
    .D(_4621_),
    .Y(_6105_)
);

FILL FILL_4__12830_ (
);

FILL FILL_4__12410_ (
);

NAND3X1 _15219_ (
    .A(_5686_),
    .B(_5694_),
    .C(_5691_),
    .Y(_5695_)
);

OAI21X1 _10774_ (
    .A(_1972_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .C(_1973_),
    .Y(_1953_[10])
);

FILL FILL_0__10489_ (
);

FILL FILL_0__8083_ (
);

DFFSR _10354_ (
    .Q(\datapath_1.regfile_1.regOut[27] [28]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_1693_[28])
);

FILL FILL_0__10069_ (
);

FILL SFILL43960x67050 (
);

FILL FILL_3__11823_ (
);

FILL FILL_3__11403_ (
);

FILL FILL_4__6916_ (
);

FILL FILL_2__10816_ (
);

FILL FILL_2__9882_ (
);

FILL FILL_2__9462_ (
);

FILL FILL_0__11850_ (
);

FILL FILL_2__9042_ (
);

FILL FILL_3__14295_ (
);

FILL FILL_0__11430_ (
);

FILL FILL_0__11010_ (
);

FILL FILL_4__9388_ (
);

FILL FILL112360x71050 (
);

FILL FILL_2__13288_ (
);

FILL FILL_5__14622_ (
);

FILL FILL_5__14202_ (
);

DFFSR _8922_ (
    .Q(\datapath_1.regfile_1.regOut[16] [4]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_978_[4])
);

NAND2X1 _8502_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_825_)
);

FILL FILL_4__13615_ (
);

FILL SFILL64040x80050 (
);

OAI21X1 _11979_ (
    .A(_3026_),
    .B(IorD_bF$buf1),
    .C(_3027_),
    .Y(_1_[30])
);

FILL FILL_0__9288_ (
);

INVX1 _11559_ (
    .A(_2276_),
    .Y(_2668_)
);

OAI21X1 _11139_ (
    .A(_2251_),
    .B(_2252_),
    .C(_2257_),
    .Y(_2258_)
);

FILL SFILL3720x15050 (
);

FILL FILL_3__12608_ (
);

FILL FILL_1__13642_ (
);

FILL FILL_1__13222_ (
);

FILL FILL_4__16087_ (
);

FILL SFILL43960x22050 (
);

FILL FILL112280x78050 (
);

FILL FILL_1_BUFX2_insert500 (
);

FILL FILL_1_BUFX2_insert501 (
);

FILL FILL_0__12635_ (
);

DFFSR _12920_ (
    .Q(\datapath_1.a [1]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_3555_[1])
);

FILL FILL_1_BUFX2_insert502 (
);

FILL FILL_1_BUFX2_insert503 (
);

NAND2X1 _12500_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [20]),
    .Y(_3400_)
);

FILL FILL_0__12215_ (
);

FILL FILL_1_BUFX2_insert504 (
);

FILL FILL_1_BUFX2_insert505 (
);

FILL FILL_1_BUFX2_insert506 (
);

FILL FILL_5__8252_ (
);

FILL FILL_1_BUFX2_insert507 (
);

FILL FILL_1_BUFX2_insert508 (
);

FILL FILL_1_BUFX2_insert509 (
);

OAI22X1 _15392_ (
    .A(_5863_),
    .B(_5545__bF$buf1),
    .C(_5485__bF$buf4),
    .D(_4381_),
    .Y(_5864_)
);

FILL FILL_5__15827_ (
);

FILL FILL_5__15407_ (
);

DFFSR _9707_ (
    .Q(\datapath_1.regfile_1.regOut[22] [21]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_1368_[21])
);

FILL FILL_3__16021_ (
);

FILL FILL_5__10962_ (
);

FILL FILL_5__10542_ (
);

FILL FILL_5__10122_ (
);

FILL FILL_1__8244_ (
);

FILL SFILL104520x39050 (
);

FILL FILL_2__15854_ (
);

FILL FILL_2__15434_ (
);

FILL FILL_2__15014_ (
);

FILL SFILL24280x60050 (
);

FILL FILL_1__14847_ (
);

FILL FILL_1__14427_ (
);

FILL FILL_1__14007_ (
);

FILL FILL_3__9531_ (
);

FILL FILL_3__9111_ (
);

NOR2X1 _13705_ (
    .A(_4208_),
    .B(_4211_),
    .Y(_4212_)
);

FILL SFILL104120x25050 (
);

FILL FILL112280x33050 (
);

FILL FILL_5__9877_ (
);

FILL FILL_5__9037_ (
);

AOI22X1 _16177_ (
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .B(_5577_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_6629_)
);

FILL FILL_1__9869_ (
);

FILL FILL_5__11747_ (
);

FILL FILL_3__12781_ (
);

FILL FILL_5__11327_ (
);

FILL FILL_3__12361_ (
);

FILL FILL_1__9029_ (
);

FILL FILL_2__16219_ (
);

FILL FILL_4__7874_ (
);

FILL FILL_4__7454_ (
);

FILL FILL_4__7034_ (
);

FILL FILL_2__11774_ (
);

FILL FILL_2__11354_ (
);

INVX1 _8099_ (
    .A(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_617_)
);

FILL FILL_1__10767_ (
);

FILL FILL_2_CLKBUF1_insert220 (
);

FILL FILL_2_CLKBUF1_insert221 (
);

FILL FILL_2_CLKBUF1_insert222 (
);

FILL FILL_2_CLKBUF1_insert223 (
);

FILL FILL_5__15580_ (
);

FILL FILL_2_CLKBUF1_insert224 (
);

FILL FILL_5__15160_ (
);

NAND2X1 _9880_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1520_)
);

FILL FILL_0__7354_ (
);

DFFSR _9460_ (
    .Q(\datapath_1.regfile_1.regOut[20] [30]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_1238_[30])
);

INVX1 _9040_ (
    .A(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_1102_)
);

FILL FILL_4__14993_ (
);

FILL FILL_4__14573_ (
);

FILL FILL_4__14153_ (
);

AOI22X1 _12097_ (
    .A(\datapath_1.ALUResult [27]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3119_)
);

FILL FILL_3__13986_ (
);

FILL FILL_2__8733_ (
);

FILL FILL_0__10701_ (
);

FILL FILL_3__13566_ (
);

FILL FILL_2__8313_ (
);

FILL FILL_3__13146_ (
);

FILL FILL_1__14180_ (
);

FILL FILL_4__8659_ (
);

FILL FILL_4__8239_ (
);

FILL FILL_2__12979_ (
);

FILL FILL_0__13593_ (
);

FILL FILL_2__12139_ (
);

FILL SFILL33880x27050 (
);

FILL FILL_0__13173_ (
);

FILL FILL_4__9600_ (
);

FILL FILL_2__13920_ (
);

FILL FILL_5__16365_ (
);

FILL FILL_2__13500_ (
);

FILL FILL_0__8979_ (
);

FILL FILL_0__8139_ (
);

FILL FILL_5__11080_ (
);

FILL FILL_4__15778_ (
);

FILL FILL_1__12913_ (
);

FILL FILL_4__15358_ (
);

FILL FILL_2__16392_ (
);

FILL FILL_4__10493_ (
);

FILL FILL_0__9920_ (
);

FILL FILL_2__9938_ (
);

FILL FILL_0__11906_ (
);

FILL FILL_0__9500_ (
);

FILL FILL_2__9518_ (
);

FILL FILL_1__15385_ (
);

FILL FILL_5__7943_ (
);

FILL FILL_5__7103_ (
);

FILL FILL_0__14798_ (
);

FILL FILL_0__14378_ (
);

INVX1 _14663_ (
    .A(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_5150_)
);

NOR2X1 _14243_ (
    .A(_4723_),
    .B(_4738_),
    .Y(_4739_)
);

FILL FILL_3__15712_ (
);

FILL FILL_1__7935_ (
);

FILL FILL_2__14705_ (
);

FILL FILL_5__12285_ (
);

FILL SFILL84120x72050 (
);

FILL FILL_4__11698_ (
);

FILL FILL_4__11278_ (
);

FILL FILL_5__8728_ (
);

NAND3X1 _15868_ (
    .A(\datapath_1.regfile_1.regOut[4] [20]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf2),
    .Y(_6328_)
);

FILL SFILL23800x68050 (
);

INVX1 _15448_ (
    .A(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_5919_)
);

NOR2X1 _15028_ (
    .A(_5507_),
    .B(_5488_),
    .Y(_5508_)
);

FILL FILL_0__10298_ (
);

DFFSR _10583_ (
    .Q(\datapath_1.regfile_1.regOut[29] [1]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_1823_[1])
);

NAND2X1 _10163_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1668_)
);

FILL SFILL23880x25050 (
);

FILL FILL_3__11632_ (
);

FILL FILL_3__11212_ (
);

FILL FILL_0__16104_ (
);

FILL FILL_2__10625_ (
);

FILL FILL_2__9271_ (
);

FILL SFILL39000x39050 (
);

FILL FILL112440x2050 (
);

FILL FILL112360x7050 (
);

FILL FILL_2__13097_ (
);

FILL FILL_5__14851_ (
);

FILL FILL_5_BUFX2_insert90 (
);

FILL FILL_5__14431_ (
);

FILL FILL_5_BUFX2_insert91 (
);

FILL FILL_5__14011_ (
);

FILL FILL_5_BUFX2_insert92 (
);

NAND2X1 _8731_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_937_)
);

FILL FILL_5_BUFX2_insert93 (
);

NAND2X1 _8311_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .Y(_782_)
);

FILL FILL_5_BUFX2_insert94 (
);

FILL FILL_5_BUFX2_insert95 (
);

FILL FILL_4__13844_ (
);

FILL FILL_5_BUFX2_insert96 (
);

FILL FILL_4__13424_ (
);

FILL FILL_5_BUFX2_insert97 (
);

FILL FILL_5_BUFX2_insert98 (
);

FILL FILL_4__13004_ (
);

FILL FILL_5_BUFX2_insert99 (
);

FILL FILL_0__9097_ (
);

FILL FILL_3__7194_ (
);

OAI21X1 _11788_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(_2151_),
    .C(_2879_),
    .Y(_2881_)
);

OAI21X1 _11368_ (
    .A(_2320_),
    .B(_2347__bF$buf2),
    .C(_2484_),
    .Y(_2485_)
);

FILL SFILL23800x23050 (
);

FILL FILL_3__12837_ (
);

FILL FILL_1__13871_ (
);

FILL FILL_3__12417_ (
);

FILL FILL_1__13451_ (
);

FILL FILL_1__13031_ (
);

FILL SFILL84040x34050 (
);

FILL FILL_0__12864_ (
);

FILL FILL_0__12444_ (
);

FILL SFILL84840x17050 (
);

FILL FILL_0__12024_ (
);

FILL FILL_5__8481_ (
);

FILL FILL_5__8061_ (
);

FILL SFILL74200x4050 (
);

FILL FILL_5__15636_ (
);

FILL FILL_5__15216_ (
);

INVX1 _9936_ (
    .A(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_1557_)
);

FILL FILL_3__16250_ (
);

INVX1 _9516_ (
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_1338_)
);

FILL FILL_1__8893_ (
);

FILL FILL_5__10771_ (
);

FILL FILL_1__8473_ (
);

FILL FILL_4__14629_ (
);

FILL FILL_2__15663_ (
);

FILL FILL_4__14209_ (
);

FILL FILL_2__15243_ (
);

FILL FILL_3__8399_ (
);

FILL SFILL13800x66050 (
);

FILL FILL_1__14656_ (
);

FILL FILL_1__14236_ (
);

FILL FILL_3__9760_ (
);

FILL FILL_0__13649_ (
);

AOI21X1 _13934_ (
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .B(_4102_),
    .C(_4435_),
    .Y(_4436_)
);

FILL FILL_3__9340_ (
);

FILL FILL_0__13229_ (
);

OAI22X1 _13514_ (
    .A(_3890_),
    .B(_4024_),
    .C(_4023_),
    .D(_3931__bF$buf3),
    .Y(_4025_)
);

FILL FILL_5__9266_ (
);

FILL SFILL53960x19050 (
);

FILL FILL_5__11976_ (
);

FILL FILL_1__9678_ (
);

FILL FILL_5__11556_ (
);

FILL FILL_3__12590_ (
);

FILL FILL_1__9258_ (
);

FILL FILL_5__11136_ (
);

FILL FILL_3__12170_ (
);

FILL FILL_2__16028_ (
);

FILL FILL_4__7683_ (
);

FILL FILL_4__10969_ (
);

FILL FILL_4__10549_ (
);

BUFX2 BUFX2_insert1084 (
    .A(rst),
    .Y(rst_hier0_bF$buf9)
);

BUFX2 BUFX2_insert1085 (
    .A(rst),
    .Y(rst_hier0_bF$buf8)
);

FILL FILL_4__10129_ (
);

FILL FILL_2__11583_ (
);

BUFX2 BUFX2_insert1086 (
    .A(rst),
    .Y(rst_hier0_bF$buf7)
);

FILL FILL_2__11163_ (
);

BUFX2 BUFX2_insert1087 (
    .A(rst),
    .Y(rst_hier0_bF$buf6)
);

BUFX2 BUFX2_insert1088 (
    .A(rst),
    .Y(rst_hier0_bF$buf5)
);

BUFX2 BUFX2_insert1089 (
    .A(rst),
    .Y(rst_hier0_bF$buf4)
);

FILL SFILL13800x21050 (
);

FILL FILL_1__10996_ (
);

FILL FILL_1__10576_ (
);

FILL FILL_1__10156_ (
);

FILL FILL_4__11910_ (
);

INVX1 _14719_ (
    .A(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_5205_)
);

FILL SFILL74040x32050 (
);

FILL FILL_0__7583_ (
);

FILL FILL_0__7163_ (
);

FILL FILL_1_CLKBUF1_insert210 (
);

FILL FILL_3__10903_ (
);

FILL FILL_1_CLKBUF1_insert211 (
);

FILL FILL_1_CLKBUF1_insert212 (
);

FILL FILL_1_CLKBUF1_insert213 (
);

FILL FILL_4__14382_ (
);

FILL FILL_1_CLKBUF1_insert214 (
);

FILL FILL_1_CLKBUF1_insert215 (
);

FILL FILL_1_CLKBUF1_insert216 (
);

FILL FILL_1_CLKBUF1_insert217 (
);

FILL FILL_1_CLKBUF1_insert218 (
);

FILL FILL_2__8962_ (
);

FILL FILL_0__10930_ (
);

FILL FILL_3__13795_ (
);

FILL FILL_1_CLKBUF1_insert219 (
);

FILL FILL_0__10510_ (
);

FILL FILL_2__8122_ (
);

FILL FILL_3__13375_ (
);

FILL FILL_4__8888_ (
);

FILL FILL_4__8468_ (
);

FILL FILL112360x66050 (
);

FILL FILL_2__12788_ (
);

FILL FILL_2__12368_ (
);

FILL FILL_5__13702_ (
);

FILL FILL_3__6885_ (
);

FILL FILL_5__16174_ (
);

FILL FILL_0__8788_ (
);

FILL FILL_0__8368_ (
);

NAND2X1 _10639_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1904_)
);

DFFSR _10219_ (
    .Q(\datapath_1.regfile_1.regOut[26] [21]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1628_[21])
);

FILL FILL_1__12722_ (
);

FILL FILL_4__15587_ (
);

FILL FILL_1__12302_ (
);

FILL FILL_4__15167_ (
);

FILL SFILL43960x17050 (
);

FILL FILL_2__9747_ (
);

FILL FILL_0__11715_ (
);

FILL FILL_1__15194_ (
);

FILL FILL_5__7752_ (
);

FILL FILL_5__7332_ (
);

INVX1 _14892_ (
    .A(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_5374_)
);

FILL SFILL108920x35050 (
);

NAND3X1 _14472_ (
    .A(_4961_),
    .B(_4962_),
    .C(_4958_),
    .Y(_4963_)
);

FILL FILL_0__14187_ (
);

INVX1 _14052_ (
    .A(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_4552_)
);

FILL FILL_5__14907_ (
);

FILL FILL_3__15941_ (
);

FILL FILL112360x21050 (
);

FILL FILL_3__15521_ (
);

FILL FILL_3__15101_ (
);

FILL FILL_1__7744_ (
);

FILL FILL_1__7324_ (
);

FILL FILL_2__14934_ (
);

FILL FILL_2__14514_ (
);

FILL SFILL64040x30050 (
);

FILL FILL_5__12094_ (
);

FILL FILL_1__13927_ (
);

FILL FILL_1__13507_ (
);

FILL SFILL84360x6050 (
);

FILL FILL_4__11087_ (
);

FILL FILL_3__8611_ (
);

FILL FILL112280x28050 (
);

FILL FILL_1__16399_ (
);

FILL FILL_5__8957_ (
);

FILL FILL_5__8117_ (
);

OAI22X1 _15677_ (
    .A(_5466__bF$buf0),
    .B(_6141_),
    .C(_4684_),
    .D(_5483__bF$buf3),
    .Y(_6142_)
);

NAND3X1 _15257_ (
    .A(_5726_),
    .B(_5732_),
    .C(_5722_),
    .Y(_5733_)
);

FILL FILL_3__16306_ (
);

NAND2X1 _10392_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1780_)
);

FILL SFILL83640x8050 (
);

FILL FILL_5__10827_ (
);

FILL FILL_5__10407_ (
);

FILL FILL_3__11861_ (
);

FILL FILL_1__8529_ (
);

FILL FILL_1__8109_ (
);

FILL FILL_3__11441_ (
);

FILL FILL_3__11021_ (
);

FILL FILL_2__15719_ (
);

FILL FILL_4__6954_ (
);

FILL FILL_0__16333_ (
);

FILL FILL_5__13299_ (
);

FILL FILL_2__10434_ (
);

FILL SFILL54040x73050 (
);

FILL FILL_2__9080_ (
);

FILL FILL_2__10014_ (
);

INVX1 _7599_ (
    .A(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_365_)
);

INVX1 _7179_ (
    .A(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_146_)
);

FILL FILL_5__14660_ (
);

FILL FILL_5__14240_ (
);

FILL FILL_0__6854_ (
);

NAND2X1 _8960_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1049_)
);

DFFSR _8540_ (
    .Q(\datapath_1.regfile_1.regOut[13] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_783_[6])
);

INVX1 _8120_ (
    .A(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_631_)
);

FILL FILL_6__12619_ (
);

FILL FILL_4__13653_ (
);

FILL FILL_4__13233_ (
);

AOI21X1 _11597_ (
    .A(_2424_),
    .B(_2703_),
    .C(_2692_),
    .Y(_2704_)
);

NOR2X1 _11177_ (
    .A(_2295_),
    .B(_2294_),
    .Y(_2296_)
);

FILL FILL_2__7813_ (
);

FILL FILL_3__12646_ (
);

FILL FILL_1__13680_ (
);

FILL FILL_3__12226_ (
);

FILL FILL_1__13260_ (
);

FILL FILL_4__7739_ (
);

FILL FILL_4__7319_ (
);

FILL FILL_2__11639_ (
);

FILL FILL_2__11219_ (
);

FILL FILL_0__12253_ (
);

FILL FILL_6__16032_ (
);

FILL FILL_5__15865_ (
);

FILL FILL_5__15445_ (
);

FILL FILL_5__15025_ (
);

INVX1 _9745_ (
    .A(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_1450_)
);

FILL FILL_0__7219_ (
);

DFFSR _9325_ (
    .Q(\datapath_1.regfile_1.regOut[19] [23]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_1173_[23])
);

FILL FILL_5__10580_ (
);

FILL FILL_5__10160_ (
);

FILL FILL_4__14858_ (
);

FILL FILL_2__15892_ (
);

FILL FILL_4__14438_ (
);

FILL FILL_4__14018_ (
);

FILL FILL_2__15472_ (
);

FILL FILL_2__15052_ (
);

FILL FILL_1__14885_ (
);

FILL FILL_1__14465_ (
);

FILL FILL_1__14045_ (
);

FILL FILL_0__13878_ (
);

INVX1 _13743_ (
    .A(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_4249_)
);

FILL FILL_0__13458_ (
);

OAI21X1 _13323_ (
    .A(\datapath_1.a3 [4]),
    .B(_3852_),
    .C(_3848_),
    .Y(_3853_)
);

FILL FILL_0__13038_ (
);

FILL FILL_5__9495_ (
);

FILL SFILL44040x71050 (
);

FILL FILL_6__12372_ (
);

FILL SFILL8120x72050 (
);

FILL FILL_5__11785_ (
);

FILL FILL_1__9487_ (
);

FILL FILL_5__11365_ (
);

FILL FILL_2__16257_ (
);

FILL FILL_4__7492_ (
);

FILL FILL_4__7072_ (
);

FILL FILL_4__10778_ (
);

FILL FILL_4__10358_ (
);

FILL FILL_2__11392_ (
);

FILL FILL_5__7808_ (
);

FILL FILL_1__10385_ (
);

INVX1 _14948_ (
    .A(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_5429_)
);

AOI22X1 _14528_ (
    .A(\datapath_1.regfile_1.regOut[27] [22]),
    .B(_4129_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_5018_)
);

NOR2X1 _14108_ (
    .A(_4606_),
    .B(_3971__bF$buf2),
    .Y(_4607_)
);

FILL SFILL84520x36050 (
);

FILL FILL_6__13577_ (
);

FILL FILL_4__14191_ (
);

FILL FILL_0__15604_ (
);

FILL FILL_2__8771_ (
);

FILL FILL_2__8351_ (
);

FILL FILL_4__8697_ (
);

FILL FILL_4__8277_ (
);

FILL SFILL53640x7050 (
);

FILL FILL_2__12597_ (
);

FILL FILL_2__12177_ (
);

FILL FILL_5__13931_ (
);

FILL FILL_5__13511_ (
);

NAND2X1 _7811_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_466_)
);

FILL FILL_4__12504_ (
);

FILL FILL_6__9984_ (
);

FILL FILL_0__8597_ (
);

DFFSR _10868_ (
    .Q(\datapath_1.regfile_1.regOut[31] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_1953_[30])
);

FILL SFILL23800x18050 (
);

INVX1 _10448_ (
    .A(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_1817_)
);

INVX1 _10028_ (
    .A(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_1598_)
);

FILL FILL_3__11917_ (
);

FILL FILL_1__12951_ (
);

FILL FILL_4__15396_ (
);

FILL FILL_1__12531_ (
);

FILL FILL_1__12111_ (
);

FILL FILL_2__9976_ (
);

FILL FILL_0__11944_ (
);

FILL FILL_2__9556_ (
);

FILL FILL_2__9136_ (
);

FILL FILL_3__14389_ (
);

FILL FILL_0__11524_ (
);

FILL FILL_0__11104_ (
);

FILL SFILL104360x5050 (
);

FILL FILL_5__7981_ (
);

FILL FILL_5__7561_ (
);

FILL SFILL74120x65050 (
);

OAI22X1 _14281_ (
    .A(_3959_),
    .B(_4775_),
    .C(_3954__bF$buf2),
    .D(_4774_),
    .Y(_4776_)
);

FILL FILL_5__14716_ (
);

FILL FILL_3__15750_ (
);

FILL FILL_3__15330_ (
);

FILL FILL_1__7973_ (
);

FILL FILL_1__7553_ (
);

FILL FILL_4__13709_ (
);

FILL FILL_2__14743_ (
);

FILL FILL_2__14323_ (
);

FILL SFILL109320x20050 (
);

FILL FILL_3__7479_ (
);

FILL FILL_3__7059_ (
);

FILL FILL_1__13736_ (
);

FILL FILL_1__13316_ (
);

FILL FILL_3__8840_ (
);

FILL FILL_0__12729_ (
);

FILL FILL_3__8000_ (
);

FILL FILL_0__12309_ (
);

FILL FILL_5__8766_ (
);

FILL FILL_5__8346_ (
);

OAI22X1 _15486_ (
    .A(_4440_),
    .B(_5548__bF$buf4),
    .C(_5489__bF$buf3),
    .D(_4438_),
    .Y(_5956_)
);

OAI22X1 _15066_ (
    .A(_5544__bF$buf3),
    .B(_5543_),
    .C(_5545__bF$buf1),
    .D(_3922_),
    .Y(_5546_)
);

FILL SFILL74120x20050 (
);

FILL FILL_3__16115_ (
);

FILL FILL_5__10636_ (
);

FILL FILL_1__8758_ (
);

FILL FILL_1__8338_ (
);

FILL FILL_3__11670_ (
);

FILL FILL_3__11250_ (
);

FILL FILL_2__15948_ (
);

FILL FILL_2__15528_ (
);

FILL FILL_2__15108_ (
);

FILL FILL_0__16142_ (
);

FILL FILL_2__10663_ (
);

FILL FILL_2__10243_ (
);

FILL FILL_3__9625_ (
);

FILL FILL_3_BUFX2_insert410 (
);

FILL FILL_3_BUFX2_insert411 (
);

FILL FILL_3_BUFX2_insert412 (
);

FILL FILL_3_BUFX2_insert413 (
);

FILL FILL_3_BUFX2_insert414 (
);

FILL FILL_3_BUFX2_insert415 (
);

FILL FILL_3_BUFX2_insert416 (
);

FILL FILL_3_BUFX2_insert417 (
);

FILL FILL_3_BUFX2_insert418 (
);

FILL FILL_6__12428_ (
);

FILL FILL_4__13882_ (
);

FILL FILL_3_BUFX2_insert419 (
);

FILL FILL_4__13462_ (
);

FILL FILL_4__13042_ (
);

FILL SFILL64120x63050 (
);

FILL FILL_2__7622_ (
);

FILL FILL_3__12875_ (
);

FILL FILL_2__7202_ (
);

FILL FILL_3__12455_ (
);

FILL FILL_3__12035_ (
);

FILL FILL_4__7968_ (
);

FILL FILL_4__7548_ (
);

FILL FILL_2__11868_ (
);

FILL FILL_2__11448_ (
);

FILL FILL_0__12482_ (
);

FILL FILL_2__11028_ (
);

FILL FILL_0__12062_ (
);

FILL SFILL89240x3050 (
);

FILL SFILL23720x1050 (
);

FILL FILL_5__15674_ (
);

FILL FILL_0__7868_ (
);

FILL FILL_5__15254_ (
);

FILL SFILL113880x74050 (
);

INVX1 _9974_ (
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_1626_)
);

FILL FILL_0__7448_ (
);

OAI21X1 _9554_ (
    .A(_1362_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1363_),
    .Y(_1303_[30])
);

OAI21X1 _9134_ (
    .A(_1143_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .C(_1144_),
    .Y(_1108_[18])
);

FILL FILL_1__8091_ (
);

FILL FILL_1__11802_ (
);

FILL FILL_4__14667_ (
);

FILL FILL_4__14247_ (
);

FILL FILL_2__15281_ (
);

FILL FILL_2__8827_ (
);

FILL FILL_1__14694_ (
);

FILL FILL_1__14274_ (
);

FILL FILL_0_BUFX2_insert540 (
);

FILL FILL_0_BUFX2_insert541 (
);

FILL FILL_0_BUFX2_insert542 (
);

FILL FILL_0_BUFX2_insert543 (
);

FILL FILL_0_BUFX2_insert544 (
);

AOI22X1 _13972_ (
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .B(_3894_),
    .C(_3995__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_4474_)
);

FILL FILL_0__13687_ (
);

FILL FILL_0__13267_ (
);

FILL FILL_0_BUFX2_insert545 (
);

INVX1 _13552_ (
    .A(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_4062_)
);

FILL FILL_0_BUFX2_insert546 (
);

OAI21X1 _13132_ (
    .A(_3718_),
    .B(PCEn_bF$buf0),
    .C(_3719_),
    .Y(_3685_[17])
);

FILL FILL112360x16050 (
);

FILL FILL_0_BUFX2_insert547 (
);

FILL FILL_3__14601_ (
);

FILL FILL_0_BUFX2_insert548 (
);

FILL FILL_0_BUFX2_insert549 (
);

FILL FILL_5__16039_ (
);

FILL SFILL64040x25050 (
);

FILL FILL_5__11594_ (
);

FILL FILL_5__11174_ (
);

FILL FILL_1__9296_ (
);

FILL FILL_2__16066_ (
);

FILL FILL_4__10167_ (
);

FILL FILL_1__15899_ (
);

FILL SFILL54120x61050 (
);

FILL FILL_1__15479_ (
);

FILL FILL_1__15059_ (
);

FILL FILL_5__7617_ (
);

FILL SFILL113880x4050 (
);

FILL FILL_1__10194_ (
);

OAI22X1 _14757_ (
    .A(_5240_),
    .B(_3916_),
    .C(_3983__bF$buf2),
    .D(_5241_),
    .Y(_5242_)
);

INVX1 _14337_ (
    .A(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_4831_)
);

FILL FILL_3__15806_ (
);

FILL FILL_1__16000_ (
);

FILL FILL_3__10941_ (
);

FILL FILL_1__7609_ (
);

FILL FILL_3__10521_ (
);

FILL FILL_0__15833_ (
);

FILL FILL_0__15413_ (
);

FILL SFILL54040x68050 (
);

FILL FILL_2__8580_ (
);

FILL FILL_5__12379_ (
);

FILL FILL_4__8086_ (
);

FILL FILL_5__13740_ (
);

FILL FILL_5__13320_ (
);

INVX1 _7620_ (
    .A(\datapath_1.regfile_1.regOut[6] [26]),
    .Y(_379_)
);

INVX1 _7200_ (
    .A(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_160_)
);

FILL FILL_1__11399_ (
);

FILL FILL_4__12733_ (
);

FILL FILL_4__12313_ (
);

INVX1 _10677_ (
    .A(\datapath_1.regfile_1.regOut[30] [21]),
    .Y(_1929_)
);

INVX1 _10257_ (
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_1710_)
);

FILL FILL_3__11726_ (
);

FILL FILL_1__12760_ (
);

FILL FILL_3__11306_ (
);

FILL FILL_1__12340_ (
);

FILL FILL_2__9785_ (
);

FILL FILL_0__11753_ (
);

FILL FILL_2__9365_ (
);

FILL FILL_3__14198_ (
);

FILL FILL_0__11333_ (
);

FILL SFILL54040x23050 (
);

FILL FILL_5__7370_ (
);

FILL FILL_6__15112_ (
);

FILL FILL_5__14945_ (
);

INVX1 _14090_ (
    .A(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_4589_)
);

FILL FILL_5__14525_ (
);

FILL FILL_5__14105_ (
);

INVX1 _8825_ (
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_979_)
);

OAI21X1 _8405_ (
    .A(_779_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_780_),
    .Y(_718_[31])
);

FILL SFILL79240x72050 (
);

FILL FILL_1__7362_ (
);

FILL FILL_4__13938_ (
);

FILL FILL_2__14972_ (
);

FILL FILL_4__13518_ (
);

FILL FILL_2__14552_ (
);

FILL FILL_2__14132_ (
);

FILL FILL_3__7288_ (
);

FILL FILL_1__13965_ (
);

FILL FILL_1__13545_ (
);

FILL SFILL59240x2050 (
);

FILL FILL_1__13125_ (
);

FILL SFILL59160x7050 (
);

FILL FILL_0__12958_ (
);

INVX1 _12823_ (
    .A(\datapath_1.a [0]),
    .Y(_3618_)
);

INVX1 _12403_ (
    .A(ALUOut[20]),
    .Y(_3334_)
);

FILL FILL_0__12118_ (
);

FILL FILL_5__8995_ (
);

FILL FILL_5__8575_ (
);

FILL SFILL44040x66050 (
);

NOR3X1 _15295_ (
    .A(_5760_),
    .B(_5751_),
    .C(_5769_),
    .Y(_5770_)
);

FILL FILL_3__16344_ (
);

FILL FILL_1__8987_ (
);

FILL FILL_1__8567_ (
);

FILL FILL_5__10445_ (
);

FILL FILL_1__8147_ (
);

FILL FILL_5__10025_ (
);

FILL FILL_2__15757_ (
);

FILL FILL_2__15337_ (
);

FILL FILL_4__6992_ (
);

FILL FILL_0__16371_ (
);

FILL FILL_2__10892_ (
);

FILL FILL_2__10052_ (
);

FILL FILL_3__9854_ (
);

FILL FILL_3__9014_ (
);

NOR2X1 _13608_ (
    .A(_4116_),
    .B(_3954__bF$buf1),
    .Y(_4117_)
);

FILL FILL_0__6892_ (
);

FILL FILL_4__13691_ (
);

FILL FILL_4__13271_ (
);

FILL FILL_2__7851_ (
);

FILL FILL_2__7431_ (
);

FILL FILL_3__12264_ (
);

FILL FILL_4__7357_ (
);

FILL FILL_2__11677_ (
);

FILL FILL_2__11257_ (
);

FILL FILL_0__12291_ (
);

FILL FILL_5__15483_ (
);

FILL FILL_5__15063_ (
);

FILL FILL_0__7677_ (
);

OAI21X1 _9783_ (
    .A(_1474_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .C(_1475_),
    .Y(_1433_[21])
);

OAI21X1 _9363_ (
    .A(_1255_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .C(_1256_),
    .Y(_1238_[9])
);

FILL FILL_4__14896_ (
);

FILL FILL_4__14476_ (
);

FILL FILL_1__11611_ (
);

FILL FILL_4__14056_ (
);

FILL FILL_2__15090_ (
);

FILL FILL_2__8636_ (
);

FILL FILL_3__13889_ (
);

FILL FILL_3__13469_ (
);

FILL FILL_2__8216_ (
);

FILL FILL_1__14083_ (
);

INVX1 _13781_ (
    .A(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_4287_)
);

FILL FILL_0__13496_ (
);

NOR2X1 _13361_ (
    .A(_3874_),
    .B(_3876_),
    .Y(\datapath_1.regfile_1.regEn [28])
);

FILL FILL_3__14830_ (
);

FILL FILL_3__14410_ (
);

FILL FILL_4__9923_ (
);

FILL FILL_4__9503_ (
);

FILL FILL_2__13823_ (
);

FILL FILL_2__13403_ (
);

FILL FILL_5__16268_ (
);

FILL FILL_3__6979_ (
);

FILL FILL_2__16295_ (
);

FILL FILL_4__10396_ (
);

FILL SFILL69160x32050 (
);

FILL FILL_3__7500_ (
);

FILL FILL_0__9403_ (
);

FILL FILL_0__11809_ (
);

FILL FILL_1__15288_ (
);

FILL FILL_5__7846_ (
);

FILL FILL_5__7426_ (
);

FILL FILL_4__16202_ (
);

NAND3X1 _14986_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5461_),
    .C(_5465_),
    .Y(_5466_)
);

INVX1 _14566_ (
    .A(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_5055_)
);

AOI22X1 _14146_ (
    .A(_3894_),
    .B(\datapath_1.regfile_1.regOut[28] [14]),
    .C(\datapath_1.regfile_1.regOut[3] [14]),
    .D(_3942__bF$buf2),
    .Y(_4644_)
);

FILL SFILL28920x4050 (
);

FILL FILL_3__15615_ (
);

FILL FILL_1__7838_ (
);

FILL FILL_1__7418_ (
);

FILL FILL_3__10750_ (
);

FILL SFILL28840x9050 (
);

FILL FILL_2__14608_ (
);

FILL SFILL99320x64050 (
);

FILL FILL_0__15642_ (
);

FILL FILL_0__15222_ (
);

FILL FILL_5__12188_ (
);

FILL SFILL8760x5050 (
);

FILL FILL_3__8705_ (
);

FILL SFILL59160x75050 (
);

FILL SFILL68680x6050 (
);

FILL FILL_4__12962_ (
);

FILL SFILL64120x58050 (
);

FILL FILL_4__12122_ (
);

INVX1 _10486_ (
    .A(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_1886_)
);

OAI21X1 _10066_ (
    .A(_1622_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .C(_1623_),
    .Y(_1563_[30])
);

FILL FILL_3__11955_ (
);

FILL FILL_3__11535_ (
);

FILL FILL_3__11115_ (
);

FILL FILL_0__16007_ (
);

FILL FILL_2__10948_ (
);

FILL FILL_2__10528_ (
);

FILL FILL_0__11982_ (
);

FILL FILL_2__9594_ (
);

FILL FILL_0__11562_ (
);

FILL FILL_2__10108_ (
);

FILL FILL_0__11142_ (
);

FILL FILL_6__15761_ (
);

FILL FILL_5__14754_ (
);

FILL FILL_0__6948_ (
);

FILL FILL_5__14334_ (
);

OAI21X1 _8634_ (
    .A(_891_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .C(_892_),
    .Y(_848_[22])
);

FILL SFILL59160x30050 (
);

OAI21X1 _8214_ (
    .A(_672_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_673_),
    .Y(_653_[10])
);

FILL FILL_1__7591_ (
);

FILL FILL_1__7171_ (
);

FILL FILL_4__13747_ (
);

FILL FILL_4__13327_ (
);

FILL FILL_2__14781_ (
);

FILL FILL_2__14361_ (
);

FILL FILL_3__7097_ (
);

FILL SFILL64120x13050 (
);

FILL FILL_1__13774_ (
);

FILL FILL_1__13354_ (
);

FILL FILL_0__12767_ (
);

OAI21X1 _12632_ (
    .A(_3466_),
    .B(vdd),
    .C(_3467_),
    .Y(_3425_[21])
);

FILL FILL_0__12347_ (
);

FILL SFILL89320x62050 (
);

NAND3X1 _12212_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3197_)
);

FILL FILL_5__8384_ (
);

FILL FILL_6__11681_ (
);

FILL FILL_5__15959_ (
);

FILL FILL_5__15539_ (
);

FILL FILL_5__15119_ (
);

FILL FILL_3__16153_ (
);

DFFSR _9839_ (
    .Q(\datapath_1.regfile_1.regOut[23] [25]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_1433_[25])
);

FILL SFILL18760x82050 (
);

NAND2X1 _9419_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1294_)
);

FILL FILL_5__10674_ (
);

FILL FILL_5__10254_ (
);

FILL FILL_1__8376_ (
);

FILL FILL_2__15986_ (
);

FILL FILL_2__15566_ (
);

FILL FILL_2__15146_ (
);

FILL FILL_0__16180_ (
);

FILL SFILL89240x69050 (
);

FILL FILL_2__10281_ (
);

FILL SFILL54120x56050 (
);

FILL FILL_1__14979_ (
);

FILL FILL_1__14559_ (
);

FILL FILL_1__14139_ (
);

FILL FILL_3__9663_ (
);

NOR2X1 _13837_ (
    .A(_4341_),
    .B(_4338_),
    .Y(_4342_)
);

FILL FILL_3__9243_ (
);

INVX1 _13417_ (
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_3929_)
);

FILL FILL_1__15920_ (
);

FILL FILL_1__15500_ (
);

FILL FILL_5__9169_ (
);

FILL FILL_4__13080_ (
);

FILL FILL_0__14913_ (
);

FILL FILL_5__11879_ (
);

FILL FILL_5__11459_ (
);

FILL FILL_3__12493_ (
);

FILL FILL_5__11039_ (
);

FILL FILL_2__7240_ (
);

FILL FILL_3__12073_ (
);

FILL FILL_4__7586_ (
);

FILL FILL_4__7166_ (
);

FILL FILL_2__11486_ (
);

FILL FILL_2__11066_ (
);

FILL FILL_5__12400_ (
);

FILL FILL_1__10899_ (
);

FILL SFILL54120x11050 (
);

FILL FILL_1__10059_ (
);

FILL FILL_4__11813_ (
);

FILL FILL_5__15292_ (
);

FILL FILL_0__7486_ (
);

OAI21X1 _9592_ (
    .A(_1431_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1432_),
    .Y(_1368_[0])
);

FILL FILL_0__7066_ (
);

NAND2X1 _9172_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1170_)
);

FILL FILL_3__10806_ (
);

FILL SFILL18680x44050 (
);

FILL FILL_1__11840_ (
);

FILL FILL_4__14285_ (
);

FILL FILL_1__11420_ (
);

FILL FILL_1__11000_ (
);

FILL FILL_2__8865_ (
);

FILL FILL_0__10833_ (
);

FILL FILL_2__8445_ (
);

FILL FILL_3__13698_ (
);

FILL FILL_3__13278_ (
);

FILL FILL_0__10413_ (
);

FILL FILL111960x73050 (
);

FILL SFILL54040x18050 (
);

FILL FILL_0_BUFX2_insert920 (
);

FILL FILL_5__6870_ (
);

FILL FILL_0_BUFX2_insert921 (
);

FILL FILL_0_BUFX2_insert922 (
);

FILL FILL_0_BUFX2_insert923 (
);

FILL FILL_0_BUFX2_insert924 (
);

OAI22X1 _13590_ (
    .A(_3944__bF$buf2),
    .B(_4097_),
    .C(_4098_),
    .D(_3955__bF$buf3),
    .Y(_4099_)
);

FILL FILL_0_BUFX2_insert925 (
);

NAND2X1 _13170_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_pcsrc.dout [30]),
    .Y(_3745_)
);

FILL FILL_0_BUFX2_insert926 (
);

FILL FILL_5__13605_ (
);

FILL FILL_0_BUFX2_insert927 (
);

FILL FILL_0_BUFX2_insert928 (
);

DFFSR _7905_ (
    .Q(\datapath_1.regfile_1.regOut[8] [11]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_458_[11])
);

FILL FILL_0_BUFX2_insert929 (
);

FILL SFILL79240x67050 (
);

FILL FILL_1__6862_ (
);

FILL FILL_4__9732_ (
);

FILL FILL_2__13632_ (
);

FILL FILL_2__13212_ (
);

FILL FILL_5__16077_ (
);

FILL FILL_6__9658_ (
);

FILL FILL_1__12625_ (
);

FILL FILL_1__12205_ (
);

FILL FILL_0__9632_ (
);

NAND2X1 _11903_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[5]),
    .Y(_2977_)
);

FILL FILL_0__9212_ (
);

FILL FILL_0__11618_ (
);

FILL FILL_1__15097_ (
);

FILL FILL_5__7235_ (
);

FILL FILL_4__16011_ (
);

FILL FILL_6__10532_ (
);

INVX1 _14795_ (
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_5279_)
);

AOI22X1 _14375_ (
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .B(_4246_),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_4868_)
);

FILL FILL_3__15844_ (
);

FILL FILL_3__15424_ (
);

FILL FILL_3__15004_ (
);

FILL FILL_1__7227_ (
);

FILL FILL_6_BUFX2_insert301 (
);

FILL FILL_2__14837_ (
);

FILL SFILL79240x22050 (
);

FILL FILL_2__14417_ (
);

FILL FILL_0__15871_ (
);

FILL FILL_0__15451_ (
);

FILL FILL_0__15031_ (
);

FILL FILL_6_BUFX2_insert306 (
);

FILL FILL_3__8514_ (
);

FILL SFILL109400x48050 (
);

FILL FILL_6__11737_ (
);

FILL FILL_4__12771_ (
);

FILL SFILL44040x16050 (
);

FILL FILL_4__12351_ (
);

FILL FILL_3__16209_ (
);

OAI21X1 _10295_ (
    .A(_1734_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .C(_1735_),
    .Y(_1693_[21])
);

FILL FILL_2__6931_ (
);

FILL FILL_3__11764_ (
);

FILL FILL_5__9801_ (
);

FILL FILL_3__11344_ (
);

FILL SFILL69240x65050 (
);

FILL FILL_4__6857_ (
);

FILL FILL_0__16236_ (
);

NAND3X1 _16101_ (
    .A(_6550_),
    .B(_6551_),
    .C(_6554_),
    .Y(_6555_)
);

FILL FILL_2__10757_ (
);

FILL FILL_0__11791_ (
);

FILL FILL_0__11371_ (
);

FILL FILL_3__9719_ (
);

FILL FILL_5__14983_ (
);

FILL FILL_5__14563_ (
);

FILL FILL_5__14143_ (
);

OAI21X1 _8863_ (
    .A(_1003_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1004_),
    .Y(_978_[13])
);

OAI21X1 _8443_ (
    .A(_784_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .C(_785_),
    .Y(_783_[1])
);

DFFSR _8023_ (
    .Q(\datapath_1.regfile_1.regOut[9] [1]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_523_[1])
);

FILL FILL_4__13976_ (
);

FILL FILL_4__13556_ (
);

FILL FILL_2__14590_ (
);

FILL FILL_4__13136_ (
);

FILL FILL_2__14170_ (
);

FILL FILL_2__7716_ (
);

FILL FILL_3__12969_ (
);

FILL FILL_3__12129_ (
);

FILL FILL_1__13583_ (
);

FILL FILL_1__13163_ (
);

FILL FILL_0__12996_ (
);

FILL FILL_0__12576_ (
);

OAI21X1 _12861_ (
    .A(_3578_),
    .B(vdd),
    .C(_3579_),
    .Y(_3555_[12])
);

OAI21X1 _12441_ (
    .A(_3423_),
    .B(vdd),
    .C(_3424_),
    .Y(_3360_[0])
);

FILL FILL_0__12156_ (
);

AOI22X1 _12021_ (
    .A(\datapath_1.ALUResult [8]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3062_)
);

FILL FILL_3__13910_ (
);

FILL FILL_6__16355_ (
);

FILL FILL_5__8193_ (
);

FILL FILL_5_BUFX2_insert320 (
);

FILL FILL_5_BUFX2_insert321 (
);

FILL FILL_2__12903_ (
);

FILL FILL_5__15768_ (
);

FILL FILL_5_BUFX2_insert322 (
);

FILL FILL_5__15348_ (
);

FILL FILL_3__16382_ (
);

FILL FILL_5_BUFX2_insert323 (
);

FILL FILL_5_BUFX2_insert324 (
);

NAND2X1 _9648_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1406_)
);

NAND2X1 _9228_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1187_)
);

FILL FILL_5_BUFX2_insert325 (
);

FILL FILL_5_BUFX2_insert326 (
);

FILL FILL_5__10063_ (
);

FILL FILL_5_BUFX2_insert327 (
);

FILL FILL_1__8185_ (
);

FILL FILL_5_BUFX2_insert328 (
);

FILL FILL_2__15795_ (
);

FILL FILL_5_BUFX2_insert329 (
);

FILL FILL_2__15375_ (
);

FILL SFILL38760x36050 (
);

FILL SFILL69160x27050 (
);

FILL FILL_0__8903_ (
);

FILL FILL_1__14788_ (
);

FILL FILL_1__14368_ (
);

FILL FILL_5__6926_ (
);

FILL FILL_4__15702_ (
);

FILL FILL_3__9892_ (
);

FILL FILL_3__9472_ (
);

INVX8 _13646_ (
    .A(_3982__bF$buf0),
    .Y(_4154_)
);

NOR2X1 _13226_ (
    .A(_3768_),
    .B(_3762_),
    .Y(_3769_)
);

FILL FILL_5__9398_ (
);

FILL FILL_1__6918_ (
);

FILL FILL_6__12275_ (
);

FILL SFILL99320x59050 (
);

FILL FILL_0__14722_ (
);

FILL FILL_0__14302_ (
);

FILL FILL_5__11688_ (
);

FILL FILL_5__11268_ (
);

FILL SFILL28760x79050 (
);

FILL FILL_2__11295_ (
);

FILL FILL_2_BUFX2_insert450 (
);

FILL FILL_2_BUFX2_insert451 (
);

FILL FILL_1__10288_ (
);

FILL FILL_2_BUFX2_insert452 (
);

FILL FILL_2_BUFX2_insert453 (
);

FILL FILL_2_BUFX2_insert454 (
);

FILL FILL_4__11622_ (
);

FILL FILL_2_BUFX2_insert455 (
);

FILL FILL_4__11202_ (
);

FILL FILL_2_BUFX2_insert456 (
);

FILL FILL_0__7295_ (
);

FILL FILL_2_BUFX2_insert457 (
);

FILL FILL_2_BUFX2_insert458 (
);

FILL FILL_6__8262_ (
);

FILL FILL_2_BUFX2_insert459 (
);

FILL FILL_3__10615_ (
);

FILL FILL_0_CLKBUF1_insert150 (
);

FILL FILL_0_CLKBUF1_insert151 (
);

FILL FILL_4__14094_ (
);

FILL FILL_0__15927_ (
);

FILL FILL_0_CLKBUF1_insert152 (
);

FILL FILL_0__15507_ (
);

FILL FILL_0_CLKBUF1_insert153 (
);

FILL FILL_0_CLKBUF1_insert154 (
);

FILL FILL_0_CLKBUF1_insert155 (
);

FILL FILL_0_CLKBUF1_insert156 (
);

FILL SFILL99320x14050 (
);

FILL FILL_0_CLKBUF1_insert157 (
);

FILL FILL_2__8254_ (
);

FILL FILL_0__10642_ (
);

FILL FILL_0_CLKBUF1_insert158 (
);

FILL FILL_3__13087_ (
);

FILL FILL_0_CLKBUF1_insert159 (
);

FILL FILL_6__14421_ (
);

FILL FILL_6__14001_ (
);

FILL FILL_5__13834_ (
);

FILL SFILL89400x50050 (
);

FILL FILL_5__13414_ (
);

FILL SFILL28760x34050 (
);

FILL SFILL59160x25050 (
);

OAI21X1 _7714_ (
    .A(_420_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_421_),
    .Y(_393_[14])
);

FILL FILL_4__9541_ (
);

FILL FILL_4__9121_ (
);

FILL FILL_4__12827_ (
);

FILL FILL_4__12407_ (
);

FILL FILL_2__13861_ (
);

FILL FILL_2__13441_ (
);

FILL FILL_2__13021_ (
);

FILL FILL_6__9467_ (
);

FILL FILL_1__12854_ (
);

FILL FILL_1__12434_ (
);

FILL FILL_4__15299_ (
);

FILL FILL_1__12014_ (
);

FILL SFILL28360x20050 (
);

FILL FILL_2__9879_ (
);

FILL FILL_0__9861_ (
);

FILL FILL_0__11847_ (
);

FILL SFILL89320x57050 (
);

FILL FILL_2__9039_ (
);

FILL FILL_0__9021_ (
);

FILL FILL_0__11427_ (
);

OAI21X1 _11712_ (
    .A(_2376_),
    .B(_2380_),
    .C(_2390_),
    .Y(_2811_)
);

FILL FILL_0__11007_ (
);

FILL FILL_5__7884_ (
);

FILL FILL_5__7464_ (
);

FILL FILL_4__16240_ (
);

FILL FILL_5__7044_ (
);

NOR2X1 _14184_ (
    .A(_4680_),
    .B(_3977__bF$buf4),
    .Y(_4681_)
);

FILL FILL_5__14619_ (
);

FILL FILL_3__15653_ (
);

FILL SFILL18760x77050 (
);

FILL FILL_3__15233_ (
);

DFFSR _8919_ (
    .Q(\datapath_1.regfile_1.regOut[16] [1]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_978_[1])
);

FILL FILL_1__7876_ (
);

FILL SFILL113880x19050 (
);

FILL FILL_1__7456_ (
);

FILL FILL_1__7036_ (
);

FILL FILL_2__14646_ (
);

FILL FILL_0__15680_ (
);

FILL FILL_2__14226_ (
);

FILL FILL_0__15260_ (
);

FILL SFILL89720x26050 (
);

FILL FILL_1__13639_ (
);

FILL FILL_1__13219_ (
);

FILL FILL_1_BUFX2_insert470 (
);

FILL FILL_1_BUFX2_insert471 (
);

FILL FILL_3__8743_ (
);

FILL FILL_3__8323_ (
);

FILL FILL_1_BUFX2_insert472 (
);

NAND2X1 _12917_ (
    .A(vdd),
    .B(\datapath_1.rd1 [31]),
    .Y(_3617_)
);

FILL FILL_1_BUFX2_insert473 (
);

FILL FILL_1_BUFX2_insert474 (
);

FILL SFILL33960x52050 (
);

FILL FILL_1_BUFX2_insert475 (
);

FILL FILL_1_BUFX2_insert476 (
);

FILL FILL_5__8249_ (
);

FILL FILL_1_BUFX2_insert477 (
);

FILL SFILL89320x12050 (
);

FILL FILL_1_BUFX2_insert478 (
);

FILL FILL_1_BUFX2_insert479 (
);

FILL FILL_4__12580_ (
);

NOR2X1 _15389_ (
    .A(_5860_),
    .B(_5853_),
    .Y(_5861_)
);

FILL FILL_4__12160_ (
);

FILL FILL_3__16018_ (
);

FILL FILL_5__10959_ (
);

FILL FILL_5__10539_ (
);

FILL FILL_3__11993_ (
);

FILL FILL_5__9610_ (
);

FILL FILL_3__11573_ (
);

FILL FILL_5__10119_ (
);

FILL FILL_3__11153_ (
);

FILL SFILL18760x32050 (
);

INVX1 _16330_ (
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_6774_)
);

FILL FILL_0__16045_ (
);

FILL FILL_2__10566_ (
);

FILL FILL_2__10146_ (
);

FILL FILL_0__11180_ (
);

FILL FILL_5__11900_ (
);

FILL FILL_1__9602_ (
);

FILL SFILL89240x19050 (
);

FILL FILL_3__9528_ (
);

FILL FILL_3__9108_ (
);

FILL FILL_5__14792_ (
);

FILL FILL_0__6986_ (
);

FILL FILL_5__14372_ (
);

FILL FILL_6__7953_ (
);

DFFSR _8672_ (
    .Q(\datapath_1.regfile_1.regOut[14] [10]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_848_[10])
);

NAND2X1 _8252_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_699_)
);

FILL SFILL18680x39050 (
);

FILL FILL_1__10920_ (
);

FILL FILL_4__13785_ (
);

FILL FILL_4__13365_ (
);

FILL FILL_1__10500_ (
);

FILL FILL_2__7945_ (
);

FILL FILL_3__12778_ (
);

FILL FILL111960x68050 (
);

FILL FILL_3__12358_ (
);

FILL FILL_2__7105_ (
);

FILL FILL_1__13392_ (
);

DFFSR _12670_ (
    .Q(\datapath_1.Data [7]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3425_[7])
);

FILL FILL_0__12385_ (
);

NAND3X1 _12250_ (
    .A(_3224_),
    .B(_3225_),
    .C(_3226_),
    .Y(\datapath_1.alu_1.ALUInB [8])
);

FILL FILL_2_CLKBUF1_insert190 (
);

FILL FILL_2_CLKBUF1_insert191 (
);

FILL FILL_2_CLKBUF1_insert192 (
);

FILL FILL_5__15997_ (
);

FILL FILL_2_CLKBUF1_insert193 (
);

FILL FILL_2__12712_ (
);

FILL FILL_5__15577_ (
);

FILL FILL_2_CLKBUF1_insert194 (
);

FILL FILL_5__15157_ (
);

FILL FILL_2_CLKBUF1_insert195 (
);

FILL FILL_6__8738_ (
);

FILL FILL_3__16191_ (
);

NAND2X1 _9877_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1518_)
);

FILL FILL_2_CLKBUF1_insert196 (
);

DFFSR _9457_ (
    .Q(\datapath_1.regfile_1.regOut[20] [27]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_1238_[27])
);

INVX1 _9037_ (
    .A(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_1100_)
);

FILL FILL_2_CLKBUF1_insert197 (
);

FILL FILL_2_CLKBUF1_insert198 (
);

FILL FILL_5__10292_ (
);

FILL FILL_2_CLKBUF1_insert199 (
);

FILL FILL_1__11705_ (
);

FILL FILL_2__15184_ (
);

FILL SFILL114440x80050 (
);

FILL FILL_0__8712_ (
);

FILL FILL_1__14597_ (
);

FILL FILL_1__14177_ (
);

FILL FILL_4__15931_ (
);

FILL FILL_4__15511_ (
);

FILL FILL_6_BUFX2_insert1073 (
);

INVX1 _13875_ (
    .A(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_4379_)
);

FILL FILL_3__9281_ (
);

NAND3X1 _13455_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3903_),
    .C(_3919_),
    .Y(_3967_)
);

INVX1 _13035_ (
    .A(_2_[28]),
    .Y(_3675_)
);

FILL FILL_3__14924_ (
);

FILL FILL_3__14504_ (
);

FILL FILL_2__13917_ (
);

FILL FILL_0__14951_ (
);

FILL FILL_0__14531_ (
);

FILL FILL_0__14111_ (
);

FILL FILL_5__11497_ (
);

FILL FILL_5__11077_ (
);

FILL FILL_2__16389_ (
);

FILL FILL_0__9917_ (
);

FILL SFILL114760x56050 (
);

FILL FILL_4__11851_ (
);

FILL FILL_4__11431_ (
);

FILL FILL_4__11011_ (
);

FILL FILL_3__15709_ (
);

FILL FILL_1__16323_ (
);

FILL FILL_3__10424_ (
);

FILL FILL_3__10004_ (
);

FILL FILL_0__15736_ (
);

FILL FILL_0__15316_ (
);

OAI22X1 _15601_ (
    .A(_5478__bF$buf3),
    .B(_6067_),
    .C(_4585_),
    .D(_5530__bF$buf1),
    .Y(_6068_)
);

FILL FILL_2__8483_ (
);

FILL FILL_0__10871_ (
);

FILL FILL_2__8063_ (
);

FILL FILL_0__10451_ (
);

FILL FILL_0__10031_ (
);

FILL SFILL100200x5050 (
);

FILL FILL_5__13643_ (
);

FILL FILL_5__13223_ (
);

OAI21X1 _7943_ (
    .A(_532_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_533_),
    .Y(_523_[5])
);

DFFSR _7523_ (
    .Q(\datapath_1.regfile_1.regOut[5] [13]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_263_[13])
);

NAND2X1 _7103_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_116_)
);

FILL FILL_4__9770_ (
);

FILL FILL_4__9350_ (
);

FILL FILL_4__12636_ (
);

FILL FILL_2__13670_ (
);

FILL FILL_4__12216_ (
);

FILL FILL_2__13250_ (
);

FILL FILL_3__11629_ (
);

FILL FILL_3__11209_ (
);

FILL FILL_1__12243_ (
);

FILL FILL_0__9670_ (
);

FILL SFILL69240x15050 (
);

FILL FILL_0__9250_ (
);

INVX1 _11941_ (
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3002_)
);

FILL FILL_2__9268_ (
);

FILL FILL_0__11656_ (
);

FILL FILL_0__11236_ (
);

OAI21X1 _11521_ (
    .A(_2631_),
    .B(_2278_),
    .C(_2410_),
    .Y(_2632_)
);

NOR2X1 _11101_ (
    .A(_2217_),
    .B(_2219_),
    .Y(_2220_)
);

FILL FILL_5__7693_ (
);

FILL FILL_6__10150_ (
);

FILL FILL_5__14848_ (
);

FILL FILL_3__15882_ (
);

FILL FILL_5__14428_ (
);

FILL FILL_5__14008_ (
);

FILL FILL_3__15462_ (
);

NAND2X1 _8728_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_935_)
);

FILL FILL_3__15042_ (
);

DFFSR _8308_ (
    .Q(\datapath_1.regfile_1.regOut[11] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_653_[30])
);

FILL FILL_1__7685_ (
);

FILL FILL_2__14875_ (
);

FILL FILL_2__14455_ (
);

FILL FILL_2__14035_ (
);

FILL FILL_1__13868_ (
);

FILL FILL_1__13448_ (
);

FILL FILL_1__13028_ (
);

FILL FILL_3__8972_ (
);

FILL SFILL59240x58050 (
);

NAND2X1 _12726_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[10]),
    .Y(_3510_)
);

FILL FILL_3__8132_ (
);

NAND3X1 _12306_ (
    .A(_3266_),
    .B(_3267_),
    .C(_3268_),
    .Y(\datapath_1.alu_1.ALUInB [22])
);

FILL FILL_5__8898_ (
);

FILL FILL_5__8478_ (
);

FILL FILL_5__8058_ (
);

INVX1 _15198_ (
    .A(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_5675_)
);

FILL FILL_0__13802_ (
);

FILL FILL_3__16247_ (
);

FILL FILL_5__10768_ (
);

FILL SFILL3800x35050 (
);

FILL FILL_3__11382_ (
);

FILL FILL_4__6895_ (
);

FILL FILL_0__16274_ (
);

FILL FILL_2__10795_ (
);

FILL FILL_2__10375_ (
);

FILL FILL_1__9411_ (
);

FILL FILL_3__9757_ (
);

FILL FILL_3__9337_ (
);

FILL FILL_4__10702_ (
);

FILL FILL_5__14181_ (
);

NAND2X1 _8481_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_811_)
);

NAND2X1 _8061_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_592_)
);

FILL FILL_4__13594_ (
);

FILL FILL_4__13174_ (
);

FILL FILL_2__7754_ (
);

FILL FILL_3__12587_ (
);

FILL FILL_2__7334_ (
);

FILL FILL_3__12167_ (
);

FILL FILL_0__12194_ (
);

FILL SFILL89400x45050 (
);

FILL FILL_5__12914_ (
);

FILL FILL_4__8621_ (
);

FILL FILL_4__8201_ (
);

FILL FILL_4__11907_ (
);

FILL FILL_5_BUFX2_insert700 (
);

FILL FILL_5_BUFX2_insert701 (
);

FILL FILL_5__15386_ (
);

FILL FILL_5_BUFX2_insert702 (
);

FILL FILL_2__12521_ (
);

FILL FILL_2__12101_ (
);

FILL FILL_5_BUFX2_insert703 (
);

FILL FILL_5_BUFX2_insert704 (
);

DFFSR _9686_ (
    .Q(\datapath_1.regfile_1.regOut[22] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_1368_[0])
);

FILL FILL_5_BUFX2_insert705 (
);

INVX1 _9266_ (
    .A(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_1212_)
);

FILL FILL_1_CLKBUF1_insert180 (
);

FILL FILL_5_BUFX2_insert706 (
);

FILL FILL_1_CLKBUF1_insert181 (
);

FILL FILL_5_BUFX2_insert707 (
);

FILL FILL_1__11934_ (
);

FILL FILL_4__14799_ (
);

FILL FILL_5_BUFX2_insert708 (
);

FILL FILL_1_CLKBUF1_insert182 (
);

FILL FILL_5_BUFX2_insert709 (
);

FILL FILL_1_CLKBUF1_insert183 (
);

FILL FILL_4__14379_ (
);

FILL FILL_1__11514_ (
);

FILL FILL_1_CLKBUF1_insert184 (
);

FILL FILL_1_CLKBUF1_insert185 (
);

FILL FILL_1_CLKBUF1_insert186 (
);

FILL FILL_1_CLKBUF1_insert187 (
);

FILL FILL_2__8959_ (
);

FILL FILL_1_CLKBUF1_insert188 (
);

FILL FILL_0__10927_ (
);

FILL FILL_0__8521_ (
);

FILL FILL_1_CLKBUF1_insert189 (
);

FILL FILL_0__10507_ (
);

FILL FILL_2__8119_ (
);

FILL FILL_0__8101_ (
);

FILL FILL_5__6964_ (
);

FILL FILL_4__15740_ (
);

FILL FILL_4__15320_ (
);

FILL FILL_3__9090_ (
);

NAND3X1 _13684_ (
    .A(_4190_),
    .B(_4191_),
    .C(_4189_),
    .Y(_4192_)
);

FILL FILL_0__13399_ (
);

OR2X2 _13264_ (
    .A(_3796_),
    .B(_3806_),
    .Y(_3807_)
);

FILL FILL_2__9900_ (
);

FILL FILL_3__14733_ (
);

FILL FILL_3__14313_ (
);

FILL FILL_1__6956_ (
);

FILL FILL_4__9406_ (
);

FILL SFILL94280x51050 (
);

FILL FILL_2__13726_ (
);

FILL FILL_2__13306_ (
);

FILL FILL_0__14760_ (
);

FILL FILL_0__14340_ (
);

FILL FILL_1__12719_ (
);

FILL FILL_2__16198_ (
);

FILL FILL_4__10299_ (
);

FILL FILL_3__7823_ (
);

FILL FILL_0__9726_ (
);

FILL FILL_5__7749_ (
);

FILL FILL_5__7329_ (
);

FILL FILL_2_BUFX2_insert830 (
);

FILL FILL_4__16105_ (
);

FILL FILL_2_BUFX2_insert831 (
);

FILL FILL_2_BUFX2_insert832 (
);

FILL FILL_6__10626_ (
);

FILL FILL_2_BUFX2_insert833 (
);

AOI22X1 _14889_ (
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .B(_4246_),
    .C(_4115_),
    .D(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_5371_)
);

NOR2X1 _14469_ (
    .A(_4959_),
    .B(_3977__bF$buf3),
    .Y(_4960_)
);

FILL FILL_2_BUFX2_insert834 (
);

FILL FILL_4__11660_ (
);

FILL FILL_2_BUFX2_insert835 (
);

INVX1 _14049_ (
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_4549_)
);

FILL FILL_4__11240_ (
);

FILL FILL_2_BUFX2_insert836 (
);

FILL FILL_3__15938_ (
);

FILL FILL_3__15518_ (
);

FILL FILL_2_BUFX2_insert837 (
);

FILL FILL_2_BUFX2_insert838 (
);

FILL FILL_2_BUFX2_insert839 (
);

FILL FILL_1__16132_ (
);

FILL SFILL79400x43050 (
);

FILL FILL_3__10653_ (
);

FILL SFILL18760x27050 (
);

FILL FILL_3__10233_ (
);

FILL FILL_0__15965_ (
);

FILL FILL_0__15545_ (
);

INVX1 _15830_ (
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_6291_)
);

OAI22X1 _15410_ (
    .A(_5463__bF$buf3),
    .B(_5881_),
    .C(_5880_),
    .D(_5504__bF$buf1),
    .Y(_5882_)
);

FILL FILL_0__15125_ (
);

FILL FILL_0__10680_ (
);

FILL FILL_0__10260_ (
);

FILL FILL_3__8608_ (
);

FILL FILL_5__13872_ (
);

FILL FILL_5__13452_ (
);

FILL FILL_5__13032_ (
);

NAND2X1 _7752_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_447_)
);

NAND2X1 _7332_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_228_)
);

FILL FILL_4__12865_ (
);

FILL FILL_4__12445_ (
);

FILL FILL_4__12025_ (
);

FILL FILL_6__9085_ (
);

NAND2X1 _10389_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1778_)
);

FILL FILL_3__11858_ (
);

FILL FILL_1__12892_ (
);

FILL FILL_3__11438_ (
);

FILL FILL_1__12472_ (
);

FILL FILL_3__11018_ (
);

FILL FILL_1__12052_ (
);

FILL FILL_0__11885_ (
);

FILL FILL_2__9497_ (
);

FILL FILL_0__11465_ (
);

AND2X2 _11750_ (
    .A(_2376_),
    .B(_2503_),
    .Y(_2846_)
);

FILL FILL_0__11045_ (
);

AOI21X1 _11330_ (
    .A(_2447_),
    .B(_2440_),
    .C(_2448_),
    .Y(_2449_)
);

FILL SFILL79720x19050 (
);

FILL FILL_6__15664_ (
);

FILL SFILL110120x67050 (
);

FILL FILL_5__7082_ (
);

FILL FILL_5__14657_ (
);

FILL SFILL59880x6050 (
);

FILL FILL_3__15691_ (
);

FILL FILL_5__14237_ (
);

FILL FILL_6__7818_ (
);

FILL FILL_3__15271_ (
);

NAND2X1 _8957_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1047_)
);

DFFSR _8537_ (
    .Q(\datapath_1.regfile_1.regOut[13] [3]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_783_[3])
);

INVX1 _8117_ (
    .A(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_629_)
);

FILL FILL_1__7494_ (
);

FILL FILL_1__7074_ (
);

FILL FILL_2__14684_ (
);

FILL SFILL114440x75050 (
);

FILL FILL_2__14264_ (
);

FILL FILL_1__13677_ (
);

FILL FILL_1__13257_ (
);

FILL FILL111960x18050 (
);

FILL FILL_1_BUFX2_insert850 (
);

FILL FILL_3__8781_ (
);

FILL FILL_1_BUFX2_insert851 (
);

FILL FILL_1_BUFX2_insert852 (
);

FILL FILL_3__8361_ (
);

NAND2X1 _12955_ (
    .A(vdd),
    .B(\datapath_1.rd2 [1]),
    .Y(_3622_)
);

FILL FILL_1_BUFX2_insert853 (
);

DFFSR _12535_ (
    .Q(ALUOut[0]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3360_[0])
);

FILL FILL_1_BUFX2_insert854 (
);

INVX1 _12115_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3194_)
);

FILL FILL_1_BUFX2_insert855 (
);

FILL FILL_1_BUFX2_insert856 (
);

FILL FILL_1_BUFX2_insert857 (
);

FILL FILL_1_BUFX2_insert858 (
);

FILL FILL_1_BUFX2_insert859 (
);

FILL FILL_6__11584_ (
);

FILL FILL_0__13611_ (
);

FILL FILL_3__16056_ (
);

FILL FILL_5__10997_ (
);

FILL FILL_5__10577_ (
);

FILL FILL_1__8699_ (
);

FILL FILL_5__10157_ (
);

FILL FILL_3__11191_ (
);

FILL FILL_2__15889_ (
);

FILL FILL_2__15469_ (
);

FILL SFILL69320x48050 (
);

FILL FILL_2__15049_ (
);

FILL FILL_0__16083_ (
);

FILL FILL_2__10184_ (
);

FILL SFILL114440x30050 (
);

FILL FILL_1__9640_ (
);

FILL FILL_1__9220_ (
);

FILL FILL_2__16410_ (
);

FILL FILL_3__9986_ (
);

FILL SFILL13560x74050 (
);

FILL FILL_4__10931_ (
);

FILL FILL_3__9146_ (
);

FILL FILL_4__10511_ (
);

FILL FILL_1__15823_ (
);

FILL FILL_1__15403_ (
);

DFFSR _8290_ (
    .Q(\datapath_1.regfile_1.regOut[11] [12]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_653_[12])
);

FILL FILL_6__12789_ (
);

FILL FILL_0__14816_ (
);

FILL FILL_2__7983_ (
);

FILL FILL_2__7563_ (
);

BUFX2 BUFX2_insert520 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf87)
);

BUFX2 BUFX2_insert521 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf86)
);

FILL FILL_3__12396_ (
);

BUFX2 BUFX2_insert522 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf85)
);

BUFX2 BUFX2_insert523 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf84)
);

BUFX2 BUFX2_insert524 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf83)
);

FILL FILL_6__13730_ (
);

BUFX2 BUFX2_insert525 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf82)
);

FILL FILL_4__7489_ (
);

BUFX2 BUFX2_insert526 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf81)
);

FILL FILL_4__7069_ (
);

BUFX2 BUFX2_insert527 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf80)
);

BUFX2 BUFX2_insert528 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf79)
);

FILL FILL_2__11389_ (
);

BUFX2 BUFX2_insert529 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf78)
);

FILL FILL_5__12723_ (
);

FILL FILL_5__12303_ (
);

FILL FILL_4__8850_ (
);

FILL FILL_4__8010_ (
);

FILL FILL_4__11716_ (
);

FILL FILL_2__12750_ (
);

FILL FILL_5__15195_ (
);

FILL FILL_2__12330_ (
);

FILL FILL_6__8356_ (
);

INVX1 _9495_ (
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_1324_)
);

DFFSR _9075_ (
    .Q(\datapath_1.regfile_1.regOut[17] [29]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_1043_[29])
);

FILL FILL_3__10709_ (
);

FILL FILL_1__11743_ (
);

FILL FILL_4__14188_ (
);

FILL FILL_1__11323_ (
);

FILL FILL_2__8768_ (
);

FILL FILL_0__8750_ (
);

FILL FILL_0__8330_ (
);

FILL FILL_2__8348_ (
);

FILL FILL_0__10316_ (
);

DFFSR _10601_ (
    .Q(\datapath_1.regfile_1.regOut[29] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1823_[19])
);

FILL FILL_0_BUFX2_insert40 (
);

FILL FILL_0_BUFX2_insert41 (
);

FILL FILL_0_BUFX2_insert42 (
);

FILL FILL_0_BUFX2_insert43 (
);

FILL FILL_0_BUFX2_insert44 (
);

FILL FILL_0_BUFX2_insert45 (
);

FILL FILL_0_BUFX2_insert46 (
);

FILL FILL_0_BUFX2_insert47 (
);

AOI21X1 _13493_ (
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .B(_4001__bF$buf1),
    .C(_4003_),
    .Y(_4004_)
);

FILL FILL_0_BUFX2_insert48 (
);

DFFSR _13073_ (
    .Q(_2_[26]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3620_[26])
);

FILL FILL_5__13928_ (
);

FILL FILL_0_BUFX2_insert49 (
);

FILL FILL_3__14962_ (
);

FILL FILL_5__13508_ (
);

FILL FILL_3__14542_ (
);

NAND2X1 _7808_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_464_)
);

FILL FILL_3__14122_ (
);

FILL FILL_4_BUFX2_insert360 (
);

FILL FILL_4__9635_ (
);

FILL FILL_4_BUFX2_insert361 (
);

FILL FILL_4__9215_ (
);

FILL FILL_4_BUFX2_insert362 (
);

FILL FILL_2__13955_ (
);

FILL FILL_4_BUFX2_insert363 (
);

FILL FILL_4_BUFX2_insert364 (
);

FILL FILL_2__13535_ (
);

FILL FILL_4_BUFX2_insert365 (
);

FILL FILL_2__13115_ (
);

FILL FILL_4_BUFX2_insert366 (
);

FILL FILL_4_BUFX2_insert367 (
);

FILL FILL_4_BUFX2_insert368 (
);

FILL FILL_4_BUFX2_insert369 (
);

FILL FILL_1__12528_ (
);

FILL FILL_1__12108_ (
);

FILL FILL_0__9535_ (
);

FILL FILL_3__7632_ (
);

FILL FILL_0__9115_ (
);

FILL FILL_3__7212_ (
);

AOI21X1 _11806_ (
    .A(_2368_),
    .B(_2363_),
    .C(_2458_),
    .Y(_2898_)
);

FILL FILL_5__7978_ (
);

FILL SFILL104360x35050 (
);

FILL FILL_5__7558_ (
);

FILL FILL_4__16334_ (
);

INVX1 _14698_ (
    .A(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_5184_)
);

OAI22X1 _14278_ (
    .A(_3982__bF$buf2),
    .B(_4771_),
    .C(_3971__bF$buf3),
    .D(_4772_),
    .Y(_4773_)
);

FILL FILL_3__15747_ (
);

FILL FILL_3__15327_ (
);

FILL FILL_1__16361_ (
);

FILL FILL_3__10882_ (
);

FILL FILL_3__10042_ (
);

FILL FILL_0__15774_ (
);

FILL FILL_0__15354_ (
);

FILL FILL_1__8911_ (
);

FILL FILL_3__8837_ (
);

FILL FILL_5__13681_ (
);

FILL FILL_5__13261_ (
);

FILL FILL_6__6842_ (
);

NAND2X1 _7981_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_559_)
);

FILL FILL112440x41050 (
);

NAND2X1 _7561_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_340_)
);

DFFSR _7141_ (
    .Q(\datapath_1.regfile_1.regOut[2] [15]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_68_[15])
);

FILL FILL_4__12254_ (
);

DFFSR _10198_ (
    .Q(\datapath_1.regfile_1.regOut[26] [0]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_1628_[0])
);

FILL SFILL114520x6050 (
);

FILL FILL_3__11667_ (
);

FILL FILL_3__11247_ (
);

FILL SFILL108600x41050 (
);

FILL FILL_1__12281_ (
);

DFFSR _16424_ (
    .Q(\datapath_1.regfile_1.regOut[0] [7]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_6769_[7])
);

FILL FILL_0__16139_ (
);

NAND2X1 _16004_ (
    .A(_6455_),
    .B(_6460_),
    .Y(_6461_)
);

FILL FILL_0__11694_ (
);

FILL FILL_0__11274_ (
);

FILL SFILL113800x8050 (
);

FILL FILL_3_BUFX2_insert380 (
);

FILL FILL_4__7701_ (
);

FILL FILL_3_BUFX2_insert381 (
);

FILL FILL_3_BUFX2_insert382 (
);

FILL FILL_5__14886_ (
);

FILL FILL_5__14466_ (
);

FILL FILL_3_BUFX2_insert383 (
);

FILL FILL_2__11601_ (
);

FILL FILL_5__14046_ (
);

FILL FILL_3_BUFX2_insert384 (
);

INVX1 _8766_ (
    .A(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_960_)
);

FILL FILL_3_BUFX2_insert385 (
);

FILL FILL_6__7627_ (
);

FILL FILL_3__15080_ (
);

FILL FILL_3_BUFX2_insert386 (
);

INVX1 _8346_ (
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_741_)
);

FILL FILL_3_BUFX2_insert387 (
);

FILL FILL_3_BUFX2_insert388 (
);

FILL FILL_4__13879_ (
);

FILL FILL_3_BUFX2_insert389 (
);

FILL FILL_4__13459_ (
);

FILL FILL_2__14493_ (
);

FILL FILL_4__13039_ (
);

FILL FILL_2__14073_ (
);

FILL FILL_0__7601_ (
);

FILL FILL_2__7619_ (
);

FILL FILL_1__13486_ (
);

FILL FILL_4__14820_ (
);

FILL FILL_4__14400_ (
);

FILL FILL_3__8590_ (
);

FILL FILL_0__12899_ (
);

INVX1 _12764_ (
    .A(\datapath_1.PCJump [25]),
    .Y(_3535_)
);

FILL FILL_0__12479_ (
);

NAND2X1 _12344_ (
    .A(\datapath_1.Data [0]),
    .B(MemToReg_bF$buf5),
    .Y(_3359_)
);

FILL FILL_0__12059_ (
);

FILL FILL_3__13813_ (
);

FILL FILL_6__16258_ (
);

FILL FILL_5__8096_ (
);

FILL FILL_4__8906_ (
);

FILL SFILL94280x46050 (
);

FILL FILL_0__13840_ (
);

FILL FILL_0__13420_ (
);

FILL FILL_3__16285_ (
);

FILL FILL_0__13000_ (
);

FILL FILL_5__10386_ (
);

FILL FILL_1__8088_ (
);

FILL FILL_2__15698_ (
);

FILL FILL_2__15278_ (
);

FILL FILL_3__6903_ (
);

FILL FILL_4__15605_ (
);

FILL FILL_3__9795_ (
);

OAI22X1 _13969_ (
    .A(_3884__bF$buf3),
    .B(_4469_),
    .C(_3955__bF$buf4),
    .D(_4470_),
    .Y(_4471_)
);

FILL FILL_3__9375_ (
);

INVX1 _13549_ (
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_4059_)
);

OAI21X1 _13129_ (
    .A(_3716_),
    .B(PCEn_bF$buf1),
    .C(_3717_),
    .Y(_3685_[16])
);

FILL FILL_4__10320_ (
);

FILL FILL_1__15632_ (
);

FILL FILL_1__15212_ (
);

FILL FILL_6__12598_ (
);

FILL FILL_0__14625_ (
);

INVX1 _14910_ (
    .A(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_5392_)
);

FILL FILL_0__14205_ (
);

FILL FILL_2__7372_ (
);

FILL FILL_4__7298_ (
);

FILL FILL_2__11198_ (
);

FILL SFILL33160x14050 (
);

FILL FILL_5__12952_ (
);

FILL FILL_5__12532_ (
);

FILL SFILL33800x7050 (
);

FILL FILL_5__12112_ (
);

FILL SFILL8680x63050 (
);

FILL FILL_4__11945_ (
);

FILL SFILL74280x7050 (
);

FILL FILL_4__11525_ (
);

FILL SFILL109560x80050 (
);

FILL FILL_4__11105_ (
);

FILL SFILL23240x50050 (
);

FILL FILL_0__7198_ (
);

FILL FILL_3__10938_ (
);

FILL FILL_1__11972_ (
);

FILL FILL_3__10518_ (
);

FILL FILL_1__11552_ (
);

FILL SFILL105160x79050 (
);

FILL FILL_1__11132_ (
);

FILL SFILL84280x44050 (
);

FILL FILL_2__8997_ (
);

FILL FILL_2__8577_ (
);

FILL FILL_0__10965_ (
);

NAND2X1 _10830_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_2011_)
);

FILL FILL_0__10545_ (
);

FILL FILL_0__10125_ (
);

NAND2X1 _10410_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1792_)
);

FILL FILL_6__14324_ (
);

FILL FILL_5__13737_ (
);

FILL FILL_5__13317_ (
);

FILL FILL_3__14771_ (
);

FILL FILL_3__14351_ (
);

FILL SFILL8600x61050 (
);

INVX1 _7617_ (
    .A(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_377_)
);

FILL FILL_1__6994_ (
);

FILL FILL_4__9864_ (
);

FILL FILL_4__9024_ (
);

FILL FILL_2__13764_ (
);

FILL FILL_2__13344_ (
);

FILL FILL_1__12757_ (
);

FILL FILL_1__12337_ (
);

FILL FILL_3__7861_ (
);

FILL FILL_0__9764_ (
);

FILL FILL_0__9344_ (
);

FILL FILL_3__7441_ (
);

INVX2 _11615_ (
    .A(_2257_),
    .Y(_2720_)
);

FILL FILL_5__7367_ (
);

FILL FILL_4__16143_ (
);

FILL SFILL13640x62050 (
);

INVX1 _14087_ (
    .A(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_4586_)
);

FILL FILL_3__15976_ (
);

FILL FILL_3__15556_ (
);

FILL FILL_3__15136_ (
);

FILL SFILL109480x42050 (
);

FILL FILL_1__16170_ (
);

FILL FILL_1__7359_ (
);

FILL FILL_3__10691_ (
);

FILL FILL_3__10271_ (
);

FILL FILL_2__14969_ (
);

FILL FILL_2__14549_ (
);

FILL FILL_2__14129_ (
);

FILL FILL_0__15583_ (
);

FILL SFILL74680x56050 (
);

FILL FILL_0__15163_ (
);

FILL SFILL114440x25050 (
);

FILL FILL_1__8720_ (
);

FILL FILL_2__15910_ (
);

FILL FILL_3__8646_ (
);

FILL FILL_3__8226_ (
);

FILL FILL_5__13490_ (
);

DFFSR _7790_ (
    .Q(\datapath_1.regfile_1.regOut[7] [24]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_393_[24])
);

FILL FILL_1__14903_ (
);

INVX1 _7370_ (
    .A(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_253_)
);

FILL FILL_4__12483_ (
);

FILL FILL_4__12063_ (
);

FILL FILL_5__9933_ (
);

FILL FILL_3__11896_ (
);

FILL FILL_5__9513_ (
);

FILL FILL_3__11476_ (
);

FILL FILL_3__11056_ (
);

FILL FILL_1__12090_ (
);

FILL FILL_4__6989_ (
);

FILL FILL_0__16368_ (
);

OAI21X1 _16233_ (
    .A(_5524__bF$buf3),
    .B(_5347_),
    .C(_6683_),
    .Y(_6684_)
);

FILL FILL_2__10889_ (
);

FILL FILL_2__10049_ (
);

FILL FILL_0__11083_ (
);

FILL FILL_1__9925_ (
);

FILL FILL_5__11803_ (
);

FILL FILL_1__9505_ (
);

FILL FILL_4__7930_ (
);

FILL FILL_2__11830_ (
);

FILL FILL_5__14695_ (
);

FILL FILL_0__6889_ (
);

FILL FILL_5__14275_ (
);

FILL FILL_2__11410_ (
);

FILL SFILL74200x40050 (
);

INVX1 _8995_ (
    .A(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_1072_)
);

INVX1 _8575_ (
    .A(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_853_)
);

FILL FILL_6__7436_ (
);

DFFSR _8155_ (
    .Q(\datapath_1.regfile_1.regOut[10] [5]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_588_[5])
);

FILL FILL_1__10823_ (
);

FILL FILL_4__13688_ (
);

FILL FILL_4__13268_ (
);

FILL FILL_1__10403_ (
);

FILL FILL_2__7848_ (
);

FILL FILL_0__7830_ (
);

FILL FILL_2__7428_ (
);

FILL FILL_1__13295_ (
);

INVX1 _12993_ (
    .A(_2_[14]),
    .Y(_3647_)
);

INVX1 _12573_ (
    .A(\datapath_1.Data [2]),
    .Y(_3428_)
);

FILL FILL_0__12288_ (
);

OAI21X1 _12153_ (
    .A(_3154_),
    .B(ALUSrcA_bF$buf2),
    .C(_3155_),
    .Y(\datapath_1.alu_1.ALUInA [12])
);

FILL FILL_3__13622_ (
);

FILL FILL_4__8715_ (
);

FILL FILL_2__12615_ (
);

FILL FILL_3__16094_ (
);

FILL FILL_5__10195_ (
);

FILL FILL_1__11608_ (
);

FILL FILL_2__15087_ (
);

FILL FILL_5__16001_ (
);

FILL FILL_0__8615_ (
);

FILL FILL_4__15834_ (
);

FILL FILL_4__15414_ (
);

OAI22X1 _13778_ (
    .A(_4283_),
    .B(_3935__bF$buf3),
    .C(_3924__bF$buf3),
    .D(_4282_),
    .Y(_4284_)
);

NAND2X1 _13358_ (
    .A(RegWrite_bF$buf0),
    .B(_3873_),
    .Y(_3874_)
);

FILL FILL_3__14827_ (
);

FILL FILL_3__14407_ (
);

FILL FILL_1__15861_ (
);

FILL FILL_1__15441_ (
);

FILL FILL112040x67050 (
);

FILL FILL_1__15021_ (
);

FILL FILL_0__14854_ (
);

FILL FILL_0__14434_ (
);

FILL FILL_0__14014_ (
);

BUFX2 BUFX2_insert900 (
    .A(_5552_),
    .Y(_5552__bF$buf2)
);

FILL SFILL68920x60050 (
);

FILL FILL_2__7181_ (
);

BUFX2 BUFX2_insert901 (
    .A(_5552_),
    .Y(_5552__bF$buf1)
);

BUFX2 BUFX2_insert902 (
    .A(_5552_),
    .Y(_5552__bF$buf0)
);

BUFX2 BUFX2_insert903 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf7)
);

BUFX2 BUFX2_insert904 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf6)
);

BUFX2 BUFX2_insert905 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf5)
);

BUFX2 BUFX2_insert906 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf4)
);

BUFX2 BUFX2_insert907 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf3)
);

BUFX2 BUFX2_insert908 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf2)
);

BUFX2 BUFX2_insert909 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf1)
);

FILL FILL_5__12761_ (
);

FILL FILL_5__12341_ (
);

FILL FILL112440x36050 (
);

FILL FILL_4__11754_ (
);

FILL FILL_4__11334_ (
);

FILL FILL_1__16226_ (
);

FILL FILL_3__10747_ (
);

FILL FILL_1__11781_ (
);

FILL FILL_1__11361_ (
);

FILL FILL112040x22050 (
);

OAI22X1 _15924_ (
    .A(_4956_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf2),
    .D(_4953_),
    .Y(_6383_)
);

FILL FILL_0__15639_ (
);

FILL FILL_0__15219_ (
);

NAND3X1 _15504_ (
    .A(_5970_),
    .B(_5972_),
    .C(_5969_),
    .Y(_5973_)
);

FILL FILL_0__10774_ (
);

FILL FILL_2__8386_ (
);

FILL FILL_6__14973_ (
);

FILL FILL_5__13966_ (
);

FILL FILL_5__13546_ (
);

FILL FILL_3__14580_ (
);

FILL FILL_5__13126_ (
);

INVX1 _7846_ (
    .A(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_489_)
);

FILL FILL_3__14160_ (
);

INVX1 _7426_ (
    .A(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_270_)
);

DFFSR _7006_ (
    .Q(\datapath_1.regfile_1.regOut[1] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_3_[8])
);

FILL FILL_4_BUFX2_insert740 (
);

FILL FILL_4_BUFX2_insert741 (
);

FILL FILL_4__9673_ (
);

FILL FILL_4__9253_ (
);

FILL FILL_4_BUFX2_insert742 (
);

FILL FILL_4__12959_ (
);

FILL FILL_2__13993_ (
);

FILL FILL_4_BUFX2_insert743 (
);

FILL FILL_4_BUFX2_insert744 (
);

FILL FILL_4__12119_ (
);

FILL FILL_2__13573_ (
);

FILL FILL_2__13153_ (
);

FILL FILL_4_BUFX2_insert745 (
);

FILL FILL_4_BUFX2_insert746 (
);

FILL FILL_4_BUFX2_insert747 (
);

FILL FILL_4_BUFX2_insert748 (
);

FILL FILL_4_BUFX2_insert749 (
);

FILL FILL_1__12986_ (
);

FILL FILL_1__12146_ (
);

FILL FILL_4__13900_ (
);

FILL FILL_0__9993_ (
);

FILL FILL_3__7670_ (
);

FILL FILL_0__11979_ (
);

OAI21X1 _11844_ (
    .A(_2931_),
    .B(gnd),
    .C(_2344__bF$buf0),
    .Y(_2932_)
);

FILL FILL_3__7250_ (
);

FILL FILL_0__11559_ (
);

FILL FILL_0__9153_ (
);

NOR2X1 _11424_ (
    .A(_2537_),
    .B(_2539_),
    .Y(_2540_)
);

FILL FILL_0__11139_ (
);

OR2X2 _11004_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2123_)
);

FILL FILL_5__7596_ (
);

FILL FILL_5__7176_ (
);

FILL FILL_4__16372_ (
);

FILL FILL_3__15785_ (
);

FILL FILL_3__15365_ (
);

FILL FILL_0__12500_ (
);

FILL FILL_1__7588_ (
);

FILL FILL_1__7168_ (
);

FILL FILL_2__14778_ (
);

FILL FILL_2__14358_ (
);

FILL FILL_0__15392_ (
);

FILL SFILL13640x2050 (
);

FILL SFILL23720x52050 (
);

FILL FILL_3__8875_ (
);

FILL FILL_3__8455_ (
);

OAI21X1 _12629_ (
    .A(_3464_),
    .B(vdd),
    .C(_3465_),
    .Y(_3425_[20])
);

NAND2X1 _12209_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [31]),
    .Y(_3193_)
);

FILL FILL_1__14712_ (
);

FILL SFILL94200x39050 (
);

FILL FILL_4__12292_ (
);

FILL FILL_0__13705_ (
);

FILL FILL_2__6872_ (
);

FILL FILL_5__9742_ (
);

FILL FILL_3__11285_ (
);

FILL FILL_0__16177_ (
);

OAI22X1 _16042_ (
    .A(_5549__bF$buf2),
    .B(_5123_),
    .C(_5466__bF$buf0),
    .D(_5120_),
    .Y(_6498_)
);

FILL FILL_2__10698_ (
);

FILL FILL_2__10278_ (
);

FILL FILL_1__9734_ (
);

FILL FILL_5__11612_ (
);

FILL SFILL8680x58050 (
);

FILL FILL_6__15091_ (
);

FILL FILL_3_BUFX2_insert760 (
);

FILL FILL_3_BUFX2_insert761 (
);

FILL SFILL109560x75050 (
);

FILL FILL_3_BUFX2_insert762 (
);

FILL FILL_3_BUFX2_insert763 (
);

FILL FILL_3_BUFX2_insert764 (
);

FILL FILL_5__14084_ (
);

FILL FILL_1__15917_ (
);

FILL FILL_3_BUFX2_insert765 (
);

FILL FILL_3_BUFX2_insert766 (
);

OAI21X1 _8384_ (
    .A(_765_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .C(_766_),
    .Y(_718_[24])
);

FILL FILL_3_BUFX2_insert767 (
);

FILL FILL_3_BUFX2_insert768 (
);

FILL FILL_3_BUFX2_insert769 (
);

FILL FILL_1__10632_ (
);

FILL FILL_4__13497_ (
);

FILL SFILL84280x39050 (
);

FILL FILL_2__7237_ (
);

FILL SFILL23640x14050 (
);

INVX1 _12382_ (
    .A(ALUOut[13]),
    .Y(_3320_)
);

FILL FILL_0__12097_ (
);

FILL FILL_3__13851_ (
);

FILL SFILL8600x56050 (
);

FILL FILL_3__13431_ (
);

FILL FILL_3__13011_ (
);

FILL FILL_4__8524_ (
);

FILL FILL_4__8104_ (
);

FILL SFILL8680x13050 (
);

FILL FILL_2__12844_ (
);

FILL SFILL13720x50050 (
);

FILL FILL_2__12424_ (
);

FILL FILL_5__15289_ (
);

FILL FILL_2__12004_ (
);

DFFSR _9589_ (
    .Q(\datapath_1.regfile_1.regOut[21] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1303_[31])
);

NAND2X1 _9169_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1168_)
);

FILL FILL_1__11837_ (
);

FILL FILL_1__11417_ (
);

FILL SFILL84200x37050 (
);

FILL FILL_0__8844_ (
);

FILL FILL_5__16230_ (
);

FILL FILL_3__6941_ (
);

FILL FILL_0__8004_ (
);

FILL FILL_5__6867_ (
);

FILL FILL_0_BUFX2_insert890 (
);

FILL FILL_0_BUFX2_insert891 (
);

FILL FILL_4__15643_ (
);

FILL FILL_0_BUFX2_insert892 (
);

FILL FILL_4__15223_ (
);

FILL FILL_0_BUFX2_insert893 (
);

FILL FILL_0_BUFX2_insert894 (
);

FILL SFILL13640x57050 (
);

OAI22X1 _13587_ (
    .A(_3947__bF$buf1),
    .B(_4095_),
    .C(_3909_),
    .D(_4094_),
    .Y(_4096_)
);

FILL FILL_0_BUFX2_insert895 (
);

NAND2X1 _13167_ (
    .A(PCEn_bF$buf6),
    .B(\datapath_1.mux_pcsrc.dout [29]),
    .Y(_3743_)
);

FILL FILL_0_BUFX2_insert896 (
);

FILL FILL_0_BUFX2_insert897 (
);

FILL FILL_2__9803_ (
);

FILL FILL_3__14636_ (
);

FILL FILL_0_BUFX2_insert898 (
);

FILL SFILL109480x37050 (
);

FILL FILL_1__15670_ (
);

FILL FILL_3__14216_ (
);

FILL FILL_0_BUFX2_insert899 (
);

FILL FILL_1__15250_ (
);

FILL FILL_1__6859_ (
);

FILL FILL_4__9729_ (
);

FILL SFILL8600x11050 (
);

FILL FILL_2__13629_ (
);

FILL SFILL19320x78050 (
);

FILL FILL_2__13209_ (
);

FILL FILL_0__14663_ (
);

FILL FILL_0__14243_ (
);

FILL FILL_1__7800_ (
);

FILL FILL_3__7726_ (
);

FILL FILL_0__9629_ (
);

FILL FILL_3__7306_ (
);

FILL FILL_0__9209_ (
);

FILL FILL_5__12990_ (
);

FILL FILL_5__12570_ (
);

FILL SFILL74280x37050 (
);

FILL FILL_5__12150_ (
);

BUFX2 _6870_ (
    .A(_2_[0]),
    .Y(memoryWriteData[0])
);

FILL FILL_4__16008_ (
);

FILL FILL_4__11983_ (
);

FILL FILL_4__11563_ (
);

FILL FILL_6__10109_ (
);

FILL FILL_4__11143_ (
);

FILL SFILL13640x12050 (
);

FILL FILL_1__16035_ (
);

FILL FILL_3__10976_ (
);

FILL FILL_6_BUFX2_insert270 (
);

FILL FILL_3__10556_ (
);

FILL FILL_3__10136_ (
);

FILL FILL_1__11590_ (
);

FILL FILL_1__11170_ (
);

FILL FILL_0__15868_ (
);

AOI22X1 _15733_ (
    .A(_5557_),
    .B(\datapath_1.regfile_1.regOut[17] [17]),
    .C(\datapath_1.regfile_1.regOut[18] [17]),
    .D(_5558_),
    .Y(_6196_)
);

FILL FILL_0__15448_ (
);

NOR3X1 _15313_ (
    .A(_4259_),
    .B(_5459__bF$buf0),
    .C(_5519_),
    .Y(_5787_)
);

FILL FILL_0__15028_ (
);

FILL FILL_6_BUFX2_insert275 (
);

FILL SFILL38840x61050 (
);

FILL FILL_2__8195_ (
);

FILL FILL_0__10163_ (
);

BUFX2 BUFX2_insert50 (
    .A(_3893_),
    .Y(_3893__bF$buf0)
);

BUFX2 BUFX2_insert51 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf7 )
);

BUFX2 BUFX2_insert52 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf6 )
);

BUFX2 BUFX2_insert53 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf5 )
);

BUFX2 BUFX2_insert54 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf4 )
);

BUFX2 BUFX2_insert55 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf3 )
);

BUFX2 BUFX2_insert56 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf2 )
);

BUFX2 BUFX2_insert57 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf1 )
);

FILL FILL_2__10910_ (
);

FILL FILL_5__13775_ (
);

FILL SFILL74200x35050 (
);

FILL FILL_5__13355_ (
);

BUFX2 BUFX2_insert58 (
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf0 )
);

FILL SFILL13560x19050 (
);

BUFX2 BUFX2_insert59 (
    .A(_5463_),
    .Y(_5463__bF$buf3)
);

DFFSR _7655_ (
    .Q(\datapath_1.regfile_1.regOut[6] [17]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_328_[17])
);

OAI21X1 _7235_ (
    .A(_182_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_183_),
    .Y(_133_[25])
);

FILL FILL_4__9482_ (
);

FILL FILL_4__12768_ (
);

FILL FILL_4__12348_ (
);

FILL FILL_2__13382_ (
);

FILL FILL_2__6928_ (
);

FILL FILL_0__6910_ (
);

FILL FILL_1__12375_ (
);

FILL SFILL99480x41050 (
);

FILL FILL_0__9382_ (
);

FILL FILL_0__11788_ (
);

FILL FILL_0__11368_ (
);

INVX1 _11653_ (
    .A(_2395_),
    .Y(_2756_)
);

NOR2X1 _11233_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2352_)
);

FILL FILL_3__12702_ (
);

FILL FILL_6__15567_ (
);

FILL SFILL104440x18050 (
);

FILL FILL_6__15147_ (
);

FILL FILL_4__16181_ (
);

FILL SFILL64200x78050 (
);

FILL FILL_3__15594_ (
);

FILL FILL_3__15174_ (
);

FILL FILL112120x55050 (
);

FILL FILL_2__14587_ (
);

FILL FILL_2__14167_ (
);

FILL FILL_5__15921_ (
);

FILL FILL_5__15501_ (
);

OAI21X1 _9801_ (
    .A(_1486_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .C(_1487_),
    .Y(_1433_[27])
);

FILL FILL_4__14914_ (
);

OAI21X1 _12858_ (
    .A(_3576_),
    .B(vdd),
    .C(_3577_),
    .Y(_3555_[11])
);

FILL FILL_3__8264_ (
);

OAI21X1 _12438_ (
    .A(_3356_),
    .B(MemToReg_bF$buf6),
    .C(_3357_),
    .Y(\datapath_1.mux_wd3.dout [31])
);

NAND3X1 _12018_ (
    .A(_3057_),
    .B(_3058_),
    .C(_3059_),
    .Y(\datapath_1.mux_pcsrc.dout [7])
);

FILL FILL_3__13907_ (
);

FILL FILL_1__14941_ (
);

FILL FILL_1__14521_ (
);

FILL FILL_1__14101_ (
);

FILL FILL_6__11487_ (
);

FILL FILL_5_BUFX2_insert290 (
);

FILL FILL_6__11067_ (
);

FILL FILL_5_BUFX2_insert291 (
);

FILL FILL_5_BUFX2_insert292 (
);

FILL FILL_0__13934_ (
);

FILL FILL_3__16379_ (
);

FILL FILL_0__13514_ (
);

FILL FILL_5_BUFX2_insert293 (
);

FILL FILL_5_BUFX2_insert294 (
);

FILL FILL_5_BUFX2_insert295 (
);

FILL FILL_5_BUFX2_insert296 (
);

FILL SFILL33800x42050 (
);

FILL FILL_5__9551_ (
);

FILL FILL_5_BUFX2_insert297 (
);

FILL SFILL64200x33050 (
);

FILL FILL_5__9131_ (
);

FILL FILL_5_BUFX2_insert298 (
);

FILL FILL_3__11094_ (
);

FILL FILL_5_BUFX2_insert299 (
);

FILL FILL_5_BUFX2_insert1084 (
);

FILL FILL112120x10050 (
);

FILL FILL_5_BUFX2_insert1085 (
);

OAI22X1 _16271_ (
    .A(_6720_),
    .B(_5518__bF$buf3),
    .C(_5478__bF$buf3),
    .D(_6719_),
    .Y(_6721_)
);

FILL FILL_5_BUFX2_insert1086 (
);

FILL FILL_5_BUFX2_insert1087 (
);

FILL FILL_5_BUFX2_insert1088 (
);

FILL FILL_5_BUFX2_insert1089 (
);

FILL FILL_5__11841_ (
);

FILL FILL_1__9543_ (
);

FILL FILL_5__11421_ (
);

FILL FILL_1__9123_ (
);

FILL FILL_5__11001_ (
);

FILL FILL_3__9889_ (
);

FILL FILL_2__16313_ (
);

FILL FILL_3__9469_ (
);

FILL FILL_4__10834_ (
);

FILL FILL_4__10414_ (
);

FILL FILL_1__15726_ (
);

OAI21X1 _8193_ (
    .A(_658_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .C(_659_),
    .Y(_653_[3])
);

FILL FILL_1__15306_ (
);

FILL SFILL113960x44050 (
);

FILL FILL_1__10441_ (
);

FILL FILL_1__10021_ (
);

FILL FILL_0__14719_ (
);

FILL FILL_2__7886_ (
);

FILL FILL_2__7466_ (
);

FILL FILL_3__12299_ (
);

FILL FILL_2__7046_ (
);

FILL FILL_6__13633_ (
);

NAND2X1 _12191_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.a [25]),
    .Y(_3181_)
);

FILL FILL_5__12626_ (
);

FILL FILL_3__13660_ (
);

FILL FILL_5__12206_ (
);

FILL FILL_3__13240_ (
);

INVX1 _6926_ (
    .A(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_18_)
);

FILL FILL_4__8753_ (
);

FILL FILL_4__8333_ (
);

FILL FILL_4__11619_ (
);

FILL FILL_2__12653_ (
);

FILL FILL_5__15098_ (
);

FILL FILL_2__12233_ (
);

NAND2X1 _9398_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1280_)
);

FILL FILL_1__11646_ (
);

FILL FILL_1__11226_ (
);

FILL FILL_0__8653_ (
);

FILL FILL_0__10639_ (
);

NOR2X1 _10924_ (
    .A(_2060_),
    .B(_2057_),
    .Y(_2062_)
);

FILL FILL_0__8233_ (
);

INVX1 _10504_ (
    .A(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_1834_)
);

FILL FILL_4__15872_ (
);

FILL FILL_4__15452_ (
);

FILL FILL_4__15032_ (
);

INVX1 _13396_ (
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_3908_)
);

FILL FILL_2__9612_ (
);

FILL FILL_3__14865_ (
);

FILL FILL_3__14445_ (
);

FILL FILL_3__14025_ (
);

FILL FILL_4__9538_ (
);

FILL FILL_4__9118_ (
);

FILL FILL_2__13858_ (
);

FILL FILL_2__13438_ (
);

FILL FILL_0__14892_ (
);

FILL FILL_0__14472_ (
);

FILL FILL_2__13018_ (
);

FILL FILL_0__14052_ (
);

FILL SFILL23720x47050 (
);

FILL FILL_0__9858_ (
);

FILL FILL_3__7955_ (
);

FILL FILL_3__7115_ (
);

FILL FILL_0__9018_ (
);

AOI22X1 _11709_ (
    .A(_2392_),
    .B(_2481__bF$buf3),
    .C(_2478_),
    .D(_2171_),
    .Y(_2808_)
);

FILL FILL_4__16237_ (
);

FILL FILL_4__11792_ (
);

FILL FILL_4__11372_ (
);

FILL SFILL23320x33050 (
);

FILL FILL_1__16264_ (
);

FILL FILL_5__8822_ (
);

FILL FILL_3__10785_ (
);

FILL FILL_5__8402_ (
);

FILL FILL_3__10365_ (
);

FILL FILL_0__15677_ (
);

INVX1 _15962_ (
    .A(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_6420_)
);

FILL FILL_0__15257_ (
);

NAND3X1 _15542_ (
    .A(_6005_),
    .B(_6006_),
    .C(_6009_),
    .Y(_6010_)
);

INVX1 _15122_ (
    .A(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_5601_)
);

FILL FILL_0__10392_ (
);

FILL FILL_5__13584_ (
);

FILL FILL_5__13164_ (
);

OAI21X1 _7884_ (
    .A(_513_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_514_),
    .Y(_458_[28])
);

OAI21X1 _7464_ (
    .A(_294_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_295_),
    .Y(_263_[16])
);

OAI21X1 _7044_ (
    .A(_75_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .C(_76_),
    .Y(_68_[4])
);

FILL FILL_4__12997_ (
);

FILL FILL_4__9291_ (
);

FILL FILL_4__12577_ (
);

FILL FILL_4__12157_ (
);

FILL FILL_5__9607_ (
);

FILL FILL_1__12184_ (
);

INVX1 _16327_ (
    .A(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_6772_)
);

NAND2X1 _11882_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [16]),
    .Y(_2965_)
);

FILL FILL_0__11597_ (
);

FILL FILL_0__11177_ (
);

INVX1 _11462_ (
    .A(_2302_),
    .Y(_2577_)
);

XOR2X1 _11042_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2161_)
);

FILL FILL_3__12511_ (
);

FILL FILL_4__7604_ (
);

FILL SFILL13720x45050 (
);

FILL FILL_2__11924_ (
);

FILL FILL_5__14789_ (
);

FILL FILL_5__14369_ (
);

FILL FILL_2__11504_ (
);

DFFSR _8669_ (
    .Q(\datapath_1.regfile_1.regOut[14] [7]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_848_[7])
);

NAND2X1 _8249_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_697_)
);

FILL FILL_1__10917_ (
);

FILL SFILL64200x50 (
);

FILL FILL_2__14396_ (
);

FILL FILL_5__15730_ (
);

FILL FILL_5__15310_ (
);

FILL FILL_0__7504_ (
);

OAI21X1 _9610_ (
    .A(_1379_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .C(_1380_),
    .Y(_1368_[6])
);

FILL FILL_1__13389_ (
);

FILL FILL_4__14723_ (
);

FILL FILL_4__14303_ (
);

FILL FILL_3__8493_ (
);

DFFSR _12667_ (
    .Q(\datapath_1.Data [4]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[4])
);

FILL FILL_3__8073_ (
);

NAND3X1 _12247_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3224_)
);

FILL FILL_3__13716_ (
);

FILL FILL_1__14750_ (
);

FILL FILL_1__14330_ (
);

FILL FILL_2__12709_ (
);

FILL FILL_0__13743_ (
);

FILL FILL_0__13323_ (
);

FILL FILL_3__16188_ (
);

FILL FILL_5__10289_ (
);

FILL FILL_5__9780_ (
);

FILL FILL_5__9360_ (
);

NOR2X1 _16080_ (
    .A(_6534_),
    .B(_6533_),
    .Y(_6535_)
);

FILL FILL_0__8709_ (
);

FILL FILL_1__9772_ (
);

FILL FILL_5__11650_ (
);

FILL FILL_1__9352_ (
);

FILL FILL_5__11230_ (
);

FILL FILL_4__15928_ (
);

FILL FILL_4__15508_ (
);

FILL FILL_2__16122_ (
);

FILL FILL_3__9278_ (
);

FILL FILL_4__10643_ (
);

FILL FILL_1__15955_ (
);

FILL FILL_1__15535_ (
);

FILL FILL_1__15115_ (
);

FILL FILL_1__10670_ (
);

FILL FILL_1__10250_ (
);

FILL FILL_0__14948_ (
);

INVX1 _14813_ (
    .A(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_5297_)
);

FILL FILL_0__14528_ (
);

FILL FILL_0__14108_ (
);

FILL SFILL38840x56050 (
);

FILL FILL_2__7695_ (
);

FILL FILL_6__13022_ (
);

FILL FILL_5__12855_ (
);

FILL FILL_5__12435_ (
);

FILL FILL_5__12015_ (
);

FILL FILL_4__8982_ (
);

FILL FILL_4__8142_ (
);

FILL FILL_4__11848_ (
);

FILL FILL_2__12882_ (
);

FILL FILL_4__11428_ (
);

FILL FILL_2__12462_ (
);

FILL FILL_4__11008_ (
);

FILL FILL_2__12042_ (
);

FILL SFILL43400x25050 (
);

FILL FILL112200x43050 (
);

FILL FILL_1__11875_ (
);

FILL SFILL99480x36050 (
);

FILL FILL_1__11455_ (
);

FILL FILL_1__11035_ (
);

FILL FILL_0__8882_ (
);

FILL FILL_0__8462_ (
);

FILL SFILL3480x55050 (
);

DFFSR _10733_ (
    .Q(\datapath_1.regfile_1.regOut[30] [23]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1888_[23])
);

FILL FILL_0__10448_ (
);

FILL FILL_0__10028_ (
);

OAI21X1 _10313_ (
    .A(_1746_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1747_),
    .Y(_1693_[27])
);

FILL SFILL38840x11050 (
);

FILL FILL_4__15681_ (
);

FILL FILL_6__14227_ (
);

FILL FILL_4__15261_ (
);

FILL FILL_2__9421_ (
);

FILL FILL_3__14674_ (
);

FILL FILL_3__14254_ (
);

FILL FILL_2__9001_ (
);

FILL FILL_1__6897_ (
);

FILL FILL_4__9767_ (
);

FILL FILL_4__9347_ (
);

FILL FILL_2__13667_ (
);

FILL FILL_2__13247_ (
);

FILL FILL_0__14281_ (
);

FILL SFILL89480x79050 (
);

FILL SFILL64840x4050 (
);

FILL FILL_3__7764_ (
);

FILL FILL_0__9667_ (
);

INVX1 _11938_ (
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3000_)
);

FILL FILL_3__7344_ (
);

FILL FILL_0__9247_ (
);

INVX1 _11518_ (
    .A(_2237_),
    .Y(_2629_)
);

FILL SFILL28840x54050 (
);

FILL FILL_1__13601_ (
);

FILL FILL_4__16046_ (
);

FILL SFILL89080x65050 (
);

FILL FILL_4__11181_ (
);

FILL FILL_3__15879_ (
);

FILL FILL_3__15459_ (
);

FILL FILL_3__15039_ (
);

FILL FILL_1__16073_ (
);

FILL SFILL33800x37050 (
);

FILL SFILL64200x28050 (
);

FILL FILL_5__8631_ (
);

FILL FILL_3__10174_ (
);

FILL FILL_5__8211_ (
);

FILL FILL_6_BUFX2_insert654 (
);

AOI22X1 _15771_ (
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_6233_)
);

FILL FILL_0__15486_ (
);

OAI22X1 _15351_ (
    .A(_5526__bF$buf0),
    .B(_4333_),
    .C(_4317_),
    .D(_5527__bF$buf0),
    .Y(_5824_)
);

FILL FILL_0__15066_ (
);

FILL FILL_3__16400_ (
);

FILL FILL_6_BUFX2_insert659 (
);

FILL FILL_5__10921_ (
);

FILL FILL_1__8623_ (
);

FILL FILL_5__10501_ (
);

FILL FILL_1__8203_ (
);

FILL FILL_2__15813_ (
);

FILL FILL_3__8969_ (
);

FILL FILL_3__8129_ (
);

FILL FILL_5__13393_ (
);

OAI21X1 _7693_ (
    .A(_406_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_407_),
    .Y(_393_[7])
);

FILL FILL_1__14806_ (
);

DFFSR _7273_ (
    .Q(\datapath_1.regfile_1.regOut[3] [19]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_133_[19])
);

FILL SFILL113960x39050 (
);

FILL FILL_4__12386_ (
);

FILL FILL_3__9910_ (
);

FILL FILL_2__6966_ (
);

FILL SFILL89080x20050 (
);

FILL FILL_3__11799_ (
);

FILL FILL_5__9416_ (
);

FILL FILL_3__11379_ (
);

INVX1 _16136_ (
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_6589_)
);

OAI21X1 _11691_ (
    .A(_2764_),
    .B(_2165_),
    .C(_2462__bF$buf3),
    .Y(_2791_)
);

AOI21X1 _11271_ (
    .A(_2387_),
    .B(_2389_),
    .C(_2385_),
    .Y(_2390_)
);

FILL FILL_5__11706_ (
);

FILL FILL_3__12740_ (
);

FILL FILL_1__9408_ (
);

FILL FILL_3__12320_ (
);

FILL FILL_4__7833_ (
);

FILL FILL_5__14598_ (
);

FILL FILL_2__11733_ (
);

FILL FILL_5__14178_ (
);

FILL FILL_2__11313_ (
);

NAND2X1 _8898_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1028_)
);

NAND2X1 _8478_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_809_)
);

NAND2X1 _8058_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_590_)
);

FILL FILL_1__10306_ (
);

FILL FILL_0__7733_ (
);

FILL FILL_0__7313_ (
);

FILL FILL_4__14952_ (
);

FILL FILL_4__14532_ (
);

FILL SFILL54200x26050 (
);

FILL FILL_4__14112_ (
);

NAND2X1 _12896_ (
    .A(vdd),
    .B(\datapath_1.rd1 [24]),
    .Y(_3603_)
);

NAND2X1 _12476_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [12]),
    .Y(_3384_)
);

NAND3X1 _12056_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3034__bF$buf1),
    .Y(_3088_)
);

FILL FILL_3__13945_ (
);

FILL FILL_3__13525_ (
);

FILL FILL_3__13105_ (
);

FILL FILL_4__8618_ (
);

FILL FILL_5_BUFX2_insert670 (
);

FILL FILL_5_BUFX2_insert671 (
);

FILL FILL_5_BUFX2_insert672 (
);

FILL FILL_2__12518_ (
);

FILL FILL_0__13972_ (
);

FILL FILL_5_BUFX2_insert673 (
);

FILL FILL_0__13552_ (
);

FILL FILL_5_BUFX2_insert674 (
);

FILL FILL_0__13132_ (
);

FILL FILL_5_BUFX2_insert675 (
);

FILL FILL_5_BUFX2_insert676 (
);

FILL FILL_5_BUFX2_insert677 (
);

FILL FILL_5_BUFX2_insert678 (
);

FILL FILL_5_BUFX2_insert679 (
);

FILL FILL_5__16324_ (
);

FILL FILL_0__8518_ (
);

FILL FILL_1__9161_ (
);

FILL FILL_4__15737_ (
);

FILL FILL_4__15317_ (
);

FILL FILL_2__16351_ (
);

FILL FILL_3__9087_ (
);

FILL FILL_4__10872_ (
);

FILL FILL_4__10452_ (
);

FILL FILL_4__10032_ (
);

FILL FILL_1__15764_ (
);

FILL FILL_1__15344_ (
);

FILL FILL_0__14757_ (
);

INVX1 _14622_ (
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_5110_)
);

FILL FILL_0__14337_ (
);

INVX1 _14202_ (
    .A(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_4699_)
);

FILL FILL_2__7084_ (
);

FILL FILL_5__12244_ (
);

OAI21X1 _6964_ (
    .A(_42_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_43_),
    .Y(_3_[20])
);

FILL FILL_4__8371_ (
);

FILL FILL_4__11657_ (
);

FILL SFILL48920x46050 (
);

FILL SFILL99320x1050 (
);

FILL FILL_4__11237_ (
);

FILL FILL_2__12271_ (
);

FILL FILL_1__16129_ (
);

FILL FILL_1__11684_ (
);

FILL FILL_1__11264_ (
);

NOR3X1 _15827_ (
    .A(_5515__bF$buf3),
    .B(_6287_),
    .C(_5521__bF$buf3),
    .Y(_6288_)
);

OAI22X1 _15407_ (
    .A(_5878_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf1),
    .D(_4371_),
    .Y(_5879_)
);

FILL FILL_0__10677_ (
);

NAND2X1 _10962_ (
    .A(_2063_),
    .B(_2093_),
    .Y(_2094_)
);

FILL FILL_0__8271_ (
);

OAI21X1 _10542_ (
    .A(_1858_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1859_),
    .Y(_1823_[18])
);

FILL FILL_0__10257_ (
);

OAI21X1 _10122_ (
    .A(_1639_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1640_),
    .Y(_1628_[6])
);

FILL FILL_6__14876_ (
);

FILL FILL_4__15490_ (
);

FILL FILL_4__15070_ (
);

FILL FILL_5__13869_ (
);

FILL SFILL88600x28050 (
);

FILL FILL_5__13449_ (
);

FILL FILL_2__9650_ (
);

FILL FILL_2__9230_ (
);

FILL FILL_3__14483_ (
);

FILL FILL_5__13029_ (
);

FILL FILL_3__14063_ (
);

NAND2X1 _7749_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_445_)
);

NAND2X1 _7329_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_226_)
);

FILL FILL_4__9996_ (
);

FILL FILL_4__9156_ (
);

FILL SFILL109400x9050 (
);

FILL FILL_2__13896_ (
);

FILL FILL_2__13476_ (
);

FILL FILL_0__14090_ (
);

FILL FILL_5__14810_ (
);

FILL FILL_1__12889_ (
);

FILL FILL_1__12469_ (
);

FILL FILL_1__12049_ (
);

FILL FILL_4__13803_ (
);

FILL SFILL3640x81050 (
);

FILL FILL_0__9896_ (
);

FILL FILL_3__7993_ (
);

FILL FILL_0__9476_ (
);

FILL FILL_3__7573_ (
);

OAI21X1 _11747_ (
    .A(_2841_),
    .B(_2480_),
    .C(_2842_),
    .Y(_2843_)
);

AOI21X1 _11327_ (
    .A(_2300_),
    .B(_2296_),
    .C(_2294_),
    .Y(_2446_)
);

FILL FILL_1__13830_ (
);

FILL FILL_5__7499_ (
);

FILL FILL_5__7079_ (
);

FILL FILL_1__13410_ (
);

FILL FILL_4__16275_ (
);

FILL FILL_6__10796_ (
);

FILL FILL_3__15688_ (
);

FILL FILL_0__12823_ (
);

FILL FILL_0__12403_ (
);

FILL FILL_3__15268_ (
);

FILL FILL_5__8860_ (
);

FILL FILL_5__8440_ (
);

FILL FILL_5__8020_ (
);

FILL FILL_0__15295_ (
);

NAND3X1 _15580_ (
    .A(_6041_),
    .B(_6042_),
    .C(_6046_),
    .Y(_6047_)
);

NOR2X1 _15160_ (
    .A(_5637_),
    .B(_5635_),
    .Y(_5638_)
);

FILL SFILL38920x44050 (
);

FILL FILL_1__8852_ (
);

FILL FILL_5__10310_ (
);

FILL FILL_1__8012_ (
);

FILL FILL_2__15622_ (
);

FILL FILL_2__15202_ (
);

FILL FILL_3__8778_ (
);

FILL FILL_3__8358_ (
);

FILL FILL_1__14615_ (
);

NAND2X1 _7082_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_102_)
);

FILL FILL_4__12195_ (
);

FILL FILL_0__13608_ (
);

FILL FILL_5__9645_ (
);

FILL FILL_5__9225_ (
);

FILL FILL_3__11188_ (
);

OAI21X1 _16365_ (
    .A(_6796_),
    .B(gnd),
    .C(_6797_),
    .Y(_6769_[14])
);

FILL SFILL3560x43050 (
);

FILL FILL_5__11935_ (
);

INVX1 _11080_ (
    .A(_2198_),
    .Y(_2199_)
);

FILL FILL_1__9637_ (
);

FILL FILL_5__11515_ (
);

FILL FILL_1__9217_ (
);

FILL FILL_2__16407_ (
);

FILL FILL_4__7222_ (
);

FILL FILL_4__10928_ (
);

FILL FILL_4__10508_ (
);

FILL FILL_2__11962_ (
);

FILL FILL_2__11542_ (
);

FILL FILL_3_CLKBUF1_insert200 (
);

FILL FILL_2__11122_ (
);

FILL FILL_3_CLKBUF1_insert201 (
);

FILL FILL_3_CLKBUF1_insert202 (
);

DFFSR _8287_ (
    .Q(\datapath_1.regfile_1.regOut[11] [9]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_653_[9])
);

FILL FILL_3_CLKBUF1_insert203 (
);

FILL FILL112200x38050 (
);

FILL FILL_3_CLKBUF1_insert204 (
);

FILL SFILL83880x46050 (
);

FILL FILL_3_CLKBUF1_insert205 (
);

FILL FILL_1__10955_ (
);

FILL FILL_1__10535_ (
);

FILL FILL_3_CLKBUF1_insert206 (
);

FILL FILL_3_CLKBUF1_insert207 (
);

FILL FILL_1__10115_ (
);

FILL FILL_3_CLKBUF1_insert208 (
);

FILL FILL_3_CLKBUF1_insert209 (
);

FILL SFILL38040x23050 (
);

FILL FILL_0__7962_ (
);

FILL FILL_0__7542_ (
);

BUFX2 BUFX2_insert490 (
    .A(_3983_),
    .Y(_3983__bF$buf3)
);

FILL SFILL24600x34050 (
);

BUFX2 BUFX2_insert491 (
    .A(_3983_),
    .Y(_3983__bF$buf2)
);

FILL FILL_0__7122_ (
);

BUFX2 BUFX2_insert492 (
    .A(_3983_),
    .Y(_3983__bF$buf1)
);

BUFX2 BUFX2_insert493 (
    .A(_3983_),
    .Y(_3983__bF$buf0)
);

FILL SFILL73960x82050 (
);

BUFX2 BUFX2_insert494 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf113)
);

BUFX2 BUFX2_insert495 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf112)
);

FILL FILL_4__14761_ (
);

BUFX2 BUFX2_insert496 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf111)
);

FILL FILL_4__14341_ (
);

BUFX2 BUFX2_insert497 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf110)
);

FILL SFILL69240x5050 (
);

BUFX2 BUFX2_insert498 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf109)
);

BUFX2 BUFX2_insert499 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf108)
);

FILL SFILL43960x1050 (
);

AOI22X1 _12285_ (
    .A(_2_[17]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3253_)
);

FILL FILL_2__8501_ (
);

FILL FILL_3__13754_ (
);

FILL FILL_3__13334_ (
);

FILL FILL_4__8847_ (
);

FILL FILL_4__8007_ (
);

FILL FILL_2__12747_ (
);

FILL FILL_0__13781_ (
);

FILL FILL_2__12327_ (
);

FILL FILL_0__13361_ (
);

FILL FILL_3__6844_ (
);

FILL FILL_0__8747_ (
);

FILL FILL_5__16133_ (
);

FILL FILL_0__8327_ (
);

FILL FILL_1__9390_ (
);

FILL SFILL28840x49050 (
);

FILL FILL_4__15966_ (
);

FILL FILL_4__15546_ (
);

FILL FILL_4__15126_ (
);

FILL FILL_2__16160_ (
);

FILL FILL_4__10681_ (
);

FILL FILL_4__10261_ (
);

FILL FILL_3__14959_ (
);

FILL FILL_1__15993_ (
);

FILL FILL_3__14539_ (
);

FILL FILL_1__15573_ (
);

FILL FILL_3__14119_ (
);

FILL FILL_1__15153_ (
);

FILL FILL_5__7711_ (
);

FILL FILL_0__14986_ (
);

FILL FILL_0__14566_ (
);

INVX1 _14851_ (
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_5334_)
);

FILL FILL_0__14146_ (
);

INVX1 _14431_ (
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_4923_)
);

NOR2X1 _14011_ (
    .A(_4508_),
    .B(_4511_),
    .Y(_4512_)
);

FILL FILL_3__15900_ (
);

FILL FILL_1__7703_ (
);

FILL FILL_6__13480_ (
);

FILL FILL_3__7629_ (
);

FILL FILL_3__7209_ (
);

FILL FILL_5__12893_ (
);

FILL FILL_5__12473_ (
);

FILL FILL_5__12053_ (
);

FILL FILL_4__11886_ (
);

FILL SFILL63960x80050 (
);

FILL FILL_4__11466_ (
);

FILL SFILL94360x71050 (
);

FILL FILL_4__11046_ (
);

FILL FILL_2__12080_ (
);

FILL FILL_1__16358_ (
);

FILL FILL_3__10879_ (
);

FILL FILL_5__8916_ (
);

FILL FILL_3__10039_ (
);

FILL FILL_1__11493_ (
);

FILL FILL_1__11073_ (
);

NAND3X1 _15636_ (
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .B(_5471__bF$buf3),
    .C(_5531__bF$buf2),
    .Y(_6102_)
);

INVX4 _15216_ (
    .A(_5532__bF$buf0),
    .Y(_5692_)
);

FILL FILL_0__8080_ (
);

FILL FILL_0__10486_ (
);

FILL FILL_2__8098_ (
);

OAI21X1 _10771_ (
    .A(_1970_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .C(_1971_),
    .Y(_1953_[9])
);

FILL SFILL79160x51050 (
);

FILL FILL_0__10066_ (
);

DFFSR _10351_ (
    .Q(\datapath_1.regfile_1.regOut[27] [25]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_1693_[25])
);

FILL FILL_1__8908_ (
);

FILL FILL_3__11820_ (
);

FILL FILL_3__11400_ (
);

FILL FILL_4__6913_ (
);

FILL FILL_2__10813_ (
);

FILL FILL_5__13678_ (
);

FILL FILL_5__13258_ (
);

FILL FILL_3__14292_ (
);

NAND2X1 _7978_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_557_)
);

NAND2X1 _7558_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_338_)
);

DFFSR _7138_ (
    .Q(\datapath_1.regfile_1.regOut[2] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_68_[12])
);

FILL FILL_4__9385_ (
);

FILL SFILL18840x47050 (
);

FILL FILL_2__13285_ (
);

FILL SFILL79080x58050 (
);

FILL FILL_1__12698_ (
);

FILL FILL_1__12278_ (
);

FILL FILL_4__13612_ (
);

OAI21X1 _11976_ (
    .A(_3024_),
    .B(IorD_bF$buf2),
    .C(_3025_),
    .Y(_1_[29])
);

FILL FILL_0__9285_ (
);

AOI21X1 _11556_ (
    .A(_2229_),
    .B(_2481__bF$buf2),
    .C(_2664_),
    .Y(_2665_)
);

FILL SFILL79880x3050 (
);

INVX1 _11136_ (
    .A(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2255_)
);

FILL FILL_3__12605_ (
);

FILL FILL_4__16084_ (
);

FILL FILL111720x62050 (
);

FILL FILL_0__12632_ (
);

FILL FILL_3__15497_ (
);

FILL SFILL79480x27050 (
);

FILL FILL_3__15077_ (
);

FILL FILL_0__12212_ (
);

FILL FILL_6__16411_ (
);

FILL SFILL38920x7050 (
);

FILL FILL_5__15824_ (
);

FILL FILL_5__15404_ (
);

DFFSR _9704_ (
    .Q(\datapath_1.regfile_1.regOut[22] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_1368_[18])
);

FILL FILL_1__8661_ (
);

FILL FILL_1__8241_ (
);

FILL SFILL79080x13050 (
);

FILL FILL_4__14817_ (
);

FILL FILL_2__15851_ (
);

FILL FILL_2__15431_ (
);

FILL FILL_3__8587_ (
);

FILL FILL_2__15011_ (
);

FILL FILL_1__14844_ (
);

FILL FILL_1__14424_ (
);

FILL FILL_1__14004_ (
);

FILL FILL_0__13837_ (
);

FILL FILL_0__13417_ (
);

INVX1 _13702_ (
    .A(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_4209_)
);

FILL FILL_5__9874_ (
);

FILL FILL_5__9034_ (
);

FILL FILL_6__12331_ (
);

OAI22X1 _16174_ (
    .A(_6625_),
    .B(_5518__bF$buf2),
    .C(_5548__bF$buf2),
    .D(_5309_),
    .Y(_6626_)
);

FILL FILL_1__9866_ (
);

FILL FILL_5__11744_ (
);

FILL FILL_5__11324_ (
);

FILL FILL_1__9026_ (
);

FILL FILL_4__7871_ (
);

FILL FILL_2__16216_ (
);

FILL FILL_4__7451_ (
);

FILL FILL_4__7031_ (
);

FILL FILL_4__10317_ (
);

FILL FILL_2__11771_ (
);

FILL FILL_2__11351_ (
);

FILL FILL_1__15629_ (
);

INVX1 _8096_ (
    .A(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_615_)
);

FILL FILL_1__15209_ (
);

FILL FILL_1__10764_ (
);

NOR2X1 _14907_ (
    .A(_5388_),
    .B(_5373_),
    .Y(_5389_)
);

FILL FILL_0__7351_ (
);

FILL FILL_2__7369_ (
);

FILL SFILL114520x50050 (
);

FILL FILL_4__14990_ (
);

FILL FILL_6__13536_ (
);

FILL FILL_4__14570_ (
);

FILL FILL_4__14150_ (
);

NAND3X1 _12094_ (
    .A(_3114_),
    .B(_3115_),
    .C(_3116_),
    .Y(\datapath_1.mux_pcsrc.dout [26])
);

FILL FILL_3__13983_ (
);

FILL FILL_2__8730_ (
);

FILL FILL_5__12529_ (
);

FILL FILL_2__8310_ (
);

FILL FILL_5__12109_ (
);

FILL FILL_3__13563_ (
);

FILL FILL_3__13143_ (
);

FILL FILL_4__8656_ (
);

FILL FILL_4__8236_ (
);

FILL FILL_2__12976_ (
);

FILL SFILL69080x11050 (
);

FILL FILL_0__13590_ (
);

FILL FILL_2__12136_ (
);

FILL FILL_0__13170_ (
);

FILL FILL_1__11969_ (
);

FILL FILL_1__11549_ (
);

FILL FILL_1__11129_ (
);

FILL SFILL3640x76050 (
);

FILL FILL_0__8976_ (
);

FILL FILL_5__16362_ (
);

NAND2X1 _10827_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_2009_)
);

FILL FILL_0__8136_ (
);

NAND2X1 _10407_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1790_)
);

FILL SFILL43880x83050 (
);

FILL FILL_1__12910_ (
);

FILL FILL_4__15775_ (
);

FILL FILL_4__15355_ (
);

INVX2 _13299_ (
    .A(_3834_),
    .Y(_3835_)
);

FILL FILL_4__10490_ (
);

FILL FILL_2__9935_ (
);

FILL FILL_0__11903_ (
);

FILL FILL_3__14768_ (
);

FILL FILL_2__9515_ (
);

FILL FILL_3__14348_ (
);

FILL FILL_1__15382_ (
);

FILL FILL_5__7940_ (
);

FILL FILL_5__7100_ (
);

FILL FILL_0__14795_ (
);

FILL FILL_0__14375_ (
);

INVX1 _14660_ (
    .A(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_5147_)
);

OAI22X1 _14240_ (
    .A(_4734_),
    .B(_3955__bF$buf3),
    .C(_3924__bF$buf0),
    .D(_4735_),
    .Y(_4736_)
);

FILL SFILL38920x39050 (
);

FILL FILL_1__7932_ (
);

FILL FILL_2__14702_ (
);

FILL FILL_3__7858_ (
);

FILL FILL_3__7438_ (
);

FILL SFILL3640x31050 (
);

FILL FILL_5__12282_ (
);

FILL FILL_4__11695_ (
);

FILL FILL_4__11275_ (
);

FILL FILL_1__16167_ (
);

FILL FILL_3__10688_ (
);

FILL FILL_5__8725_ (
);

FILL FILL_3__10268_ (
);

FILL SFILL99560x19050 (
);

NAND3X1 _15865_ (
    .A(_6322_),
    .B(_6323_),
    .C(_6324_),
    .Y(_6325_)
);

OAI22X1 _15445_ (
    .A(_4404_),
    .B(_5548__bF$buf1),
    .C(_5489__bF$buf0),
    .D(_4417_),
    .Y(_5916_)
);

OAI22X1 _15025_ (
    .A(_3907_),
    .B(_5503__bF$buf1),
    .C(_5504__bF$buf4),
    .D(_3981_),
    .Y(_5505_)
);

FILL SFILL3560x38050 (
);

FILL FILL_0__10295_ (
);

NAND2X1 _10580_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1885_)
);

NAND2X1 _10160_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1666_)
);

FILL FILL_1__8717_ (
);

FILL SFILL104440x55050 (
);

FILL FILL_2__15907_ (
);

FILL FILL_0__16101_ (
);

FILL FILL_5__13487_ (
);

FILL FILL_2__10622_ (
);

DFFSR _7787_ (
    .Q(\datapath_1.regfile_1.regOut[7] [21]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_393_[21])
);

INVX1 _7367_ (
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_251_)
);

FILL SFILL33880x81050 (
);

FILL SFILL108760x63050 (
);

FILL FILL_2__13094_ (
);

FILL FILL_5_BUFX2_insert60 (
);

FILL FILL_5_BUFX2_insert61 (
);

FILL FILL_5_BUFX2_insert62 (
);

FILL FILL_5_BUFX2_insert63 (
);

FILL FILL_1__12087_ (
);

FILL FILL_5_BUFX2_insert64 (
);

FILL FILL_5_BUFX2_insert65 (
);

FILL FILL_4__13841_ (
);

FILL FILL_5_BUFX2_insert66 (
);

FILL FILL_4__13421_ (
);

FILL FILL_5_BUFX2_insert67 (
);

FILL FILL_4__13001_ (
);

FILL FILL_5_BUFX2_insert68 (
);

FILL FILL_5_BUFX2_insert69 (
);

FILL FILL_3__7191_ (
);

INVX1 _11785_ (
    .A(_2152_),
    .Y(_2878_)
);

FILL FILL_0__9094_ (
);

FILL SFILL49080x52050 (
);

NAND2X1 _11365_ (
    .A(_2319_),
    .B(_2481__bF$buf1),
    .Y(_2482_)
);

FILL FILL_3__12834_ (
);

FILL FILL_3__12414_ (
);

FILL SFILL28920x37050 (
);

FILL FILL_4__7927_ (
);

FILL FILL_4__7507_ (
);

FILL FILL_2__11827_ (
);

FILL FILL_0__12861_ (
);

FILL FILL_2__11407_ (
);

FILL FILL_0__12441_ (
);

FILL FILL_0__12021_ (
);

FILL FILL_2__14299_ (
);

FILL FILL_5__15633_ (
);

FILL FILL_5__15213_ (
);

FILL FILL_0__7827_ (
);

INVX1 _9933_ (
    .A(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_1555_)
);

INVX1 _9513_ (
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_1336_)
);

FILL FILL_1__8890_ (
);

FILL FILL_1__8470_ (
);

FILL FILL_4__14626_ (
);

FILL FILL_2__15660_ (
);

FILL FILL_4__14206_ (
);

FILL FILL_2__15240_ (
);

FILL FILL_3__8396_ (
);

FILL SFILL49000x50050 (
);

FILL FILL_3__13619_ (
);

FILL FILL_1__14653_ (
);

FILL FILL_1__14233_ (
);

FILL FILL_0__13646_ (
);

AOI22X1 _13931_ (
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .B(_3942__bF$buf3),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_4433_)
);

FILL FILL_0__13226_ (
);

NOR2X1 _13511_ (
    .A(_4018_),
    .B(_4021_),
    .Y(_4022_)
);

FILL FILL_5__9683_ (
);

FILL FILL_5__9263_ (
);

FILL FILL_5__11973_ (
);

FILL FILL_1__9675_ (
);

FILL FILL_5__11553_ (
);

FILL FILL_1__9255_ (
);

FILL FILL_5__11133_ (
);

BUFX2 BUFX2_insert1050 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf2 )
);

BUFX2 BUFX2_insert1051 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf1 )
);

FILL FILL_4__7680_ (
);

FILL FILL_2__16025_ (
);

BUFX2 BUFX2_insert1052 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf0 )
);

FILL FILL_4__10966_ (
);

BUFX2 BUFX2_insert1053 (
    .A(_4038_),
    .Y(_4038__bF$buf3)
);

FILL SFILL94360x66050 (
);

BUFX2 BUFX2_insert1054 (
    .A(_4038_),
    .Y(_4038__bF$buf2)
);

FILL FILL_4__10546_ (
);

FILL FILL_4__10126_ (
);

BUFX2 BUFX2_insert1055 (
    .A(_4038_),
    .Y(_4038__bF$buf1)
);

FILL FILL_2__11580_ (
);

BUFX2 BUFX2_insert1056 (
    .A(_4038_),
    .Y(_4038__bF$buf0)
);

FILL FILL_2__11160_ (
);

BUFX2 BUFX2_insert1057 (
    .A(_5531_),
    .Y(_5531__bF$buf4)
);

FILL FILL_1__15858_ (
);

BUFX2 BUFX2_insert1058 (
    .A(_5531_),
    .Y(_5531__bF$buf3)
);

FILL FILL_1__15438_ (
);

BUFX2 BUFX2_insert1059 (
    .A(_5531_),
    .Y(_5531__bF$buf2)
);

FILL FILL_1__15018_ (
);

FILL FILL_1__10993_ (
);

FILL FILL_1__10573_ (
);

FILL FILL_1__10153_ (
);

INVX1 _14716_ (
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_5202_)
);

FILL SFILL98680x74050 (
);

FILL FILL_0__7580_ (
);

BUFX2 BUFX2_insert870 (
    .A(_3891_),
    .Y(_3891__bF$buf1)
);

FILL FILL_2__7598_ (
);

FILL SFILL79160x46050 (
);

FILL FILL_2__7178_ (
);

BUFX2 BUFX2_insert871 (
    .A(_3891_),
    .Y(_3891__bF$buf0)
);

FILL FILL_0__7160_ (
);

BUFX2 BUFX2_insert872 (
    .A(_3947_),
    .Y(_3947__bF$buf3)
);

BUFX2 BUFX2_insert873 (
    .A(_3947_),
    .Y(_3947__bF$buf2)
);

FILL FILL_3__10900_ (
);

BUFX2 BUFX2_insert874 (
    .A(_3947_),
    .Y(_3947__bF$buf1)
);

BUFX2 BUFX2_insert875 (
    .A(_3947_),
    .Y(_3947__bF$buf0)
);

BUFX2 BUFX2_insert876 (
    .A(_5499_),
    .Y(_5499__bF$buf3)
);

BUFX2 BUFX2_insert877 (
    .A(_5499_),
    .Y(_5499__bF$buf2)
);

BUFX2 BUFX2_insert878 (
    .A(_5499_),
    .Y(_5499__bF$buf1)
);

BUFX2 BUFX2_insert879 (
    .A(_5499_),
    .Y(_5499__bF$buf0)
);

FILL FILL_5__12758_ (
);

FILL SFILL18760x2050 (
);

FILL FILL_3__13792_ (
);

FILL FILL_5__12338_ (
);

FILL FILL_3__13372_ (
);

FILL FILL_4__8885_ (
);

FILL SFILL18680x7050 (
);

FILL FILL_4__8465_ (
);

FILL FILL_2__12785_ (
);

FILL FILL_2__12365_ (
);

FILL FILL_1__11778_ (
);

FILL FILL_1__11358_ (
);

FILL FILL_5__16171_ (
);

FILL FILL_3__6882_ (
);

FILL FILL_0__8785_ (
);

FILL FILL_0__8365_ (
);

NAND2X1 _10636_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1902_)
);

DFFSR _10216_ (
    .Q(\datapath_1.regfile_1.regOut[26] [18]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_1628_[18])
);

FILL FILL_4__15584_ (
);

FILL FILL_4__15164_ (
);

FILL SFILL8760x83050 (
);

FILL FILL_2__9744_ (
);

FILL FILL_3__14997_ (
);

FILL FILL_3__14577_ (
);

FILL FILL_0__11712_ (
);

FILL FILL_3__14157_ (
);

FILL SFILL29480x62050 (
);

FILL FILL_1__15191_ (
);

FILL FILL_0__14184_ (
);

FILL FILL_5__14904_ (
);

FILL SFILL53960x73050 (
);

FILL SFILL84360x64050 (
);

FILL FILL_1__7741_ (
);

FILL FILL_1__7321_ (
);

FILL FILL_2__14931_ (
);

FILL FILL_2__14511_ (
);

FILL FILL_3__7247_ (
);

FILL FILL_5__12091_ (
);

FILL FILL_1__13924_ (
);

FILL FILL_4__16369_ (
);

FILL FILL_1__13504_ (
);

FILL FILL_4__11084_ (
);

FILL FILL_0__12917_ (
);

FILL FILL_1__16396_ (
);

FILL FILL_5__8954_ (
);

FILL FILL_3__10497_ (
);

FILL FILL_5__8114_ (
);

FILL FILL_0__15389_ (
);

OAI22X1 _15674_ (
    .A(_4670_),
    .B(_5544__bF$buf2),
    .C(_5480__bF$buf0),
    .D(_6138_),
    .Y(_6139_)
);

INVX1 _15254_ (
    .A(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_5730_)
);

FILL FILL_3__16303_ (
);

FILL FILL_5__10824_ (
);

FILL FILL_1__8526_ (
);

FILL FILL_5__10404_ (
);

FILL FILL_1__8106_ (
);

FILL FILL_2__15716_ (
);

FILL FILL_4__6951_ (
);

FILL FILL_0__16330_ (
);

FILL FILL_5__13296_ (
);

FILL FILL_2__10431_ (
);

FILL FILL_2__10011_ (
);

FILL FILL_1__14709_ (
);

FILL FILL_4_BUFX2_insert1090 (
);

INVX1 _7596_ (
    .A(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_363_)
);

INVX1 _7176_ (
    .A(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_144_)
);

FILL FILL_4_BUFX2_insert1091 (
);

FILL FILL_4_BUFX2_insert1092 (
);

FILL FILL_4_BUFX2_insert1093 (
);

FILL FILL_4__12289_ (
);

FILL FILL_3__9813_ (
);

FILL FILL_2__6869_ (
);

FILL FILL_0__6851_ (
);

FILL FILL_5__9739_ (
);

FILL SFILL114520x45050 (
);

FILL FILL_4__13650_ (
);

FILL FILL_4__13230_ (
);

NOR2X1 _16039_ (
    .A(_6492_),
    .B(_6494_),
    .Y(_6495_)
);

FILL SFILL3720x64050 (
);

OAI21X1 _11594_ (
    .A(_2700_),
    .B(_2423_),
    .C(_2263_),
    .Y(_2701_)
);

OAI21X1 _11174_ (
    .A(_2291_),
    .B(_2292_),
    .C(_2289_),
    .Y(_2293_)
);

FILL FILL_2__7810_ (
);

FILL FILL_5__11609_ (
);

FILL FILL_3__12643_ (
);

FILL SFILL43960x71050 (
);

FILL FILL_3__12223_ (
);

FILL SFILL74360x62050 (
);

FILL FILL_4__7736_ (
);

FILL FILL_4__7316_ (
);

FILL FILL_2__11636_ (
);

FILL FILL_2__11216_ (
);

FILL FILL_0__12250_ (
);

FILL SFILL114920x14050 (
);

FILL FILL_1__10629_ (
);

FILL FILL_5__15862_ (
);

FILL FILL_5__15442_ (
);

FILL FILL_5__15022_ (
);

FILL FILL_0__7636_ (
);

INVX1 _9742_ (
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_1448_)
);

FILL FILL_0__7216_ (
);

DFFSR _9322_ (
    .Q(\datapath_1.regfile_1.regOut[19] [20]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_1173_[20])
);

FILL SFILL43880x78050 (
);

FILL FILL_4__14855_ (
);

FILL FILL_4__14435_ (
);

FILL FILL_4__14015_ (
);

DFFSR _12799_ (
    .Q(\datapath_1.PCJump [10]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[8])
);

INVX1 _12379_ (
    .A(ALUOut[12]),
    .Y(_3318_)
);

FILL SFILL3560x9050 (
);

FILL FILL_3__13848_ (
);

FILL FILL_3__13428_ (
);

FILL FILL_1__14882_ (
);

FILL FILL_1__14462_ (
);

FILL FILL_3__13008_ (
);

FILL FILL_1__14042_ (
);

FILL FILL_0__13875_ (
);

FILL FILL_0__13455_ (
);

INVX8 _13740_ (
    .A(_3905__bF$buf0),
    .Y(_4246_)
);

NOR2X1 _13320_ (
    .A(_3781_),
    .B(_3850_),
    .Y(\datapath_1.regfile_1.regEn [13])
);

FILL FILL_0__13035_ (
);

FILL FILL_5__9492_ (
);

FILL FILL_5__16227_ (
);

FILL FILL_3__6938_ (
);

FILL FILL_6__9808_ (
);

FILL FILL_5__11782_ (
);

FILL FILL_1__9484_ (
);

FILL FILL_5__11362_ (
);

FILL FILL_2__16254_ (
);

FILL FILL_4__10775_ (
);

FILL FILL_1__15667_ (
);

FILL FILL_1__15247_ (
);

FILL FILL_5__7805_ (
);

FILL SFILL59000x47050 (
);

FILL FILL_1__10382_ (
);

INVX1 _14945_ (
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_5426_)
);

AOI21X1 _14525_ (
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .B(_4115_),
    .C(_5014_),
    .Y(_5015_)
);

NOR2X1 _14105_ (
    .A(_4603_),
    .B(_4600_),
    .Y(_4604_)
);

FILL FILL_0__15601_ (
);

FILL FILL_5__12987_ (
);

FILL FILL_5__12567_ (
);

FILL FILL_5__12147_ (
);

BUFX2 _6867_ (
    .A(_1_[29]),
    .Y(memoryAddress[29])
);

FILL FILL_4__8694_ (
);

FILL SFILL33880x76050 (
);

FILL FILL_4__8274_ (
);

FILL FILL_2__12594_ (
);

FILL FILL_2__12174_ (
);

FILL FILL_1__11587_ (
);

FILL FILL_1__11167_ (
);

FILL FILL_4__12501_ (
);

FILL FILL_0__8594_ (
);

FILL SFILL49080x47050 (
);

DFFSR _10865_ (
    .Q(\datapath_1.regfile_1.regOut[31] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_1953_[27])
);

FILL FILL_6__9141_ (
);

INVX1 _10445_ (
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_1815_)
);

INVX1 _10025_ (
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_1596_)
);

FILL FILL_3__11914_ (
);

FILL FILL_6__14779_ (
);

FILL FILL_4__15393_ (
);

FILL FILL_2__10907_ (
);

FILL FILL_0__11941_ (
);

FILL FILL_2__9553_ (
);

FILL FILL_2__9133_ (
);

FILL FILL_3__14386_ (
);

FILL FILL_0__11521_ (
);

FILL FILL_0__11101_ (
);

FILL FILL_6__15720_ (
);

FILL FILL_4__9899_ (
);

FILL FILL_4__9479_ (
);

FILL FILL_2__13799_ (
);

FILL FILL_2__13379_ (
);

FILL FILL_5__14713_ (
);

FILL FILL_0__6907_ (
);

FILL FILL_1__7970_ (
);

FILL FILL_1__7550_ (
);

FILL FILL_4__13706_ (
);

FILL FILL_2__14740_ (
);

FILL FILL_2__14320_ (
);

FILL FILL_0__9799_ (
);

FILL SFILL33400x60050 (
);

FILL FILL_0__9379_ (
);

FILL FILL_3__7476_ (
);

FILL FILL_3__7056_ (
);

FILL FILL_1__13733_ (
);

FILL FILL_1__13313_ (
);

FILL FILL_4__16178_ (
);

FILL FILL_6__10279_ (
);

FILL SFILL94440x54050 (
);

FILL FILL_0__12726_ (
);

FILL FILL_0__12306_ (
);

FILL FILL_5__8763_ (
);

FILL FILL_5__8343_ (
);

FILL FILL_6__11640_ (
);

FILL FILL_0__15198_ (
);

INVX1 _15483_ (
    .A(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_5953_)
);

FILL FILL_5__15918_ (
);

INVX1 _15063_ (
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_5543_)
);

FILL FILL_3__16112_ (
);

FILL FILL_5__10633_ (
);

FILL FILL_1__8755_ (
);

FILL FILL_1__8335_ (
);

FILL FILL_2__15945_ (
);

FILL FILL_2__15525_ (
);

FILL FILL_2__15105_ (
);

FILL FILL_2__10660_ (
);

FILL FILL_2__10240_ (
);

FILL FILL_1__14938_ (
);

FILL FILL_1__14518_ (
);

FILL FILL_4__12098_ (
);

FILL FILL_3__9622_ (
);

FILL FILL_5__9548_ (
);

FILL FILL_5__9128_ (
);

NAND3X1 _16268_ (
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6718_)
);

FILL FILL_5__11838_ (
);

FILL FILL_3__12872_ (
);

FILL FILL_5__11418_ (
);

FILL FILL_3__12452_ (
);

FILL SFILL54280x20050 (
);

FILL FILL_3__12032_ (
);

FILL FILL_4__7965_ (
);

FILL FILL_4__7545_ (
);

FILL FILL_4__7125_ (
);

FILL FILL_2__11865_ (
);

FILL FILL_2__11445_ (
);

FILL FILL_2__11025_ (
);

FILL FILL_1__10438_ (
);

FILL FILL_1__10018_ (
);

FILL FILL_5__15671_ (
);

FILL FILL_5__15251_ (
);

FILL FILL_0__7865_ (
);

FILL FILL_6__8832_ (
);

DFFSR _9971_ (
    .Q(\datapath_1.regfile_1.regOut[24] [29]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_1498_[29])
);

FILL FILL_0__7445_ (
);

FILL SFILL84440x52050 (
);

OAI21X1 _9551_ (
    .A(_1360_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .C(_1361_),
    .Y(_1303_[29])
);

OAI21X1 _9131_ (
    .A(_1141_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .C(_1142_),
    .Y(_1108_[17])
);

FILL FILL_4__14664_ (
);

FILL SFILL8760x78050 (
);

FILL FILL_4__14244_ (
);

NAND2X1 _12188_ (
    .A(ALUSrcA_bF$buf6),
    .B(\datapath_1.a [24]),
    .Y(_3179_)
);

FILL FILL_2__8824_ (
);

FILL FILL_3__13657_ (
);

FILL FILL_2__8404_ (
);

FILL FILL_3__13237_ (
);

FILL FILL_1__14691_ (
);

FILL FILL_1__14271_ (
);

FILL FILL_0_BUFX2_insert510 (
);

FILL FILL_0_BUFX2_insert511 (
);

FILL FILL_0_BUFX2_insert512 (
);

FILL FILL_0_BUFX2_insert513 (
);

FILL FILL_0__13684_ (
);

FILL FILL_0_BUFX2_insert514 (
);

FILL SFILL114600x78050 (
);

FILL FILL_0__13264_ (
);

FILL FILL_0_BUFX2_insert515 (
);

FILL SFILL53960x68050 (
);

FILL FILL_0_BUFX2_insert516 (
);

FILL SFILL84360x59050 (
);

FILL FILL_0_BUFX2_insert517 (
);

FILL FILL_0_BUFX2_insert518 (
);

FILL FILL_0_BUFX2_insert519 (
);

FILL FILL_5__16036_ (
);

FILL FILL_6__9617_ (
);

FILL FILL_5__11591_ (
);

FILL FILL_1__9293_ (
);

FILL FILL_5__11171_ (
);

FILL FILL_4__15869_ (
);

FILL FILL_4__15449_ (
);

FILL FILL_4__15029_ (
);

FILL FILL_2__16063_ (
);

FILL FILL_4__10164_ (
);

FILL SFILL8760x33050 (
);

FILL FILL_2__9609_ (
);

FILL SFILL13800x70050 (
);

FILL FILL_1__15896_ (
);

FILL FILL_1__15476_ (
);

FILL FILL_1__15056_ (
);

FILL FILL_5__7614_ (
);

FILL FILL_1__10191_ (
);

FILL FILL_0__14889_ (
);

FILL FILL_0__14469_ (
);

NAND3X1 _14754_ (
    .A(_5231_),
    .B(_5230_),
    .C(_5238_),
    .Y(_5239_)
);

FILL FILL_0__14049_ (
);

INVX1 _14334_ (
    .A(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_4828_)
);

FILL FILL_3__15803_ (
);

FILL SFILL114600x33050 (
);

FILL FILL_1__7606_ (
);

FILL SFILL84360x14050 (
);

FILL FILL_0__15830_ (
);

FILL FILL_0__15410_ (
);

FILL FILL_5__12376_ (
);

FILL FILL_4__11789_ (
);

FILL FILL_4__8083_ (
);

FILL FILL_4__11369_ (
);

FILL FILL_1__11396_ (
);

NOR2X1 _15959_ (
    .A(_6416_),
    .B(_6414_),
    .Y(_6417_)
);

FILL FILL_4__12730_ (
);

OAI22X1 _15539_ (
    .A(_5530__bF$buf3),
    .B(_4552_),
    .C(_4560_),
    .D(_5534__bF$buf4),
    .Y(_6007_)
);

FILL FILL_4__12310_ (
);

NOR2X1 _15119_ (
    .A(_5594_),
    .B(_5597_),
    .Y(_5598_)
);

INVX1 _10674_ (
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_1927_)
);

FILL FILL_0__10389_ (
);

INVX1 _10254_ (
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_1708_)
);

FILL SFILL43960x66050 (
);

FILL FILL_3__11723_ (
);

FILL FILL_3__11303_ (
);

FILL FILL_2__9782_ (
);

FILL FILL_0__11750_ (
);

FILL FILL_2__9362_ (
);

FILL FILL_3__14195_ (
);

FILL FILL_0__11330_ (
);

FILL FILL_4__9288_ (
);

FILL FILL112360x70050 (
);

FILL FILL_5__14942_ (
);

FILL FILL_5__14522_ (
);

FILL FILL_5__14102_ (
);

INVX1 _8822_ (
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_1041_)
);

OAI21X1 _8402_ (
    .A(_777_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .C(_778_),
    .Y(_718_[30])
);

FILL FILL_4__13935_ (
);

FILL FILL_4__13515_ (
);

NAND2X1 _11879_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [15]),
    .Y(_2963_)
);

AOI21X1 _11459_ (
    .A(_2526_),
    .B(_2522_),
    .C(_2302_),
    .Y(_2574_)
);

NOR2X1 _11039_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2157_),
    .Y(_2158_)
);

FILL FILL_3__12508_ (
);

FILL FILL_1__13962_ (
);

FILL SFILL64840x62050 (
);

FILL FILL_1__13542_ (
);

FILL FILL_1__13122_ (
);

FILL SFILL43960x21050 (
);

FILL FILL112280x77050 (
);

FILL FILL_0__12955_ (
);

DFFSR _12820_ (
    .Q(\control_1.op [3]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3490_[29])
);

FILL FILL_0__12115_ (
);

INVX1 _12400_ (
    .A(ALUOut[19]),
    .Y(_3332_)
);

FILL FILL_5__8992_ (
);

FILL FILL_6__16314_ (
);

FILL FILL_5__8572_ (
);

OAI22X1 _15292_ (
    .A(_5549__bF$buf1),
    .B(_4238_),
    .C(_5466__bF$buf1),
    .D(_4202_),
    .Y(_5767_)
);

FILL FILL_5__15727_ (
);

FILL FILL_5__15307_ (
);

FILL FILL_3__16341_ (
);

OAI21X1 _9607_ (
    .A(_1377_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .C(_1378_),
    .Y(_1368_[5])
);

FILL FILL_1__8984_ (
);

FILL FILL_5__10442_ (
);

FILL FILL_5__10022_ (
);

FILL FILL_1__8144_ (
);

FILL SFILL104520x38050 (
);

FILL FILL_2__15754_ (
);

FILL SFILL43880x28050 (
);

FILL FILL_2__15334_ (
);

FILL FILL_1__14747_ (
);

FILL FILL_1__14327_ (
);

FILL FILL_3__9851_ (
);

AOI21X1 _13605_ (
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .B(_3894_),
    .C(_4113_),
    .Y(_4114_)
);

FILL FILL_3__9011_ (
);

FILL FILL112280x32050 (
);

FILL FILL_5__9777_ (
);

FILL FILL_5__9357_ (
);

FILL FILL_6__12234_ (
);

INVX1 _16077_ (
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_6532_)
);

FILL FILL_1__9769_ (
);

FILL FILL_5__11647_ (
);

FILL FILL_5__11227_ (
);

FILL FILL_1__9349_ (
);

FILL FILL_3__12261_ (
);

FILL FILL_2__16119_ (
);

FILL FILL_4__7354_ (
);

FILL FILL_2__11674_ (
);

FILL FILL_2__11254_ (
);

FILL FILL_1__10667_ (
);

FILL FILL_1__10247_ (
);

FILL FILL_5__15480_ (
);

FILL FILL_5__15060_ (
);

FILL FILL_0__7674_ (
);

OAI21X1 _9780_ (
    .A(_1472_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .C(_1473_),
    .Y(_1433_[20])
);

OAI21X1 _9360_ (
    .A(_1253_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .C(_1254_),
    .Y(_1238_[8])
);

FILL FILL_6__8221_ (
);

FILL FILL_6__13439_ (
);

FILL FILL_4__14893_ (
);

FILL FILL_4__14473_ (
);

FILL FILL_4__14053_ (
);

FILL FILL_3__13886_ (
);

FILL FILL_2__8633_ (
);

FILL FILL_3__13466_ (
);

FILL FILL_2__8213_ (
);

FILL FILL_3__13046_ (
);

FILL FILL_1__14080_ (
);

FILL FILL_6__14800_ (
);

FILL FILL_4__8979_ (
);

FILL FILL_4__8139_ (
);

FILL FILL_2__12879_ (
);

FILL FILL_2__12459_ (
);

FILL SFILL94520x42050 (
);

FILL FILL_2__12039_ (
);

FILL FILL_0__13493_ (
);

FILL SFILL33880x26050 (
);

FILL FILL_4__9920_ (
);

FILL FILL_4__9500_ (
);

FILL FILL_2__13820_ (
);

FILL FILL_3__6976_ (
);

FILL FILL_2__13400_ (
);

FILL FILL_0__8879_ (
);

FILL FILL_5__16265_ (
);

FILL FILL_0__8459_ (
);

FILL FILL_4__15678_ (
);

FILL FILL_4__15258_ (
);

FILL FILL_2__16292_ (
);

FILL SFILL94440x49050 (
);

FILL FILL_4__10393_ (
);

FILL FILL_2__9418_ (
);

FILL FILL_0__9400_ (
);

FILL FILL_0__11806_ (
);

FILL FILL_1__15285_ (
);

FILL FILL_5__7843_ (
);

FILL FILL_5__7423_ (
);

NAND3X1 _14983_ (
    .A(_5459__bF$buf2),
    .B(_5462_),
    .C(_5461_),
    .Y(_5463_)
);

FILL FILL_0__14698_ (
);

INVX1 _14563_ (
    .A(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_5052_)
);

FILL FILL_6__10300_ (
);

FILL FILL_0__14278_ (
);

NAND3X1 _14143_ (
    .A(_4632_),
    .B(_4633_),
    .C(_4640_),
    .Y(_4641_)
);

FILL FILL_3__15612_ (
);

FILL FILL_1__7835_ (
);

FILL FILL_1__7415_ (
);

FILL FILL_2__14605_ (
);

FILL FILL_5__12185_ (
);

FILL FILL_4__11598_ (
);

FILL FILL_4__11178_ (
);

FILL FILL_3__8702_ (
);

FILL FILL_5__8628_ (
);

FILL FILL_5__8208_ (
);

NAND2X1 _15768_ (
    .A(_6225_),
    .B(_6230_),
    .Y(_6231_)
);

NAND3X1 _15348_ (
    .A(_5812_),
    .B(_5820_),
    .C(_5816_),
    .Y(_5821_)
);

DFFSR _10483_ (
    .Q(\datapath_1.regfile_1.regOut[28] [29]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1758_[29])
);

OAI21X1 _10063_ (
    .A(_1620_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .C(_1621_),
    .Y(_1563_[29])
);

FILL FILL_5__10918_ (
);

FILL SFILL23880x24050 (
);

FILL FILL_3__11952_ (
);

FILL FILL_3__11532_ (
);

FILL FILL_3__11112_ (
);

FILL SFILL4120x44050 (
);

FILL FILL_0__16004_ (
);

FILL FILL_2__10945_ (
);

FILL FILL_2__9591_ (
);

FILL FILL_2__10525_ (
);

FILL FILL_2__9171_ (
);

FILL FILL_2__10105_ (
);

FILL SFILL39000x38050 (
);

FILL FILL112440x1050 (
);

FILL FILL_4__9097_ (
);

FILL FILL112360x6050 (
);

FILL FILL_3__9907_ (
);

FILL FILL_5__14751_ (
);

FILL FILL_0__6945_ (
);

FILL FILL_5__14331_ (
);

OAI21X1 _8631_ (
    .A(_889_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .C(_890_),
    .Y(_848_[21])
);

OAI21X1 _8211_ (
    .A(_670_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_671_),
    .Y(_653_[9])
);

FILL FILL_4__13744_ (
);

FILL FILL_4__13324_ (
);

FILL SFILL18840x50 (
);

FILL FILL_3__7094_ (
);

OAI21X1 _11688_ (
    .A(_2787_),
    .B(_2788_),
    .C(_2784_),
    .Y(_2789_)
);

INVX1 _11268_ (
    .A(_2386_),
    .Y(_2387_)
);

FILL SFILL23800x22050 (
);

FILL FILL_3__12737_ (
);

FILL FILL_1__13771_ (
);

FILL FILL_3__12317_ (
);

FILL FILL_1__13351_ (
);

FILL FILL_0__12764_ (
);

FILL FILL_0__12344_ (
);

FILL FILL_5__8381_ (
);

FILL SFILL74200x3050 (
);

FILL SFILL29080x38050 (
);

FILL FILL_5__15956_ (
);

FILL FILL_5__15536_ (
);

FILL FILL_5__15116_ (
);

DFFSR _9836_ (
    .Q(\datapath_1.regfile_1.regOut[23] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_1433_[22])
);

FILL FILL_3__16150_ (
);

NAND2X1 _9416_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1292_)
);

FILL FILL_5__10671_ (
);

FILL SFILL114200x59050 (
);

FILL FILL_1__8373_ (
);

FILL FILL_5__10251_ (
);

FILL FILL_4__14949_ (
);

FILL FILL_2__15983_ (
);

FILL FILL_4__14529_ (
);

FILL FILL_2__15563_ (
);

FILL FILL_4__14109_ (
);

FILL FILL_2__15143_ (
);

FILL FILL_1__14976_ (
);

FILL FILL_1__14556_ (
);

FILL FILL_1__14136_ (
);

FILL FILL_3__9660_ (
);

FILL FILL_0__13969_ (
);

INVX1 _13834_ (
    .A(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_4339_)
);

FILL FILL_3__9240_ (
);

FILL FILL_0__13549_ (
);

OAI22X1 _13414_ (
    .A(_3922_),
    .B(_3925_),
    .C(_3924__bF$buf3),
    .D(_3923_),
    .Y(_3926_)
);

FILL FILL_0__13129_ (
);

FILL FILL_5__9166_ (
);

FILL SFILL29000x36050 (
);

FILL FILL_0__14910_ (
);

FILL FILL_5__11876_ (
);

FILL FILL_1__9998_ (
);

FILL FILL_5__11456_ (
);

FILL FILL_1__9158_ (
);

FILL FILL_3__12490_ (
);

FILL FILL_5__11036_ (
);

FILL FILL_3__12070_ (
);

FILL FILL_2__16348_ (
);

FILL FILL_4__7583_ (
);

FILL FILL_4__7163_ (
);

FILL FILL_4__10449_ (
);

FILL FILL_4__10029_ (
);

FILL FILL_2__11483_ (
);

FILL FILL_2__11063_ (
);

FILL FILL_6__7089_ (
);

FILL SFILL13800x20050 (
);

FILL FILL_1__10896_ (
);

FILL FILL_1__10056_ (
);

INVX1 _14619_ (
    .A(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_5107_)
);

FILL FILL_4__11810_ (
);

FILL SFILL74040x31050 (
);

FILL FILL_0__7483_ (
);

FILL FILL_0__7063_ (
);

FILL FILL_3__10803_ (
);

FILL FILL_4__14282_ (
);

FILL FILL_2__8862_ (
);

FILL FILL_0__10830_ (
);

FILL FILL_2__8442_ (
);

FILL FILL_3__13695_ (
);

FILL FILL_3__13275_ (
);

FILL FILL_0__10410_ (
);

FILL FILL_4__8788_ (
);

FILL FILL_4__8368_ (
);

FILL FILL112360x65050 (
);

FILL FILL_2__12268_ (
);

FILL FILL_5__13602_ (
);

DFFSR _7902_ (
    .Q(\datapath_1.regfile_1.regOut[8] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_458_[8])
);

FILL SFILL64040x74050 (
);

FILL FILL_5__16074_ (
);

NAND3X1 _10959_ (
    .A(_2084_),
    .B(_2090_),
    .C(_2072_),
    .Y(_2091_)
);

FILL FILL_0__8268_ (
);

OAI21X1 _10539_ (
    .A(_1856_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1857_),
    .Y(_1823_[17])
);

FILL FILL_6__9235_ (
);

OAI21X1 _10119_ (
    .A(_1637_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .C(_1638_),
    .Y(_1628_[5])
);

FILL FILL_1__12622_ (
);

FILL FILL_4__15487_ (
);

FILL FILL_1__12202_ (
);

FILL FILL_4__15067_ (
);

FILL SFILL43960x16050 (
);

FILL FILL_2__9647_ (
);

FILL FILL_2__9227_ (
);

NAND2X1 _11900_ (
    .A(IorD_bF$buf3),
    .B(ALUOut[4]),
    .Y(_2975_)
);

FILL FILL_0__11615_ (
);

FILL FILL_1__15094_ (
);

FILL FILL_5__7232_ (
);

FILL SFILL44600x3050 (
);

AOI22X1 _14792_ (
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .B(_4005__bF$buf3),
    .C(_3998__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_5276_)
);

INVX1 _14372_ (
    .A(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_4865_)
);

FILL FILL_0__14087_ (
);

FILL FILL_5__14807_ (
);

FILL FILL_3__15841_ (
);

FILL FILL112360x20050 (
);

FILL FILL_3__15421_ (
);

FILL FILL_3__15001_ (
);

FILL FILL_1__7224_ (
);

FILL FILL_2__14834_ (
);

FILL FILL_2__14414_ (
);

FILL FILL_1__13827_ (
);

FILL FILL_1__13407_ (
);

FILL SFILL84360x5050 (
);

FILL FILL_3__8511_ (
);

FILL FILL112280x27050 (
);

FILL FILL_1__16299_ (
);

FILL FILL_5__8857_ (
);

FILL FILL_5__8017_ (
);

OAI22X1 _15997_ (
    .A(_5478__bF$buf1),
    .B(_5066_),
    .C(_5073_),
    .D(_5485__bF$buf3),
    .Y(_6454_)
);

INVX1 _15577_ (
    .A(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_6044_)
);

OAI22X1 _15157_ (
    .A(_5472__bF$buf2),
    .B(_4059_),
    .C(_4056_),
    .D(_5526__bF$buf4),
    .Y(_5635_)
);

FILL FILL_3__16206_ (
);

OAI21X1 _10292_ (
    .A(_1732_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .C(_1733_),
    .Y(_1693_[20])
);

FILL FILL_1__8849_ (
);

FILL FILL_3__11761_ (
);

FILL FILL_5__10307_ (
);

FILL FILL_3__11341_ (
);

FILL FILL_1__8009_ (
);

FILL FILL_2__15619_ (
);

FILL FILL_4__6854_ (
);

FILL FILL_0__16233_ (
);

FILL FILL_2__10754_ (
);

NAND2X1 _7499_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_319_)
);

NAND2X1 _7079_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_100_)
);

FILL FILL_5__14980_ (
);

FILL FILL_5__14560_ (
);

FILL FILL_5__14140_ (
);

OAI21X1 _8860_ (
    .A(_1001_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .C(_1002_),
    .Y(_978_[12])
);

OAI21X1 _8440_ (
    .A(_846_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_847_),
    .Y(_783_[0])
);

NAND2X1 _8020_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_585_)
);

FILL FILL_4__13973_ (
);

FILL FILL_4__13553_ (
);

FILL FILL_4__13133_ (
);

OAI21X1 _11497_ (
    .A(_2295_),
    .B(_2347__bF$buf0),
    .C(_2609_),
    .Y(_2610_)
);

NOR2X1 _11077_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(_2195_),
    .Y(_2196_)
);

FILL FILL_2__7713_ (
);

FILL FILL_3__12966_ (
);

FILL FILL_3__12126_ (
);

FILL FILL_1__13580_ (
);

FILL FILL_1__13160_ (
);

FILL FILL_4__7219_ (
);

FILL FILL_2__11959_ (
);

FILL FILL_0__12993_ (
);

FILL FILL_2__11539_ (
);

FILL FILL_0__12573_ (
);

FILL FILL_3_CLKBUF1_insert170 (
);

FILL FILL_2__11119_ (
);

FILL FILL_0__12153_ (
);

FILL FILL_3_CLKBUF1_insert171 (
);

FILL FILL_3_CLKBUF1_insert172 (
);

FILL FILL_3_CLKBUF1_insert173 (
);

FILL FILL_3_CLKBUF1_insert174 (
);

FILL FILL_3_CLKBUF1_insert175 (
);

FILL FILL_5__8190_ (
);

FILL FILL_3_CLKBUF1_insert176 (
);

FILL FILL_3_CLKBUF1_insert177 (
);

FILL FILL_3_CLKBUF1_insert178 (
);

FILL FILL_3_CLKBUF1_insert179 (
);

FILL FILL_5__15765_ (
);

FILL FILL_2__12900_ (
);

FILL FILL_5__15345_ (
);

FILL FILL_0__7959_ (
);

FILL SFILL98840x45050 (
);

FILL FILL_0__7119_ (
);

NAND2X1 _9645_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1404_)
);

NAND2X1 _9225_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1185_)
);

FILL FILL_5__10060_ (
);

FILL FILL_1__8182_ (
);

FILL FILL_4__14758_ (
);

FILL FILL_4__14338_ (
);

FILL FILL_2__15792_ (
);

FILL FILL_2__15372_ (
);

FILL FILL_0__8900_ (
);

FILL FILL_1__14785_ (
);

FILL FILL_1__14365_ (
);

FILL FILL_5__6923_ (
);

FILL FILL_0__13778_ (
);

FILL FILL_0__13358_ (
);

OAI22X1 _13643_ (
    .A(_4149_),
    .B(_3905__bF$buf2),
    .C(_3935__bF$buf4),
    .D(_4150_),
    .Y(_4151_)
);

NAND2X1 _13223_ (
    .A(\datapath_1.a3 [4]),
    .B(_3758_),
    .Y(_3766_)
);

FILL FILL_5__9395_ (
);

FILL SFILL44040x70050 (
);

FILL FILL_1__6915_ (
);

FILL FILL_5__11685_ (
);

FILL FILL_1__9387_ (
);

FILL FILL_5__11265_ (
);

FILL FILL_2__16157_ (
);

FILL FILL_4__10678_ (
);

FILL FILL_4__10258_ (
);

FILL FILL_2__11292_ (
);

FILL FILL_5__7708_ (
);

FILL FILL_2_BUFX2_insert420 (
);

FILL FILL_2_BUFX2_insert421 (
);

FILL FILL_1__10285_ (
);

FILL FILL_2_BUFX2_insert422 (
);

INVX1 _14848_ (
    .A(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_5331_)
);

FILL FILL_2_BUFX2_insert423 (
);

FILL FILL_2_BUFX2_insert424 (
);

INVX1 _14428_ (
    .A(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_4920_)
);

INVX1 _14008_ (
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_4509_)
);

FILL FILL_2_BUFX2_insert425 (
);

FILL FILL_2_BUFX2_insert426 (
);

FILL FILL_2_BUFX2_insert427 (
);

FILL FILL_0__7292_ (
);

FILL FILL_2_BUFX2_insert428 (
);

FILL FILL_2_BUFX2_insert429 (
);

FILL FILL_0_CLKBUF1_insert120 (
);

FILL FILL_0_CLKBUF1_insert121 (
);

FILL FILL_4__14091_ (
);

FILL FILL_0__15924_ (
);

FILL FILL_0_CLKBUF1_insert122 (
);

FILL FILL_0__15504_ (
);

FILL FILL_0_CLKBUF1_insert123 (
);

FILL FILL_0_CLKBUF1_insert124 (
);

FILL FILL_0_CLKBUF1_insert125 (
);

FILL FILL_0_CLKBUF1_insert126 (
);

FILL FILL_2__8251_ (
);

FILL FILL_0_CLKBUF1_insert127 (
);

FILL FILL_3__13084_ (
);

FILL FILL_0_CLKBUF1_insert128 (
);

FILL FILL_0_CLKBUF1_insert129 (
);

FILL FILL_4__8597_ (
);

FILL SFILL84120x21050 (
);

FILL FILL_2__12497_ (
);

FILL FILL_2__12077_ (
);

FILL FILL_5__13831_ (
);

FILL FILL_5__13411_ (
);

OAI21X1 _7711_ (
    .A(_418_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .C(_419_),
    .Y(_393_[13])
);

FILL FILL_4__12824_ (
);

FILL FILL_4__12404_ (
);

FILL FILL_0__8497_ (
);

OAI21X1 _10768_ (
    .A(_1968_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .C(_1969_),
    .Y(_1953_[8])
);

FILL FILL_0__8077_ (
);

FILL SFILL23800x17050 (
);

DFFSR _10348_ (
    .Q(\datapath_1.regfile_1.regOut[27] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_1693_[22])
);

FILL FILL_3__11817_ (
);

FILL FILL_1__12851_ (
);

FILL FILL_1__12431_ (
);

FILL FILL_4__15296_ (
);

FILL FILL_1__12011_ (
);

FILL FILL_2__9876_ (
);

FILL FILL_0__11844_ (
);

FILL FILL_2__9036_ (
);

FILL FILL_3__14289_ (
);

FILL FILL_0__11424_ (
);

FILL FILL_0__11004_ (
);

FILL FILL_6__15623_ (
);

FILL FILL_5__7881_ (
);

FILL FILL_5__7461_ (
);

FILL SFILL74120x64050 (
);

FILL FILL_5__7041_ (
);

AOI22X1 _14181_ (
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .B(_4246_),
    .C(_4115_),
    .D(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_4678_)
);

FILL FILL_5__14616_ (
);

FILL FILL_3__15650_ (
);

FILL FILL_3__15230_ (
);

NAND2X1 _8916_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1040_)
);

FILL SFILL103720x1050 (
);

FILL FILL_1__7873_ (
);

FILL FILL_1__7453_ (
);

FILL FILL_1__7033_ (
);

FILL FILL_4__13609_ (
);

FILL FILL_2__14643_ (
);

FILL FILL_2__14223_ (
);

FILL FILL_3__7799_ (
);

FILL FILL_3__7379_ (
);

FILL FILL_1__13636_ (
);

FILL FILL_1__13216_ (
);

FILL FILL_1_BUFX2_insert440 (
);

FILL FILL_3__8740_ (
);

FILL FILL_1_BUFX2_insert441 (
);

FILL FILL_3__8320_ (
);

FILL FILL_0__12629_ (
);

FILL FILL_1_BUFX2_insert442 (
);

NAND2X1 _12914_ (
    .A(vdd),
    .B(\datapath_1.rd1 [30]),
    .Y(_3615_)
);

FILL FILL_1_BUFX2_insert443 (
);

FILL FILL_0__12209_ (
);

FILL FILL_1_BUFX2_insert444 (
);

FILL FILL_1_BUFX2_insert445 (
);

FILL FILL_1_BUFX2_insert446 (
);

FILL FILL_5__8246_ (
);

FILL FILL_1_BUFX2_insert447 (
);

FILL FILL_1_BUFX2_insert448 (
);

FILL FILL_1_BUFX2_insert449 (
);

FILL FILL_6__11963_ (
);

FILL FILL_6__11543_ (
);

OAI22X1 _15386_ (
    .A(_4363_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf1),
    .D(_5857_),
    .Y(_5858_)
);

FILL FILL_3__16015_ (
);

FILL FILL_5__10956_ (
);

FILL FILL_5__10536_ (
);

FILL FILL_3__11990_ (
);

FILL FILL_1__8658_ (
);

FILL FILL_5__10116_ (
);

FILL FILL_1__8238_ (
);

FILL FILL_3__11570_ (
);

FILL FILL_3__11150_ (
);

FILL FILL_2__15848_ (
);

FILL FILL_2__15428_ (
);

FILL FILL_2__15008_ (
);

FILL FILL_0__16042_ (
);

FILL FILL_2__10983_ (
);

FILL FILL_2__10563_ (
);

FILL FILL_2__10143_ (
);

FILL SFILL13800x15050 (
);

FILL FILL_3__9525_ (
);

FILL FILL_3__9105_ (
);

FILL FILL_0__6983_ (
);

FILL FILL_6__7110_ (
);

FILL FILL_6__12748_ (
);

FILL FILL_4__13782_ (
);

FILL FILL_4__13362_ (
);

FILL FILL_2__7942_ (
);

FILL FILL_3__12775_ (
);

BUFX2 BUFX2_insert110 (
    .A(IorD),
    .Y(IorD_bF$buf0)
);

FILL FILL_2__7102_ (
);

FILL FILL_3__12355_ (
);

FILL FILL_4__7868_ (
);

FILL FILL_4__7448_ (
);

FILL FILL_2__11768_ (
);

FILL FILL_2__11348_ (
);

FILL FILL_0__12382_ (
);

FILL FILL_2_CLKBUF1_insert160 (
);

FILL SFILL49000x4050 (
);

FILL FILL_2_CLKBUF1_insert161 (
);

FILL SFILL64040x69050 (
);

FILL FILL_5__15994_ (
);

FILL FILL_2_CLKBUF1_insert162 (
);

FILL SFILL89240x2050 (
);

FILL FILL_2_CLKBUF1_insert163 (
);

FILL FILL_5__15574_ (
);

FILL FILL_2_CLKBUF1_insert164 (
);

FILL FILL_5__15154_ (
);

FILL FILL_0__7348_ (
);

NAND2X1 _9874_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1516_)
);

FILL FILL_2_CLKBUF1_insert165 (
);

FILL FILL_2_CLKBUF1_insert166 (
);

DFFSR _9454_ (
    .Q(\datapath_1.regfile_1.regOut[20] [24]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1238_[24])
);

FILL FILL_6__8315_ (
);

INVX1 _9034_ (
    .A(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_1098_)
);

FILL FILL_2_CLKBUF1_insert167 (
);

FILL SFILL23640x5050 (
);

FILL FILL_2_CLKBUF1_insert168 (
);

FILL FILL_4__14987_ (
);

FILL FILL_2_CLKBUF1_insert169 (
);

FILL FILL_4__14567_ (
);

FILL FILL_1__11702_ (
);

FILL FILL_4__14147_ (
);

FILL FILL_2__15181_ (
);

FILL FILL_2__8727_ (
);

FILL FILL_1__14594_ (
);

FILL FILL_1__14174_ (
);

FILL FILL_6_BUFX2_insert1042 (
);

FILL FILL_0__13587_ (
);

NOR2X1 _13872_ (
    .A(_4375_),
    .B(_4372_),
    .Y(_4376_)
);

FILL FILL_0__13167_ (
);

INVX1 _13452_ (
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_3964_)
);

FILL FILL_6_BUFX2_insert1047 (
);

INVX1 _13032_ (
    .A(_2_[27]),
    .Y(_3673_)
);

FILL FILL112360x15050 (
);

FILL FILL_3__14921_ (
);

FILL FILL_3__14501_ (
);

FILL FILL_2__13914_ (
);

FILL FILL_5__16359_ (
);

FILL SFILL64040x24050 (
);

FILL FILL_5__11494_ (
);

FILL FILL_5__11074_ (
);

FILL FILL_1__12907_ (
);

FILL FILL_2__16386_ (
);

FILL FILL_4__10487_ (
);

FILL FILL_0__9914_ (
);

FILL FILL_4__10067_ (
);

FILL SFILL89240x73050 (
);

FILL FILL_1__15799_ (
);

FILL SFILL54120x60050 (
);

FILL FILL_1__15379_ (
);

FILL FILL_5__7937_ (
);

FILL SFILL89880x50 (
);

NAND3X1 _14657_ (
    .A(_5142_),
    .B(_5143_),
    .C(_5141_),
    .Y(_5144_)
);

OAI22X1 _14237_ (
    .A(_4732_),
    .B(_3972__bF$buf2),
    .C(_3920_),
    .D(_4731_),
    .Y(_4733_)
);

FILL FILL_3__15706_ (
);

FILL FILL_1__16320_ (
);

FILL FILL_1__7929_ (
);

FILL FILL_1__7509_ (
);

FILL FILL_3__10421_ (
);

FILL FILL_3__10001_ (
);

FILL FILL_0__15733_ (
);

FILL FILL_0__15313_ (
);

FILL FILL_5__12699_ (
);

FILL SFILL54040x67050 (
);

FILL FILL_2__8480_ (
);

FILL FILL_5__12279_ (
);

FILL FILL_2__8060_ (
);

DFFSR _6999_ (
    .Q(\datapath_1.regfile_1.regOut[1] [1]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_3_[1])
);

FILL FILL_5__13640_ (
);

FILL FILL_5__13220_ (
);

OAI21X1 _7940_ (
    .A(_530_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_531_),
    .Y(_523_[4])
);

DFFSR _7520_ (
    .Q(\datapath_1.regfile_1.regOut[5] [10]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_263_[10])
);

NAND2X1 _7100_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_114_)
);

FILL FILL_1__11299_ (
);

FILL FILL_4__12633_ (
);

FILL FILL_4__12213_ (
);

NOR2X1 _10997_ (
    .A(_2115_),
    .B(_2114_),
    .Y(_2116_)
);

NAND2X1 _10577_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1883_)
);

NAND2X1 _10157_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1664_)
);

FILL FILL_3__11626_ (
);

FILL FILL_1__12660_ (
);

FILL FILL_3__11206_ (
);

FILL FILL_1__12240_ (
);

FILL FILL_2__9685_ (
);

FILL FILL_2__10619_ (
);

FILL FILL_2__9265_ (
);

FILL FILL_0__11653_ (
);

FILL FILL_0__11233_ (
);

FILL FILL_3__14098_ (
);

FILL FILL_5__7690_ (
);

FILL SFILL54040x22050 (
);

FILL FILL_5__14845_ (
);

FILL FILL_5__14425_ (
);

FILL FILL_5__14005_ (
);

NAND2X1 _8725_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_933_)
);

DFFSR _8305_ (
    .Q(\datapath_1.regfile_1.regOut[11] [27]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_653_[27])
);

FILL SFILL79240x71050 (
);

FILL FILL_1__7682_ (
);

FILL FILL_4__13838_ (
);

FILL FILL_2__14872_ (
);

FILL FILL_4__13418_ (
);

FILL FILL_2__14452_ (
);

FILL FILL_2__14032_ (
);

FILL FILL_3__7188_ (
);

FILL FILL_1__13865_ (
);

FILL FILL_1__13445_ (
);

FILL FILL_1__13025_ (
);

FILL FILL_0__12858_ (
);

NAND2X1 _12723_ (
    .A(IRWrite_bF$buf3),
    .B(memoryOutData[9]),
    .Y(_3508_)
);

FILL FILL_0__12438_ (
);

FILL SFILL33880x2050 (
);

FILL FILL_0__12018_ (
);

NAND3X1 _12303_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3266_)
);

FILL FILL_5__8895_ (
);

FILL SFILL79160x78050 (
);

FILL FILL_6__16217_ (
);

FILL FILL_5__8475_ (
);

FILL SFILL44040x65050 (
);

FILL FILL_5__8055_ (
);

NOR2X1 _15195_ (
    .A(_5671_),
    .B(_5670_),
    .Y(_5672_)
);

FILL FILL_3__16244_ (
);

FILL FILL_5__10765_ (
);

FILL FILL_1__8887_ (
);

FILL FILL_1__8467_ (
);

FILL FILL_2__15657_ (
);

FILL FILL_2__15237_ (
);

FILL FILL_4__6892_ (
);

FILL FILL_0__16271_ (
);

FILL FILL_2__10792_ (
);

FILL FILL_2__10372_ (
);

FILL FILL_3__9754_ (
);

FILL FILL_3__9334_ (
);

NAND3X1 _13928_ (
    .A(_4429_),
    .B(_4430_),
    .C(_4428_),
    .Y(_4431_)
);

INVX1 _13508_ (
    .A(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_4019_)
);

FILL FILL_4__13591_ (
);

FILL FILL_6__12137_ (
);

FILL FILL_4__13171_ (
);

FILL SFILL44040x20050 (
);

FILL FILL_2__7751_ (
);

FILL FILL_2__7331_ (
);

FILL FILL_3__12584_ (
);

FILL FILL_3__12164_ (
);

FILL FILL_4__7677_ (
);

FILL FILL_2__11997_ (
);

FILL FILL_2__11577_ (
);

FILL FILL_2__11157_ (
);

FILL FILL_0__12191_ (
);

FILL FILL_5__12911_ (
);

FILL SFILL109800x21050 (
);

FILL FILL_4__11904_ (
);

FILL FILL_5__15383_ (
);

FILL FILL_0__7997_ (
);

FILL FILL_0__7577_ (
);

INVX1 _9683_ (
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_1429_)
);

INVX1 _9263_ (
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_1210_)
);

FILL FILL_1_CLKBUF1_insert150 (
);

FILL FILL_1_CLKBUF1_insert151 (
);

FILL FILL_4__14796_ (
);

FILL FILL_1__11931_ (
);

FILL FILL_1_CLKBUF1_insert152 (
);

FILL FILL_1_CLKBUF1_insert153 (
);

FILL FILL_4__14376_ (
);

FILL FILL_1__11511_ (
);

FILL FILL_1_CLKBUF1_insert154 (
);

FILL FILL_1_CLKBUF1_insert155 (
);

FILL FILL_1_CLKBUF1_insert156 (
);

FILL FILL_1_CLKBUF1_insert157 (
);

FILL FILL_1_CLKBUF1_insert158 (
);

FILL FILL_2__8956_ (
);

FILL FILL_0__10924_ (
);

FILL FILL_3__13789_ (
);

FILL FILL_1_CLKBUF1_insert159 (
);

FILL FILL_3__13369_ (
);

FILL FILL_0__10504_ (
);

FILL FILL_2__8116_ (
);

FILL SFILL109720x28050 (
);

FILL FILL_5__6961_ (
);

FILL SFILL74120x59050 (
);

NOR2X1 _13681_ (
    .A(_4188_),
    .B(_4185_),
    .Y(_4189_)
);

FILL FILL_0__13396_ (
);

NOR2X1 _13261_ (
    .A(\datapath_1.a3 [4]),
    .B(_3799_),
    .Y(_3804_)
);

FILL FILL_3__14730_ (
);

FILL FILL_3__14310_ (
);

FILL FILL_1__6953_ (
);

FILL FILL_4__9403_ (
);

FILL FILL_2__13723_ (
);

FILL SFILL109320x14050 (
);

FILL FILL_2__13303_ (
);

FILL FILL_5__16168_ (
);

FILL FILL_3__6879_ (
);

FILL FILL_1__12716_ (
);

FILL FILL_2__16195_ (
);

FILL FILL_4__10296_ (
);

FILL FILL_3__7820_ (
);

FILL FILL_0__9723_ (
);

FILL SFILL69160x31050 (
);

FILL FILL_0__11709_ (
);

FILL FILL_1__15188_ (
);

FILL FILL_5__7746_ (
);

FILL FILL_2_BUFX2_insert800 (
);

FILL FILL_5__7326_ (
);

FILL FILL_4__16102_ (
);

FILL FILL_2_BUFX2_insert801 (
);

FILL FILL_2_BUFX2_insert802 (
);

FILL SFILL78840x36050 (
);

FILL FILL_2_BUFX2_insert803 (
);

INVX1 _14886_ (
    .A(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_5368_)
);

OAI22X1 _14466_ (
    .A(_4956_),
    .B(_3910_),
    .C(_3944__bF$buf3),
    .D(_4955_),
    .Y(_4957_)
);

FILL FILL_2_BUFX2_insert804 (
);

FILL SFILL74120x14050 (
);

FILL FILL_2_BUFX2_insert805 (
);

NOR3X1 _14046_ (
    .A(_4542_),
    .B(_4545_),
    .C(_4540_),
    .Y(_4546_)
);

FILL FILL_3__15935_ (
);

FILL FILL_2_BUFX2_insert806 (
);

FILL SFILL28920x3050 (
);

FILL FILL_3__15515_ (
);

FILL FILL_2_BUFX2_insert807 (
);

FILL FILL_2_BUFX2_insert808 (
);

FILL FILL_2_BUFX2_insert809 (
);

FILL FILL_1__7738_ (
);

FILL FILL_3__10650_ (
);

FILL FILL_1__7318_ (
);

FILL SFILL28840x8050 (
);

FILL FILL_3__10230_ (
);

FILL FILL_6__13095_ (
);

FILL FILL_2__14928_ (
);

FILL FILL_2__14508_ (
);

FILL FILL_0__15962_ (
);

FILL SFILL99320x63050 (
);

FILL FILL_0__15542_ (
);

FILL FILL_0__15122_ (
);

FILL FILL_5__12088_ (
);

FILL SFILL8760x4050 (
);

FILL FILL_3__8605_ (
);

FILL SFILL8680x9050 (
);

FILL SFILL68840x79050 (
);

FILL FILL_4__12862_ (
);

FILL FILL_4__12442_ (
);

FILL SFILL64120x57050 (
);

FILL FILL_4__12022_ (
);

NAND2X1 _10386_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1776_)
);

FILL FILL_3__11855_ (
);

FILL FILL_3__11435_ (
);

FILL FILL_3__11015_ (
);

FILL FILL_4__6948_ (
);

FILL FILL_0__16327_ (
);

FILL FILL_2__10428_ (
);

FILL FILL_0__11882_ (
);

FILL FILL_2__9494_ (
);

FILL FILL_2__10008_ (
);

FILL FILL_0__11462_ (
);

FILL FILL_0__11042_ (
);

FILL FILL_5__14654_ (
);

FILL FILL_5__14234_ (
);

FILL FILL_0__6848_ (
);

NAND2X1 _8954_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1045_)
);

DFFSR _8534_ (
    .Q(\datapath_1.regfile_1.regOut[13] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_783_[0])
);

INVX1 _8114_ (
    .A(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_627_)
);

FILL FILL_1__7491_ (
);

FILL FILL_1__7071_ (
);

FILL FILL_4__13647_ (
);

FILL FILL_4__13227_ (
);

FILL FILL_2__14681_ (
);

FILL FILL_2__14261_ (
);

FILL FILL_2__7807_ (
);

FILL SFILL64120x12050 (
);

FILL FILL_1__13674_ (
);

FILL FILL_1__13254_ (
);

FILL FILL_1_BUFX2_insert820 (
);

FILL FILL_1_BUFX2_insert821 (
);

NAND2X1 _12952_ (
    .A(\datapath_1.rd2 [0]),
    .B(vdd),
    .Y(_3684_)
);

FILL FILL_1_BUFX2_insert822 (
);

INVX1 _12532_ (
    .A(ALUOut[31]),
    .Y(_3421_)
);

FILL FILL_1_BUFX2_insert823 (
);

FILL FILL_0__12247_ (
);

FILL SFILL89320x61050 (
);

NAND3X1 _12112_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump [31]),
    .C(_3034__bF$buf1),
    .Y(_3130_)
);

FILL FILL_1_BUFX2_insert824 (
);

FILL FILL_1_BUFX2_insert825 (
);

FILL FILL_1_BUFX2_insert826 (
);

FILL FILL_1_BUFX2_insert827 (
);

FILL FILL_1_BUFX2_insert828 (
);

FILL FILL_1_BUFX2_insert829 (
);

FILL FILL_5__15859_ (
);

FILL FILL_5__15439_ (
);

FILL FILL_5__15019_ (
);

INVX1 _9739_ (
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_1446_)
);

FILL FILL_3__16053_ (
);

FILL SFILL18760x81050 (
);

FILL SFILL64040x19050 (
);

FILL SFILL3560x50 (
);

DFFSR _9319_ (
    .Q(\datapath_1.regfile_1.regOut[19] [17]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1173_[17])
);

FILL FILL_5__10994_ (
);

FILL FILL_5__10574_ (
);

FILL FILL_1__8696_ (
);

FILL FILL_5__10154_ (
);

FILL FILL_1__8276_ (
);

FILL FILL_2__15886_ (
);

FILL FILL_2__15466_ (
);

FILL FILL_2__15046_ (
);

FILL FILL_0__16080_ (
);

FILL SFILL89240x68050 (
);

FILL FILL_2__10181_ (
);

FILL SFILL54120x55050 (
);

FILL FILL_1__14879_ (
);

FILL FILL_1__14459_ (
);

FILL FILL_1__14039_ (
);

FILL FILL_3__9983_ (
);

FILL FILL_3__9143_ (
);

NAND3X1 _13737_ (
    .A(_4242_),
    .B(_4243_),
    .C(_4241_),
    .Y(_4244_)
);

OAI21X1 _13317_ (
    .A(\datapath_1.a3 [4]),
    .B(_3837_),
    .C(_3848_),
    .Y(_3849_)
);

FILL FILL_1__15820_ (
);

FILL FILL_5__9489_ (
);

FILL FILL_1__15400_ (
);

FILL FILL_0__14813_ (
);

FILL FILL_2__7980_ (
);

FILL FILL_5__11779_ (
);

FILL FILL_2__7560_ (
);

FILL FILL_5__11359_ (
);

FILL FILL_3__12393_ (
);

FILL FILL_4__7486_ (
);

FILL FILL_4__7066_ (
);

FILL FILL_2__11386_ (
);

FILL FILL_5__12720_ (
);

FILL FILL_5__12300_ (
);

FILL FILL_1__10799_ (
);

FILL SFILL54120x10050 (
);

FILL FILL_1__10379_ (
);

FILL FILL_4__11713_ (
);

FILL FILL_5__15192_ (
);

INVX1 _9492_ (
    .A(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_1322_)
);

DFFSR _9072_ (
    .Q(\datapath_1.regfile_1.regOut[17] [26]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_1043_[26])
);

FILL FILL_3__10706_ (
);

FILL SFILL18680x43050 (
);

FILL FILL_1__11740_ (
);

FILL FILL_4__14185_ (
);

FILL FILL_1__11320_ (
);

FILL FILL_2__8765_ (
);

FILL FILL_3__13598_ (
);

FILL FILL_2__8345_ (
);

FILL FILL_0__10313_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL SFILL54040x17050 (
);

FILL FILL_0_BUFX2_insert12 (
);

FILL FILL_0_BUFX2_insert13 (
);

FILL FILL_0_BUFX2_insert14 (
);

FILL FILL_0_BUFX2_insert15 (
);

FILL FILL_0_BUFX2_insert16 (
);

INVX8 _13490_ (
    .A(_3909_),
    .Y(_4001_)
);

FILL FILL_0_BUFX2_insert17 (
);

DFFSR _13070_ (
    .Q(_2_[23]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_3620_[23])
);

FILL FILL_0_BUFX2_insert18 (
);

FILL FILL_5__13925_ (
);

FILL FILL_0_BUFX2_insert19 (
);

FILL FILL_5__13505_ (
);

NAND2X1 _7805_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_462_)
);

FILL SFILL79240x66050 (
);

FILL FILL_4_BUFX2_insert330 (
);

FILL FILL_4__9632_ (
);

FILL FILL_4_BUFX2_insert331 (
);

FILL FILL_4__12918_ (
);

FILL FILL_4_BUFX2_insert332 (
);

FILL FILL_4__9212_ (
);

FILL FILL_4_BUFX2_insert333 (
);

FILL FILL_2__13952_ (
);

FILL FILL_4_BUFX2_insert334 (
);

FILL FILL_2__13532_ (
);

FILL FILL_5__16397_ (
);

FILL FILL_2__13112_ (
);

FILL FILL_4_BUFX2_insert335 (
);

FILL FILL_4_BUFX2_insert336 (
);

FILL FILL_4_BUFX2_insert337 (
);

FILL FILL_4_BUFX2_insert338 (
);

FILL FILL_4_BUFX2_insert339 (
);

FILL FILL_1__12525_ (
);

FILL FILL_1__12105_ (
);

FILL FILL_0__9532_ (
);

FILL FILL_0__11938_ (
);

FILL FILL_0__9112_ (
);

AOI22X1 _11803_ (
    .A(_2143_),
    .B(_2481__bF$buf0),
    .C(_2341__bF$buf3),
    .D(_2144_),
    .Y(_2895_)
);

FILL FILL_0__11518_ (
);

FILL FILL_5__7975_ (
);

FILL FILL_5__7555_ (
);

FILL FILL_4__16331_ (
);

INVX1 _14695_ (
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_5181_)
);

NAND3X1 _14275_ (
    .A(_4768_),
    .B(_4769_),
    .C(_4767_),
    .Y(_4770_)
);

FILL FILL_3__15744_ (
);

FILL FILL_3__15324_ (
);

FILL FILL_1__7967_ (
);

FILL FILL_1__7547_ (
);

FILL FILL_2__14737_ (
);

FILL FILL_2__14317_ (
);

FILL FILL_0__15771_ (
);

FILL FILL_0__15351_ (
);

FILL FILL_3__8834_ (
);

FILL SFILL109400x47050 (
);

FILL SFILL44040x15050 (
);

FILL FILL_4__12251_ (
);

FILL FILL_3__16109_ (
);

INVX1 _10195_ (
    .A(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_1689_)
);

FILL FILL_3__11664_ (
);

FILL FILL_3__11244_ (
);

FILL SFILL69240x64050 (
);

DFFSR _16421_ (
    .Q(\datapath_1.regfile_1.regOut[0] [4]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_6769_[4])
);

FILL FILL_0__16136_ (
);

INVX1 _16001_ (
    .A(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_6458_)
);

FILL SFILL109000x33050 (
);

FILL FILL_2__10657_ (
);

FILL FILL_2__10237_ (
);

FILL FILL_0__11691_ (
);

FILL FILL_0__11271_ (
);

FILL FILL_6__15470_ (
);

FILL FILL_6__15050_ (
);

FILL FILL_3_BUFX2_insert350 (
);

FILL FILL_3__9619_ (
);

FILL FILL_3_BUFX2_insert351 (
);

FILL FILL_5__14883_ (
);

FILL FILL_3_BUFX2_insert352 (
);

FILL FILL_3_BUFX2_insert353 (
);

FILL FILL_5__14463_ (
);

FILL FILL_3_BUFX2_insert354 (
);

FILL FILL_5__14043_ (
);

INVX1 _8763_ (
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_958_)
);

FILL FILL_3_BUFX2_insert355 (
);

FILL FILL_3_BUFX2_insert356 (
);

INVX1 _8343_ (
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_739_)
);

FILL FILL_3_BUFX2_insert357 (
);

FILL FILL_3_BUFX2_insert358 (
);

FILL FILL_4__13876_ (
);

FILL FILL_3_BUFX2_insert359 (
);

FILL FILL_4__13456_ (
);

FILL FILL_2__14490_ (
);

FILL FILL_4__13036_ (
);

FILL FILL_2__14070_ (
);

FILL FILL_3__12869_ (
);

FILL FILL_2__7616_ (
);

FILL FILL_3__12449_ (
);

FILL FILL_3__12029_ (
);

FILL FILL_1__13483_ (
);

FILL FILL_0__12896_ (
);

INVX1 _12761_ (
    .A(\datapath_1.PCJump [24]),
    .Y(_3533_)
);

FILL FILL_0__12476_ (
);

FILL FILL_0__12056_ (
);

AOI22X1 _12341_ (
    .A(_2_[31]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3295_)
);

FILL FILL_3__13810_ (
);

FILL FILL_5__8093_ (
);

FILL FILL_4__8903_ (
);

FILL FILL_6__11390_ (
);

FILL FILL_5__15668_ (
);

FILL FILL_5__15248_ (
);

DFFSR _9968_ (
    .Q(\datapath_1.regfile_1.regOut[24] [26]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_1498_[26])
);

FILL FILL_3__16282_ (
);

OAI21X1 _9548_ (
    .A(_1358_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .C(_1359_),
    .Y(_1303_[28])
);

OAI21X1 _9128_ (
    .A(_1139_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1140_),
    .Y(_1108_[16])
);

FILL FILL_5__10383_ (
);

FILL FILL_1__8085_ (
);

FILL FILL_2__15695_ (
);

FILL FILL_2__15275_ (
);

FILL SFILL99400x51050 (
);

FILL SFILL38760x35050 (
);

FILL SFILL69160x26050 (
);

FILL FILL_3__6900_ (
);

FILL SFILL34040x13050 (
);

FILL FILL_1__14688_ (
);

FILL FILL_1__14268_ (
);

FILL FILL_0_BUFX2_insert480 (
);

FILL FILL_0_BUFX2_insert481 (
);

FILL FILL_4__15602_ (
);

FILL FILL_0_BUFX2_insert482 (
);

FILL FILL_3__9792_ (
);

FILL FILL_0_BUFX2_insert483 (
);

FILL FILL_3__9372_ (
);

OAI22X1 _13966_ (
    .A(_4466_),
    .B(_3916_),
    .C(_3983__bF$buf2),
    .D(_4467_),
    .Y(_4468_)
);

FILL FILL_0_BUFX2_insert484 (
);

FILL FILL_0_BUFX2_insert485 (
);

INVX1 _13546_ (
    .A(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_4056_)
);

OAI21X1 _13126_ (
    .A(_3714_),
    .B(PCEn_bF$buf6),
    .C(_3715_),
    .Y(_3685_[15])
);

FILL FILL_0_BUFX2_insert486 (
);

FILL FILL_0_BUFX2_insert487 (
);

FILL FILL_0_BUFX2_insert488 (
);

FILL FILL_0_BUFX2_insert489 (
);

FILL FILL_5__9298_ (
);

FILL SFILL99320x58050 (
);

FILL FILL_0__14622_ (
);

FILL FILL_0__14202_ (
);

FILL FILL_5__11588_ (
);

FILL FILL_5__11168_ (
);

FILL FILL_4__7295_ (
);

FILL SFILL28760x78050 (
);

FILL SFILL59160x69050 (
);

FILL FILL_2__11195_ (
);

FILL FILL_1__10188_ (
);

FILL FILL_4__11942_ (
);

FILL FILL_4__11522_ (
);

FILL FILL_4__11102_ (
);

FILL FILL_0__7195_ (
);

FILL FILL_1__16414_ (
);

FILL FILL_3__10935_ (
);

FILL FILL_3__10515_ (
);

FILL FILL_0__15827_ (
);

FILL FILL_0__15407_ (
);

FILL FILL_2__8994_ (
);

FILL FILL_0__10962_ (
);

FILL FILL_2__8574_ (
);

FILL SFILL99320x13050 (
);

FILL FILL_0__10542_ (
);

FILL FILL_0__10122_ (
);

FILL SFILL49640x74050 (
);

FILL FILL_5__13734_ (
);

FILL FILL_5__13314_ (
);

FILL SFILL28760x33050 (
);

FILL SFILL59160x24050 (
);

INVX1 _7614_ (
    .A(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_375_)
);

FILL FILL_1__6991_ (
);

FILL FILL_4__9861_ (
);

FILL FILL_4__9021_ (
);

FILL FILL_4__12727_ (
);

FILL FILL_2__13761_ (
);

FILL FILL_4__12307_ (
);

FILL FILL_2__13341_ (
);

FILL FILL_6__9787_ (
);

FILL FILL_1__12754_ (
);

FILL FILL_4__15199_ (
);

FILL FILL_1__12334_ (
);

FILL FILL_0__9761_ (
);

FILL FILL_2__9779_ (
);

FILL FILL_2__9359_ (
);

FILL FILL_0__11747_ (
);

FILL FILL_0__9341_ (
);

FILL SFILL89320x56050 (
);

FILL FILL_0__11327_ (
);

NOR2X1 _11612_ (
    .A(_2710_),
    .B(_2717_),
    .Y(_2718_)
);

FILL FILL_6__15526_ (
);

FILL FILL_5__7364_ (
);

FILL FILL_6__15106_ (
);

FILL FILL_4__16140_ (
);

FILL FILL_5__14939_ (
);

NOR2X1 _14084_ (
    .A(_4582_),
    .B(_4579_),
    .Y(_4583_)
);

FILL FILL_3__15973_ (
);

FILL FILL_5__14519_ (
);

FILL FILL_3__15553_ (
);

FILL SFILL18760x76050 (
);

DFFSR _8819_ (
    .Q(\datapath_1.regfile_1.regOut[15] [29]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_913_[29])
);

FILL FILL_3__15133_ (
);

FILL SFILL113880x18050 (
);

FILL FILL_1__7356_ (
);

FILL FILL_2__14966_ (
);

FILL FILL_2__14546_ (
);

FILL FILL_2__14126_ (
);

FILL FILL_0__15580_ (
);

FILL FILL_0__15160_ (
);

FILL SFILL73640x78050 (
);

FILL FILL_1__13959_ (
);

FILL FILL_1__13539_ (
);

FILL FILL_1__13119_ (
);

FILL FILL_3__8643_ (
);

DFFSR _12817_ (
    .Q(\control_1.op [0]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3490_[26])
);

FILL FILL_3__8223_ (
);

FILL FILL_5__8989_ (
);

FILL FILL_1__14900_ (
);

FILL FILL_5__8569_ (
);

FILL FILL_5__8149_ (
);

FILL SFILL89320x11050 (
);

FILL FILL_6__11446_ (
);

FILL FILL_4__12480_ (
);

FILL FILL_6__11026_ (
);

NOR2X1 _15289_ (
    .A(_5763_),
    .B(_5761_),
    .Y(_5764_)
);

FILL FILL_4__12060_ (
);

FILL FILL_3__16338_ (
);

FILL FILL_5__9930_ (
);

FILL FILL_3__11893_ (
);

FILL FILL_5__10439_ (
);

FILL FILL_5__10019_ (
);

FILL FILL_5__9510_ (
);

FILL FILL_3__11473_ (
);

FILL FILL_3__11053_ (
);

FILL SFILL18760x31050 (
);

FILL FILL_4__6986_ (
);

FILL FILL_0__16365_ (
);

NOR2X1 _16230_ (
    .A(_6679_),
    .B(_6680_),
    .Y(_6681_)
);

FILL FILL_2__10886_ (
);

FILL FILL_2__10046_ (
);

FILL FILL_0__11080_ (
);

FILL FILL_5__11800_ (
);

FILL FILL_1__9922_ (
);

FILL FILL_1__9502_ (
);

FILL SFILL89240x18050 (
);

FILL FILL_3__9848_ (
);

FILL FILL_3__9428_ (
);

FILL FILL_3__9008_ (
);

FILL FILL_5__14692_ (
);

FILL FILL_0__6886_ (
);

FILL FILL_5__14272_ (
);

INVX1 _8992_ (
    .A(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_1070_)
);

INVX1 _8572_ (
    .A(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_851_)
);

DFFSR _8152_ (
    .Q(\datapath_1.regfile_1.regOut[10] [2]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_588_[2])
);

FILL SFILL79320x54050 (
);

FILL SFILL18680x38050 (
);

FILL FILL_4__13685_ (
);

FILL FILL_1__10820_ (
);

FILL FILL_4__13265_ (
);

FILL FILL_1__10400_ (
);

FILL FILL_2__7845_ (
);

FILL FILL_2__7425_ (
);

FILL FILL111960x67050 (
);

FILL FILL_3__12258_ (
);

FILL FILL_1__13292_ (
);

INVX1 _12990_ (
    .A(_2_[13]),
    .Y(_3645_)
);

INVX1 _12570_ (
    .A(\datapath_1.Data [1]),
    .Y(_3426_)
);

FILL FILL_0__12285_ (
);

OAI21X1 _12150_ (
    .A(_3152_),
    .B(ALUSrcA_bF$buf2),
    .C(_3153_),
    .Y(\datapath_1.alu_1.ALUInA [11])
);

FILL FILL_4__8712_ (
);

FILL FILL_5__15897_ (
);

FILL FILL_2__12612_ (
);

FILL FILL_5__15477_ (
);

FILL FILL_5__15057_ (
);

FILL FILL_3__16091_ (
);

OAI21X1 _9777_ (
    .A(_1470_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1471_),
    .Y(_1433_[19])
);

OAI21X1 _9357_ (
    .A(_1251_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .C(_1252_),
    .Y(_1238_[7])
);

FILL FILL_5__10192_ (
);

FILL FILL_1__11605_ (
);

FILL FILL_2__15084_ (
);

FILL FILL_0__8612_ (
);

FILL FILL_1__14497_ (
);

FILL FILL_1__14077_ (
);

FILL FILL_4__15831_ (
);

FILL FILL_4__15411_ (
);

FILL FILL111960x22050 (
);

OAI22X1 _13775_ (
    .A(_4279_),
    .B(_3936__bF$buf3),
    .C(_3971__bF$buf4),
    .D(_4280_),
    .Y(_4281_)
);

OAI21X1 _13355_ (
    .A(_3766_),
    .B(\datapath_1.a3 [1]),
    .C(_3756_),
    .Y(_3872_)
);

FILL FILL_3__14824_ (
);

FILL FILL_3__14404_ (
);

FILL FILL_4__9917_ (
);

FILL FILL_2__13817_ (
);

FILL FILL_0__14851_ (
);

FILL FILL_0__14431_ (
);

FILL FILL_0__14011_ (
);

FILL FILL_5__11397_ (
);

FILL FILL_1__9099_ (
);

FILL FILL_2__16289_ (
);

FILL FILL_4__11751_ (
);

FILL FILL_4__11331_ (
);

FILL FILL_3__15609_ (
);

FILL FILL_6__8391_ (
);

FILL FILL_1__16223_ (
);

FILL FILL_3__10744_ (
);

FILL FILL_3__10324_ (
);

INVX1 _15921_ (
    .A(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_6380_)
);

FILL FILL_0__15636_ (
);

AOI22X1 _15501_ (
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [11]),
    .C(\datapath_1.regfile_1.regOut[11] [11]),
    .D(_5496_),
    .Y(_5970_)
);

FILL FILL_0__15216_ (
);

FILL SFILL114360x41050 (
);

FILL FILL_2__8383_ (
);

FILL FILL_0__10771_ (
);

FILL FILL_5__13963_ (
);

FILL FILL_5__13543_ (
);

FILL FILL_5__13123_ (
);

INVX1 _7843_ (
    .A(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_487_)
);

INVX1 _7423_ (
    .A(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_268_)
);

FILL FILL_4_BUFX2_insert710 (
);

DFFSR _7003_ (
    .Q(\datapath_1.regfile_1.regOut[1] [5]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_3_[5])
);

FILL FILL_4_BUFX2_insert711 (
);

FILL FILL_4__9670_ (
);

FILL FILL_4__9250_ (
);

FILL FILL_4_BUFX2_insert712 (
);

FILL FILL_4__12956_ (
);

FILL FILL_2__13990_ (
);

FILL FILL_4_BUFX2_insert713 (
);

FILL FILL_4_BUFX2_insert714 (
);

FILL FILL_4__12116_ (
);

FILL FILL_2__13570_ (
);

FILL FILL_4_BUFX2_insert715 (
);

FILL FILL_2__13150_ (
);

FILL FILL_4_BUFX2_insert716 (
);

FILL FILL_4_BUFX2_insert717 (
);

FILL FILL_4_BUFX2_insert718 (
);

FILL FILL_3__11949_ (
);

FILL FILL_4_BUFX2_insert719 (
);

FILL FILL_1__12983_ (
);

FILL FILL_3__11529_ (
);

FILL FILL_3__11109_ (
);

FILL FILL_1__12143_ (
);

FILL SFILL99000x77050 (
);

FILL FILL_0__9990_ (
);

FILL FILL_0__11976_ (
);

FILL SFILL69240x14050 (
);

FILL FILL_0__9150_ (
);

OR2X2 _11841_ (
    .A(_2929_),
    .B(_2923_),
    .Y(\datapath_1.ALUResult [1])
);

FILL FILL_2__9168_ (
);

FILL FILL_0__11556_ (
);

OAI22X1 _11421_ (
    .A(_2474_),
    .B(_2480_),
    .C(_2324_),
    .D(_2344__bF$buf0),
    .Y(_2537_)
);

FILL FILL_0__11136_ (
);

INVX1 _11001_ (
    .A(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2120_)
);

FILL FILL_5__7593_ (
);

FILL FILL_5__7173_ (
);

FILL FILL_5__14748_ (
);

FILL FILL_3__15782_ (
);

FILL FILL_5__14328_ (
);

FILL FILL_3__15362_ (
);

OAI21X1 _8628_ (
    .A(_887_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .C(_888_),
    .Y(_848_[20])
);

OAI21X1 _8208_ (
    .A(_668_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .C(_669_),
    .Y(_653_[8])
);

FILL FILL_1__7585_ (
);

FILL FILL_1__7165_ (
);

FILL FILL_2__14775_ (
);

FILL FILL_2__14355_ (
);

FILL SFILL99400x46050 (
);

FILL SFILL13720x50 (
);

FILL FILL_1__13768_ (
);

FILL FILL_1__13348_ (
);

FILL FILL_3__8872_ (
);

FILL FILL_3__8452_ (
);

OAI21X1 _12626_ (
    .A(_3462_),
    .B(vdd),
    .C(_3463_),
    .Y(_3425_[19])
);

NAND2X1 _12206_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [30]),
    .Y(_3191_)
);

FILL FILL_5__8378_ (
);

INVX4 _15098_ (
    .A(_5503__bF$buf1),
    .Y(_5577_)
);

FILL FILL_0__13702_ (
);

FILL FILL_3__16147_ (
);

FILL FILL_5__10668_ (
);

FILL FILL_5__10248_ (
);

FILL FILL_3__11282_ (
);

FILL FILL_0__16174_ (
);

FILL FILL_2__10695_ (
);

FILL FILL_2__10275_ (
);

FILL FILL_1__9731_ (
);

FILL FILL_3_BUFX2_insert730 (
);

FILL FILL_3__9657_ (
);

FILL FILL_3_BUFX2_insert731 (
);

FILL FILL_3__9237_ (
);

FILL FILL_3_BUFX2_insert732 (
);

FILL FILL_3_BUFX2_insert733 (
);

FILL FILL_3_BUFX2_insert734 (
);

FILL FILL_5__14081_ (
);

FILL SFILL89000x75050 (
);

FILL FILL_1__15914_ (
);

FILL FILL_3_BUFX2_insert735 (
);

OAI21X1 _8381_ (
    .A(_763_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .C(_764_),
    .Y(_718_[23])
);

FILL FILL_3_BUFX2_insert736 (
);

FILL SFILL59240x12050 (
);

FILL FILL_3_BUFX2_insert737 (
);

FILL SFILL85000x7050 (
);

FILL FILL_3_BUFX2_insert738 (
);

FILL FILL_3_BUFX2_insert739 (
);

FILL FILL_4__13494_ (
);

FILL FILL_0__14907_ (
);

FILL FILL_3__12487_ (
);

FILL FILL_2__7234_ (
);

FILL FILL_3__12067_ (
);

FILL FILL_0__12094_ (
);

FILL SFILL89400x44050 (
);

FILL SFILL28760x28050 (
);

FILL SFILL59160x19050 (
);

FILL FILL_6__16293_ (
);

FILL FILL_4__8521_ (
);

FILL FILL_4__11807_ (
);

FILL FILL_4__8101_ (
);

FILL FILL_2__12841_ (
);

FILL FILL_2__12421_ (
);

FILL FILL_5__15286_ (
);

FILL FILL_2__12001_ (
);

FILL FILL_6__8867_ (
);

DFFSR _9586_ (
    .Q(\datapath_1.regfile_1.regOut[21] [28]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_1303_[28])
);

NAND2X1 _9166_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1166_)
);

FILL FILL_4__14699_ (
);

FILL FILL_1__11834_ (
);

FILL FILL_4__14279_ (
);

FILL FILL_1__11414_ (
);

FILL FILL_0__8841_ (
);

FILL FILL_2__8859_ (
);

FILL FILL_0__10827_ (
);

FILL FILL_2__8439_ (
);

FILL FILL_0__10407_ (
);

FILL FILL_2__8019_ (
);

FILL FILL_0__8001_ (
);

FILL FILL_0_BUFX2_insert860 (
);

FILL FILL_5__6864_ (
);

FILL FILL_4__15640_ (
);

FILL FILL_0_BUFX2_insert861 (
);

FILL FILL_0_BUFX2_insert862 (
);

FILL FILL_4__15220_ (
);

FILL FILL_0_BUFX2_insert863 (
);

FILL FILL_0_BUFX2_insert864 (
);

FILL FILL_0__13299_ (
);

FILL FILL_0_BUFX2_insert865 (
);

AOI21X1 _13584_ (
    .A(_4070_),
    .B(_4093_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [2])
);

NAND2X1 _13164_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [28]),
    .Y(_3741_)
);

FILL FILL_0_BUFX2_insert866 (
);

FILL FILL_0_BUFX2_insert867 (
);

FILL FILL_2__9800_ (
);

FILL FILL_3__14633_ (
);

FILL FILL_0_BUFX2_insert868 (
);

FILL FILL_3__14213_ (
);

FILL FILL_0_BUFX2_insert869 (
);

FILL FILL_1__6856_ (
);

FILL FILL_4__9726_ (
);

FILL SFILL94280x50050 (
);

FILL FILL_2__13626_ (
);

FILL FILL_0__14660_ (
);

FILL FILL_0__14240_ (
);

FILL FILL_1__12619_ (
);

FILL FILL_2__16098_ (
);

FILL FILL_0__9626_ (
);

FILL FILL_3__7723_ (
);

FILL FILL_0__9206_ (
);

FILL FILL_3__7303_ (
);

FILL SFILL33960x46050 (
);

FILL FILL_5__7229_ (
);

FILL FILL_4__16005_ (
);

FILL FILL_6__10946_ (
);

FILL FILL_4__11980_ (
);

NAND3X1 _14789_ (
    .A(_5268_),
    .B(_5273_),
    .C(_5267_),
    .Y(_5274_)
);

INVX1 _14369_ (
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_4862_)
);

FILL FILL_4__11560_ (
);

FILL FILL_4__11140_ (
);

FILL FILL_3__15838_ (
);

FILL FILL_3__15418_ (
);

FILL FILL_1__16032_ (
);

FILL FILL_3__10973_ (
);

FILL SFILL79400x42050 (
);

FILL FILL_3__10553_ (
);

FILL SFILL18760x26050 (
);

FILL FILL_3__10133_ (
);

FILL SFILL49160x17050 (
);

FILL FILL_0__15865_ (
);

NAND2X1 _15730_ (
    .A(_6189_),
    .B(_6193_),
    .Y(_6194_)
);

FILL FILL_6_BUFX2_insert244 (
);

FILL FILL_0__15445_ (
);

NOR2X1 _15310_ (
    .A(_5783_),
    .B(_5777_),
    .Y(_5784_)
);

FILL FILL_0__15025_ (
);

FILL FILL_2__8192_ (
);

FILL FILL_0__10580_ (
);

FILL FILL_0__10160_ (
);

FILL FILL_6_BUFX2_insert249 (
);

BUFX2 BUFX2_insert20 (
    .A(_3955_),
    .Y(_3955__bF$buf1)
);

BUFX2 BUFX2_insert21 (
    .A(_3955_),
    .Y(_3955__bF$buf0)
);

BUFX2 BUFX2_insert22 (
    .A(_2462_),
    .Y(_2462__bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .A(_2462_),
    .Y(_2462__bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .A(_2462_),
    .Y(_2462__bF$buf1)
);

FILL FILL_3__8508_ (
);

BUFX2 BUFX2_insert25 (
    .A(_2462_),
    .Y(_2462__bF$buf0)
);

BUFX2 BUFX2_insert26 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf7 )
);

FILL FILL_5__13772_ (
);

BUFX2 BUFX2_insert27 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf6 )
);

FILL FILL_5__13352_ (
);

BUFX2 BUFX2_insert28 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf5 )
);

BUFX2 BUFX2_insert29 (
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf4 )
);

DFFSR _7652_ (
    .Q(\datapath_1.regfile_1.regOut[6] [14]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_328_[14])
);

OAI21X1 _7232_ (
    .A(_180_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .C(_181_),
    .Y(_133_[24])
);

FILL FILL_4__12765_ (
);

FILL FILL_4__12345_ (
);

OAI21X1 _10289_ (
    .A(_1730_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .C(_1731_),
    .Y(_1693_[19])
);

FILL FILL_2__6925_ (
);

FILL FILL_3__11758_ (
);

FILL FILL_3__11338_ (
);

FILL FILL_1__12372_ (
);

FILL FILL_2__9397_ (
);

FILL FILL_0__11785_ (
);

FILL FILL_0__11365_ (
);

INVX1 _11650_ (
    .A(_2378_),
    .Y(_2753_)
);

NOR2X1 _11230_ (
    .A(_2348_),
    .B(_2345_),
    .Y(_2349_)
);

FILL FILL_5__14977_ (
);

FILL FILL_5__14557_ (
);

FILL FILL_5__14137_ (
);

FILL FILL_3__15591_ (
);

FILL FILL_3__15171_ (
);

OAI21X1 _8857_ (
    .A(_999_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .C(_1000_),
    .Y(_978_[11])
);

DFFSR _8437_ (
    .Q(\datapath_1.regfile_1.regOut[12] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_718_[31])
);

NAND2X1 _8017_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_583_)
);

FILL FILL_2__14584_ (
);

FILL FILL_2__14164_ (
);

FILL FILL_1__13997_ (
);

FILL FILL_1__13577_ (
);

FILL FILL_1__13157_ (
);

FILL SFILL29640x65050 (
);

FILL FILL_4__14911_ (
);

FILL FILL_3__8261_ (
);

OAI21X1 _12855_ (
    .A(_3574_),
    .B(vdd),
    .C(_3575_),
    .Y(_3555_[10])
);

OAI21X1 _12435_ (
    .A(_3354_),
    .B(MemToReg_bF$buf4),
    .C(_3355_),
    .Y(\datapath_1.mux_wd3.dout [30])
);

NAND3X1 _12015_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[7]),
    .C(_3032__bF$buf0),
    .Y(_3057_)
);

FILL FILL_3__13904_ (
);

FILL FILL_5__8187_ (
);

FILL FILL_5_BUFX2_insert260 (
);

FILL FILL_5_BUFX2_insert261 (
);

FILL FILL_0__13931_ (
);

FILL FILL_5_BUFX2_insert262 (
);

FILL FILL_3__16376_ (
);

FILL FILL_0__13511_ (
);

FILL FILL_5_BUFX2_insert263 (
);

FILL FILL_5_BUFX2_insert264 (
);

FILL FILL_5__10897_ (
);

FILL FILL_5_BUFX2_insert265 (
);

FILL FILL_1__8599_ (
);

FILL FILL_5_BUFX2_insert266 (
);

FILL FILL_5_BUFX2_insert267 (
);

FILL FILL_5_BUFX2_insert1050 (
);

FILL FILL_5__10057_ (
);

FILL FILL_5_BUFX2_insert1051 (
);

FILL FILL_5_BUFX2_insert268 (
);

FILL FILL_3__11091_ (
);

FILL FILL_2__15789_ (
);

FILL FILL_5_BUFX2_insert1052 (
);

FILL FILL_5_BUFX2_insert269 (
);

FILL FILL_2__15369_ (
);

FILL FILL_5_BUFX2_insert1053 (
);

FILL FILL_5_BUFX2_insert1054 (
);

FILL FILL_5_BUFX2_insert1055 (
);

FILL FILL_5_BUFX2_insert1056 (
);

FILL FILL_5_BUFX2_insert1057 (
);

FILL FILL_5_BUFX2_insert1058 (
);

FILL FILL_5_BUFX2_insert1059 (
);

FILL FILL_1__9540_ (
);

FILL FILL_1__9120_ (
);

FILL FILL_2__16310_ (
);

FILL FILL_3__9886_ (
);

FILL FILL_3__9466_ (
);

FILL FILL_4__10831_ (
);

FILL FILL_4__10411_ (
);

FILL FILL_1__15723_ (
);

FILL FILL_1__15303_ (
);

OAI21X1 _8190_ (
    .A(_656_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_657_),
    .Y(_653_[2])
);

FILL FILL_0__14716_ (
);

FILL FILL_2__7883_ (
);

FILL FILL_2__7463_ (
);

FILL FILL_2__7043_ (
);

FILL FILL_3__12296_ (
);

FILL FILL_2__11289_ (
);

FILL FILL_5__12623_ (
);

FILL FILL_5__12203_ (
);

INVX1 _6923_ (
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_16_)
);

FILL FILL_2_BUFX2_insert390 (
);

FILL FILL_2_BUFX2_insert391 (
);

FILL FILL_2_BUFX2_insert392 (
);

FILL FILL_4__8750_ (
);

FILL FILL_4__8330_ (
);

FILL FILL_2_BUFX2_insert393 (
);

FILL FILL_2_BUFX2_insert394 (
);

FILL FILL_4__11616_ (
);

FILL FILL_2__12650_ (
);

FILL FILL_2_BUFX2_insert395 (
);

FILL FILL_2_BUFX2_insert396 (
);

FILL FILL_2__12230_ (
);

FILL FILL_5__15095_ (
);

FILL FILL_2_BUFX2_insert397 (
);

FILL FILL_0__7289_ (
);

FILL FILL_2_BUFX2_insert398 (
);

NAND2X1 _9395_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1278_)
);

FILL FILL_2_BUFX2_insert399 (
);

FILL FILL_1__11643_ (
);

FILL FILL_1__11223_ (
);

FILL FILL_4__14088_ (
);

FILL FILL_0__8650_ (
);

FILL FILL_0__10636_ (
);

FILL FILL_2__8248_ (
);

OAI21X1 _10921_ (
    .A(_2051_),
    .B(_2053_),
    .C(_2060_),
    .Y(_2061_)
);

FILL FILL_0__8230_ (
);

INVX1 _10501_ (
    .A(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_1832_)
);

FILL FILL_6__14835_ (
);

NAND3X1 _13393_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3904_),
    .C(_3903_),
    .Y(_3905_)
);

FILL FILL_5__13828_ (
);

FILL FILL_3__14862_ (
);

FILL FILL_5__13408_ (
);

FILL FILL_3__14442_ (
);

FILL FILL_3__14022_ (
);

OAI21X1 _7708_ (
    .A(_416_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_417_),
    .Y(_393_[12])
);

FILL FILL_4__9535_ (
);

FILL FILL_4__9115_ (
);

FILL FILL_2__13855_ (
);

FILL FILL_2__13435_ (
);

FILL FILL_2__13015_ (
);

FILL FILL_1__12848_ (
);

FILL FILL_1__12428_ (
);

FILL FILL_1__12008_ (
);

FILL FILL_3__7952_ (
);

FILL FILL_0__9855_ (
);

FILL FILL_0__9015_ (
);

FILL FILL_3__7112_ (
);

AOI21X1 _11706_ (
    .A(_2188_),
    .B(_2803_),
    .C(_2804_),
    .Y(_2805_)
);

FILL SFILL64520x5050 (
);

FILL FILL_5__7878_ (
);

FILL SFILL104360x34050 (
);

FILL FILL_5__7458_ (
);

FILL FILL_4__16234_ (
);

FILL FILL_5__7038_ (
);

FILL FILL_6__10755_ (
);

INVX1 _14598_ (
    .A(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_5086_)
);

NOR2X1 _14178_ (
    .A(_4674_),
    .B(_3983__bF$buf0),
    .Y(_4675_)
);

FILL FILL_3__15647_ (
);

FILL FILL_3__15227_ (
);

FILL FILL_1__16261_ (
);

FILL FILL112040x71050 (
);

FILL FILL_3__10782_ (
);

FILL FILL_3__10362_ (
);

FILL FILL_0__15674_ (
);

FILL FILL_0__15254_ (
);

FILL SFILL64040x9050 (
);

FILL FILL_3__8737_ (
);

FILL FILL_3__8317_ (
);

FILL FILL_5__13581_ (
);

FILL FILL_5__13161_ (
);

OAI21X1 _7881_ (
    .A(_511_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .C(_512_),
    .Y(_458_[27])
);

FILL FILL112440x40050 (
);

OAI21X1 _7461_ (
    .A(_292_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .C(_293_),
    .Y(_263_[15])
);

OAI21X1 _7041_ (
    .A(_73_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_74_),
    .Y(_68_[3])
);

FILL FILL_4__12994_ (
);

FILL FILL_4__12574_ (
);

FILL FILL_4__12154_ (
);

DFFSR _10098_ (
    .Q(\datapath_1.regfile_1.regOut[25] [28]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_1563_[28])
);

FILL FILL_3__11987_ (
);

FILL FILL_5__9604_ (
);

FILL FILL_3__11567_ (
);

FILL FILL_3__11147_ (
);

FILL FILL_1__12181_ (
);

FILL FILL_0__16039_ (
);

INVX1 _16324_ (
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_6770_)
);

FILL FILL_0__11594_ (
);

FILL FILL_0__11174_ (
);

FILL FILL_4__7601_ (
);

FILL FILL_2__11921_ (
);

FILL FILL_5__14786_ (
);

FILL FILL_5__14366_ (
);

FILL FILL_2__11501_ (
);

DFFSR _8666_ (
    .Q(\datapath_1.regfile_1.regOut[14] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_848_[4])
);

NAND2X1 _8246_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_695_)
);

FILL FILL_1__10914_ (
);

FILL FILL_4__13779_ (
);

FILL FILL_4__13359_ (
);

FILL FILL_2__14393_ (
);

FILL FILL_2__7939_ (
);

FILL FILL_0__7501_ (
);

FILL SFILL94680x59050 (
);

FILL FILL_1__13386_ (
);

FILL FILL_4__14720_ (
);

FILL FILL_4__14300_ (
);

FILL FILL_3__8490_ (
);

DFFSR _12664_ (
    .Q(\datapath_1.Data [1]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3425_[1])
);

FILL FILL_0__12379_ (
);

FILL FILL_3__8070_ (
);

NAND3X1 _12244_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [9]),
    .C(_3198__bF$buf3),
    .Y(_3222_)
);

FILL FILL_3__13713_ (
);

FILL FILL_2__12706_ (
);

FILL FILL_0__13740_ (
);

FILL FILL_0__13320_ (
);

FILL FILL_3__16185_ (
);

FILL FILL_5__10286_ (
);

FILL FILL_2__15598_ (
);

FILL FILL_2__15178_ (
);

FILL FILL_0__8706_ (
);

FILL SFILL94600x57050 (
);

FILL FILL_4__15925_ (
);

FILL FILL_4__15505_ (
);

INVX1 _13869_ (
    .A(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_4373_)
);

FILL FILL_3__9275_ (
);

FILL FILL_4__10640_ (
);

OAI22X1 _13449_ (
    .A(_3958_),
    .B(_3960_),
    .C(_3959_),
    .D(_3957_),
    .Y(_3961_)
);

INVX1 _13029_ (
    .A(_2_[26]),
    .Y(_3671_)
);

FILL FILL_3__14918_ (
);

FILL FILL_1__15952_ (
);

FILL FILL_1__15532_ (
);

FILL FILL_1__15112_ (
);

FILL SFILL34520x4050 (
);

FILL FILL_0__14945_ (
);

NOR2X1 _14810_ (
    .A(_5290_),
    .B(_5293_),
    .Y(_5294_)
);

FILL FILL_0__14525_ (
);

FILL FILL_0__14105_ (
);

FILL FILL_2__7692_ (
);

FILL SFILL39720x10050 (
);

FILL FILL_4__7198_ (
);

FILL FILL_2__11098_ (
);

FILL FILL_5__12852_ (
);

FILL FILL_5__12432_ (
);

FILL FILL_5__12012_ (
);

FILL SFILL8680x62050 (
);

FILL FILL_4__11845_ (
);

FILL SFILL74280x6050 (
);

FILL FILL_4__11425_ (
);

FILL FILL_4__11005_ (
);

FILL FILL_6__8485_ (
);

FILL FILL_0__7098_ (
);

FILL FILL_1__16317_ (
);

FILL FILL_1__11872_ (
);

FILL FILL_3__10418_ (
);

FILL FILL_1__11452_ (
);

FILL FILL_1__11032_ (
);

FILL SFILL84280x43050 (
);

FILL FILL_2__8897_ (
);

FILL FILL_2__8477_ (
);

FILL FILL_0__10445_ (
);

DFFSR _10730_ (
    .Q(\datapath_1.regfile_1.regOut[30] [20]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_1888_[20])
);

FILL FILL_2__8057_ (
);

OAI21X1 _10310_ (
    .A(_1744_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .C(_1745_),
    .Y(_1693_[26])
);

FILL FILL_0__10025_ (
);

FILL FILL_5__13637_ (
);

FILL FILL_5__13217_ (
);

FILL FILL_3__14671_ (
);

OAI21X1 _7937_ (
    .A(_528_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_529_),
    .Y(_523_[3])
);

FILL FILL_3__14251_ (
);

FILL SFILL8600x60050 (
);

DFFSR _7517_ (
    .Q(\datapath_1.regfile_1.regOut[5] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_263_[7])
);

FILL FILL_1__6894_ (
);

FILL FILL_4__9764_ (
);

FILL FILL_4__9344_ (
);

FILL FILL_2__13664_ (
);

FILL FILL_2__13244_ (
);

FILL FILL_1__12657_ (
);

FILL FILL_1__12237_ (
);

FILL SFILL53800x50050 (
);

FILL SFILL84200x41050 (
);

FILL FILL_0__9664_ (
);

FILL FILL_3__7761_ (
);

INVX1 _11935_ (
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_2998_)
);

FILL FILL_0__9244_ (
);

FILL FILL_3__7341_ (
);

NOR2X1 _11515_ (
    .A(_2619_),
    .B(_2626_),
    .Y(_2627_)
);

FILL FILL_5__7687_ (
);

FILL FILL_6__15429_ (
);

FILL FILL_6__15009_ (
);

FILL FILL_4__16043_ (
);

FILL SFILL13640x61050 (
);

FILL FILL_3__15876_ (
);

FILL FILL_3__15456_ (
);

FILL FILL_3__15036_ (
);

FILL FILL_1__16070_ (
);

FILL FILL_1__7679_ (
);

FILL FILL_3__10171_ (
);

FILL FILL_2__14869_ (
);

FILL FILL_6_BUFX2_insert623 (
);

FILL FILL_2__14449_ (
);

FILL FILL_2__14029_ (
);

FILL FILL_0__15483_ (
);

FILL FILL_0__15063_ (
);

FILL SFILL114440x24050 (
);

FILL FILL_6_BUFX2_insert628 (
);

FILL FILL_1__8620_ (
);

FILL FILL_1__8200_ (
);

FILL FILL_2__15810_ (
);

FILL FILL_3__8966_ (
);

FILL FILL_3__8126_ (
);

FILL FILL_5__13390_ (
);

OAI21X1 _7690_ (
    .A(_404_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .C(_405_),
    .Y(_393_[6])
);

FILL FILL_1__14803_ (
);

DFFSR _7270_ (
    .Q(\datapath_1.regfile_1.regOut[3] [16]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_133_[16])
);

FILL FILL_1_BUFX2_insert80 (
);

FILL FILL_1_BUFX2_insert81 (
);

FILL FILL_1_BUFX2_insert82 (
);

FILL FILL_1_BUFX2_insert83 (
);

FILL FILL_6__11349_ (
);

FILL FILL_4__12383_ (
);

FILL FILL_1_BUFX2_insert84 (
);

FILL FILL_1_BUFX2_insert85 (
);

FILL FILL_1_BUFX2_insert86 (
);

FILL FILL_1_BUFX2_insert87 (
);

FILL FILL_1_BUFX2_insert88 (
);

FILL FILL_1_BUFX2_insert89 (
);

FILL FILL_2__6963_ (
);

FILL FILL_3__11796_ (
);

FILL FILL_5__9413_ (
);

FILL FILL_3__11376_ (
);

FILL FILL_4__6889_ (
);

FILL FILL_0__16268_ (
);

AOI22X1 _16133_ (
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_6586_)
);

FILL FILL_2__10789_ (
);

FILL FILL_2__10369_ (
);

FILL FILL_5__11703_ (
);

FILL FILL_1__9405_ (
);

FILL FILL_4__7830_ (
);

FILL FILL_5__14595_ (
);

FILL FILL_2__11730_ (
);

FILL FILL_5__14175_ (
);

FILL FILL_2__11310_ (
);

NAND2X1 _8895_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1026_)
);

FILL FILL_6__7756_ (
);

NAND2X1 _8475_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_807_)
);

NAND2X1 _8055_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .Y(_652_)
);

FILL FILL_4__13588_ (
);

FILL FILL_1__10303_ (
);

FILL FILL_4__13168_ (
);

FILL FILL_0__7730_ (
);

FILL FILL_2__7748_ (
);

FILL FILL_0__7310_ (
);

FILL FILL_2__7328_ (
);

NAND2X1 _12893_ (
    .A(vdd),
    .B(\datapath_1.rd1 [23]),
    .Y(_3601_)
);

FILL FILL_0__12188_ (
);

NAND2X1 _12473_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [11]),
    .Y(_3382_)
);

FILL FILL_5__12908_ (
);

AOI22X1 _12053_ (
    .A(\datapath_1.ALUResult [16]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3086_)
);

FILL FILL_3__13942_ (
);

FILL FILL_3__13522_ (
);

FILL FILL_3__13102_ (
);

FILL FILL_4__8615_ (
);

FILL FILL_5_BUFX2_insert640 (
);

FILL FILL_5_BUFX2_insert641 (
);

FILL FILL_2__12515_ (
);

FILL FILL_5_BUFX2_insert642 (
);

FILL FILL_5_BUFX2_insert643 (
);

FILL SFILL64200x82050 (
);

FILL FILL_5_BUFX2_insert644 (
);

FILL FILL_5_BUFX2_insert645 (
);

FILL FILL_5_BUFX2_insert646 (
);

FILL FILL_5_BUFX2_insert647 (
);

FILL FILL_5_BUFX2_insert648 (
);

FILL FILL_1__11928_ (
);

FILL FILL_5_BUFX2_insert649 (
);

FILL FILL_1__11508_ (
);

FILL FILL_5__16321_ (
);

FILL FILL_0__8515_ (
);

FILL FILL_5__6958_ (
);

FILL FILL_4__15734_ (
);

FILL FILL_4__15314_ (
);

INVX1 _13678_ (
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_4186_)
);

FILL FILL_3__9084_ (
);

OAI21X1 _13258_ (
    .A(_3759_),
    .B(_3799_),
    .C(_3800_),
    .Y(_3801_)
);

FILL FILL_3__14727_ (
);

FILL FILL_3__14307_ (
);

FILL FILL_1__15761_ (
);

FILL FILL_1__15341_ (
);

FILL FILL112040x66050 (
);

FILL FILL_0__14754_ (
);

FILL FILL_0__14334_ (
);

FILL FILL_2__7081_ (
);

FILL FILL_3__7817_ (
);

FILL FILL_5__12661_ (
);

FILL FILL_5__12241_ (
);

FILL FILL112440x35050 (
);

OAI21X1 _6961_ (
    .A(_40_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_41_),
    .Y(_3_[19])
);

FILL FILL_2_BUFX2_insert770 (
);

FILL FILL_2_BUFX2_insert771 (
);

FILL FILL_2_BUFX2_insert772 (
);

FILL FILL_2_BUFX2_insert773 (
);

FILL FILL_2_BUFX2_insert774 (
);

FILL FILL_4__11654_ (
);

FILL FILL_4__11234_ (
);

FILL FILL_2_BUFX2_insert775 (
);

FILL FILL_2_BUFX2_insert776 (
);

FILL FILL_2_BUFX2_insert777 (
);

FILL FILL_2_BUFX2_insert778 (
);

FILL FILL_2_BUFX2_insert779 (
);

FILL FILL_1__16126_ (
);

FILL FILL_3__10647_ (
);

FILL FILL_1__11681_ (
);

FILL SFILL85080x42050 (
);

FILL FILL_1__11261_ (
);

FILL FILL_0__15959_ (
);

FILL FILL112040x21050 (
);

FILL FILL_0__15539_ (
);

NAND3X1 _15824_ (
    .A(_6283_),
    .B(_6284_),
    .C(_6282_),
    .Y(_6285_)
);

OAI22X1 _15404_ (
    .A(_5874_),
    .B(_5548__bF$buf0),
    .C(_5489__bF$buf1),
    .D(_5875_),
    .Y(_5876_)
);

FILL FILL_0__15119_ (
);

FILL FILL_0__10674_ (
);

FILL FILL_0__10254_ (
);

FILL FILL_5__13866_ (
);

FILL FILL_5__13446_ (
);

FILL FILL_3__14480_ (
);

FILL FILL_5__13026_ (
);

FILL FILL_3__14060_ (
);

NAND2X1 _7746_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_443_)
);

NAND2X1 _7326_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_224_)
);

FILL FILL_4__9993_ (
);

FILL FILL_4__12859_ (
);

FILL FILL_4__9153_ (
);

FILL FILL_4__12439_ (
);

FILL FILL_2__13893_ (
);

FILL FILL_4__12019_ (
);

FILL FILL_2__13473_ (
);

FILL FILL_1__12886_ (
);

FILL FILL_1__12466_ (
);

FILL FILL_1__12046_ (
);

FILL FILL_4__13800_ (
);

FILL FILL_3__7990_ (
);

FILL FILL_6_CLKBUF1_insert224 (
);

FILL FILL_0__9893_ (
);

FILL FILL_0__9473_ (
);

FILL FILL_0__11879_ (
);

FILL FILL_3__7570_ (
);

AOI21X1 _11744_ (
    .A(_2838_),
    .B(_2169_),
    .C(_2839_),
    .Y(_2840_)
);

FILL FILL_0__11459_ (
);

FILL FILL_0__11039_ (
);

NAND2X1 _11324_ (
    .A(_2296_),
    .B(_2442_),
    .Y(_2443_)
);

FILL FILL_5__7496_ (
);

FILL FILL_5__7076_ (
);

FILL FILL_4__16272_ (
);

FILL FILL_6__10373_ (
);

FILL FILL_3__15685_ (
);

FILL FILL_0__12400_ (
);

FILL FILL_3__15265_ (
);

FILL FILL_1__7488_ (
);

FILL FILL_1__7068_ (
);

FILL FILL_2__14678_ (
);

FILL FILL_2__14258_ (
);

FILL FILL_0__15292_ (
);

FILL SFILL13640x1050 (
);

FILL SFILL23720x51050 (
);

FILL FILL_1_BUFX2_insert790 (
);

FILL FILL_1_BUFX2_insert791 (
);

FILL FILL_3__8775_ (
);

FILL SFILL37960x23050 (
);

FILL FILL_3__8355_ (
);

FILL FILL_1_BUFX2_insert792 (
);

DFFSR _12949_ (
    .Q(\datapath_1.a [30]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_3555_[30])
);

INVX1 _12529_ (
    .A(ALUOut[30]),
    .Y(_3419_)
);

FILL FILL_1_BUFX2_insert793 (
);

FILL FILL_1_BUFX2_insert794 (
);

AOI22X1 _12109_ (
    .A(\datapath_1.ALUResult [30]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3128_)
);

FILL FILL_1_BUFX2_insert795 (
);

FILL FILL_1_BUFX2_insert796 (
);

FILL FILL_1__14612_ (
);

FILL FILL_1_BUFX2_insert797 (
);

FILL FILL_1_BUFX2_insert798 (
);

FILL FILL_1_BUFX2_insert799 (
);

FILL FILL_6__11998_ (
);

FILL FILL_4__12192_ (
);

FILL FILL_0__13605_ (
);

FILL FILL_5__9642_ (
);

FILL FILL_5__9222_ (
);

FILL FILL_3__11185_ (
);

FILL FILL_0__16077_ (
);

OAI21X1 _16362_ (
    .A(_6794_),
    .B(gnd),
    .C(_6795_),
    .Y(_6769_[13])
);

FILL FILL_2__10178_ (
);

FILL FILL_5__11932_ (
);

FILL FILL_1__9634_ (
);

FILL FILL_5__11512_ (
);

FILL FILL_1__9214_ (
);

FILL FILL_2__16404_ (
);

FILL FILL_4__10925_ (
);

FILL SFILL109560x74050 (
);

FILL FILL_4__10505_ (
);

FILL SFILL23240x44050 (
);

FILL FILL_6__7565_ (
);

FILL FILL_1__15817_ (
);

DFFSR _8284_ (
    .Q(\datapath_1.regfile_1.regOut[11] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_653_[6])
);

FILL FILL_1__10952_ (
);

FILL FILL_1__10532_ (
);

FILL FILL_4__13397_ (
);

FILL FILL_1__10112_ (
);

FILL SFILL84280x38050 (
);

FILL FILL_2__7977_ (
);

BUFX2 BUFX2_insert460 (
    .A(_5524_),
    .Y(_5524__bF$buf3)
);

FILL FILL_2__7557_ (
);

BUFX2 BUFX2_insert461 (
    .A(_5524_),
    .Y(_5524__bF$buf2)
);

BUFX2 BUFX2_insert462 (
    .A(_5524_),
    .Y(_5524__bF$buf1)
);

BUFX2 BUFX2_insert463 (
    .A(_5524_),
    .Y(_5524__bF$buf0)
);

BUFX2 BUFX2_insert464 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf7 )
);

BUFX2 BUFX2_insert465 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf6 )
);

BUFX2 BUFX2_insert466 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf5 )
);

BUFX2 BUFX2_insert467 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf4 )
);

BUFX2 BUFX2_insert468 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf3 )
);

BUFX2 BUFX2_insert469 (
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf2 )
);

NAND3X1 _12282_ (
    .A(_3248_),
    .B(_3249_),
    .C(_3250_),
    .Y(\datapath_1.alu_1.ALUInB [16])
);

FILL FILL_5__12717_ (
);

FILL FILL_3__13751_ (
);

FILL SFILL8600x55050 (
);

FILL FILL_3__13331_ (
);

FILL FILL_6__16196_ (
);

FILL FILL_4__8844_ (
);

FILL FILL_4__8004_ (
);

FILL SFILL8680x12050 (
);

FILL FILL_2__12744_ (
);

FILL FILL_5__15189_ (
);

FILL FILL_2__12324_ (
);

INVX1 _9489_ (
    .A(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_1320_)
);

DFFSR _9069_ (
    .Q(\datapath_1.regfile_1.regOut[17] [23]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_1043_[23])
);

FILL FILL_1__11737_ (
);

FILL FILL_1__11317_ (
);

FILL FILL_3__6841_ (
);

FILL FILL_0__8744_ (
);

FILL FILL_5__16130_ (
);

FILL FILL_0__8324_ (
);

FILL FILL_4__15963_ (
);

FILL FILL_4__15543_ (
);

FILL FILL_4__15123_ (
);

FILL SFILL13640x56050 (
);

INVX8 _13487_ (
    .A(_3960_),
    .Y(_3998_)
);

DFFSR _13067_ (
    .Q(_2_[20]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3620_[20])
);

FILL FILL_3__14956_ (
);

FILL FILL_1__15990_ (
);

FILL FILL_3__14536_ (
);

FILL FILL_1__15570_ (
);

FILL FILL_3__14116_ (
);

FILL FILL_1__15150_ (
);

FILL FILL_4__9629_ (
);

FILL FILL_4__9209_ (
);

FILL SFILL8600x10050 (
);

FILL FILL_2__13949_ (
);

FILL FILL_0__14983_ (
);

FILL FILL_2__13529_ (
);

FILL FILL_0__14563_ (
);

FILL FILL_2__13109_ (
);

FILL FILL_0__14143_ (
);

FILL FILL_1__7700_ (
);

FILL SFILL74200x79050 (
);

FILL FILL_3__7626_ (
);

FILL FILL_0__9529_ (
);

FILL FILL_3__7206_ (
);

FILL FILL_0__9109_ (
);

FILL FILL_5__12890_ (
);

FILL FILL_5__12470_ (
);

FILL FILL_5__12050_ (
);

FILL FILL_4__16328_ (
);

FILL FILL_6__10429_ (
);

FILL FILL_4__11883_ (
);

FILL FILL_4__11463_ (
);

FILL FILL_4__11043_ (
);

FILL FILL_1__16355_ (
);

FILL SFILL13640x11050 (
);

FILL FILL_3__10876_ (
);

FILL FILL_5__8913_ (
);

FILL FILL_1__11490_ (
);

FILL FILL_3__10036_ (
);

FILL FILL_1__11070_ (
);

FILL FILL_0__15768_ (
);

FILL FILL_0__15348_ (
);

OAI22X1 _15633_ (
    .A(_5480__bF$buf3),
    .B(_4653_),
    .C(_4635_),
    .D(_5499__bF$buf1),
    .Y(_6099_)
);

NOR3X1 _15213_ (
    .A(_4160_),
    .B(_5509_),
    .C(_5688_),
    .Y(_5689_)
);

FILL SFILL38840x60050 (
);

FILL FILL_2__8095_ (
);

FILL FILL_0__10063_ (
);

FILL FILL_1__8905_ (
);

FILL FILL_6__14682_ (
);

FILL FILL_6__14262_ (
);

FILL FILL_4__6910_ (
);

FILL FILL_5__13675_ (
);

FILL FILL_2__10810_ (
);

FILL SFILL74200x34050 (
);

FILL FILL_5__13255_ (
);

NAND2X1 _7975_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_555_)
);

NAND2X1 _7555_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_336_)
);

DFFSR _7135_ (
    .Q(\datapath_1.regfile_1.regOut[2] [9]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_68_[9])
);

FILL FILL_4__9382_ (
);

FILL FILL_4__12248_ (
);

FILL FILL_2__13282_ (
);

FILL FILL_1__12695_ (
);

FILL FILL_1__12275_ (
);

FILL SFILL99480x40050 (
);

DFFSR _16418_ (
    .Q(\datapath_1.regfile_1.regOut[0] [1]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_6769_[1])
);

OAI21X1 _11973_ (
    .A(_3022_),
    .B(IorD_bF$buf5),
    .C(_3023_),
    .Y(_1_[28])
);

FILL FILL_0__11688_ (
);

FILL FILL_0__9282_ (
);

OAI21X1 _11553_ (
    .A(_2660_),
    .B(_2231_),
    .C(_2470__bF$buf2),
    .Y(_2662_)
);

FILL FILL_0__11268_ (
);

FILL FILL_5_CLKBUF1_insert210 (
);

NOR2X1 _11133_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2252_)
);

FILL FILL_5_CLKBUF1_insert211 (
);

FILL FILL_3__12602_ (
);

FILL FILL_5_CLKBUF1_insert212 (
);

FILL FILL_5_CLKBUF1_insert213 (
);

FILL FILL_5_CLKBUF1_insert214 (
);

FILL FILL_4__16081_ (
);

FILL FILL_5_CLKBUF1_insert215 (
);

FILL FILL_5_CLKBUF1_insert216 (
);

FILL FILL_5_CLKBUF1_insert217 (
);

FILL FILL_5_CLKBUF1_insert218 (
);

FILL FILL_5_CLKBUF1_insert219 (
);

FILL SFILL64200x77050 (
);

FILL FILL_3__15494_ (
);

FILL FILL_3__15074_ (
);

FILL FILL112120x54050 (
);

FILL FILL_1__7297_ (
);

FILL FILL_2__14487_ (
);

FILL FILL_2__14067_ (
);

FILL FILL_5__15821_ (
);

FILL FILL_5__15401_ (
);

DFFSR _9701_ (
    .Q(\datapath_1.regfile_1.regOut[22] [15]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_1368_[15])
);

FILL FILL_4__14814_ (
);

FILL FILL_3__8584_ (
);

INVX1 _12758_ (
    .A(\datapath_1.PCJump [23]),
    .Y(_3531_)
);

NAND3X1 _12338_ (
    .A(_3290_),
    .B(_3291_),
    .C(_3292_),
    .Y(\datapath_1.alu_1.ALUInB [30])
);

FILL FILL_3__13807_ (
);

FILL FILL_1__14841_ (
);

FILL FILL_1__14421_ (
);

FILL FILL_1__14001_ (
);

FILL FILL_0__13834_ (
);

FILL FILL_0__13414_ (
);

FILL FILL_3__16279_ (
);

FILL FILL_5__9871_ (
);

FILL SFILL33800x41050 (
);

FILL SFILL89880x52050 (
);

FILL FILL_5__9031_ (
);

NOR2X1 _16171_ (
    .A(_6620_),
    .B(_6622_),
    .Y(_6623_)
);

FILL FILL_5__11741_ (
);

FILL FILL_1__9863_ (
);

FILL FILL_5__11321_ (
);

FILL FILL_1__9023_ (
);

FILL FILL_3__9789_ (
);

FILL FILL_2__16213_ (
);

FILL FILL_3__9369_ (
);

FILL FILL_4__10314_ (
);

FILL FILL_1__15626_ (
);

FILL SFILL33720x48050 (
);

FILL FILL_1__15206_ (
);

INVX1 _8093_ (
    .A(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_613_)
);

FILL FILL_1__10761_ (
);

FILL FILL_0__14619_ (
);

OAI22X1 _14904_ (
    .A(_5384_),
    .B(_3936__bF$buf1),
    .C(_3935__bF$buf0),
    .D(_5385_),
    .Y(_5386_)
);

FILL FILL_2__7366_ (
);

FILL FILL_3__12199_ (
);

NAND3X1 _12091_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[26]),
    .C(_3032__bF$buf4),
    .Y(_3114_)
);

FILL FILL_5__12526_ (
);

FILL FILL_3__13980_ (
);

FILL FILL_5__12106_ (
);

FILL FILL_3__13560_ (
);

FILL FILL_3__13140_ (
);

FILL FILL_4__8653_ (
);

FILL FILL_4__11939_ (
);

FILL FILL_4__8233_ (
);

FILL FILL_2__12973_ (
);

FILL FILL_4__11519_ (
);

FILL FILL_2__12133_ (
);

OAI21X1 _9298_ (
    .A(_1232_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1233_),
    .Y(_1173_[30])
);

FILL FILL_1__11966_ (
);

FILL FILL_1__11546_ (
);

FILL FILL_1__11126_ (
);

FILL FILL_0__8973_ (
);

FILL FILL_0__10959_ (
);

FILL FILL_0__10539_ (
);

FILL FILL_0__8133_ (
);

NAND2X1 _10824_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_2007_)
);

FILL FILL_6__9100_ (
);

NAND2X1 _10404_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1788_)
);

FILL FILL_0__10119_ (
);

FILL FILL_5__6996_ (
);

FILL FILL_6__14738_ (
);

FILL FILL_4__15772_ (
);

FILL FILL_4__15352_ (
);

NAND2X1 _13296_ (
    .A(_3832_),
    .B(_3828_),
    .Y(_3833_)
);

FILL FILL_2__9932_ (
);

FILL FILL_2__9512_ (
);

FILL FILL_0__11900_ (
);

FILL FILL_3__14765_ (
);

FILL FILL_3__14345_ (
);

FILL FILL_1__6988_ (
);

FILL FILL_4__9858_ (
);

FILL FILL_4__9018_ (
);

FILL FILL_2__13758_ (
);

FILL FILL_2__13338_ (
);

FILL FILL_0__14792_ (
);

FILL FILL_0__14372_ (
);

FILL SFILL23720x46050 (
);

FILL FILL_3__7855_ (
);

FILL FILL_0__9758_ (
);

FILL FILL_3__7435_ (
);

FILL FILL_0__9338_ (
);

NAND3X1 _11609_ (
    .A(_2692_),
    .B(_2424_),
    .C(_2703_),
    .Y(_2715_)
);

FILL FILL_4__16137_ (
);

FILL FILL_6__10238_ (
);

FILL FILL_4__11692_ (
);

FILL FILL_4__11272_ (
);

FILL SFILL23320x32050 (
);

FILL FILL_1__16164_ (
);

FILL FILL_3__10685_ (
);

FILL FILL_5__8722_ (
);

FILL FILL_3__10265_ (
);

FILL FILL_0__15997_ (
);

AOI21X1 _15862_ (
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .B(_5649_),
    .C(_6321_),
    .Y(_6322_)
);

FILL FILL_0__15577_ (
);

INVX1 _15442_ (
    .A(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_5913_)
);

FILL FILL_0__15157_ (
);

OAI22X1 _15022_ (
    .A(_5498_),
    .B(_5501_),
    .C(_5499__bF$buf1),
    .D(_3957_),
    .Y(_5502_)
);

FILL FILL_0__10292_ (
);

FILL FILL_1__8714_ (
);

FILL FILL_2__15904_ (
);

FILL SFILL109560x69050 (
);

FILL FILL_5__13484_ (
);

DFFSR _7784_ (
    .Q(\datapath_1.regfile_1.regOut[7] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_393_[18])
);

INVX1 _7364_ (
    .A(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_249_)
);

FILL FILL_4__12897_ (
);

FILL FILL_4__12477_ (
);

FILL FILL_4__12057_ (
);

FILL FILL_2__13091_ (
);

FILL FILL_5_BUFX2_insert30 (
);

FILL FILL_5_BUFX2_insert31 (
);

FILL FILL_5__9927_ (
);

FILL FILL_5__9507_ (
);

FILL FILL_5_BUFX2_insert32 (
);

FILL FILL_5_BUFX2_insert33 (
);

FILL FILL_5_BUFX2_insert34 (
);

FILL FILL_1__12084_ (
);

FILL FILL_5_BUFX2_insert35 (
);

FILL FILL_5_BUFX2_insert36 (
);

INVX1 _16227_ (
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_6678_)
);

FILL FILL_5_BUFX2_insert37 (
);

FILL FILL_5_BUFX2_insert38 (
);

FILL FILL_5_BUFX2_insert39 (
);

FILL FILL_0__9091_ (
);

OAI21X1 _11782_ (
    .A(_2863_),
    .B(_2558_),
    .C(_2470__bF$buf3),
    .Y(_2876_)
);

FILL FILL_0__11497_ (
);

INVX1 _11362_ (
    .A(_2320_),
    .Y(_2479_)
);

FILL FILL_0__11077_ (
);

FILL FILL_1__9919_ (
);

FILL FILL_3__12831_ (
);

FILL FILL_3__12411_ (
);

FILL FILL_4__7504_ (
);

FILL FILL_4_CLKBUF1_insert200 (
);

FILL SFILL13720x44050 (
);

FILL FILL_4_CLKBUF1_insert201 (
);

FILL FILL_2__11824_ (
);

FILL FILL_5__14689_ (
);

FILL FILL_4_CLKBUF1_insert202 (
);

FILL FILL_5__14269_ (
);

FILL FILL_2__11404_ (
);

FILL FILL_4_CLKBUF1_insert203 (
);

INVX1 _8989_ (
    .A(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_1068_)
);

INVX1 _8569_ (
    .A(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_849_)
);

FILL FILL_4_CLKBUF1_insert204 (
);

FILL FILL_4_CLKBUF1_insert205 (
);

OAI21X1 _8149_ (
    .A(_649_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_650_),
    .Y(_588_[31])
);

FILL FILL_4_CLKBUF1_insert206 (
);

FILL FILL_4_CLKBUF1_insert207 (
);

FILL FILL_4_CLKBUF1_insert208 (
);

FILL FILL_1__10817_ (
);

FILL FILL_4_CLKBUF1_insert209 (
);

FILL FILL_2__14296_ (
);

FILL FILL_5__15630_ (
);

FILL FILL_0__7824_ (
);

FILL FILL_5__15210_ (
);

INVX1 _9930_ (
    .A(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_1553_)
);

INVX1 _9510_ (
    .A(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_1334_)
);

FILL FILL_1__13289_ (
);

FILL FILL_4__14623_ (
);

FILL FILL_4__14203_ (
);

INVX1 _12987_ (
    .A(_2_[12]),
    .Y(_3643_)
);

FILL FILL_3__8393_ (
);

INVX1 _12567_ (
    .A(\datapath_1.Data [0]),
    .Y(_3488_)
);

OAI21X1 _12147_ (
    .A(_3150_),
    .B(ALUSrcA_bF$buf0),
    .C(_3151_),
    .Y(\datapath_1.alu_1.ALUInA [10])
);

FILL FILL_3__13616_ (
);

FILL FILL_1__14650_ (
);

FILL FILL_1__14230_ (
);

FILL FILL_0_BUFX2_insert100 (
);

FILL FILL_4__8709_ (
);

FILL FILL_0_BUFX2_insert101 (
);

FILL FILL_0_BUFX2_insert102 (
);

FILL FILL_2__12609_ (
);

FILL FILL_0_BUFX2_insert103 (
);

FILL FILL_0__13643_ (
);

FILL FILL_0_BUFX2_insert104 (
);

FILL FILL_0__13223_ (
);

FILL FILL_0_BUFX2_insert105 (
);

FILL FILL_3__16088_ (
);

FILL FILL_0_BUFX2_insert106 (
);

FILL SFILL48840x12050 (
);

FILL FILL_0_BUFX2_insert107 (
);

FILL FILL_5__10189_ (
);

FILL FILL_0_BUFX2_insert108 (
);

FILL FILL_5__9680_ (
);

FILL FILL_0_BUFX2_insert109 (
);

FILL FILL_5__9260_ (
);

FILL FILL_5__16415_ (
);

FILL FILL_0__8609_ (
);

FILL FILL_5__11970_ (
);

FILL FILL_1__9672_ (
);

FILL FILL_5__11550_ (
);

FILL FILL_1__9252_ (
);

FILL FILL_5__11130_ (
);

FILL FILL_4__15828_ (
);

FILL FILL_4__15408_ (
);

BUFX2 BUFX2_insert1020 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf6 )
);

BUFX2 BUFX2_insert1021 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf5 )
);

BUFX2 BUFX2_insert1022 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf4 )
);

FILL FILL_2__16022_ (
);

FILL FILL_3__9598_ (
);

FILL FILL_4__10963_ (
);

BUFX2 BUFX2_insert1023 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf3 )
);

BUFX2 BUFX2_insert1024 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf2 )
);

FILL FILL_4__10543_ (
);

BUFX2 BUFX2_insert1025 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf1 )
);

FILL FILL_4__10123_ (
);

BUFX2 BUFX2_insert1026 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf0 )
);

FILL FILL_1__15855_ (
);

BUFX2 BUFX2_insert1027 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf7 )
);

FILL FILL_6__7183_ (
);

BUFX2 BUFX2_insert1028 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf6 )
);

FILL FILL_1__15435_ (
);

BUFX2 BUFX2_insert1029 (
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf5 )
);

FILL FILL_1__15015_ (
);

FILL FILL_1__10990_ (
);

FILL FILL_1__10570_ (
);

FILL FILL_1__10150_ (
);

FILL FILL_0__14848_ (
);

AOI22X1 _14713_ (
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .B(_4102_),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_5199_)
);

FILL FILL_0__14428_ (
);

FILL FILL_0__14008_ (
);

FILL SFILL38840x55050 (
);

FILL FILL_2__7595_ (
);

BUFX2 BUFX2_insert840 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf2 )
);

BUFX2 BUFX2_insert841 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf1 )
);

FILL FILL_2__7175_ (
);

BUFX2 BUFX2_insert842 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf0 )
);

BUFX2 BUFX2_insert843 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf4 )
);

BUFX2 BUFX2_insert844 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf3 )
);

BUFX2 BUFX2_insert845 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf2 )
);

BUFX2 BUFX2_insert846 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf1 )
);

BUFX2 BUFX2_insert847 (
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf0 )
);

BUFX2 BUFX2_insert848 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf7 )
);

BUFX2 BUFX2_insert849 (
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf6 )
);

FILL SFILL74200x29050 (
);

FILL FILL_5__12755_ (
);

FILL FILL_5__12335_ (
);

FILL FILL_4__8882_ (
);

FILL FILL_4__8462_ (
);

FILL FILL_4__11748_ (
);

FILL FILL_2__12782_ (
);

FILL FILL_4__11328_ (
);

FILL FILL_2__12362_ (
);

FILL FILL112200x42050 (
);

FILL FILL_1__11775_ (
);

FILL SFILL99480x35050 (
);

FILL FILL_1__11355_ (
);

NAND3X1 _15918_ (
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6377_)
);

FILL FILL_0__8782_ (
);

FILL FILL_0__10768_ (
);

FILL FILL_0__8362_ (
);

FILL SFILL3480x54050 (
);

NAND2X1 _10633_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1900_)
);

DFFSR _10213_ (
    .Q(\datapath_1.regfile_1.regOut[26] [15]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1628_[15])
);

FILL FILL_4__15581_ (
);

FILL FILL_4__15161_ (
);

FILL FILL_2__9741_ (
);

FILL FILL_3__14994_ (
);

FILL FILL_3__14574_ (
);

FILL FILL_3__14154_ (
);

FILL FILL112120x49050 (
);

FILL FILL_4_BUFX2_insert680 (
);

FILL FILL_4_BUFX2_insert681 (
);

FILL FILL_4__9667_ (
);

FILL FILL_4_BUFX2_insert682 (
);

FILL FILL_4__9247_ (
);

FILL FILL_2__13987_ (
);

FILL FILL_4_BUFX2_insert683 (
);

FILL FILL_4_BUFX2_insert684 (
);

FILL FILL_2__13567_ (
);

FILL FILL_2__13147_ (
);

FILL FILL_4_BUFX2_insert685 (
);

FILL FILL_0__14181_ (
);

FILL FILL_4_BUFX2_insert686 (
);

FILL FILL_4_BUFX2_insert687 (
);

FILL FILL_5__14901_ (
);

FILL FILL_4_BUFX2_insert688 (
);

FILL FILL_4_BUFX2_insert689 (
);

FILL FILL_0__9987_ (
);

FILL FILL_0__9147_ (
);

FILL FILL_3__7244_ (
);

NAND2X1 _11838_ (
    .A(_2926_),
    .B(_2920_),
    .Y(_2927_)
);

OAI21X1 _11418_ (
    .A(_2476_),
    .B(_2477_),
    .C(_2534_),
    .Y(\datapath_1.ALUResult [29])
);

FILL FILL_1__13921_ (
);

FILL SFILL28840x53050 (
);

FILL FILL_4__16366_ (
);

FILL FILL_1__13501_ (
);

FILL SFILL24120x31050 (
);

FILL FILL_4__11081_ (
);

FILL FILL_3__15779_ (
);

FILL FILL_0__12914_ (
);

FILL FILL_3__15359_ (
);

FILL FILL_1__16393_ (
);

FILL SFILL33800x36050 (
);

FILL FILL_5__8951_ (
);

FILL SFILL64200x27050 (
);

FILL FILL_5__8531_ (
);

FILL FILL_3__10494_ (
);

FILL FILL_5__8111_ (
);

FILL FILL_0__15386_ (
);

INVX1 _15671_ (
    .A(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_6136_)
);

INVX1 _15251_ (
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_5727_)
);

FILL FILL_3__16300_ (
);

FILL FILL_5__10821_ (
);

FILL FILL_5__10401_ (
);

FILL FILL_1__8523_ (
);

FILL FILL_1__8103_ (
);

FILL FILL_2__15713_ (
);

FILL FILL_3__8869_ (
);

FILL SFILL89480x33050 (
);

FILL FILL_3__8449_ (
);

FILL FILL_5__13293_ (
);

FILL FILL_1__14706_ (
);

FILL FILL_4_BUFX2_insert1060 (
);

INVX1 _7593_ (
    .A(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_361_)
);

FILL FILL_4_BUFX2_insert1061 (
);

INVX1 _7173_ (
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_142_)
);

FILL FILL_4_BUFX2_insert1062 (
);

FILL FILL_4_BUFX2_insert1063 (
);

FILL SFILL113960x38050 (
);

FILL FILL_4_BUFX2_insert1064 (
);

FILL FILL_4__12286_ (
);

FILL FILL_4_BUFX2_insert1065 (
);

FILL FILL_4_BUFX2_insert1066 (
);

FILL FILL_3__9810_ (
);

FILL FILL_4_BUFX2_insert1067 (
);

FILL FILL_4_BUFX2_insert1068 (
);

FILL FILL_4_BUFX2_insert1069 (
);

FILL FILL_2__6866_ (
);

FILL FILL_5__9736_ (
);

FILL FILL_3__11699_ (
);

FILL FILL_3__11279_ (
);

OAI21X1 _16036_ (
    .A(_5530__bF$buf3),
    .B(_6490_),
    .C(_6491_),
    .Y(_6492_)
);

OAI22X1 _11591_ (
    .A(_2246_),
    .B(_2347__bF$buf1),
    .C(_2245_),
    .D(_2346_),
    .Y(_2698_)
);

NAND2X1 _11171_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2290_)
);

FILL FILL_1__9728_ (
);

FILL FILL_5__11606_ (
);

FILL FILL_3__12640_ (
);

FILL FILL_3__12220_ (
);

FILL FILL_4__7733_ (
);

FILL FILL_4__7313_ (
);

FILL FILL_5__14498_ (
);

FILL FILL_2__11633_ (
);

FILL FILL_2__11213_ (
);

FILL FILL_5__14078_ (
);

DFFSR _8798_ (
    .Q(\datapath_1.regfile_1.regOut[15] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_913_[8])
);

OAI21X1 _8378_ (
    .A(_761_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .C(_762_),
    .Y(_718_[22])
);

FILL FILL_6__7239_ (
);

FILL FILL_1__10626_ (
);

FILL SFILL18840x51050 (
);

FILL FILL_0__7633_ (
);

FILL FILL_0__7213_ (
);

FILL FILL_1__13098_ (
);

FILL FILL_4__14852_ (
);

FILL FILL_4__14432_ (
);

FILL FILL_4__14012_ (
);

DFFSR _12796_ (
    .Q(\aluControl_1.inst [5]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3490_[5])
);

INVX1 _12376_ (
    .A(ALUOut[11]),
    .Y(_3316_)
);

FILL FILL_3__13845_ (
);

FILL FILL_3__13425_ (
);

FILL FILL_3__13005_ (
);

FILL FILL_4__8518_ (
);

FILL FILL_2__12838_ (
);

FILL FILL_0__13872_ (
);

FILL FILL_2__12418_ (
);

FILL FILL_0__13452_ (
);

FILL FILL_0__13032_ (
);

FILL FILL_5__16224_ (
);

FILL FILL_3__6935_ (
);

FILL FILL_0__8838_ (
);

FILL FILL_1__9481_ (
);

FILL FILL_4__15637_ (
);

FILL FILL_4__15217_ (
);

FILL FILL_2__16251_ (
);

FILL FILL_4__10772_ (
);

FILL FILL_1__15664_ (
);

FILL FILL_1__15244_ (
);

FILL FILL_5__7802_ (
);

AOI21X1 _14942_ (
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .B(_3894_),
    .C(_5422_),
    .Y(_5423_)
);

FILL FILL_0__14657_ (
);

FILL FILL_0__14237_ (
);

AOI21X1 _14522_ (
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .B(_3995__bF$buf3),
    .C(_5011_),
    .Y(_5012_)
);

INVX1 _14102_ (
    .A(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_4601_)
);

FILL FILL_6__13991_ (
);

FILL FILL_6__13151_ (
);

FILL FILL_5__12984_ (
);

FILL FILL_5__12144_ (
);

BUFX2 _6864_ (
    .A(_1_[26]),
    .Y(memoryAddress[26])
);

FILL SFILL69080x60050 (
);

FILL FILL_4__8271_ (
);

FILL FILL_4__11977_ (
);

FILL FILL_4__11557_ (
);

FILL FILL_2__12591_ (
);

FILL FILL_4__11137_ (
);

FILL FILL_2__12171_ (
);

FILL FILL_1__16449_ (
);

FILL FILL_1__16029_ (
);

FILL FILL_1__11584_ (
);

FILL FILL_1__11164_ (
);

INVX1 _15727_ (
    .A(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_6191_)
);

OAI22X1 _15307_ (
    .A(_4279_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf1),
    .D(_4253_),
    .Y(_5781_)
);

FILL FILL_0__8591_ (
);

FILL FILL_0__10997_ (
);

DFFSR _10862_ (
    .Q(\datapath_1.regfile_1.regOut[31] [24]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_1953_[24])
);

FILL FILL_0__10577_ (
);

FILL FILL_2__8189_ (
);

INVX1 _10442_ (
    .A(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_1813_)
);

FILL FILL_0__10157_ (
);

INVX1 _10022_ (
    .A(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_1594_)
);

FILL FILL_3__11911_ (
);

FILL FILL_4__15390_ (
);

FILL SFILL13720x39050 (
);

FILL FILL_2__10904_ (
);

FILL FILL_5__13769_ (
);

FILL FILL_2__9550_ (
);

FILL FILL_5__13349_ (
);

FILL FILL_3__14383_ (
);

FILL FILL_2__9130_ (
);

FILL SFILL93480x78050 (
);

FILL SFILL109560x19050 (
);

DFFSR _7649_ (
    .Q(\datapath_1.regfile_1.regOut[6] [11]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_328_[11])
);

OAI21X1 _7229_ (
    .A(_178_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .C(_179_),
    .Y(_133_[23])
);

FILL FILL_4__9896_ (
);

FILL FILL_4__9476_ (
);

FILL FILL_2__13796_ (
);

FILL FILL_2__13376_ (
);

FILL FILL_5__14710_ (
);

FILL FILL_0__6904_ (
);

FILL FILL_1__12789_ (
);

FILL FILL_1__12369_ (
);

FILL FILL_4__13703_ (
);

FILL SFILL3640x80050 (
);

FILL FILL_0__9796_ (
);

FILL FILL_3__7893_ (
);

FILL FILL_0__9376_ (
);

FILL FILL_3__7473_ (
);

FILL FILL_3__7053_ (
);

OAI21X1 _11647_ (
    .A(_2344__bF$buf1),
    .B(_2402_),
    .C(_2347__bF$buf1),
    .Y(_2750_)
);

NAND2X1 _11227_ (
    .A(_2340_),
    .B(_2343_),
    .Y(_2346_)
);

FILL SFILL59480x72050 (
);

FILL FILL_1__13730_ (
);

FILL FILL_1__13310_ (
);

FILL FILL_4__16175_ (
);

FILL FILL_0__12723_ (
);

FILL FILL_3__15588_ (
);

FILL FILL_3__15168_ (
);

FILL FILL_0__12303_ (
);

FILL FILL_5__8760_ (
);

FILL FILL_5__8340_ (
);

FILL FILL_0__15195_ (
);

AOI21X1 _15480_ (
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .B(_5481_),
    .C(_5949_),
    .Y(_5950_)
);

FILL FILL_5__15915_ (
);

NOR2X1 _15060_ (
    .A(_3933_),
    .B(_5539__bF$buf4),
    .Y(_5540_)
);

FILL FILL_1__8752_ (
);

FILL FILL_5__10630_ (
);

FILL FILL_1__8332_ (
);

FILL FILL_4__14908_ (
);

FILL FILL_2__15942_ (
);

FILL FILL_2__15522_ (
);

FILL FILL_2__15102_ (
);

FILL FILL_3__8258_ (
);

FILL FILL_1__14935_ (
);

FILL FILL_1__14515_ (
);

FILL FILL_4__12095_ (
);

FILL FILL_0__13928_ (
);

FILL FILL_0__13508_ (
);

FILL FILL_5__9545_ (
);

FILL FILL_5__9125_ (
);

FILL FILL_3__11088_ (
);

NOR3X1 _16265_ (
    .A(_5375_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6715_)
);

FILL SFILL3560x42050 (
);

FILL FILL_5__11835_ (
);

FILL FILL_5__11415_ (
);

FILL FILL_1__9537_ (
);

FILL FILL_1__9117_ (
);

FILL FILL_4__7962_ (
);

FILL FILL_2__16307_ (
);

FILL FILL_4__7542_ (
);

FILL FILL_4__10828_ (
);

FILL FILL_4__7122_ (
);

FILL FILL_4__10408_ (
);

FILL FILL_2__11862_ (
);

FILL FILL_2__11442_ (
);

FILL FILL_2__11022_ (
);

FILL FILL_6__7048_ (
);

OAI21X1 _8187_ (
    .A(_654_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_655_),
    .Y(_653_[1])
);

FILL FILL112200x37050 (
);

FILL FILL_1__10435_ (
);

FILL SFILL49480x70050 (
);

FILL FILL_1__10015_ (
);

FILL FILL_0__7862_ (
);

FILL FILL_0__7442_ (
);

FILL FILL_4__14661_ (
);

FILL FILL_4__14241_ (
);

NAND2X1 _12185_ (
    .A(ALUSrcA_bF$buf6),
    .B(\datapath_1.a [23]),
    .Y(_3177_)
);

FILL FILL_3__13654_ (
);

FILL FILL_2__8401_ (
);

FILL FILL_3__13234_ (
);

FILL FILL_6__16099_ (
);

FILL FILL_4__8747_ (
);

FILL FILL_4__8327_ (
);

FILL FILL_2__12647_ (
);

FILL FILL_0__13681_ (
);

FILL FILL_2__12227_ (
);

FILL FILL_0__13261_ (
);

FILL FILL_6_BUFX2_insert81 (
);

FILL FILL_5__16033_ (
);

FILL FILL_0__8647_ (
);

FILL FILL_0__8227_ (
);

NAND2X1 _10918_ (
    .A(\control_1.reg_state.dout [1]),
    .B(\control_1.reg_state.dout [0]),
    .Y(_2060_)
);

FILL FILL_1__9290_ (
);

FILL FILL_6_BUFX2_insert86 (
);

FILL SFILL28840x48050 (
);

FILL FILL_4__15866_ (
);

FILL FILL_4__15446_ (
);

FILL FILL_4__15026_ (
);

FILL FILL_2__16060_ (
);

FILL SFILL73480x74050 (
);

FILL FILL_4__10581_ (
);

FILL FILL_4__10161_ (
);

FILL FILL_3__14859_ (
);

FILL FILL_2__9606_ (
);

FILL FILL_1__15893_ (
);

FILL FILL_3__14439_ (
);

FILL FILL_3__14019_ (
);

FILL FILL_1__15473_ (
);

FILL FILL_1__15053_ (
);

FILL FILL_5__7611_ (
);

FILL FILL_0__14886_ (
);

FILL FILL_0__14466_ (
);

INVX1 _14751_ (
    .A(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_5236_)
);

FILL FILL_0__14046_ (
);

NOR2X1 _14331_ (
    .A(_4821_),
    .B(_4824_),
    .Y(_4825_)
);

FILL FILL_3__15800_ (
);

FILL FILL_1__7603_ (
);

FILL FILL_3__7949_ (
);

FILL FILL_3__7109_ (
);

FILL FILL_5__12373_ (
);

FILL FILL_4__8080_ (
);

FILL FILL_4__11786_ (
);

FILL FILL_4__11366_ (
);

FILL SFILL94360x70050 (
);

FILL FILL_1__16258_ (
);

FILL FILL_3__10779_ (
);

FILL FILL_3__10359_ (
);

FILL FILL_1__11393_ (
);

OAI22X1 _15956_ (
    .A(_5495__bF$buf3),
    .B(_5023_),
    .C(_5526__bF$buf2),
    .D(_5034_),
    .Y(_6414_)
);

AOI21X1 _15536_ (
    .A(_5980_),
    .B(_6004_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [11])
);

INVX1 _15116_ (
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_5595_)
);

INVX1 _10671_ (
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_1925_)
);

FILL FILL_0__10386_ (
);

INVX1 _10251_ (
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_1706_)
);

FILL FILL_6__14585_ (
);

FILL FILL_3__11720_ (
);

FILL FILL_6__14165_ (
);

FILL FILL_3__11300_ (
);

FILL FILL_5__13998_ (
);

FILL FILL_5__13578_ (
);

FILL FILL_5__13158_ (
);

FILL FILL_3__14192_ (
);

OAI21X1 _7878_ (
    .A(_509_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_510_),
    .Y(_458_[26])
);

OAI21X1 _7458_ (
    .A(_290_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_291_),
    .Y(_263_[14])
);

OAI21X1 _7038_ (
    .A(_71_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_72_),
    .Y(_68_[2])
);

FILL FILL_4__9285_ (
);

FILL SFILL18840x46050 (
);

FILL FILL_1__12598_ (
);

FILL FILL_1__12178_ (
);

FILL FILL_4__13932_ (
);

FILL FILL_4__13512_ (
);

NAND2X1 _11876_ (
    .A(RegDst),
    .B(\datapath_1.PCJump [14]),
    .Y(_2961_)
);

NAND3X1 _11456_ (
    .A(_2470__bF$buf2),
    .B(_2557_),
    .C(_2571_),
    .Y(_2572_)
);

INVX1 _11036_ (
    .A(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2155_)
);

FILL FILL_3__12505_ (
);

FILL FILL_2__11918_ (
);

FILL FILL_0__12952_ (
);

FILL FILL_3__15397_ (
);

FILL FILL_0__12532_ (
);

FILL SFILL63880x41050 (
);

FILL FILL_0__12112_ (
);

FILL SFILL38920x6050 (
);

FILL FILL_5__15724_ (
);

FILL FILL_5__15304_ (
);

OAI21X1 _9604_ (
    .A(_1375_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1376_),
    .Y(_1368_[4])
);

FILL FILL_1__8981_ (
);

FILL FILL_1__8141_ (
);

FILL FILL_4__14717_ (
);

FILL FILL_2__15751_ (
);

FILL FILL_2__15331_ (
);

FILL FILL_3__8487_ (
);

FILL FILL_3__8067_ (
);

FILL FILL_1__14744_ (
);

FILL FILL_1__14324_ (
);

FILL FILL_0__13737_ (
);

FILL FILL_0__13317_ (
);

NOR2X1 _13602_ (
    .A(_4110_),
    .B(_4107_),
    .Y(_4111_)
);

FILL FILL_5__9774_ (
);

FILL SFILL109240x38050 (
);

FILL FILL_5__9354_ (
);

AOI21X1 _16074_ (
    .A(\datapath_1.regfile_1.regOut[30] [25]),
    .B(_5481_),
    .C(_6528_),
    .Y(_6529_)
);

FILL FILL_1__9766_ (
);

FILL FILL_5__11644_ (
);

FILL FILL_1__9346_ (
);

FILL FILL_5__11224_ (
);

FILL FILL_2__16116_ (
);

FILL FILL_4__7351_ (
);

FILL FILL_4__10637_ (
);

FILL FILL_2__11671_ (
);

FILL FILL_2__11251_ (
);

FILL FILL_1__15949_ (
);

FILL FILL_1__15529_ (
);

FILL FILL_1__15109_ (
);

FILL FILL_1__10664_ (
);

FILL FILL_1__10244_ (
);

INVX1 _14807_ (
    .A(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_5291_)
);

FILL FILL_2__7689_ (
);

FILL FILL_0__7671_ (
);

FILL FILL_0__7251_ (
);

FILL FILL_4__14890_ (
);

FILL FILL_4__14470_ (
);

FILL FILL_4__14050_ (
);

FILL FILL_5__12849_ (
);

FILL FILL_2__8630_ (
);

FILL FILL_3__13883_ (
);

FILL FILL_5__12429_ (
);

FILL FILL_3__13463_ (
);

FILL FILL_5__12009_ (
);

FILL FILL_2__8210_ (
);

FILL FILL_3__13043_ (
);

FILL FILL_4__8976_ (
);

FILL FILL_4__8136_ (
);

FILL FILL_2__12876_ (
);

FILL SFILL69080x10050 (
);

FILL FILL_2__12456_ (
);

FILL FILL_0__13490_ (
);

FILL FILL_2__12036_ (
);

FILL FILL_1__11869_ (
);

FILL FILL_1__11449_ (
);

FILL FILL_1__11029_ (
);

FILL SFILL3640x75050 (
);

FILL FILL_3__6973_ (
);

FILL FILL_0__8876_ (
);

FILL FILL_5__16262_ (
);

FILL FILL_0__8456_ (
);

DFFSR _10727_ (
    .Q(\datapath_1.regfile_1.regOut[30] [17]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_1888_[17])
);

OAI21X1 _10307_ (
    .A(_1742_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .C(_1743_),
    .Y(_1693_[25])
);

FILL SFILL43880x82050 (
);

FILL FILL_5__6899_ (
);

FILL FILL_4__15675_ (
);

FILL FILL_4__15255_ (
);

DFFSR _13199_ (
    .Q(\datapath_1.mux_iord.din0 [24]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3685_[24])
);

FILL FILL_4__10390_ (
);

FILL FILL_2__9415_ (
);

FILL FILL_0__11803_ (
);

FILL FILL_3__14668_ (
);

FILL FILL_3__14248_ (
);

FILL FILL_1__15282_ (
);

FILL FILL_5__7840_ (
);

FILL FILL_5__7420_ (
);

FILL SFILL59080x53050 (
);

INVX2 _14980_ (
    .A(\datapath_1.PCJump [23]),
    .Y(_5460_)
);

FILL FILL_0__14695_ (
);

AOI22X1 _14560_ (
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .B(_4225_),
    .C(_4129_),
    .D(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_5049_)
);

FILL FILL_0__14275_ (
);

INVX1 _14140_ (
    .A(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_4638_)
);

FILL SFILL38920x38050 (
);

FILL FILL_1__7832_ (
);

FILL FILL_2__14602_ (
);

FILL FILL_3__7758_ (
);

FILL FILL_3__7338_ (
);

FILL SFILL3640x30050 (
);

FILL FILL_5__12182_ (
);

FILL FILL_4__11595_ (
);

FILL FILL_4__11175_ (
);

FILL FILL_1__16067_ (
);

FILL FILL_5__8625_ (
);

FILL FILL_5__8205_ (
);

FILL FILL_3__10168_ (
);

FILL FILL_6_BUFX2_insert592 (
);

FILL SFILL59000x51050 (
);

FILL FILL_6__11922_ (
);

OAI21X1 _15765_ (
    .A(_6226_),
    .B(_5535__bF$buf1),
    .C(_6227_),
    .Y(_6228_)
);

FILL FILL_6__11502_ (
);

OAI22X1 _15345_ (
    .A(_5530__bF$buf2),
    .B(_5817_),
    .C(_5532__bF$buf3),
    .D(_4298_),
    .Y(_5818_)
);

FILL FILL_6_BUFX2_insert597 (
);

FILL SFILL3560x37050 (
);

DFFSR _10480_ (
    .Q(\datapath_1.regfile_1.regOut[28] [26]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_1758_[26])
);

FILL FILL_0__10195_ (
);

FILL FILL_5__10915_ (
);

OAI21X1 _10060_ (
    .A(_1618_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .C(_1619_),
    .Y(_1563_[28])
);

FILL FILL_1__8617_ (
);

FILL FILL_2__15807_ (
);

FILL FILL_0__16001_ (
);

FILL FILL_2__10942_ (
);

FILL FILL_5__13387_ (
);

FILL FILL_2__10522_ (
);

FILL FILL_2__10102_ (
);

OAI21X1 _7687_ (
    .A(_402_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .C(_403_),
    .Y(_393_[5])
);

DFFSR _7267_ (
    .Q(\datapath_1.regfile_1.regOut[3] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_133_[13])
);

FILL FILL_4__9094_ (
);

FILL SFILL33880x80050 (
);

FILL FILL_3__9904_ (
);

FILL SFILL38040x17050 (
);

FILL FILL_0__6942_ (
);

FILL FILL_6__12707_ (
);

FILL FILL_4__13741_ (
);

FILL FILL_4__13321_ (
);

FILL FILL_3__7091_ (
);

OAI21X1 _11685_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(_2183_),
    .C(_2164_),
    .Y(_2786_)
);

INVX1 _11265_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .Y(_2384_)
);

FILL FILL_3__12734_ (
);

FILL FILL_3__12314_ (
);

FILL SFILL28920x36050 (
);

FILL FILL_4__7827_ (
);

FILL FILL_2__11727_ (
);

FILL FILL_0__12761_ (
);

FILL FILL_2__11307_ (
);

FILL FILL_0__12341_ (
);

FILL FILL_2__14199_ (
);

FILL FILL_5__15953_ (
);

FILL FILL_5__15533_ (
);

FILL FILL_0__7727_ (
);

FILL FILL_5__15113_ (
);

FILL FILL_0__7307_ (
);

DFFSR _9833_ (
    .Q(\datapath_1.regfile_1.regOut[23] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_1433_[19])
);

NAND2X1 _9413_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1290_)
);

FILL FILL_1__8370_ (
);

FILL FILL_4__14946_ (
);

FILL FILL_2__15980_ (
);

FILL FILL_4__14526_ (
);

FILL FILL_2__15560_ (
);

FILL FILL_4__14106_ (
);

FILL FILL_2__15140_ (
);

FILL SFILL73960x31050 (
);

FILL SFILL89560x16050 (
);

FILL FILL_3__13939_ (
);

FILL FILL_1__14973_ (
);

FILL FILL_3__13519_ (
);

FILL FILL_1__14553_ (
);

FILL FILL_1__14133_ (
);

FILL SFILL28440x29050 (
);

FILL FILL_0__13966_ (
);

INVX1 _13831_ (
    .A(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_4336_)
);

FILL FILL_0__13546_ (
);

FILL FILL_0__13126_ (
);

INVX1 _13411_ (
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_3923_)
);

FILL FILL_5__9163_ (
);

FILL FILL_5__16318_ (
);

FILL FILL_1__9995_ (
);

FILL FILL_5__11873_ (
);

FILL FILL_5__11453_ (
);

FILL FILL_5__11033_ (
);

FILL FILL_1__9155_ (
);

FILL FILL_2__16345_ (
);

FILL FILL_4__7580_ (
);

FILL SFILL79560x59050 (
);

FILL FILL_4__7160_ (
);

FILL SFILL94360x65050 (
);

FILL FILL_4__10446_ (
);

FILL FILL_4__10026_ (
);

FILL FILL_2__11480_ (
);

FILL FILL_2__11060_ (
);

FILL FILL_1__15758_ (
);

FILL FILL_1__15338_ (
);

FILL FILL_1__10893_ (
);

FILL FILL_1__10053_ (
);

NOR2X1 _14616_ (
    .A(_5100_),
    .B(_5103_),
    .Y(_5104_)
);

FILL FILL_2__7498_ (
);

FILL FILL_0__7480_ (
);

FILL SFILL79160x45050 (
);

FILL FILL_2__7078_ (
);

FILL FILL_0__7060_ (
);

FILL FILL_3__10800_ (
);

FILL FILL_5__12658_ (
);

FILL SFILL18760x1050 (
);

FILL FILL_5__12238_ (
);

FILL FILL_3__13692_ (
);

FILL FILL_3__13272_ (
);

OAI21X1 _6958_ (
    .A(_38_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .C(_39_),
    .Y(_3_[18])
);

FILL FILL_4__8785_ (
);

FILL SFILL18680x6050 (
);

FILL FILL_4__8365_ (
);

FILL FILL_2__12265_ (
);

FILL SFILL94360x20050 (
);

FILL FILL_1__11678_ (
);

FILL FILL_1__11258_ (
);

FILL FILL_5__16071_ (
);

NAND3X1 _10956_ (
    .A(_2079_),
    .B(_2088_),
    .C(_2083_),
    .Y(\control_1.next [1])
);

FILL FILL_0__8265_ (
);

OAI21X1 _10536_ (
    .A(_1854_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .C(_1855_),
    .Y(_1823_[16])
);

OAI21X1 _10116_ (
    .A(_1635_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .C(_1636_),
    .Y(_1628_[4])
);

FILL FILL_4__15484_ (
);

FILL FILL_4__15064_ (
);

FILL SFILL8760x82050 (
);

FILL FILL_2__9644_ (
);

FILL FILL_3__14897_ (
);

FILL FILL_3__14477_ (
);

FILL FILL_2__9224_ (
);

FILL FILL_0__11612_ (
);

FILL FILL_3__14057_ (
);

FILL FILL_1__15091_ (
);

FILL FILL_0__14084_ (
);

FILL SFILL114600x82050 (
);

FILL FILL_5__14804_ (
);

FILL SFILL84360x63050 (
);

FILL SFILL63480x22050 (
);

FILL FILL_1__7221_ (
);

FILL FILL_6_CLKBUF1_insert193 (
);

FILL FILL_2__14831_ (
);

FILL FILL_2__14411_ (
);

FILL FILL_3__7987_ (
);

FILL FILL_3__7567_ (
);

FILL FILL_6_CLKBUF1_insert198 (
);

FILL FILL_1__13824_ (
);

FILL FILL_1__13404_ (
);

FILL FILL_4__16269_ (
);

FILL SFILL53880x79050 (
);

FILL FILL_1__16296_ (
);

FILL FILL_5__8854_ (
);

FILL FILL_3__10397_ (
);

FILL FILL_5__8014_ (
);

NAND2X1 _15994_ (
    .A(_6445_),
    .B(_6450_),
    .Y(_6451_)
);

FILL FILL_0__15289_ (
);

AOI22X1 _15574_ (
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_6041_)
);

OAI22X1 _15154_ (
    .A(_5631_),
    .B(_5545__bF$buf3),
    .C(_5466__bF$buf1),
    .D(_4063_),
    .Y(_5632_)
);

FILL FILL_3__16203_ (
);

FILL FILL_1__8846_ (
);

FILL FILL_5__10304_ (
);

FILL FILL_1__8006_ (
);

FILL FILL_2__15616_ (
);

FILL FILL_4__6851_ (
);

FILL FILL_0__16230_ (
);

FILL FILL_2__10751_ (
);

FILL FILL_1__14609_ (
);

NAND2X1 _7496_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_317_)
);

NAND2X1 _7076_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_98_)
);

FILL FILL_4__12189_ (
);

FILL FILL_5__9639_ (
);

FILL FILL_5__9219_ (
);

FILL FILL_4__13970_ (
);

OAI21X1 _16359_ (
    .A(_6792_),
    .B(gnd),
    .C(_6793_),
    .Y(_6769_[12])
);

FILL FILL_4__13550_ (
);

FILL FILL_4__13130_ (
);

NAND2X1 _11494_ (
    .A(_2296_),
    .B(_2478_),
    .Y(_2607_)
);

FILL FILL_5__11929_ (
);

OAI21X1 _11074_ (
    .A(_2191_),
    .B(_2192_),
    .C(_2188_),
    .Y(_2193_)
);

FILL FILL_3__12963_ (
);

FILL FILL_5__11509_ (
);

FILL FILL_2__7710_ (
);

FILL SFILL43960x70050 (
);

FILL FILL_3__12123_ (
);

FILL FILL_4__7636_ (
);

FILL FILL_4__7216_ (
);

FILL FILL_2__11956_ (
);

FILL FILL_0__12990_ (
);

FILL FILL_2__11536_ (
);

FILL FILL_0__12570_ (
);

FILL FILL_3_CLKBUF1_insert140 (
);

FILL FILL_2__11116_ (
);

FILL FILL_3_CLKBUF1_insert141 (
);

FILL FILL_0__12150_ (
);

FILL FILL_3_CLKBUF1_insert142 (
);

FILL FILL_3_CLKBUF1_insert143 (
);

FILL FILL_3_CLKBUF1_insert144 (
);

FILL FILL_1__10949_ (
);

FILL FILL_3_CLKBUF1_insert145 (
);

FILL FILL_1__10529_ (
);

FILL FILL_3_CLKBUF1_insert146 (
);

FILL FILL_3_CLKBUF1_insert147 (
);

FILL FILL_1__10109_ (
);

FILL FILL_3_CLKBUF1_insert148 (
);

FILL FILL_3_CLKBUF1_insert149 (
);

FILL FILL_5__15762_ (
);

FILL FILL_5__15342_ (
);

FILL FILL_0__7956_ (
);

FILL FILL_0__7116_ (
);

NAND2X1 _9642_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1402_)
);

NAND2X1 _9222_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1183_)
);

FILL SFILL43880x77050 (
);

FILL FILL_4__14755_ (
);

FILL FILL_4__14335_ (
);

NAND2X1 _12699_ (
    .A(IRWrite_bF$buf1),
    .B(memoryOutData[1]),
    .Y(_3492_)
);

NAND3X1 _12279_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3248_)
);

FILL FILL_2__8915_ (
);

FILL SFILL3560x8050 (
);

FILL FILL_3__13748_ (
);

FILL FILL_3__13328_ (
);

FILL FILL_1__14782_ (
);

FILL FILL_1__14362_ (
);

FILL FILL_5__6920_ (
);

FILL SFILL59080x48050 (
);

FILL FILL112280x81050 (
);

FILL FILL_0__13775_ (
);

FILL FILL_0__13355_ (
);

OAI22X1 _13640_ (
    .A(_4146_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf3),
    .D(_4147_),
    .Y(_4148_)
);

INVX2 _13220_ (
    .A(\datapath_1.a3 [1]),
    .Y(_3763_)
);

FILL FILL_5__9392_ (
);

FILL FILL_1__6912_ (
);

FILL FILL_3__6838_ (
);

FILL FILL_5__16127_ (
);

FILL SFILL3640x25050 (
);

FILL FILL_5__11682_ (
);

FILL FILL_1__9384_ (
);

FILL FILL_5__11262_ (
);

FILL FILL_2__16154_ (
);

FILL FILL_4__10675_ (
);

FILL FILL_4__10255_ (
);

FILL FILL_1__15987_ (
);

FILL FILL_1__15567_ (
);

FILL FILL_1__15147_ (
);

FILL FILL_5__7705_ (
);

FILL FILL_1__10282_ (
);

NOR2X1 _14845_ (
    .A(_5327_),
    .B(_5324_),
    .Y(_5328_)
);

INVX1 _14425_ (
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_4917_)
);

INVX1 _14005_ (
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_4506_)
);

FILL FILL_6__13894_ (
);

FILL FILL_6__13474_ (
);

FILL SFILL104440x49050 (
);

FILL FILL_0__15921_ (
);

FILL FILL_0__15501_ (
);

FILL FILL_5__12887_ (
);

FILL FILL_5__12467_ (
);

FILL FILL_5__12047_ (
);

FILL FILL_3__13081_ (
);

FILL FILL_4__8594_ (
);

FILL SFILL33880x75050 (
);

FILL FILL_2__12494_ (
);

FILL FILL_2__12074_ (
);

FILL FILL_1__11487_ (
);

FILL FILL_1__11067_ (
);

FILL FILL_4__12401_ (
);

FILL FILL_6__9881_ (
);

FILL FILL_0__8494_ (
);

FILL SFILL49080x46050 (
);

OAI21X1 _10765_ (
    .A(_1966_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1967_),
    .Y(_1953_[7])
);

FILL FILL_0__8074_ (
);

DFFSR _10345_ (
    .Q(\datapath_1.regfile_1.regOut[27] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1693_[19])
);

FILL FILL_3__11814_ (
);

FILL FILL_4__15293_ (
);

FILL FILL_4__6907_ (
);

FILL FILL_2__10807_ (
);

FILL FILL_2__9873_ (
);

FILL FILL_0__11841_ (
);

FILL FILL_3__14286_ (
);

FILL FILL_0__11421_ (
);

FILL FILL_2__9033_ (
);

FILL FILL_0__11001_ (
);

FILL FILL_4__9799_ (
);

FILL FILL_4__9379_ (
);

FILL FILL_2__13699_ (
);

FILL FILL_2__13279_ (
);

FILL FILL_5__14613_ (
);

NAND2X1 _8913_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1038_)
);

FILL FILL_1__7870_ (
);

FILL FILL_1__7450_ (
);

FILL FILL_1__7030_ (
);

FILL FILL_4__13606_ (
);

FILL FILL_2__14640_ (
);

FILL FILL_2__14220_ (
);

FILL SFILL49000x44050 (
);

FILL FILL_0__9279_ (
);

FILL FILL_3__7376_ (
);

FILL FILL_5_CLKBUF1_insert180 (
);

FILL FILL_5_CLKBUF1_insert181 (
);

FILL FILL_5_CLKBUF1_insert182 (
);

FILL FILL_1__13633_ (
);

FILL FILL_5_CLKBUF1_insert183 (
);

FILL FILL_1__13213_ (
);

FILL FILL_5_CLKBUF1_insert184 (
);

FILL FILL_4__16078_ (
);

FILL FILL_5_CLKBUF1_insert185 (
);

FILL FILL_5_CLKBUF1_insert186 (
);

FILL FILL_5_CLKBUF1_insert187 (
);

FILL FILL_5_CLKBUF1_insert188 (
);

FILL FILL_1_BUFX2_insert410 (
);

FILL FILL_1_BUFX2_insert411 (
);

FILL FILL_5_CLKBUF1_insert189 (
);

NAND2X1 _12911_ (
    .A(vdd),
    .B(\datapath_1.rd1 [29]),
    .Y(_3613_)
);

FILL FILL_0__12626_ (
);

FILL FILL_1_BUFX2_insert412 (
);

FILL FILL_1_BUFX2_insert413 (
);

FILL FILL_0__12206_ (
);

FILL FILL_1_BUFX2_insert414 (
);

FILL FILL_1_BUFX2_insert415 (
);

FILL FILL_1_BUFX2_insert416 (
);

FILL FILL_6_BUFX2_insert971 (
);

FILL FILL_1_BUFX2_insert417 (
);

FILL FILL_5__8243_ (
);

FILL FILL_1_BUFX2_insert418 (
);

FILL FILL_1_BUFX2_insert419 (
);

AOI22X1 _15383_ (
    .A(_5565__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [8]),
    .C(\datapath_1.regfile_1.regOut[5] [8]),
    .D(_5700_),
    .Y(_5855_)
);

FILL FILL_0__15098_ (
);

FILL FILL_6_BUFX2_insert976 (
);

FILL FILL_5__15818_ (
);

FILL SFILL23880x73050 (
);

FILL FILL_3__16012_ (
);

FILL FILL_5__10953_ (
);

FILL FILL_1__8655_ (
);

FILL FILL_5__10533_ (
);

FILL FILL_5__10113_ (
);

FILL FILL_1__8235_ (
);

FILL FILL_2__15845_ (
);

FILL FILL_2__15425_ (
);

FILL FILL_2__15005_ (
);

FILL FILL_2__10980_ (
);

FILL FILL_2__10560_ (
);

FILL FILL_2__10140_ (
);

FILL FILL_1__14838_ (
);

FILL FILL_1__14418_ (
);

FILL FILL_3__9522_ (
);

FILL FILL_3__9102_ (
);

FILL FILL_0__6980_ (
);

FILL FILL_5__9868_ (
);

FILL FILL_5__9028_ (
);

OAI22X1 _16168_ (
    .A(_5478__bF$buf0),
    .B(_6619_),
    .C(_5552__bF$buf2),
    .D(_5312_),
    .Y(_6620_)
);

FILL FILL_5__11738_ (
);

FILL FILL_3__12772_ (
);

FILL FILL_5__11318_ (
);

FILL FILL_3__12352_ (
);

FILL FILL_4__7865_ (
);

FILL FILL_4__7445_ (
);

FILL FILL_2__11765_ (
);

FILL FILL111800x44050 (
);

FILL FILL_2__11345_ (
);

FILL SFILL94360x15050 (
);

FILL FILL_1__10758_ (
);

FILL FILL_2_CLKBUF1_insert130 (
);

FILL FILL_2_CLKBUF1_insert131 (
);

FILL FILL_5__15991_ (
);

FILL FILL_2_CLKBUF1_insert132 (
);

FILL FILL_2_CLKBUF1_insert133 (
);

FILL FILL_5__15571_ (
);

FILL FILL_0__7765_ (
);

FILL FILL_2_CLKBUF1_insert134 (
);

FILL FILL_5__15151_ (
);

NAND2X1 _9871_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1514_)
);

FILL FILL_2_CLKBUF1_insert135 (
);

FILL FILL_0__7345_ (
);

DFFSR _9451_ (
    .Q(\datapath_1.regfile_1.regOut[20] [21]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_1238_[21])
);

FILL FILL_2_CLKBUF1_insert136 (
);

INVX1 _9031_ (
    .A(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_1096_)
);

FILL FILL_2_CLKBUF1_insert137 (
);

FILL FILL_2_CLKBUF1_insert138 (
);

FILL FILL_4__14984_ (
);

FILL FILL_2_CLKBUF1_insert139 (
);

FILL FILL_4__14564_ (
);

FILL SFILL8760x77050 (
);

FILL FILL_4__14144_ (
);

NAND3X1 _12088_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [25]),
    .C(_3034__bF$buf4),
    .Y(_3112_)
);

FILL FILL_3__13977_ (
);

FILL FILL_2__8724_ (
);

FILL FILL_3__13557_ (
);

FILL FILL_1__14591_ (
);

FILL FILL_3__13137_ (
);

FILL FILL_1__14171_ (
);

FILL FILL_6_BUFX2_insert1012 (
);

FILL FILL_5_BUFX2_insert990 (
);

FILL FILL_5_BUFX2_insert991 (
);

FILL FILL_5_BUFX2_insert992 (
);

FILL FILL_5_BUFX2_insert993 (
);

FILL FILL_0__13584_ (
);

FILL FILL_5_BUFX2_insert994 (
);

FILL FILL_0__13164_ (
);

FILL SFILL53960x67050 (
);

FILL FILL_5_BUFX2_insert995 (
);

FILL FILL_6_BUFX2_insert1017 (
);

FILL SFILL84360x58050 (
);

FILL FILL_5_BUFX2_insert996 (
);

FILL FILL_5_BUFX2_insert997 (
);

FILL FILL_5_BUFX2_insert998 (
);

FILL FILL_5_BUFX2_insert999 (
);

FILL SFILL29080x42050 (
);

FILL FILL_2__13911_ (
);

FILL FILL_5__16356_ (
);

FILL FILL_6__9937_ (
);

FILL FILL_5__11491_ (
);

FILL FILL_5__11071_ (
);

FILL FILL_1__12904_ (
);

FILL FILL_4__15769_ (
);

FILL FILL_4__15349_ (
);

FILL FILL_2__16383_ (
);

FILL FILL_0__9911_ (
);

FILL FILL_4__10064_ (
);

FILL FILL_2__9929_ (
);

FILL SFILL8760x32050 (
);

FILL FILL_2__9509_ (
);

FILL FILL_1__15796_ (
);

FILL FILL_1__15376_ (
);

FILL FILL_5__7934_ (
);

FILL FILL_6__10811_ (
);

FILL FILL_0__14789_ (
);

FILL FILL_0__14369_ (
);

NOR2X1 _14654_ (
    .A(_5137_),
    .B(_5140_),
    .Y(_5141_)
);

NOR2X1 _14234_ (
    .A(_4726_),
    .B(_4729_),
    .Y(_4730_)
);

FILL FILL_3__15703_ (
);

FILL SFILL114600x32050 (
);

FILL FILL_1__7926_ (
);

FILL SFILL53960x22050 (
);

FILL FILL_1__7506_ (
);

FILL SFILL84360x13050 (
);

FILL FILL_0__15730_ (
);

FILL FILL_0__15310_ (
);

FILL FILL_5__12696_ (
);

FILL FILL_5__12276_ (
);

NAND2X1 _6996_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_65_)
);

FILL FILL_4__11689_ (
);

FILL FILL_4__11269_ (
);

FILL FILL_5__8719_ (
);

FILL FILL_1__11296_ (
);

NAND2X1 _15859_ (
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .B(_5971_),
    .Y(_6319_)
);

FILL FILL_4__12630_ (
);

AOI21X1 _15439_ (
    .A(\datapath_1.regfile_1.regOut[30] [9]),
    .B(_5481_),
    .C(_5909_),
    .Y(_5910_)
);

NAND3X1 _15019_ (
    .A(_5459__bF$buf0),
    .B(_5477_),
    .C(_5461_),
    .Y(_5499_)
);

FILL FILL_4__12210_ (
);

INVX1 _10994_ (
    .A(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2113_)
);

NAND2X1 _10574_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1881_)
);

FILL FILL_6__9270_ (
);

FILL FILL_0__10289_ (
);

NAND2X1 _10154_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1662_)
);

FILL FILL_3_BUFX2_insert1070 (
);

FILL FILL_3_BUFX2_insert1071 (
);

FILL SFILL43960x65050 (
);

FILL FILL_3_BUFX2_insert1072 (
);

FILL FILL_3__11623_ (
);

FILL FILL_3_BUFX2_insert1073 (
);

FILL FILL_6__14068_ (
);

FILL FILL_3__11203_ (
);

FILL FILL_2__10616_ (
);

FILL FILL_2__9682_ (
);

FILL FILL_2__9262_ (
);

FILL FILL_0__11650_ (
);

FILL FILL_0__11230_ (
);

FILL FILL_3__14095_ (
);

FILL SFILL104200x61050 (
);

FILL FILL_2__13088_ (
);

FILL FILL_5__14842_ (
);

FILL FILL_5__14422_ (
);

FILL FILL_5__14002_ (
);

NAND2X1 _8722_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_931_)
);

DFFSR _8302_ (
    .Q(\datapath_1.regfile_1.regOut[11] [24]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_653_[24])
);

FILL FILL_4__13835_ (
);

FILL FILL_4__13415_ (
);

FILL FILL_0__9088_ (
);

OAI22X1 _11779_ (
    .A(_2861_),
    .B(_2346_),
    .C(_2347__bF$buf2),
    .D(_2139_),
    .Y(_2873_)
);

FILL FILL_3__7185_ (
);

AND2X2 _11359_ (
    .A(_2475_),
    .B(_2452_),
    .Y(_2476_)
);

FILL SFILL3720x13050 (
);

FILL FILL_3__12828_ (
);

FILL FILL_3__12408_ (
);

FILL FILL_1__13862_ (
);

FILL FILL_1__13442_ (
);

FILL FILL_1__13022_ (
);

FILL SFILL43960x20050 (
);

FILL FILL112280x76050 (
);

FILL FILL_4_CLKBUF1_insert170 (
);

FILL FILL_4_CLKBUF1_insert171 (
);

FILL FILL_0__12855_ (
);

FILL FILL_4_CLKBUF1_insert172 (
);

NAND2X1 _12720_ (
    .A(IRWrite_bF$buf5),
    .B(memoryOutData[8]),
    .Y(_3506_)
);

FILL FILL_4_CLKBUF1_insert173 (
);

FILL FILL_0__12435_ (
);

FILL FILL_0__12015_ (
);

NAND3X1 _12300_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf1),
    .Y(_3264_)
);

FILL FILL_4_CLKBUF1_insert174 (
);

FILL FILL_4_CLKBUF1_insert175 (
);

FILL FILL_5__8892_ (
);

FILL FILL_4_CLKBUF1_insert176 (
);

FILL FILL_5__8472_ (
);

FILL FILL_4_CLKBUF1_insert177 (
);

FILL FILL_4_CLKBUF1_insert178 (
);

FILL FILL_4_CLKBUF1_insert179 (
);

NOR2X1 _15192_ (
    .A(_5665_),
    .B(_5668_),
    .Y(_5669_)
);

FILL FILL_5__15627_ (
);

FILL FILL_5__15207_ (
);

FILL FILL_3__16241_ (
);

INVX1 _9927_ (
    .A(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_1551_)
);

INVX1 _9507_ (
    .A(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_1332_)
);

FILL FILL_5__10762_ (
);

FILL FILL_1__8884_ (
);

FILL FILL_1__8464_ (
);

FILL FILL_2__15654_ (
);

FILL SFILL43880x27050 (
);

FILL FILL_2__15234_ (
);

FILL FILL_1__14647_ (
);

FILL FILL_1__14227_ (
);

FILL FILL_3__9751_ (
);

NOR2X1 _13925_ (
    .A(_4424_),
    .B(_4427_),
    .Y(_4428_)
);

INVX1 _13505_ (
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_4016_)
);

FILL FILL112280x31050 (
);

FILL FILL_5__9677_ (
);

FILL FILL_5__9257_ (
);

NAND2X1 _16397_ (
    .A(gnd),
    .B(gnd),
    .Y(_6819_)
);

FILL FILL_5__11967_ (
);

FILL FILL_1__9669_ (
);

FILL FILL_5__11547_ (
);

FILL FILL_3__12581_ (
);

FILL FILL_1__9249_ (
);

FILL FILL_5__11127_ (
);

FILL FILL_3__12161_ (
);

FILL FILL_2__16019_ (
);

FILL FILL_4__7674_ (
);

FILL FILL_2__11994_ (
);

FILL FILL_2__11574_ (
);

FILL FILL_2__11154_ (
);

FILL FILL_1__10567_ (
);

FILL FILL_1__10147_ (
);

FILL FILL_4__11901_ (
);

FILL FILL_5__15380_ (
);

FILL FILL_0__7994_ (
);

FILL FILL_6__8961_ (
);

FILL FILL_0__7574_ (
);

INVX1 _9680_ (
    .A(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_1427_)
);

INVX1 _9260_ (
    .A(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_1208_)
);

FILL FILL_1_CLKBUF1_insert120 (
);

FILL FILL_1_CLKBUF1_insert121 (
);

FILL FILL_4__14793_ (
);

FILL FILL_1_CLKBUF1_insert122 (
);

FILL FILL_1_CLKBUF1_insert123 (
);

FILL FILL_4__14373_ (
);

FILL FILL_1_CLKBUF1_insert124 (
);

FILL FILL_1_CLKBUF1_insert125 (
);

FILL FILL_1_CLKBUF1_insert126 (
);

FILL FILL_1_CLKBUF1_insert127 (
);

FILL FILL_1_CLKBUF1_insert128 (
);

FILL FILL_2__8953_ (
);

FILL FILL_0__10921_ (
);

FILL FILL_3__13786_ (
);

FILL FILL_2__8533_ (
);

FILL FILL_1_CLKBUF1_insert129 (
);

FILL FILL_3__13366_ (
);

FILL FILL_2__8113_ (
);

FILL FILL_0__10501_ (
);

FILL FILL_4__8879_ (
);

FILL FILL_4__8459_ (
);

FILL FILL_2__12779_ (
);

FILL FILL_2__12359_ (
);

FILL FILL_0__13393_ (
);

FILL SFILL33880x25050 (
);

FILL FILL_1__6950_ (
);

FILL FILL_4__9400_ (
);

FILL SFILL18600x48050 (
);

FILL FILL_2__13720_ (
);

FILL SFILL49000x39050 (
);

FILL FILL_2__13300_ (
);

FILL FILL_5__16165_ (
);

FILL FILL_0__8779_ (
);

FILL FILL_3__6876_ (
);

FILL FILL_0__8359_ (
);

FILL FILL_6__9746_ (
);

FILL FILL_4__15998_ (
);

FILL FILL_1__12713_ (
);

FILL FILL_4__15578_ (
);

FILL FILL_4__15158_ (
);

FILL FILL_2__16192_ (
);

FILL SFILL94440x48050 (
);

FILL FILL_4__10293_ (
);

FILL FILL_2__9738_ (
);

FILL FILL_0__9720_ (
);

FILL FILL_0__9300_ (
);

FILL FILL_0__11706_ (
);

FILL FILL_1__15185_ (
);

FILL FILL_6__15905_ (
);

FILL FILL_5__7743_ (
);

FILL FILL_5__7323_ (
);

FILL FILL_0__14598_ (
);

INVX1 _14883_ (
    .A(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_5365_)
);

OAI22X1 _14463_ (
    .A(_3949_),
    .B(_4953_),
    .C(_3966__bF$buf0),
    .D(_4952_),
    .Y(_4954_)
);

FILL FILL_0__14178_ (
);

FILL SFILL23880x68050 (
);

INVX1 _14043_ (
    .A(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_4543_)
);

FILL FILL_3__15932_ (
);

FILL FILL_3__15512_ (
);

FILL FILL_1__7735_ (
);

FILL FILL_1__7315_ (
);

FILL FILL_2__14925_ (
);

FILL FILL_2__14505_ (
);

FILL FILL_5__12085_ (
);

FILL FILL_1__13918_ (
);

FILL SFILL105080x62050 (
);

FILL FILL_4__11498_ (
);

FILL FILL_4__11078_ (
);

FILL FILL_3__8602_ (
);

FILL FILL_5__8528_ (
);

FILL FILL_5__8108_ (
);

NOR2X1 _15668_ (
    .A(_6132_),
    .B(_6125_),
    .Y(_6133_)
);

FILL FILL_6__11405_ (
);

FILL SFILL23800x66050 (
);

INVX1 _15248_ (
    .A(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_5724_)
);

NAND2X1 _10383_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1774_)
);

FILL FILL_5__10818_ (
);

FILL FILL_3__11852_ (
);

FILL FILL_3__11432_ (
);

FILL FILL_3__11012_ (
);

FILL FILL_4__6945_ (
);

FILL FILL_0__16324_ (
);

FILL FILL_2__10425_ (
);

FILL FILL_2__9491_ (
);

FILL FILL_2__10005_ (
);

FILL SFILL39000x37050 (
);

FILL FILL112360x5050 (
);

FILL FILL_3__9807_ (
);

FILL FILL_5__14651_ (
);

FILL FILL_0__6845_ (
);

FILL FILL_5__14231_ (
);

NAND2X1 _8951_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .Y(_1107_)
);

INVX1 _8531_ (
    .A(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_844_)
);

INVX1 _8111_ (
    .A(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_625_)
);

FILL FILL_4__13644_ (
);

FILL FILL_4__13224_ (
);

NAND3X1 _11588_ (
    .A(_2264_),
    .B(_2691_),
    .C(_2694_),
    .Y(_2695_)
);

INVX1 _11168_ (
    .A(_2286_),
    .Y(_2287_)
);

FILL SFILL23800x21050 (
);

FILL FILL_2__7804_ (
);

FILL FILL_3__12637_ (
);

FILL FILL_1__13671_ (
);

FILL FILL_3__12217_ (
);

FILL FILL_1__13251_ (
);

FILL FILL_0__12244_ (
);

FILL SFILL74200x2050 (
);

FILL FILL_5__15856_ (
);

FILL FILL_5__15436_ (
);

FILL FILL_5__15016_ (
);

INVX1 _9736_ (
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_1444_)
);

FILL FILL_3__16050_ (
);

DFFSR _9316_ (
    .Q(\datapath_1.regfile_1.regOut[19] [14]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_1173_[14])
);

FILL FILL_5__10991_ (
);

FILL FILL_5__10571_ (
);

FILL SFILL114200x58050 (
);

FILL FILL_5__10151_ (
);

FILL FILL_1__8273_ (
);

FILL FILL_4__14849_ (
);

FILL FILL_2__15883_ (
);

FILL FILL_4__14429_ (
);

FILL FILL_4__14009_ (
);

FILL FILL_2__15463_ (
);

FILL FILL_2__15043_ (
);

FILL FILL_3__8199_ (
);

FILL FILL_1__14876_ (
);

FILL FILL_1__14456_ (
);

FILL FILL_1__14036_ (
);

FILL FILL_3__9980_ (
);

FILL FILL_0__13869_ (
);

FILL FILL_0__13449_ (
);

FILL FILL_3__9140_ (
);

NOR2X1 _13734_ (
    .A(_4240_),
    .B(_4237_),
    .Y(_4241_)
);

NOR2X1 _13314_ (
    .A(_3846_),
    .B(_3781_),
    .Y(\datapath_1.regfile_1.regEn [11])
);

FILL FILL_0__13029_ (
);

FILL FILL_5__9486_ (
);

FILL SFILL114600x27050 (
);

FILL SFILL53960x17050 (
);

FILL FILL_0__14810_ (
);

FILL FILL_5__11776_ (
);

FILL FILL_1__9898_ (
);

FILL FILL_5__11356_ (
);

FILL FILL_1__9478_ (
);

FILL FILL_3__12390_ (
);

FILL FILL_2__16248_ (
);

FILL FILL_4__7483_ (
);

FILL FILL_4__7063_ (
);

FILL FILL_4__10769_ (
);

FILL FILL_2__11383_ (
);

FILL FILL_1__10796_ (
);

FILL FILL_1__10376_ (
);

NAND3X1 _14939_ (
    .A(_5411_),
    .B(_5412_),
    .C(_5419_),
    .Y(_5420_)
);

NOR2X1 _14519_ (
    .A(_5005_),
    .B(_5008_),
    .Y(_5009_)
);

FILL FILL_4__11710_ (
);

FILL FILL_3__10703_ (
);

FILL FILL_4__14182_ (
);

FILL FILL_2__8762_ (
);

FILL FILL_3__13595_ (
);

FILL FILL_2__8342_ (
);

FILL FILL_0__10310_ (
);

FILL FILL_4__8268_ (
);

FILL FILL112360x64050 (
);

FILL FILL_2__12588_ (
);

FILL FILL_2__12168_ (
);

FILL FILL_5__13922_ (
);

FILL FILL_5__13502_ (
);

NAND2X1 _7802_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_460_)
);

FILL FILL_4_BUFX2_insert300 (
);

FILL FILL_4_BUFX2_insert301 (
);

FILL FILL_4_BUFX2_insert302 (
);

FILL FILL_4__12915_ (
);

FILL FILL_4_BUFX2_insert303 (
);

FILL SFILL64040x73050 (
);

FILL FILL_4_BUFX2_insert304 (
);

FILL FILL_5__16394_ (
);

FILL FILL_0__8588_ (
);

FILL FILL_4_BUFX2_insert305 (
);

DFFSR _10859_ (
    .Q(\datapath_1.regfile_1.regOut[31] [21]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1953_[21])
);

FILL FILL_4_BUFX2_insert306 (
);

FILL FILL_4_BUFX2_insert307 (
);

INVX1 _10439_ (
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_1811_)
);

INVX1 _10019_ (
    .A(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_1592_)
);

FILL FILL_4_BUFX2_insert308 (
);

FILL FILL_3__11908_ (
);

FILL FILL_4_BUFX2_insert309 (
);

FILL FILL_4__15387_ (
);

FILL FILL_1__12522_ (
);

FILL FILL_1__12102_ (
);

FILL SFILL43960x15050 (
);

FILL FILL_2__9547_ (
);

FILL FILL_0__11935_ (
);

FILL SFILL68360x81050 (
);

FILL FILL_2__9127_ (
);

INVX1 _11800_ (
    .A(_2892_),
    .Y(\datapath_1.ALUResult [5])
);

FILL FILL_0__11515_ (
);

FILL FILL_5__7972_ (
);

FILL FILL_5__7552_ (
);

AOI21X1 _14692_ (
    .A(_5155_),
    .B(_5178_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [25])
);

FILL SFILL108920x33050 (
);

NOR2X1 _14272_ (
    .A(_4763_),
    .B(_4766_),
    .Y(_4767_)
);

FILL FILL_5__14707_ (
);

FILL FILL_3__15741_ (
);

FILL FILL_3__15321_ (
);

FILL FILL_1__7964_ (
);

FILL FILL_1__7544_ (
);

FILL FILL_1__7124_ (
);

FILL FILL_2__14734_ (
);

FILL FILL_2__14314_ (
);

FILL FILL_1__13727_ (
);

FILL FILL_1__13307_ (
);

FILL SFILL84360x4050 (
);

FILL FILL_3__8831_ (
);

FILL FILL112280x26050 (
);

FILL FILL_1__16199_ (
);

FILL FILL_5__8757_ (
);

FILL FILL_5__8337_ (
);

INVX1 _15897_ (
    .A(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_6356_)
);

AOI21X1 _15477_ (
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .B(_5567_),
    .C(_5946_),
    .Y(_5947_)
);

NOR2X1 _15057_ (
    .A(_5536_),
    .B(_5533_),
    .Y(_5537_)
);

FILL FILL_3__16106_ (
);

INVX1 _10192_ (
    .A(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_1687_)
);

FILL FILL_5__10627_ (
);

FILL FILL_1__8749_ (
);

FILL FILL_1__8329_ (
);

FILL FILL_3__11661_ (
);

FILL FILL_3__11241_ (
);

FILL FILL_2__15939_ (
);

FILL FILL_2__15519_ (
);

FILL FILL_0__16133_ (
);

FILL FILL_2__10654_ (
);

FILL FILL_5__13099_ (
);

FILL FILL_2__10234_ (
);

FILL SFILL54040x71050 (
);

DFFSR _7399_ (
    .Q(\datapath_1.regfile_1.regOut[4] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_198_[17])
);

FILL FILL_3__9616_ (
);

FILL FILL_3_BUFX2_insert320 (
);

FILL FILL_3_BUFX2_insert321 (
);

FILL FILL_3_BUFX2_insert322 (
);

FILL FILL_5__14880_ (
);

FILL FILL_5__14460_ (
);

FILL FILL_3_BUFX2_insert323 (
);

FILL FILL_5__14040_ (
);

FILL FILL_3_BUFX2_insert324 (
);

INVX1 _8760_ (
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_956_)
);

FILL FILL_6__7621_ (
);

FILL FILL_3_BUFX2_insert325 (
);

FILL FILL_3_BUFX2_insert326 (
);

INVX1 _8340_ (
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_737_)
);

FILL FILL_3_BUFX2_insert327 (
);

FILL FILL_3_BUFX2_insert328 (
);

FILL FILL_4__13873_ (
);

FILL FILL_3_BUFX2_insert329 (
);

FILL FILL_4__13453_ (
);

FILL FILL_4__13033_ (
);

OAI21X1 _11397_ (
    .A(_2397_),
    .B(_2398_),
    .C(_2208_),
    .Y(_2514_)
);

FILL FILL_2__7613_ (
);

FILL FILL_3__12866_ (
);

FILL FILL_3__12446_ (
);

FILL FILL_3__12026_ (
);

FILL FILL_1__13480_ (
);

FILL FILL_4__7959_ (
);

FILL FILL_4__7119_ (
);

FILL FILL_2__11859_ (
);

FILL FILL_0__12893_ (
);

FILL FILL_2__11439_ (
);

FILL FILL_0__12473_ (
);

FILL FILL_2__11019_ (
);

FILL FILL_0__12053_ (
);

FILL FILL_6__16252_ (
);

FILL FILL_5__8090_ (
);

FILL FILL_4__8900_ (
);

FILL FILL_5__15665_ (
);

FILL FILL_5__15245_ (
);

FILL FILL_0__7859_ (
);

DFFSR _9965_ (
    .Q(\datapath_1.regfile_1.regOut[24] [23]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_1498_[23])
);

FILL FILL_0__7439_ (
);

FILL FILL_6__8826_ (
);

FILL SFILL98840x44050 (
);

OAI21X1 _9545_ (
    .A(_1356_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .C(_1357_),
    .Y(_1303_[27])
);

OAI21X1 _9125_ (
    .A(_1137_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .C(_1138_),
    .Y(_1108_[15])
);

FILL FILL_5__10380_ (
);

FILL FILL_1__8082_ (
);

FILL FILL_4__14658_ (
);

FILL FILL_4__14238_ (
);

FILL FILL_2__15692_ (
);

FILL FILL_2__15272_ (
);

FILL FILL_1__14685_ (
);

FILL FILL_1__14265_ (
);

FILL FILL_0_BUFX2_insert450 (
);

FILL FILL_0_BUFX2_insert451 (
);

FILL FILL_0_BUFX2_insert452 (
);

FILL FILL_0_BUFX2_insert453 (
);

FILL FILL_0_BUFX2_insert454 (
);

FILL FILL_0__13678_ (
);

NAND3X1 _13963_ (
    .A(_4463_),
    .B(_4464_),
    .C(_4462_),
    .Y(_4465_)
);

FILL FILL_0__13258_ (
);

FILL FILL_0_BUFX2_insert455 (
);

AOI22X1 _13543_ (
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .B(_3942__bF$buf0),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_4053_)
);

FILL FILL_0_BUFX2_insert456 (
);

OAI21X1 _13123_ (
    .A(_3712_),
    .B(PCEn_bF$buf1),
    .C(_3713_),
    .Y(_3685_[14])
);

FILL FILL_0_BUFX2_insert457 (
);

FILL FILL_0_BUFX2_insert458 (
);

FILL FILL_5__9295_ (
);

FILL FILL_0_BUFX2_insert459 (
);

FILL SFILL79160x82050 (
);

FILL FILL_6__12172_ (
);

FILL FILL_5__11585_ (
);

FILL FILL_1__9287_ (
);

FILL FILL_5__11165_ (
);

FILL FILL_2__16057_ (
);

FILL FILL_4__10998_ (
);

FILL FILL_4__7292_ (
);

FILL FILL_4__10578_ (
);

FILL FILL_4__10158_ (
);

FILL FILL_2__11192_ (
);

FILL FILL_5__7608_ (
);

FILL FILL_1__10185_ (
);

FILL FILL_6__10905_ (
);

INVX1 _14748_ (
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_5233_)
);

INVX1 _14328_ (
    .A(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_4822_)
);

FILL FILL_0__7192_ (
);

FILL FILL_1__16411_ (
);

FILL SFILL23880x18050 (
);

FILL FILL_3__10932_ (
);

FILL FILL_6__13797_ (
);

FILL FILL_3__10512_ (
);

FILL FILL_6__13377_ (
);

FILL FILL_0__15824_ (
);

FILL FILL_0__15404_ (
);

FILL FILL_2__8991_ (
);

FILL FILL_2__8571_ (
);

FILL FILL_4__8497_ (
);

FILL FILL_4__8077_ (
);

FILL FILL_2__12397_ (
);

FILL FILL_5__13731_ (
);

FILL FILL_5__13311_ (
);

INVX1 _7611_ (
    .A(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_373_)
);

FILL FILL_4__12724_ (
);

FILL FILL_4__12304_ (
);

FILL FILL_0__8397_ (
);

INVX1 _10668_ (
    .A(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_1923_)
);

FILL FILL_6__9364_ (
);

FILL SFILL23800x16050 (
);

INVX1 _10248_ (
    .A(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_1704_)
);

FILL FILL_3__11717_ (
);

FILL FILL_1__12751_ (
);

FILL FILL_4__15196_ (
);

FILL FILL_1__12331_ (
);

FILL FILL_2__9776_ (
);

FILL FILL_2__9356_ (
);

FILL FILL_0__11744_ (
);

FILL FILL_3__14189_ (
);

FILL FILL_0__11324_ (
);

FILL FILL_5__7361_ (
);

FILL SFILL74120x63050 (
);

FILL FILL_5__14936_ (
);

INVX1 _14081_ (
    .A(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_4580_)
);

FILL FILL_3__15970_ (
);

FILL FILL_5__14516_ (
);

FILL FILL_3__15550_ (
);

DFFSR _8816_ (
    .Q(\datapath_1.regfile_1.regOut[15] [26]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_913_[26])
);

FILL FILL_3__15130_ (
);

FILL FILL_1__7353_ (
);

FILL FILL_4__13929_ (
);

FILL FILL_2__14963_ (
);

FILL FILL_4__13509_ (
);

FILL FILL_2__14543_ (
);

FILL FILL_2__14123_ (
);

FILL FILL_3__7699_ (
);

FILL FILL_1__13956_ (
);

FILL FILL_1__13536_ (
);

FILL FILL_1__13116_ (
);

FILL FILL_3__8640_ (
);

DFFSR _12814_ (
    .Q(\datapath_1.PCJump [25]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3490_[23])
);

FILL FILL_3__8220_ (
);

FILL FILL_0__12529_ (
);

FILL FILL_0__12109_ (
);

FILL FILL_5__8986_ (
);

FILL FILL_5__8566_ (
);

FILL FILL_5__8146_ (
);

OAI22X1 _15286_ (
    .A(_5472__bF$buf2),
    .B(_4213_),
    .C(_4222_),
    .D(_5526__bF$buf4),
    .Y(_5761_)
);

FILL FILL_3__16335_ (
);

FILL FILL_1__8978_ (
);

FILL FILL_5__10436_ (
);

FILL FILL_3__11890_ (
);

FILL FILL_5__10016_ (
);

FILL FILL_1__8138_ (
);

FILL FILL_3__11470_ (
);

FILL SFILL74440x39050 (
);

FILL FILL_3__11050_ (
);

FILL FILL_2__15748_ (
);

FILL FILL_2__15328_ (
);

FILL FILL_4__6983_ (
);

FILL FILL_0__16362_ (
);

FILL SFILL38680x51050 (
);

FILL FILL_2__10883_ (
);

FILL FILL_2__10043_ (
);

FILL SFILL13800x14050 (
);

FILL FILL_3__9425_ (
);

FILL FILL_3__9005_ (
);

FILL FILL_0__6883_ (
);

FILL FILL_4__13682_ (
);

FILL FILL_4__13262_ (
);

FILL FILL_2__7842_ (
);

FILL FILL_2__7422_ (
);

FILL FILL_3__12255_ (
);

FILL FILL_4__7348_ (
);

FILL FILL112360x59050 (
);

FILL FILL_2__11668_ (
);

FILL FILL_2__11248_ (
);

FILL FILL_0__12282_ (
);

FILL SFILL49000x3050 (
);

FILL SFILL64040x68050 (
);

FILL FILL_5__15894_ (
);

FILL SFILL89240x1050 (
);

FILL FILL_5__15474_ (
);

FILL SFILL88920x4050 (
);

FILL FILL_5__15054_ (
);

FILL FILL_6__8635_ (
);

FILL FILL_0__7248_ (
);

OAI21X1 _9774_ (
    .A(_1468_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1469_),
    .Y(_1433_[18])
);

OAI21X1 _9354_ (
    .A(_1249_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1250_),
    .Y(_1238_[6])
);

FILL FILL_4__14887_ (
);

FILL FILL_4__14467_ (
);

FILL FILL_1__11602_ (
);

FILL FILL_4__14047_ (
);

FILL FILL_2__15081_ (
);

FILL FILL_2__8627_ (
);

FILL FILL_2__8207_ (
);

FILL FILL_1__14494_ (
);

FILL FILL_1__14074_ (
);

NAND3X1 _13772_ (
    .A(_4276_),
    .B(_4277_),
    .C(_4275_),
    .Y(_4278_)
);

FILL FILL_0__13487_ (
);

NOR2X1 _13352_ (
    .A(_3798_),
    .B(_3865_),
    .Y(\datapath_1.regfile_1.regEn [26])
);

FILL FILL112360x14050 (
);

FILL FILL_3__14821_ (
);

FILL FILL_3__14401_ (
);

FILL FILL_4__9914_ (
);

FILL FILL_2__13814_ (
);

FILL FILL_5__16259_ (
);

FILL SFILL64040x23050 (
);

FILL FILL_5__11394_ (
);

FILL FILL_1__9096_ (
);

FILL FILL_2__16286_ (
);

FILL FILL_4__10387_ (
);

FILL SFILL89240x72050 (
);

FILL FILL_1__15699_ (
);

FILL FILL_1__15279_ (
);

FILL FILL_5__7837_ (
);

FILL FILL_5__7417_ (
);

FILL SFILL113880x2050 (
);

NOR2X1 _14977_ (
    .A(_5457_),
    .B(_5445_),
    .Y(_5458_)
);

AOI22X1 _14557_ (
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .B(_4005__bF$buf3),
    .C(_3950__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_5046_)
);

INVX1 _14137_ (
    .A(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_4635_)
);

FILL FILL_3__15606_ (
);

FILL FILL_1__16220_ (
);

FILL FILL_1__7829_ (
);

FILL FILL_3__10321_ (
);

FILL FILL_0__15633_ (
);

FILL FILL_0__15213_ (
);

FILL FILL_5__12599_ (
);

FILL SFILL54040x66050 (
);

FILL FILL_2__8380_ (
);

FILL FILL_5__12179_ (
);

BUFX2 _6899_ (
    .A(_2_[29]),
    .Y(memoryWriteData[29])
);

FILL FILL_5__13960_ (
);

FILL FILL_5__13540_ (
);

FILL FILL_5__13120_ (
);

INVX1 _7840_ (
    .A(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_485_)
);

FILL SFILL58360x74050 (
);

INVX1 _7420_ (
    .A(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_266_)
);

FILL FILL_1__11199_ (
);

DFFSR _7000_ (
    .Q(\datapath_1.regfile_1.regOut[1] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_3_[2])
);

FILL FILL_4__12953_ (
);

FILL FILL_4__12533_ (
);

FILL FILL_4__12113_ (
);

INVX2 _10897_ (
    .A(\control_1.reg_state.dout [2]),
    .Y(_2046_)
);

DFFSR _10477_ (
    .Q(\datapath_1.regfile_1.regOut[28] [23]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_1758_[23])
);

OAI21X1 _10057_ (
    .A(_1616_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .C(_1617_),
    .Y(_1563_[27])
);

FILL FILL_3__11946_ (
);

FILL FILL_1__12980_ (
);

FILL FILL_3__11526_ (
);

FILL FILL_3__11106_ (
);

FILL FILL_1__12140_ (
);

FILL FILL_2__10939_ (
);

FILL FILL_0__11973_ (
);

FILL FILL_2__10519_ (
);

FILL FILL_2__9165_ (
);

FILL FILL_0__11553_ (
);

FILL FILL_0__11133_ (
);

FILL SFILL58760x43050 (
);

FILL FILL_5__7590_ (
);

FILL FILL_6__15332_ (
);

FILL SFILL54040x21050 (
);

FILL FILL_5__7170_ (
);

FILL FILL_5__14745_ (
);

FILL FILL_0__6939_ (
);

FILL FILL_5__14325_ (
);

OAI21X1 _8625_ (
    .A(_885_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_886_),
    .Y(_848_[19])
);

OAI21X1 _8205_ (
    .A(_666_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .C(_667_),
    .Y(_653_[7])
);

FILL FILL_1__7582_ (
);

FILL FILL_1__7162_ (
);

FILL FILL_4__13738_ (
);

FILL FILL_4__13318_ (
);

FILL FILL_2__14772_ (
);

FILL FILL_2__14352_ (
);

FILL FILL_3__7088_ (
);

FILL FILL_1__13765_ (
);

FILL FILL_1__13345_ (
);

FILL SFILL109480x50 (
);

FILL FILL_0__12758_ (
);

OAI21X1 _12623_ (
    .A(_3460_),
    .B(vdd),
    .C(_3461_),
    .Y(_3425_[18])
);

FILL FILL_0__12338_ (
);

FILL SFILL33880x1050 (
);

NAND2X1 _12203_ (
    .A(ALUSrcA_bF$buf6),
    .B(\datapath_1.a [29]),
    .Y(_3189_)
);

FILL FILL_5__8375_ (
);

FILL SFILL44040x64050 (
);

OAI22X1 _15095_ (
    .A(_3991_),
    .B(_5539__bF$buf2),
    .C(_5469__bF$buf2),
    .D(_4011_),
    .Y(_5574_)
);

FILL FILL_3__16144_ (
);

FILL SFILL8120x65050 (
);

FILL FILL_5__10665_ (
);

FILL FILL_1__8787_ (
);

FILL FILL_1__8367_ (
);

FILL FILL_5__10245_ (
);

FILL FILL_2__15977_ (
);

FILL FILL_2__15557_ (
);

FILL FILL_2__15137_ (
);

FILL FILL_0__16171_ (
);

FILL FILL_2__10692_ (
);

FILL FILL_2__10272_ (
);

FILL SFILL44440x33050 (
);

FILL FILL_3__9654_ (
);

FILL FILL_3_BUFX2_insert700 (
);

INVX1 _13828_ (
    .A(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_4333_)
);

FILL FILL_3_BUFX2_insert701 (
);

FILL FILL_3__9234_ (
);

NAND2X1 _13408_ (
    .A(_3919_),
    .B(_3917_),
    .Y(_3920_)
);

FILL FILL_3_BUFX2_insert702 (
);

FILL FILL_3_BUFX2_insert703 (
);

FILL FILL_3_BUFX2_insert704 (
);

FILL FILL_1__15911_ (
);

FILL FILL_3_BUFX2_insert705 (
);

FILL FILL_3_BUFX2_insert706 (
);

FILL FILL_3_BUFX2_insert707 (
);

FILL FILL_3_BUFX2_insert708 (
);

FILL FILL_6__12877_ (
);

FILL SFILL109400x51050 (
);

FILL FILL_3_BUFX2_insert709 (
);

FILL FILL_4__13491_ (
);

FILL FILL_0__14904_ (
);

FILL FILL_2__7231_ (
);

FILL FILL_3__12484_ (
);

FILL FILL_3__12064_ (
);

FILL FILL_4__7997_ (
);

FILL FILL_4__7577_ (
);

FILL FILL_2__11897_ (
);

FILL FILL_2__11477_ (
);

FILL FILL_2__11057_ (
);

FILL FILL_0__12091_ (
);

FILL FILL_4__11804_ (
);

FILL FILL_5__15283_ (
);

FILL FILL_0__7477_ (
);

FILL FILL_0__7057_ (
);

FILL FILL_6__8444_ (
);

DFFSR _9583_ (
    .Q(\datapath_1.regfile_1.regOut[21] [25]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_1303_[25])
);

NAND2X1 _9163_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1164_)
);

FILL FILL_4__14696_ (
);

FILL FILL_1__11831_ (
);

FILL FILL_4__14276_ (
);

FILL FILL_1__11411_ (
);

FILL SFILL69160x75050 (
);

FILL FILL_2__8856_ (
);

FILL FILL_0__10824_ (
);

FILL FILL_3__13689_ (
);

FILL FILL_3__13269_ (
);

FILL FILL_0__10404_ (
);

FILL FILL_2__8016_ (
);

FILL FILL_5__6861_ (
);

FILL FILL_0_BUFX2_insert830 (
);

FILL FILL_0_BUFX2_insert831 (
);

FILL FILL_0_BUFX2_insert832 (
);

FILL FILL_0_BUFX2_insert833 (
);

FILL FILL_0_BUFX2_insert834 (
);

FILL FILL_0__13296_ (
);

FILL FILL_0_BUFX2_insert835 (
);

AOI22X1 _13581_ (
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .B(_4090_),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_4091_)
);

FILL FILL_0_BUFX2_insert836 (
);

NAND2X1 _13161_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_pcsrc.dout [27]),
    .Y(_3739_)
);

FILL FILL_0_BUFX2_insert837 (
);

FILL FILL_0_BUFX2_insert838 (
);

FILL FILL_3__14630_ (
);

FILL FILL_3__14210_ (
);

FILL FILL_0_BUFX2_insert839 (
);

FILL FILL_1__6853_ (
);

FILL FILL_4__9723_ (
);

FILL FILL_2__13623_ (
);

FILL FILL_5__16068_ (
);

FILL FILL_6__9229_ (
);

FILL FILL_1__12616_ (
);

FILL FILL_2__16095_ (
);

FILL FILL_4__10196_ (
);

FILL FILL_3__7720_ (
);

FILL FILL_0__9623_ (
);

FILL SFILL69160x30050 (
);

FILL FILL_3__7300_ (
);

FILL FILL_0__11609_ (
);

FILL FILL_1__15088_ (
);

FILL FILL_5__7226_ (
);

FILL FILL_4__16002_ (
);

FILL SFILL78840x35050 (
);

INVX1 _14786_ (
    .A(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_5271_)
);

NOR2X1 _14366_ (
    .A(_4858_),
    .B(_4855_),
    .Y(_4859_)
);

FILL SFILL74120x13050 (
);

FILL FILL_3__15835_ (
);

FILL SFILL28920x2050 (
);

FILL FILL_3__15415_ (
);

FILL FILL_3__10970_ (
);

FILL FILL_3__10550_ (
);

FILL FILL_1__7218_ (
);

FILL SFILL28840x7050 (
);

FILL FILL_3__10130_ (
);

FILL FILL_2__14828_ (
);

FILL FILL_2__14408_ (
);

FILL FILL_0__15862_ (
);

FILL SFILL99320x62050 (
);

FILL FILL_0__15442_ (
);

FILL FILL_0__15022_ (
);

FILL SFILL28760x82050 (
);

FILL SFILL8760x3050 (
);

FILL FILL_3__8505_ (
);

FILL SFILL59160x73050 (
);

FILL SFILL68680x4050 (
);

FILL SFILL38280x32050 (
);

FILL SFILL8680x8050 (
);

FILL SFILL68840x78050 (
);

FILL FILL_4__12762_ (
);

FILL FILL_6__11308_ (
);

FILL FILL_4__12342_ (
);

FILL SFILL64120x56050 (
);

OAI21X1 _10286_ (
    .A(_1728_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1729_),
    .Y(_1693_[18])
);

FILL FILL_2__6922_ (
);

FILL FILL_3__11755_ (
);

FILL FILL_3__11335_ (
);

FILL FILL_4__6848_ (
);

FILL FILL_0__16227_ (
);

FILL FILL_2__10748_ (
);

FILL FILL_2__9394_ (
);

FILL FILL_0__11782_ (
);

FILL FILL_0__11362_ (
);

FILL FILL_6__15981_ (
);

FILL FILL_5__14974_ (
);

FILL FILL_5__14554_ (
);

FILL FILL_5__14134_ (
);

FILL FILL_6__7715_ (
);

OAI21X1 _8854_ (
    .A(_997_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_998_),
    .Y(_978_[10])
);

DFFSR _8434_ (
    .Q(\datapath_1.regfile_1.regOut[12] [28]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_718_[28])
);

NAND2X1 _8014_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_581_)
);

FILL FILL_4__13967_ (
);

FILL FILL_4__13547_ (
);

FILL FILL_2__14581_ (
);

FILL FILL_4__13127_ (
);

FILL FILL_2__14161_ (
);

FILL FILL_2__7707_ (
);

FILL SFILL64120x11050 (
);

FILL FILL_1__13994_ (
);

FILL FILL_1__13574_ (
);

FILL FILL_1__13154_ (
);

FILL FILL_0__12987_ (
);

FILL FILL_0__12567_ (
);

OAI21X1 _12852_ (
    .A(_3572_),
    .B(vdd),
    .C(_3573_),
    .Y(_3555_[9])
);

OAI21X1 _12432_ (
    .A(_3352_),
    .B(MemToReg_bF$buf7),
    .C(_3353_),
    .Y(\datapath_1.mux_wd3.dout [29])
);

FILL FILL_0__12147_ (
);

FILL SFILL89320x60050 (
);

NAND3X1 _12012_ (
    .A(PCSource_1_bF$buf2),
    .B(\aluControl_1.inst [4]),
    .C(_3034__bF$buf4),
    .Y(_3055_)
);

FILL FILL_3__13901_ (
);

FILL FILL_5__8184_ (
);

FILL FILL_5_BUFX2_insert230 (
);

FILL FILL_5__15759_ (
);

FILL FILL_5_BUFX2_insert231 (
);

FILL FILL_5__15339_ (
);

FILL FILL_5_BUFX2_insert232 (
);

FILL FILL_5_BUFX2_insert233 (
);

FILL FILL_3__16373_ (
);

NAND2X1 _9639_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1400_)
);

FILL FILL_5_BUFX2_insert234 (
);

FILL SFILL18760x80050 (
);

FILL SFILL64040x18050 (
);

NAND2X1 _9219_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1181_)
);

FILL FILL_5__10894_ (
);

FILL FILL_5_BUFX2_insert235 (
);

FILL FILL_5_BUFX2_insert236 (
);

FILL FILL_1__8596_ (
);

FILL FILL_5_BUFX2_insert1020 (
);

FILL FILL_5__10054_ (
);

FILL FILL_5_BUFX2_insert237 (
);

FILL FILL_5_BUFX2_insert238 (
);

FILL FILL_5_BUFX2_insert1021 (
);

FILL FILL_5_BUFX2_insert1022 (
);

FILL FILL_5_BUFX2_insert239 (
);

FILL FILL_2__15786_ (
);

FILL FILL_2__15366_ (
);

FILL FILL_5_BUFX2_insert1023 (
);

FILL FILL_5_BUFX2_insert1024 (
);

FILL FILL_5_BUFX2_insert1025 (
);

FILL FILL_5_BUFX2_insert1026 (
);

FILL FILL_5_BUFX2_insert1027 (
);

FILL FILL_5_BUFX2_insert1028 (
);

FILL SFILL54120x54050 (
);

FILL FILL_5_BUFX2_insert1029 (
);

FILL FILL_1__14779_ (
);

FILL FILL_1__14359_ (
);

FILL FILL_5__6917_ (
);

FILL FILL_3__9883_ (
);

FILL FILL_3__9463_ (
);

AOI21X1 _13637_ (
    .A(_4120_),
    .B(_4145_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [3])
);

FILL FILL_3__9043_ (
);

INVX1 _13217_ (
    .A(_3759_),
    .Y(_3760_)
);

FILL FILL_1__15720_ (
);

FILL FILL_5__9389_ (
);

FILL FILL_1__15300_ (
);

FILL FILL_1__6909_ (
);

FILL FILL_0__14713_ (
);

FILL FILL_2__7880_ (
);

FILL FILL_5__11679_ (
);

FILL FILL_2__7460_ (
);

FILL FILL_5__11259_ (
);

FILL FILL_2__7040_ (
);

FILL FILL_3__12293_ (
);

FILL FILL_2__11286_ (
);

FILL FILL_5__12620_ (
);

FILL FILL_5__12200_ (
);

INVX1 _6920_ (
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_14_)
);

FILL SFILL89240x22050 (
);

FILL FILL_1__10699_ (
);

FILL FILL_2_BUFX2_insert360 (
);

FILL FILL_1__10279_ (
);

FILL FILL_2_BUFX2_insert361 (
);

FILL FILL_2_BUFX2_insert362 (
);

FILL FILL_2_BUFX2_insert363 (
);

FILL FILL_4__11613_ (
);

FILL FILL_2_BUFX2_insert364 (
);

FILL FILL_2_BUFX2_insert365 (
);

FILL FILL_2_BUFX2_insert366 (
);

FILL FILL_5__15092_ (
);

FILL FILL_0__7286_ (
);

FILL FILL_2_BUFX2_insert367 (
);

FILL FILL_2_BUFX2_insert368 (
);

NAND2X1 _9392_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1276_)
);

FILL FILL_2_BUFX2_insert369 (
);

FILL SFILL18680x42050 (
);

FILL FILL_1__11640_ (
);

FILL FILL_1__11220_ (
);

FILL FILL_4__14085_ (
);

FILL FILL_0__15918_ (
);

FILL SFILL79640x79050 (
);

FILL FILL_2__8245_ (
);

FILL FILL_0__10633_ (
);

FILL FILL_3__13498_ (
);

FILL FILL111960x71050 (
);

FILL SFILL54040x16050 (
);

NAND2X1 _13390_ (
    .A(_3898_),
    .B(_3901_),
    .Y(_3902_)
);

FILL FILL_5__13825_ (
);

FILL FILL_5__13405_ (
);

OAI21X1 _7705_ (
    .A(_414_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_415_),
    .Y(_393_[11])
);

FILL SFILL79240x65050 (
);

FILL FILL_2_BUFX2_insert1084 (
);

FILL FILL_4__9532_ (
);

FILL FILL_2_BUFX2_insert1085 (
);

FILL FILL_2_BUFX2_insert1086 (
);

FILL FILL_4__9112_ (
);

FILL FILL_2_BUFX2_insert1087 (
);

FILL FILL_2__13852_ (
);

FILL FILL_2__13432_ (
);

FILL FILL_2_BUFX2_insert1088 (
);

FILL FILL_5__16297_ (
);

FILL FILL_2_BUFX2_insert1089 (
);

FILL FILL_2__13012_ (
);

FILL FILL_6__9038_ (
);

FILL FILL_1__12845_ (
);

FILL FILL_1__12425_ (
);

FILL FILL_1__12005_ (
);

FILL FILL_0__9852_ (
);

FILL FILL_0__11838_ (
);

FILL FILL_0__11418_ (
);

FILL FILL_0__9012_ (
);

OAI21X1 _11703_ (
    .A(_2801_),
    .B(_2509_),
    .C(_2800_),
    .Y(_2802_)
);

FILL FILL_5__7875_ (
);

FILL SFILL44040x59050 (
);

FILL FILL_5__7455_ (
);

FILL FILL_4__16231_ (
);

FILL FILL_5__7035_ (
);

NAND2X1 _14595_ (
    .A(_5083_),
    .B(_5076_),
    .Y(_5084_)
);

INVX1 _14175_ (
    .A(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_4672_)
);

FILL FILL_3__15644_ (
);

FILL FILL_3__15224_ (
);

FILL FILL_1__7867_ (
);

FILL FILL_1__7447_ (
);

FILL FILL_2__14637_ (
);

FILL SFILL79240x20050 (
);

FILL FILL_0__15671_ (
);

FILL FILL_2__14217_ (
);

FILL FILL_0__15251_ (
);

FILL FILL_1_BUFX2_insert380 (
);

FILL FILL_1_BUFX2_insert381 (
);

FILL FILL_3__8734_ (
);

NAND2X1 _12908_ (
    .A(vdd),
    .B(\datapath_1.rd1 [28]),
    .Y(_3611_)
);

FILL FILL_1_BUFX2_insert382 (
);

FILL FILL_3__8314_ (
);

FILL FILL_1_BUFX2_insert383 (
);

FILL SFILL8520x29050 (
);

FILL FILL_1_BUFX2_insert384 (
);

FILL FILL_1_BUFX2_insert385 (
);

FILL FILL_1_BUFX2_insert386 (
);

FILL FILL_1_BUFX2_insert387 (
);

FILL FILL_1_BUFX2_insert388 (
);

FILL SFILL109400x46050 (
);

FILL FILL_6__11957_ (
);

FILL FILL_1_BUFX2_insert389 (
);

FILL FILL_4__12991_ (
);

FILL FILL_4__12571_ (
);

FILL FILL_4__12151_ (
);

FILL FILL_3__16009_ (
);

DFFSR _10095_ (
    .Q(\datapath_1.regfile_1.regOut[25] [25]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_1563_[25])
);

FILL FILL_3__11984_ (
);

FILL FILL_5__9601_ (
);

FILL FILL_3__11564_ (
);

FILL FILL_3__11144_ (
);

FILL SFILL69240x63050 (
);

FILL FILL_0__16036_ (
);

INVX1 _16321_ (
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_6832_)
);

FILL FILL_2__10977_ (
);

FILL FILL_2__10557_ (
);

FILL FILL_2__10137_ (
);

FILL FILL_0__11591_ (
);

FILL FILL_0__11171_ (
);

FILL FILL_3__9939_ (
);

FILL FILL_3__9519_ (
);

FILL FILL_5__14783_ (
);

FILL FILL_5__14363_ (
);

FILL FILL_0__6977_ (
);

DFFSR _8663_ (
    .Q(\datapath_1.regfile_1.regOut[14] [1]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_848_[1])
);

NAND2X1 _8243_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_693_)
);

FILL SFILL38760x79050 (
);

FILL FILL_1__10911_ (
);

FILL FILL_4__13776_ (
);

FILL FILL_4__13356_ (
);

FILL SFILL34040x57050 (
);

FILL FILL_2__14390_ (
);

FILL FILL_2__7936_ (
);

FILL FILL_3__12769_ (
);

FILL FILL_3__12349_ (
);

FILL FILL_1__13383_ (
);

NAND2X1 _12661_ (
    .A(vdd),
    .B(memoryOutData[31]),
    .Y(_3487_)
);

FILL FILL_0__12376_ (
);

AOI22X1 _12241_ (
    .A(_2_[6]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf0),
    .D(\aluControl_1.inst [4]),
    .Y(_3220_)
);

FILL FILL_3__13710_ (
);

FILL FILL_6__16155_ (
);

FILL FILL_5__15988_ (
);

FILL FILL_2__12703_ (
);

FILL FILL_5__15568_ (
);

FILL FILL_5__15148_ (
);

NAND2X1 _9868_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1512_)
);

FILL FILL_3__16182_ (
);

DFFSR _9448_ (
    .Q(\datapath_1.regfile_1.regOut[20] [18]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_1238_[18])
);

INVX1 _9028_ (
    .A(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_1094_)
);

FILL FILL_5__10283_ (
);

FILL FILL_2__15595_ (
);

FILL FILL_2__15175_ (
);

FILL SFILL99400x50050 (
);

FILL SFILL69160x25050 (
);

FILL FILL_0__8703_ (
);

FILL FILL_1__14588_ (
);

FILL FILL_1__14168_ (
);

FILL FILL_4__15922_ (
);

FILL FILL_4__15502_ (
);

INVX1 _13866_ (
    .A(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_4370_)
);

FILL FILL_3__9272_ (
);

INVX1 _13446_ (
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_3958_)
);

INVX1 _13026_ (
    .A(_2_[25]),
    .Y(_3669_)
);

FILL FILL_3__14915_ (
);

FILL FILL_6__12495_ (
);

FILL FILL_6__12075_ (
);

FILL FILL_2__13908_ (
);

FILL SFILL99320x57050 (
);

FILL FILL_0__14942_ (
);

FILL FILL_0__14522_ (
);

FILL FILL_0__14102_ (
);

FILL FILL_5__11488_ (
);

FILL FILL_5__11068_ (
);

FILL FILL_4__7195_ (
);

FILL SFILL28760x77050 (
);

FILL FILL_0__9908_ (
);

FILL SFILL59160x68050 (
);

FILL FILL_2__11095_ (
);

FILL SFILL83640x79050 (
);

FILL FILL_4__11842_ (
);

FILL FILL_4__11422_ (
);

FILL FILL_4__11002_ (
);

FILL FILL_0__7095_ (
);

FILL FILL_1__16314_ (
);

FILL FILL_3__10835_ (
);

FILL FILL_3__10415_ (
);

FILL FILL_0__15727_ (
);

FILL FILL_0__15307_ (
);

FILL FILL_2__8894_ (
);

FILL FILL_2__8474_ (
);

FILL SFILL99320x12050 (
);

FILL FILL_0__10442_ (
);

FILL FILL_2__8054_ (
);

FILL FILL_0__10022_ (
);

FILL FILL_6__14641_ (
);

FILL FILL_6__14221_ (
);

FILL FILL_5__13634_ (
);

FILL FILL_5__13214_ (
);

FILL SFILL28760x32050 (
);

OAI21X1 _7934_ (
    .A(_526_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_527_),
    .Y(_523_[2])
);

DFFSR _7514_ (
    .Q(\datapath_1.regfile_1.regOut[5] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_263_[4])
);

FILL FILL_1__6891_ (
);

FILL FILL_4__9761_ (
);

FILL FILL_4__9341_ (
);

FILL FILL_4__12627_ (
);

FILL FILL_2__13661_ (
);

FILL FILL_4__12207_ (
);

FILL FILL_2__13241_ (
);

FILL FILL_1__12654_ (
);

FILL FILL_1__12234_ (
);

FILL FILL_4__15099_ (
);

FILL FILL_0__9661_ (
);

FILL FILL_2__9679_ (
);

INVX1 _11932_ (
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_2996_)
);

FILL FILL_0__9241_ (
);

FILL FILL_2__9259_ (
);

FILL FILL_0__11647_ (
);

FILL FILL_0__11227_ (
);

NOR2X1 _11512_ (
    .A(_2442_),
    .B(_2603_),
    .Y(_2624_)
);

FILL FILL_5__7684_ (
);

FILL FILL_4__16040_ (
);

FILL FILL_6__10981_ (
);

FILL FILL_5__14839_ (
);

FILL FILL_5__14419_ (
);

FILL FILL_3__15873_ (
);

FILL FILL_3__15453_ (
);

FILL SFILL18760x75050 (
);

NAND2X1 _8719_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_929_)
);

FILL FILL_3__15033_ (
);

FILL FILL_1__7676_ (
);

FILL FILL_2__14866_ (
);

FILL FILL_2__14446_ (
);

FILL FILL_2__14026_ (
);

FILL FILL_0__15480_ (
);

FILL FILL_0__15060_ (
);

FILL SFILL73640x77050 (
);

FILL SFILL54120x49050 (
);

FILL FILL_1__13859_ (
);

FILL FILL_1__13439_ (
);

FILL FILL_1__13019_ (
);

FILL FILL_3__8963_ (
);

NAND2X1 _12717_ (
    .A(IRWrite_bF$buf7),
    .B(memoryOutData[7]),
    .Y(_3504_)
);

FILL FILL_3__8123_ (
);

FILL FILL_5__8889_ (
);

FILL FILL_1__14800_ (
);

FILL FILL_5__8469_ (
);

FILL FILL_1_BUFX2_insert50 (
);

FILL FILL_1_BUFX2_insert51 (
);

FILL FILL_1_BUFX2_insert52 (
);

FILL FILL_1_BUFX2_insert53 (
);

INVX1 _15189_ (
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_5666_)
);

FILL FILL_4__12380_ (
);

FILL FILL_1_BUFX2_insert54 (
);

FILL FILL_1_BUFX2_insert55 (
);

FILL FILL_1_BUFX2_insert56 (
);

FILL FILL_1_BUFX2_insert57 (
);

FILL FILL_3__16238_ (
);

FILL FILL_1_BUFX2_insert58 (
);

FILL FILL_1_BUFX2_insert59 (
);

FILL FILL_2__6960_ (
);

FILL FILL_5__10759_ (
);

FILL FILL_3__11793_ (
);

FILL FILL_3__11373_ (
);

FILL FILL_5__9410_ (
);

FILL SFILL18760x30050 (
);

FILL FILL_4__6886_ (
);

FILL FILL_0__16265_ (
);

AOI22X1 _16130_ (
    .A(_5649_),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .C(\datapath_1.regfile_1.regOut[21] [27]),
    .D(_5685_),
    .Y(_6583_)
);

FILL FILL_2__10786_ (
);

FILL FILL_2__10366_ (
);

FILL FILL_5__11700_ (
);

FILL FILL_1__9402_ (
);

FILL SFILL89240x17050 (
);

FILL FILL_3__9748_ (
);

FILL FILL_5__14592_ (
);

FILL FILL_5__14172_ (
);

NAND2X1 _8892_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1024_)
);

NAND2X1 _8472_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_805_)
);

DFFSR _8052_ (
    .Q(\datapath_1.regfile_1.regOut[9] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_523_[30])
);

FILL SFILL79320x53050 (
);

FILL SFILL18680x37050 (
);

FILL FILL_4__13585_ (
);

FILL FILL_1__10300_ (
);

FILL FILL_4__13165_ (
);

FILL FILL_3__12998_ (
);

FILL FILL_2__7745_ (
);

FILL FILL_3__12578_ (
);

FILL FILL_2__7325_ (
);

FILL FILL111960x66050 (
);

FILL FILL_3__12158_ (
);

NAND2X1 _12890_ (
    .A(vdd),
    .B(\datapath_1.rd1 [22]),
    .Y(_3599_)
);

FILL FILL_0__12185_ (
);

NAND2X1 _12470_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [10]),
    .Y(_3380_)
);

NAND3X1 _12050_ (
    .A(_3081_),
    .B(_3082_),
    .C(_3083_),
    .Y(\datapath_1.mux_pcsrc.dout [15])
);

FILL FILL_5__12905_ (
);

FILL FILL_4__8612_ (
);

FILL FILL_5_BUFX2_insert610 (
);

FILL FILL_5__15797_ (
);

FILL FILL_5_BUFX2_insert611 (
);

FILL FILL_5__15377_ (
);

FILL FILL_2__12512_ (
);

FILL FILL_5_BUFX2_insert612 (
);

FILL FILL_5_BUFX2_insert613 (
);

INVX1 _9677_ (
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_1425_)
);

FILL FILL_5_BUFX2_insert614 (
);

FILL FILL_6__8118_ (
);

FILL FILL_5_BUFX2_insert615 (
);

INVX1 _9257_ (
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_1206_)
);

FILL FILL_5_BUFX2_insert616 (
);

FILL FILL_5_BUFX2_insert617 (
);

FILL FILL_1__11925_ (
);

FILL FILL_5_BUFX2_insert618 (
);

FILL FILL_5_BUFX2_insert619 (
);

FILL FILL_1__11505_ (
);

FILL FILL_0__10918_ (
);

FILL FILL_0__8512_ (
);

FILL FILL_1__14397_ (
);

FILL FILL_5__6955_ (
);

FILL FILL_4__15731_ (
);

FILL FILL_4__15311_ (
);

FILL FILL111960x21050 (
);

INVX1 _13675_ (
    .A(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_4183_)
);

FILL FILL_3__9081_ (
);

NAND2X1 _13255_ (
    .A(\datapath_1.a3 [4]),
    .B(RegWrite_bF$buf0),
    .Y(_3798_)
);

FILL FILL_3__14724_ (
);

FILL FILL_3__14304_ (
);

FILL FILL_1__6947_ (
);

FILL FILL_2__13717_ (
);

FILL FILL_0__14751_ (
);

FILL FILL_0__14331_ (
);

FILL FILL_5__11297_ (
);

FILL FILL_2__16189_ (
);

FILL FILL_3__7814_ (
);

FILL FILL_2_BUFX2_insert740 (
);

FILL FILL_2_BUFX2_insert741 (
);

FILL FILL_2_BUFX2_insert742 (
);

FILL FILL_2_BUFX2_insert743 (
);

FILL FILL_2_BUFX2_insert744 (
);

FILL FILL_4__11651_ (
);

FILL FILL_2_BUFX2_insert745 (
);

FILL FILL_4__11231_ (
);

FILL FILL_3__15929_ (
);

FILL FILL_2_BUFX2_insert746 (
);

FILL FILL_3__15509_ (
);

FILL FILL_2_BUFX2_insert747 (
);

FILL FILL_2_BUFX2_insert748 (
);

FILL FILL_2_BUFX2_insert749 (
);

FILL FILL_1__16123_ (
);

FILL FILL_3__10644_ (
);

FILL SFILL69240x58050 (
);

FILL SFILL69720x20050 (
);

FILL FILL_0__15956_ (
);

FILL FILL_0__15536_ (
);

AOI21X1 _15821_ (
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .B(_5606_),
    .C(_6281_),
    .Y(_6282_)
);

OAI22X1 _15401_ (
    .A(_4346_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf0),
    .D(_5872_),
    .Y(_5873_)
);

FILL FILL_0__15116_ (
);

FILL FILL_0__10671_ (
);

FILL FILL_0__10251_ (
);

FILL FILL_5__13863_ (
);

FILL FILL_5__13443_ (
);

FILL FILL_5__13023_ (
);

NAND2X1 _7743_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_441_)
);

NAND2X1 _7323_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_222_)
);

FILL FILL_4__9990_ (
);

FILL FILL_4__9150_ (
);

FILL FILL_4__12856_ (
);

FILL FILL_4__12436_ (
);

FILL FILL_2__13890_ (
);

FILL FILL_4__12016_ (
);

FILL FILL_2__13470_ (
);

FILL FILL_3__11849_ (
);

FILL FILL_1__12883_ (
);

FILL FILL_3__11429_ (
);

FILL FILL_1__12463_ (
);

FILL FILL_3__11009_ (
);

FILL FILL_1__12043_ (
);

FILL SFILL99000x76050 (
);

FILL FILL_0__9890_ (
);

FILL FILL_2__9488_ (
);

FILL FILL_0__11876_ (
);

FILL FILL_0__9470_ (
);

FILL SFILL69240x13050 (
);

OAI21X1 _11741_ (
    .A(_2827_),
    .B(_2828_),
    .C(_2837_),
    .Y(\datapath_1.ALUResult [9])
);

FILL FILL_0__11456_ (
);

FILL FILL_0__11036_ (
);

NOR2X1 _11321_ (
    .A(_2289_),
    .B(_2439_),
    .Y(_2440_)
);

FILL FILL_5__7493_ (
);

FILL FILL_5__7073_ (
);

FILL SFILL93720x24050 (
);

FILL FILL_5__14648_ (
);

FILL SFILL3800x78050 (
);

FILL FILL_3__15682_ (
);

FILL FILL_5__14228_ (
);

DFFSR _8948_ (
    .Q(\datapath_1.regfile_1.regOut[16] [30]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_978_[30])
);

FILL FILL_3__15262_ (
);

INVX1 _8528_ (
    .A(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_842_)
);

INVX1 _8108_ (
    .A(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_623_)
);

FILL FILL_1__7485_ (
);

FILL FILL_1__7065_ (
);

FILL FILL_2__14675_ (
);

FILL FILL_2__14255_ (
);

FILL SFILL19160x60050 (
);

FILL FILL_1__13668_ (
);

FILL FILL_1__13248_ (
);

FILL FILL_1_BUFX2_insert760 (
);

FILL FILL_3__8772_ (
);

FILL FILL_1_BUFX2_insert761 (
);

FILL FILL_3__8352_ (
);

FILL FILL_1_BUFX2_insert762 (
);

DFFSR _12946_ (
    .Q(\datapath_1.a [27]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_3555_[27])
);

INVX1 _12526_ (
    .A(ALUOut[29]),
    .Y(_3417_)
);

FILL FILL_1_BUFX2_insert763 (
);

FILL FILL_1_BUFX2_insert764 (
);

NAND3X1 _12106_ (
    .A(_3123_),
    .B(_3124_),
    .C(_3125_),
    .Y(\datapath_1.mux_pcsrc.dout [29])
);

FILL FILL_1_BUFX2_insert765 (
);

FILL FILL_1_BUFX2_insert766 (
);

FILL FILL_5__8698_ (
);

FILL SFILL38360x15050 (
);

FILL FILL_1_BUFX2_insert767 (
);

FILL FILL_1_BUFX2_insert768 (
);

FILL FILL_1_BUFX2_insert769 (
);

FILL FILL_0__13602_ (
);

FILL FILL_3__16047_ (
);

FILL FILL_5__10988_ (
);

FILL FILL_5__10568_ (
);

FILL FILL_5__10148_ (
);

FILL FILL_3__11182_ (
);

FILL FILL_0__16074_ (
);

FILL FILL_2__10175_ (
);

FILL FILL_1__9631_ (
);

FILL SFILL104280x45050 (
);

FILL FILL_1__9211_ (
);

FILL FILL_2__16401_ (
);

FILL FILL_3__9977_ (
);

FILL FILL_3__9557_ (
);

FILL FILL_4__10922_ (
);

FILL FILL_3__9137_ (
);

FILL FILL_4__10502_ (
);

FILL FILL_1__15814_ (
);

DFFSR _8281_ (
    .Q(\datapath_1.regfile_1.regOut[11] [3]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_653_[3])
);

FILL SFILL59240x11050 (
);

FILL FILL_4__13394_ (
);

FILL FILL_0__14807_ (
);

FILL FILL_2__7974_ (
);

FILL FILL_2__7554_ (
);

BUFX2 BUFX2_insert430 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf7 )
);

BUFX2 BUFX2_insert431 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf6 )
);

FILL FILL_3__12387_ (
);

BUFX2 BUFX2_insert432 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf5 )
);

BUFX2 BUFX2_insert433 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf4 )
);

BUFX2 BUFX2_insert434 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf3 )
);

FILL FILL_6__13301_ (
);

BUFX2 BUFX2_insert435 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf2 )
);

BUFX2 BUFX2_insert436 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf1 )
);

BUFX2 BUFX2_insert437 (
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf0 )
);

FILL SFILL49640x68050 (
);

BUFX2 BUFX2_insert438 (
    .A(_5565_),
    .Y(_5565__bF$buf3)
);

BUFX2 BUFX2_insert439 (
    .A(_5565_),
    .Y(_5565__bF$buf2)
);

FILL FILL_5__12714_ (
);

FILL SFILL28760x27050 (
);

FILL SFILL59160x18050 (
);

FILL FILL_4__8841_ (
);

FILL FILL_4__11707_ (
);

FILL FILL_4__8001_ (
);

FILL FILL_2__12741_ (
);

FILL FILL_5__15186_ (
);

FILL FILL_2__12321_ (
);

INVX1 _9486_ (
    .A(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_1318_)
);

DFFSR _9066_ (
    .Q(\datapath_1.regfile_1.regOut[17] [20]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_1043_[20])
);

FILL FILL_4__14599_ (
);

FILL FILL_1__11734_ (
);

FILL FILL_4__14179_ (
);

FILL FILL_1__11314_ (
);

FILL FILL_0__8741_ (
);

FILL FILL_2__8759_ (
);

FILL FILL_0__8321_ (
);

FILL FILL_2__8339_ (
);

FILL FILL_0__10307_ (
);

FILL FILL_4__15960_ (
);

FILL FILL_4__15540_ (
);

FILL FILL_4__15120_ (
);

INVX8 _13484_ (
    .A(_3925_),
    .Y(_3995_)
);

DFFSR _13064_ (
    .Q(_2_[17]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3620_[17])
);

FILL FILL_5__13919_ (
);

FILL FILL_3__14953_ (
);

FILL FILL_3__14533_ (
);

FILL FILL_3__14113_ (
);

FILL FILL_4_BUFX2_insert270 (
);

FILL FILL_4__9626_ (
);

FILL FILL_4_BUFX2_insert271 (
);

FILL FILL_4__9206_ (
);

FILL FILL_4_BUFX2_insert272 (
);

FILL FILL_4_BUFX2_insert273 (
);

FILL FILL_2__13946_ (
);

FILL FILL_4_BUFX2_insert274 (
);

FILL FILL_0__14980_ (
);

FILL FILL_2__13526_ (
);

FILL FILL_0__14560_ (
);

FILL FILL_2__13106_ (
);

FILL FILL_4_BUFX2_insert275 (
);

FILL FILL_0__14140_ (
);

FILL FILL_4_BUFX2_insert276 (
);

FILL FILL_4_BUFX2_insert277 (
);

FILL FILL_4_BUFX2_insert278 (
);

FILL FILL_4_BUFX2_insert279 (
);

FILL FILL_1__12519_ (
);

FILL FILL_0__9526_ (
);

FILL FILL_3__7623_ (
);

FILL FILL_3__7203_ (
);

FILL FILL_0__9106_ (
);

FILL SFILL33960x45050 (
);

FILL FILL_5__7969_ (
);

FILL FILL_5__7549_ (
);

FILL FILL_4__16325_ (
);

FILL FILL_4__11880_ (
);

AOI22X1 _14689_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [25]),
    .C(\datapath_1.regfile_1.regOut[18] [25]),
    .D(_4135_),
    .Y(_5176_)
);

INVX1 _14269_ (
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_4764_)
);

FILL FILL_4__11460_ (
);

FILL FILL_4__11040_ (
);

FILL FILL_3__15738_ (
);

FILL FILL_3__15318_ (
);

FILL FILL_1__16352_ (
);

FILL FILL_5__8910_ (
);

FILL FILL_3__10873_ (
);

FILL FILL_3__10453_ (
);

FILL FILL_3__10033_ (
);

FILL FILL_0__15765_ (
);

FILL FILL_0__15345_ (
);

NOR3X1 _15630_ (
    .A(_5515__bF$buf3),
    .B(_4656_),
    .C(_5521__bF$buf3),
    .Y(_6096_)
);

AOI22X1 _15210_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [4]),
    .C(\datapath_1.regfile_1.regOut[22] [4]),
    .D(_5650_),
    .Y(_5686_)
);

FILL FILL_2__8092_ (
);

FILL FILL_0__10060_ (
);

FILL FILL_1__8902_ (
);

FILL FILL_3__8828_ (
);

FILL FILL_5__13672_ (
);

FILL FILL_5__13252_ (
);

NAND2X1 _7972_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_553_)
);

NAND2X1 _7552_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_334_)
);

FILL SFILL79320x48050 (
);

DFFSR _7132_ (
    .Q(\datapath_1.regfile_1.regOut[2] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_68_[6])
);

FILL FILL_4__12245_ (
);

INVX1 _10189_ (
    .A(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_1685_)
);

FILL FILL_3__11658_ (
);

FILL FILL_3__11238_ (
);

FILL FILL_1__12272_ (
);

NAND2X1 _16415_ (
    .A(gnd),
    .B(gnd),
    .Y(_6831_)
);

OAI21X1 _11970_ (
    .A(_3020_),
    .B(IorD_bF$buf1),
    .C(_3021_),
    .Y(_1_[27])
);

FILL FILL_0__11685_ (
);

FILL FILL_2__9297_ (
);

FILL FILL_0__11265_ (
);

AOI21X1 _11550_ (
    .A(_2567_),
    .B(_2408_),
    .C(_2427_),
    .Y(_2659_)
);

OAI21X1 _11130_ (
    .A(_2239_),
    .B(_2241_),
    .C(_2248_),
    .Y(_2249_)
);

FILL FILL_6__15884_ (
);

FILL FILL_3_BUFX2_insert290 (
);

FILL FILL_3_BUFX2_insert291 (
);

FILL FILL_3_BUFX2_insert292 (
);

FILL FILL_5__14877_ (
);

FILL FILL_5__14457_ (
);

FILL FILL_3_BUFX2_insert293 (
);

FILL FILL_3_BUFX2_insert294 (
);

FILL FILL_5__14037_ (
);

FILL FILL_3__15491_ (
);

FILL FILL_3_BUFX2_insert295 (
);

INVX1 _8757_ (
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_954_)
);

FILL FILL_3__15071_ (
);

FILL FILL_3_BUFX2_insert296 (
);

INVX1 _8337_ (
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_735_)
);

FILL FILL_3_BUFX2_insert297 (
);

FILL FILL_1__7294_ (
);

FILL FILL_3_BUFX2_insert298 (
);

FILL FILL_3_BUFX2_insert299 (
);

FILL FILL_2__14484_ (
);

FILL SFILL114440x73050 (
);

FILL FILL_2__14064_ (
);

FILL FILL_1__13897_ (
);

FILL FILL_1__13477_ (
);

FILL FILL_4__14811_ (
);

FILL FILL_3__8581_ (
);

INVX1 _12755_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_3529_)
);

NAND3X1 _12335_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3290_)
);

FILL FILL_3__13804_ (
);

FILL FILL_5__8087_ (
);

FILL FILL_6__11384_ (
);

FILL FILL_0__13831_ (
);

FILL FILL_0__13411_ (
);

FILL FILL_3__16276_ (
);

FILL FILL_5__10797_ (
);

FILL FILL_5__10377_ (
);

FILL FILL_1__8499_ (
);

FILL FILL_1__8079_ (
);

FILL FILL_2__15689_ (
);

FILL FILL_2__15269_ (
);

FILL FILL_1__9860_ (
);

FILL FILL_1__9020_ (
);

FILL FILL_2__16210_ (
);

FILL FILL_3__9786_ (
);

FILL FILL_3__9366_ (
);

FILL FILL_4__10311_ (
);

FILL FILL_1__15623_ (
);

INVX1 _8090_ (
    .A(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_611_)
);

FILL FILL_1__15203_ (
);

FILL FILL_0__14616_ (
);

OAI21X1 _14901_ (
    .A(_5381_),
    .B(_3931__bF$buf1),
    .C(_5382_),
    .Y(_5383_)
);

FILL FILL_2__7363_ (
);

FILL FILL_3__12196_ (
);

FILL FILL_6__13950_ (
);

FILL FILL_6__13110_ (
);

FILL FILL_4__7289_ (
);

FILL FILL_2__11189_ (
);

FILL FILL_5__12523_ (
);

FILL FILL_5__12103_ (
);

FILL FILL_4__8650_ (
);

FILL FILL_4__8230_ (
);

FILL FILL_4__11936_ (
);

FILL FILL_4__11516_ (
);

FILL FILL_2__12970_ (
);

FILL FILL_2__12130_ (
);

FILL FILL_0__7189_ (
);

OAI21X1 _9295_ (
    .A(_1230_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .C(_1231_),
    .Y(_1173_[29])
);

FILL FILL_1__16408_ (
);

FILL FILL_3__10929_ (
);

FILL FILL_3__10509_ (
);

FILL FILL_1__11963_ (
);

FILL FILL_1__11543_ (
);

FILL FILL_1__11123_ (
);

FILL FILL_0__8970_ (
);

FILL FILL_2__8988_ (
);

FILL SFILL104360x78050 (
);

FILL FILL_0__10956_ (
);

FILL FILL_2__8568_ (
);

FILL FILL_0__10536_ (
);

FILL FILL_2__8148_ (
);

NAND2X1 _10821_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_2005_)
);

FILL FILL_0__8130_ (
);

FILL FILL_0__10116_ (
);

NAND2X1 _10401_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1786_)
);

FILL FILL_5__6993_ (
);

NOR2X1 _13293_ (
    .A(_3781_),
    .B(_3830_),
    .Y(\datapath_1.regfile_1.regEn [6])
);

FILL FILL_5__13728_ (
);

FILL FILL_5__13308_ (
);

FILL FILL_3__14762_ (
);

FILL FILL_3__14342_ (
);

INVX1 _7608_ (
    .A(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_371_)
);

FILL FILL_1__6985_ (
);

FILL FILL_4__9855_ (
);

FILL FILL_4__9015_ (
);

FILL FILL_2__13755_ (
);

FILL FILL_2__13335_ (
);

FILL FILL_1__12748_ (
);

FILL FILL_1__12328_ (
);

FILL FILL_0__9755_ (
);

FILL FILL_3__7852_ (
);

FILL FILL_3__7432_ (
);

FILL FILL_0__9335_ (
);

OAI21X1 _11606_ (
    .A(_2692_),
    .B(_2344__bF$buf2),
    .C(_2711_),
    .Y(_2712_)
);

FILL SFILL104360x33050 (
);

FILL FILL_5__7358_ (
);

FILL FILL_4__16134_ (
);

NAND2X1 _14498_ (
    .A(_4988_),
    .B(_4981_),
    .Y(_4989_)
);

INVX1 _14078_ (
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_4577_)
);

FILL FILL_3__15967_ (
);

FILL FILL_3__15547_ (
);

FILL FILL_3__15127_ (
);

FILL FILL_1__16161_ (
);

FILL FILL_3__10682_ (
);

FILL FILL_3__10262_ (
);

FILL SFILL108680x41050 (
);

FILL SFILL64120x3050 (
);

FILL FILL_0__15994_ (
);

FILL SFILL63800x6050 (
);

FILL FILL_0__15574_ (
);

FILL FILL_0__15154_ (
);

FILL FILL_1__8711_ (
);

FILL FILL_2__15901_ (
);

FILL FILL_3__8637_ (
);

FILL FILL_3__8217_ (
);

FILL FILL_5__13481_ (
);

DFFSR _7781_ (
    .Q(\datapath_1.regfile_1.regOut[7] [15]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_393_[15])
);

INVX1 _7361_ (
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_247_)
);

FILL FILL_4__12894_ (
);

FILL FILL_4__12474_ (
);

FILL FILL_4__12054_ (
);

FILL FILL_3__11887_ (
);

FILL FILL_5__9924_ (
);

FILL FILL_5__9504_ (
);

FILL FILL_3__11467_ (
);

FILL FILL_3__11047_ (
);

FILL FILL_1__12081_ (
);

FILL SFILL114440x9050 (
);

FILL FILL_0__16359_ (
);

INVX1 _16224_ (
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_6675_)
);

FILL FILL_0__11494_ (
);

FILL SFILL89400x38050 (
);

FILL FILL_0__11074_ (
);

FILL FILL_1__9916_ (
);

FILL FILL_4__7501_ (
);

FILL FILL_2__11821_ (
);

FILL FILL_5__14686_ (
);

FILL FILL_5__14266_ (
);

FILL FILL_2__11401_ (
);

INVX1 _8986_ (
    .A(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_1066_)
);

INVX1 _8566_ (
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_911_)
);

OAI21X1 _8146_ (
    .A(_647_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_648_),
    .Y(_588_[30])
);

FILL FILL_1__10814_ (
);

FILL FILL_4__13679_ (
);

FILL FILL_4__13259_ (
);

FILL FILL_2__14293_ (
);

FILL FILL_0__7821_ (
);

FILL FILL_2__7839_ (
);

FILL FILL_2__7419_ (
);

FILL FILL_1__13286_ (
);

FILL FILL_4__14620_ (
);

FILL FILL_4__14200_ (
);

FILL FILL_0__12699_ (
);

FILL FILL_3__8390_ (
);

INVX1 _12984_ (
    .A(_2_[11]),
    .Y(_3641_)
);

DFFSR _12564_ (
    .Q(ALUOut[29]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[29])
);

FILL FILL_0__12279_ (
);

OAI21X1 _12144_ (
    .A(_3148_),
    .B(ALUSrcA_bF$buf0),
    .C(_3149_),
    .Y(\datapath_1.alu_1.ALUInA [9])
);

FILL FILL_3__13613_ (
);

FILL FILL_6__16058_ (
);

FILL FILL_4__8706_ (
);

FILL SFILL94280x44050 (
);

FILL FILL_2__12606_ (
);

FILL FILL_0__13640_ (
);

FILL FILL_0__13220_ (
);

FILL FILL_3__16085_ (
);

FILL FILL_5__10186_ (
);

FILL FILL_2__15498_ (
);

FILL FILL_2__15078_ (
);

FILL FILL_5__16412_ (
);

FILL FILL_0__8606_ (
);

FILL FILL_4__15825_ (
);

FILL FILL_4__15405_ (
);

FILL FILL_3__9595_ (
);

FILL FILL_4__10960_ (
);

NOR3X1 _13769_ (
    .A(_4271_),
    .B(_4274_),
    .C(_4269_),
    .Y(_4275_)
);

INVX1 _13349_ (
    .A(_3862_),
    .Y(_3868_)
);

FILL FILL_4__10540_ (
);

FILL FILL_4__10120_ (
);

FILL FILL_3__14818_ (
);

FILL FILL_1__15852_ (
);

FILL FILL_1__15432_ (
);

FILL FILL_1__15012_ (
);

FILL SFILL115160x34050 (
);

FILL FILL_0__14845_ (
);

INVX1 _14710_ (
    .A(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_5196_)
);

FILL FILL_0__14425_ (
);

FILL FILL_0__14005_ (
);

FILL FILL_2__7592_ (
);

BUFX2 BUFX2_insert810 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf6 )
);

BUFX2 BUFX2_insert811 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf5 )
);

FILL FILL_2__7172_ (
);

BUFX2 BUFX2_insert812 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf4 )
);

BUFX2 BUFX2_insert813 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf3 )
);

BUFX2 BUFX2_insert814 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf2 )
);

BUFX2 BUFX2_insert815 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf1 )
);

BUFX2 BUFX2_insert816 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf0 )
);

FILL FILL_4__7098_ (
);

BUFX2 BUFX2_insert817 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf4 )
);

BUFX2 BUFX2_insert818 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf3 )
);

BUFX2 BUFX2_insert819 (
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf2 )
);

FILL FILL_5__12752_ (
);

FILL FILL_5__12332_ (
);

FILL SFILL33800x5050 (
);

FILL SFILL8680x61050 (
);

FILL FILL_4__11745_ (
);

FILL SFILL74280x5050 (
);

FILL FILL_4__11325_ (
);

FILL FILL_1__16217_ (
);

FILL FILL_3__10318_ (
);

FILL FILL_1__11772_ (
);

FILL FILL_1__11352_ (
);

OAI22X1 _15915_ (
    .A(_6373_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf3),
    .D(_4945_),
    .Y(_6374_)
);

FILL FILL_0__10765_ (
);

FILL FILL_2__8377_ (
);

NAND2X1 _10630_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1898_)
);

DFFSR _10210_ (
    .Q(\datapath_1.regfile_1.regOut[26] [12]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_1628_[12])
);

FILL FILL_6__14544_ (
);

FILL FILL_6__14124_ (
);

FILL FILL_5__13957_ (
);

FILL FILL_3__14991_ (
);

FILL FILL_5__13537_ (
);

FILL FILL_3__14571_ (
);

FILL FILL_5__13117_ (
);

FILL FILL_3__14151_ (
);

INVX1 _7837_ (
    .A(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_483_)
);

INVX1 _7417_ (
    .A(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_264_)
);

FILL FILL_4_BUFX2_insert650 (
);

FILL FILL_4__9664_ (
);

FILL FILL_4_BUFX2_insert651 (
);

FILL FILL_4_BUFX2_insert652 (
);

FILL FILL_4__9244_ (
);

FILL FILL_4_BUFX2_insert653 (
);

FILL FILL_2__13984_ (
);

FILL SFILL114440x68050 (
);

FILL FILL_4_BUFX2_insert654 (
);

FILL FILL_2__13564_ (
);

FILL FILL_2__13144_ (
);

FILL FILL_4_BUFX2_insert655 (
);

FILL FILL_4_BUFX2_insert656 (
);

FILL FILL_4_BUFX2_insert657 (
);

FILL FILL_4_BUFX2_insert658 (
);

FILL FILL_4_BUFX2_insert659 (
);

FILL FILL_1__12977_ (
);

FILL FILL_1__12137_ (
);

FILL SFILL84200x40050 (
);

FILL FILL_0__9984_ (
);

FILL FILL_0__9144_ (
);

AOI21X1 _11835_ (
    .A(_2920_),
    .B(_2542_),
    .C(_2458_),
    .Y(_2924_)
);

FILL FILL_3__7241_ (
);

OAI21X1 _11415_ (
    .A(_2451_),
    .B(_2486_),
    .C(_2462__bF$buf2),
    .Y(_2532_)
);

FILL FILL_5__7587_ (
);

FILL FILL_5__7167_ (
);

FILL FILL_4__16363_ (
);

FILL FILL_6__10884_ (
);

FILL SFILL13640x60050 (
);

FILL FILL_0__12911_ (
);

FILL FILL_3__15776_ (
);

FILL FILL_3__15356_ (
);

FILL FILL_1__16390_ (
);

FILL SFILL109480x40050 (
);

FILL FILL_1__7999_ (
);

FILL FILL_1__7579_ (
);

FILL FILL_1__7159_ (
);

FILL FILL_3__10491_ (
);

FILL FILL_2__14769_ (
);

FILL FILL_2__14349_ (
);

FILL FILL_0__15383_ (
);

FILL SFILL114440x23050 (
);

FILL FILL_1__8520_ (
);

FILL FILL_1__8100_ (
);

FILL FILL_2__15710_ (
);

FILL FILL_3__8866_ (
);

FILL FILL_3__8446_ (
);

FILL FILL_5__13290_ (
);

FILL SFILL74280x40050 (
);

INVX1 _7590_ (
    .A(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_359_)
);

FILL FILL_1__14703_ (
);

FILL FILL_4_BUFX2_insert1030 (
);

INVX1 _7170_ (
    .A(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_140_)
);

FILL FILL_4_BUFX2_insert1031 (
);

FILL FILL_4_BUFX2_insert1032 (
);

FILL FILL_4_BUFX2_insert1033 (
);

FILL FILL_4_BUFX2_insert1034 (
);

FILL FILL_4_BUFX2_insert1035 (
);

FILL FILL_4__12283_ (
);

FILL FILL_4_BUFX2_insert1036 (
);

FILL FILL_4_BUFX2_insert1037 (
);

FILL FILL_4_BUFX2_insert1038 (
);

FILL FILL_4_BUFX2_insert1039 (
);

FILL FILL_2__6863_ (
);

FILL FILL_5__9733_ (
);

FILL FILL_3__11696_ (
);

FILL FILL_3__11276_ (
);

FILL SFILL74600x52050 (
);

FILL FILL_0__16168_ (
);

NAND2X1 _16033_ (
    .A(_6488_),
    .B(_6483_),
    .Y(_6489_)
);

FILL FILL_2__10689_ (
);

FILL FILL_2__10269_ (
);

FILL FILL_1__9725_ (
);

FILL FILL_5__11603_ (
);

FILL FILL_3_BUFX2_insert670 (
);

FILL FILL_4__7730_ (
);

FILL FILL_4__7310_ (
);

FILL FILL_3_BUFX2_insert671 (
);

FILL FILL_3_BUFX2_insert672 (
);

FILL FILL_5__14495_ (
);

FILL FILL_3_BUFX2_insert673 (
);

FILL FILL_2__11630_ (
);

FILL FILL_5__14075_ (
);

FILL FILL_3_BUFX2_insert674 (
);

FILL FILL_2__11210_ (
);

FILL FILL_1__15908_ (
);

FILL FILL_3_BUFX2_insert675 (
);

DFFSR _8795_ (
    .Q(\datapath_1.regfile_1.regOut[15] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_913_[5])
);

OAI21X1 _8375_ (
    .A(_759_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_760_),
    .Y(_718_[21])
);

FILL FILL_3_BUFX2_insert676 (
);

FILL FILL_3_BUFX2_insert677 (
);

FILL FILL_3_BUFX2_insert678 (
);

FILL FILL_3_BUFX2_insert679 (
);

FILL FILL_1__10623_ (
);

FILL FILL_4__13488_ (
);

FILL FILL_0__7630_ (
);

FILL FILL_2__7228_ (
);

FILL FILL_0__7210_ (
);

FILL FILL_1__13095_ (
);

DFFSR _12793_ (
    .Q(\aluControl_1.inst [2]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3490_[2])
);

FILL SFILL43720x54050 (
);

FILL FILL_0__12088_ (
);

INVX1 _12373_ (
    .A(ALUOut[10]),
    .Y(_3314_)
);

FILL FILL_3__13842_ (
);

FILL FILL_3__13422_ (
);

FILL FILL_3__13002_ (
);

FILL FILL_4__8515_ (
);

FILL FILL_2__12835_ (
);

FILL FILL_2__12415_ (
);

FILL SFILL64200x81050 (
);

FILL FILL_1__11828_ (
);

FILL FILL_1__11408_ (
);

FILL FILL_5__16221_ (
);

FILL FILL_0__8835_ (
);

FILL FILL_3__6932_ (
);

FILL FILL_6__9802_ (
);

FILL SFILL104360x28050 (
);

FILL FILL_5__6858_ (
);

FILL FILL_4__15634_ (
);

FILL FILL_4__15214_ (
);

NOR2X1 _13998_ (
    .A(_4498_),
    .B(_4488_),
    .Y(_4499_)
);

NOR2X1 _13578_ (
    .A(_4084_),
    .B(_4087_),
    .Y(_4088_)
);

NAND2X1 _13158_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [26]),
    .Y(_3737_)
);

FILL FILL_3__14627_ (
);

FILL FILL_1__15661_ (
);

FILL FILL_3__14207_ (
);

FILL FILL_1__15241_ (
);

FILL FILL112040x65050 (
);

FILL FILL_0__14654_ (
);

FILL FILL_0__14234_ (
);

FILL FILL_3__7717_ (
);

FILL FILL_5__12981_ (
);

FILL FILL_5__12141_ (
);

FILL FILL112440x34050 (
);

BUFX2 _6861_ (
    .A(_1_[23]),
    .Y(memoryAddress[23])
);

FILL FILL_4__11974_ (
);

FILL FILL_4__11554_ (
);

FILL FILL_4__11134_ (
);

FILL FILL_1__16026_ (
);

FILL FILL_3__10967_ (
);

FILL FILL_3__10547_ (
);

FILL FILL_3__10127_ (
);

FILL FILL_1__11581_ (
);

FILL FILL_1__11161_ (
);

FILL FILL_0__15859_ (
);

FILL FILL112040x20050 (
);

OAI22X1 _15724_ (
    .A(_6186_),
    .B(_5545__bF$buf0),
    .C(_5530__bF$buf2),
    .D(_6187_),
    .Y(_6188_)
);

FILL FILL_0__15439_ (
);

AOI22X1 _15304_ (
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_5778_)
);

FILL FILL_0__15019_ (
);

FILL FILL_0__10994_ (
);

FILL FILL_0__10574_ (
);

FILL FILL_2__8186_ (
);

FILL FILL_0__10154_ (
);

FILL FILL_2__10901_ (
);

FILL FILL_5__13766_ (
);

FILL FILL_5__13346_ (
);

FILL FILL_3__14380_ (
);

DFFSR _7646_ (
    .Q(\datapath_1.regfile_1.regOut[6] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_328_[8])
);

OAI21X1 _7226_ (
    .A(_176_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_177_),
    .Y(_133_[22])
);

FILL FILL_4__9893_ (
);

FILL FILL_4__9473_ (
);

FILL FILL_4__12759_ (
);

FILL FILL_2__13793_ (
);

FILL FILL_4__12339_ (
);

FILL FILL_2__13373_ (
);

FILL FILL_0__6901_ (
);

FILL FILL_2__6919_ (
);

FILL FILL_1__12786_ (
);

FILL FILL_1__12366_ (
);

FILL FILL_4__13700_ (
);

FILL FILL_3__7890_ (
);

FILL FILL_0__9793_ (
);

FILL FILL_3__7470_ (
);

FILL FILL_0__11779_ (
);

FILL FILL_0__9373_ (
);

FILL FILL_3__7050_ (
);

FILL FILL_0__11359_ (
);

OAI21X1 _11644_ (
    .A(_2161_),
    .B(_2745_),
    .C(_2746_),
    .Y(_2747_)
);

NOR2X1 _11224_ (
    .A(gnd),
    .B(ALUControl[2]),
    .Y(_2343_)
);

FILL FILL_4__16172_ (
);

FILL SFILL94280x39050 (
);

FILL FILL_0__12720_ (
);

FILL FILL_3__15585_ (
);

FILL FILL_0__12300_ (
);

FILL FILL_3__15165_ (
);

FILL FILL_2__14998_ (
);

FILL FILL_2__14578_ (
);

FILL FILL_2__14158_ (
);

FILL FILL_0__15192_ (
);

FILL FILL_5__15912_ (
);

FILL SFILL13560x5050 (
);

FILL FILL_4__14905_ (
);

FILL FILL_3__8255_ (
);

OAI21X1 _12849_ (
    .A(_3570_),
    .B(vdd),
    .C(_3571_),
    .Y(_3555_[8])
);

OAI21X1 _12429_ (
    .A(_3350_),
    .B(MemToReg_bF$buf5),
    .C(_3351_),
    .Y(\datapath_1.mux_wd3.dout [28])
);

AOI22X1 _12009_ (
    .A(\datapath_1.ALUResult [5]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3053_)
);

FILL FILL_1__14932_ (
);

FILL FILL_1__14512_ (
);

FILL SFILL94200x37050 (
);

FILL FILL_4__12092_ (
);

FILL FILL_0__13925_ (
);

FILL FILL_0__13505_ (
);

FILL SFILL4360x48050 (
);

FILL FILL_5__9542_ (
);

FILL FILL_5__9122_ (
);

FILL FILL_3__11085_ (
);

FILL FILL_0__16397_ (
);

AOI21X1 _16262_ (
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .B(_5649_),
    .C(_6711_),
    .Y(_6712_)
);

FILL SFILL79000x17050 (
);

FILL FILL_2__10498_ (
);

FILL FILL_5__11832_ (
);

FILL FILL_1__9534_ (
);

FILL FILL_5__11412_ (
);

FILL FILL_1__9114_ (
);

FILL SFILL8680x56050 (
);

FILL FILL_2__16304_ (
);

FILL FILL_4__10825_ (
);

FILL SFILL109560x73050 (
);

FILL FILL_4__10405_ (
);

FILL FILL_6__7885_ (
);

FILL FILL_1__15717_ (
);

OAI21X1 _8184_ (
    .A(_716_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_717_),
    .Y(_653_[0])
);

FILL FILL_4__13297_ (
);

FILL FILL_1__10432_ (
);

FILL FILL_1__10012_ (
);

FILL SFILL84280x37050 (
);

FILL FILL_2__7877_ (
);

FILL FILL_2__7457_ (
);

FILL FILL_2__7037_ (
);

NAND2X1 _12182_ (
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [22]),
    .Y(_3175_)
);

FILL FILL_5__12617_ (
);

FILL FILL_3__13651_ (
);

FILL SFILL8600x54050 (
);

FILL FILL_3__13231_ (
);

INVX1 _6917_ (
    .A(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_12_)
);

FILL FILL_4__8744_ (
);

FILL FILL_4__8324_ (
);

FILL FILL_2__12644_ (
);

FILL FILL_2__12224_ (
);

FILL FILL_5__15089_ (
);

NAND2X1 _9389_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1274_)
);

FILL FILL_1__11637_ (
);

FILL FILL_1__11217_ (
);

FILL FILL_6_BUFX2_insert50 (
);

FILL SFILL23560x19050 (
);

FILL FILL_5__16450_ (
);

FILL FILL_5__16030_ (
);

FILL FILL_0__8644_ (
);

NOR2X1 _10915_ (
    .A(_2058_),
    .B(_2051_),
    .Y(PCSource[1])
);

FILL FILL_0__8224_ (
);

FILL FILL_6_BUFX2_insert55 (
);

FILL FILL_4__15863_ (
);

FILL FILL_4__15443_ (
);

FILL FILL_4__15023_ (
);

FILL SFILL13640x55050 (
);

NAND2X1 _13387_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3899_)
);

FILL FILL_3__14856_ (
);

FILL FILL_2__9603_ (
);

FILL FILL_1__15890_ (
);

FILL FILL_3__14436_ (
);

FILL FILL_3__14016_ (
);

FILL FILL_1__15470_ (
);

FILL FILL_1__15050_ (
);

FILL FILL_4__9529_ (
);

FILL FILL_4__9109_ (
);

FILL FILL_2__13849_ (
);

FILL FILL_2__13429_ (
);

FILL FILL_0__14883_ (
);

FILL FILL_0__14463_ (
);

FILL FILL_2__13009_ (
);

FILL FILL_0__14043_ (
);

FILL SFILL13240x41050 (
);

FILL FILL_1__7600_ (
);

FILL FILL_3__7946_ (
);

FILL FILL_0__9849_ (
);

FILL FILL_0__9429_ (
);

FILL FILL_0__9009_ (
);

FILL FILL_3__7106_ (
);

FILL FILL_5__12790_ (
);

FILL FILL_5__12370_ (
);

FILL SFILL74280x35050 (
);

FILL FILL_4__16228_ (
);

FILL FILL_4__11783_ (
);

FILL FILL_4__11363_ (
);

FILL SFILL34520x51050 (
);

FILL FILL_1__16255_ (
);

FILL FILL_3__10776_ (
);

FILL FILL_1__11390_ (
);

FILL FILL_0__15668_ (
);

OAI22X1 _15953_ (
    .A(_5485__bF$buf1),
    .B(_6410_),
    .C(_5483__bF$buf2),
    .D(_4998_),
    .Y(_6411_)
);

FILL FILL_0__15248_ (
);

NOR2X1 _15533_ (
    .A(_5999_),
    .B(_6001_),
    .Y(_6002_)
);

NAND2X1 _15113_ (
    .A(_5588_),
    .B(_5591_),
    .Y(_5592_)
);

FILL FILL_0__10383_ (
);

FILL FILL_5__13995_ (
);

FILL SFILL43800x42050 (
);

FILL FILL_5__13575_ (
);

FILL SFILL74200x33050 (
);

FILL FILL_5__13155_ (
);

OAI21X1 _7875_ (
    .A(_507_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .C(_508_),
    .Y(_458_[25])
);

OAI21X1 _7455_ (
    .A(_288_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .C(_289_),
    .Y(_263_[13])
);

OAI21X1 _7035_ (
    .A(_69_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .C(_70_),
    .Y(_68_[1])
);

FILL FILL_4__12988_ (
);

FILL FILL_4__9282_ (
);

FILL FILL_4__12568_ (
);

FILL FILL_4__12148_ (
);

FILL FILL_1__12595_ (
);

FILL FILL_1__12175_ (
);

NAND2X1 _16318_ (
    .A(_6766_),
    .B(_6761_),
    .Y(_6767_)
);

NAND2X1 _11873_ (
    .A(\datapath_1.PCJump [13]),
    .B(RegDst),
    .Y(_2959_)
);

FILL FILL_0__11588_ (
);

FILL FILL_0__11168_ (
);

AOI21X1 _11453_ (
    .A(_2407_),
    .B(_2565_),
    .C(_2568_),
    .Y(_2569_)
);

NOR2X1 _11033_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(_2151_),
    .Y(_2152_)
);

FILL FILL_6__15787_ (
);

FILL FILL_6__15367_ (
);

FILL FILL_3__12502_ (
);

FILL SFILL104440x16050 (
);

FILL FILL_2__11915_ (
);

FILL SFILL64200x76050 (
);

FILL FILL_3__15394_ (
);

FILL FILL112120x53050 (
);

FILL FILL_1__7197_ (
);

FILL FILL_1__10908_ (
);

FILL FILL_2__14387_ (
);

FILL FILL_5__15721_ (
);

FILL FILL_5__15301_ (
);

OAI21X1 _9601_ (
    .A(_1373_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1374_),
    .Y(_1368_[3])
);

FILL FILL_4__14714_ (
);

FILL FILL_3__8484_ (
);

NAND2X1 _12658_ (
    .A(vdd),
    .B(memoryOutData[30]),
    .Y(_3485_)
);

FILL FILL_3__8064_ (
);

NAND3X1 _12238_ (
    .A(_3215_),
    .B(_3216_),
    .C(_3217_),
    .Y(\datapath_1.alu_1.ALUInB [5])
);

FILL FILL_3__13707_ (
);

FILL FILL_1__14741_ (
);

FILL FILL_1__14321_ (
);

FILL FILL_6__11287_ (
);

FILL FILL_0__13734_ (
);

FILL FILL_0__13314_ (
);

FILL FILL_3__16179_ (
);

FILL FILL_5__9771_ (
);

FILL SFILL33800x40050 (
);

FILL FILL_5__9351_ (
);

FILL SFILL64200x31050 (
);

INVX1 _16071_ (
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_6526_)
);

FILL FILL_1__9763_ (
);

FILL FILL_5__11641_ (
);

FILL FILL112440x29050 (
);

FILL FILL_1__9343_ (
);

FILL FILL_5__11221_ (
);

FILL FILL_4__15919_ (
);

FILL FILL_2__16113_ (
);

FILL FILL_3__9269_ (
);

FILL FILL_4__10634_ (
);

FILL FILL_6__7694_ (
);

FILL FILL_1__15946_ (
);

FILL FILL_1__15526_ (
);

FILL SFILL33720x47050 (
);

FILL FILL_1__15106_ (
);

FILL FILL_1__10661_ (
);

FILL FILL_1__10241_ (
);

FILL FILL_0__14939_ (
);

INVX1 _14804_ (
    .A(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_5288_)
);

FILL FILL_0__14519_ (
);

FILL FILL_2__7686_ (
);

FILL FILL_3__12099_ (
);

FILL FILL_6__13853_ (
);

FILL FILL_5__12846_ (
);

FILL FILL_3__13880_ (
);

FILL FILL_5__12426_ (
);

FILL FILL_3__13460_ (
);

FILL FILL_5__12006_ (
);

FILL FILL_3__13040_ (
);

FILL FILL_4__8973_ (
);

FILL FILL_4__8133_ (
);

FILL FILL_4__11839_ (
);

FILL FILL_2__12873_ (
);

FILL FILL_4__11419_ (
);

FILL FILL_2__12453_ (
);

FILL FILL_2__12033_ (
);

DFFSR _9198_ (
    .Q(\datapath_1.regfile_1.regOut[18] [24]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_1108_[24])
);

FILL FILL_1__11866_ (
);

FILL FILL_1__11446_ (
);

FILL FILL_1__11026_ (
);

FILL FILL_3__6970_ (
);

FILL FILL_0__8873_ (
);

FILL FILL_0__8453_ (
);

FILL FILL_6__9420_ (
);

DFFSR _10724_ (
    .Q(\datapath_1.regfile_1.regOut[30] [14]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1888_[14])
);

FILL FILL_0__10439_ (
);

OAI21X1 _10304_ (
    .A(_1740_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1741_),
    .Y(_1693_[24])
);

FILL FILL_0__10019_ (
);

FILL FILL_5__6896_ (
);

FILL FILL_4__15672_ (
);

FILL FILL_4__15252_ (
);

DFFSR _13196_ (
    .Q(\datapath_1.mux_iord.din0 [21]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3685_[21])
);

FILL FILL_2__9412_ (
);

FILL FILL_0__11800_ (
);

FILL FILL_3__14665_ (
);

FILL FILL_3__14245_ (
);

FILL FILL_1__6888_ (
);

FILL FILL_4__9758_ (
);

FILL FILL_4__9338_ (
);

FILL FILL_2__13658_ (
);

FILL FILL_2__13238_ (
);

FILL FILL_0__14692_ (
);

FILL FILL_0__14272_ (
);

FILL SFILL23720x45050 (
);

FILL FILL_3__7755_ (
);

FILL FILL_0__9658_ (
);

FILL FILL_3__7335_ (
);

INVX1 _11929_ (
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_2994_)
);

FILL FILL_0__9238_ (
);

AOI22X1 _11509_ (
    .A(_2300_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf0),
    .D(_2301_),
    .Y(_2621_)
);

FILL FILL_4__16037_ (
);

FILL FILL_6__10558_ (
);

FILL FILL_4__11592_ (
);

FILL FILL_4__11172_ (
);

FILL SFILL109640x61050 (
);

FILL FILL_1__16064_ (
);

FILL FILL_5__8622_ (
);

FILL FILL_3__10165_ (
);

FILL FILL_5__8202_ (
);

FILL FILL_6_BUFX2_insert561 (
);

FILL FILL_0__15897_ (
);

NOR2X1 _15762_ (
    .A(_6223_),
    .B(_6224_),
    .Y(_6225_)
);

FILL FILL_0__15477_ (
);

NOR2X1 _15342_ (
    .A(_4306_),
    .B(_5535__bF$buf4),
    .Y(_5815_)
);

FILL FILL_0__15057_ (
);

FILL SFILL48520x80050 (
);

FILL FILL_6_BUFX2_insert567 (
);

FILL FILL_0__10192_ (
);

FILL FILL_5__10912_ (
);

FILL FILL_1__8614_ (
);

FILL FILL_2__15804_ (
);

FILL FILL_5__13384_ (
);

FILL FILL_6__6965_ (
);

OAI21X1 _7684_ (
    .A(_400_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_401_),
    .Y(_393_[4])
);

DFFSR _7264_ (
    .Q(\datapath_1.regfile_1.regOut[3] [10]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_133_[10])
);

FILL FILL_4__9091_ (
);

FILL FILL_4__12377_ (
);

FILL FILL_3__9901_ (
);

FILL FILL_2__6957_ (
);

FILL FILL_5__9407_ (
);

OAI22X1 _16127_ (
    .A(_5480__bF$buf2),
    .B(_5254_),
    .C(_5523_),
    .D(_5265_),
    .Y(_6580_)
);

OAI21X1 _11682_ (
    .A(_2398_),
    .B(_2347__bF$buf3),
    .C(_2782_),
    .Y(_2783_)
);

FILL FILL_0__11397_ (
);

NAND2X1 _11262_ (
    .A(_2171_),
    .B(_2172_),
    .Y(_2381_)
);

FILL SFILL8600x49050 (
);

FILL FILL_3__12731_ (
);

FILL FILL_3__12311_ (
);

FILL FILL_4__7824_ (
);

FILL FILL_5__14589_ (
);

FILL FILL_2__11724_ (
);

FILL FILL_5__14169_ (
);

FILL FILL_2__11304_ (
);

NAND2X1 _8889_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1022_)
);

NAND2X1 _8469_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_803_)
);

FILL SFILL109560x23050 (
);

DFFSR _8049_ (
    .Q(\datapath_1.regfile_1.regOut[9] [27]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_523_[27])
);

FILL SFILL53800x39050 (
);

FILL FILL_2__14196_ (
);

FILL FILL_5__15950_ (
);

FILL FILL_5__15530_ (
);

FILL FILL_0__7724_ (
);

FILL FILL_5__15110_ (
);

DFFSR _9830_ (
    .Q(\datapath_1.regfile_1.regOut[23] [16]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1433_[16])
);

FILL FILL_0__7304_ (
);

NAND2X1 _9410_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1288_)
);

FILL FILL_6__13909_ (
);

FILL FILL_4__14943_ (
);

FILL FILL_4__14523_ (
);

FILL FILL_4__14103_ (
);

NAND2X1 _12887_ (
    .A(vdd),
    .B(\datapath_1.rd1 [21]),
    .Y(_3597_)
);

NAND2X1 _12467_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [9]),
    .Y(_3378_)
);

NAND3X1 _12047_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[15]),
    .C(_3032__bF$buf4),
    .Y(_3081_)
);

FILL FILL_3__13936_ (
);

FILL FILL_1__14970_ (
);

FILL FILL_3__13516_ (
);

FILL FILL_1__14550_ (
);

FILL FILL_1__14130_ (
);

FILL FILL_4__8609_ (
);

FILL FILL_5_BUFX2_insert580 (
);

FILL FILL_5_BUFX2_insert581 (
);

FILL FILL_5_BUFX2_insert582 (
);

FILL FILL_2__12509_ (
);

FILL FILL_0__13963_ (
);

FILL FILL_5_BUFX2_insert583 (
);

FILL FILL_0__13543_ (
);

FILL FILL_5_BUFX2_insert584 (
);

FILL FILL_0__13123_ (
);

FILL FILL_5_BUFX2_insert585 (
);

FILL FILL_5_BUFX2_insert586 (
);

FILL FILL_5_BUFX2_insert587 (
);

FILL FILL_5_BUFX2_insert588 (
);

FILL FILL_5__9160_ (
);

FILL FILL_5_BUFX2_insert589 (
);

FILL FILL_5__16315_ (
);

FILL FILL_0__8509_ (
);

FILL FILL_1__9992_ (
);

FILL FILL_5__11870_ (
);

FILL FILL_5__11450_ (
);

FILL FILL_1__9152_ (
);

FILL FILL_5__11030_ (
);

FILL FILL_4__15728_ (
);

FILL FILL_4__15308_ (
);

FILL FILL_2__16342_ (
);

FILL FILL_3__9498_ (
);

FILL FILL_3__9078_ (
);

FILL FILL_4__10443_ (
);

FILL FILL_4__10023_ (
);

FILL SFILL99480x79050 (
);

FILL FILL_1__15755_ (
);

FILL FILL_1__15335_ (
);

FILL FILL_1__10890_ (
);

FILL FILL_1__10050_ (
);

FILL FILL_0__14748_ (
);

INVX1 _14613_ (
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_5101_)
);

FILL FILL_0__14328_ (
);

FILL FILL_2__7495_ (
);

FILL FILL_2__7075_ (
);

FILL SFILL74200x28050 (
);

FILL FILL_5__12655_ (
);

FILL FILL_5__12235_ (
);

OAI21X1 _6955_ (
    .A(_36_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .C(_37_),
    .Y(_3_[17])
);

FILL SFILL38440x40050 (
);

FILL FILL_4__8782_ (
);

FILL FILL_4__8362_ (
);

FILL FILL_4__11648_ (
);

FILL FILL_4__11228_ (
);

FILL FILL_2__12262_ (
);

FILL FILL112200x41050 (
);

FILL FILL_1__11675_ (
);

FILL SFILL99480x34050 (
);

FILL FILL_1__11255_ (
);

AOI22X1 _15818_ (
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .B(_5577_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_6279_)
);

INVX1 _10953_ (
    .A(_2085_),
    .Y(_2086_)
);

FILL FILL_0__8262_ (
);

FILL FILL_0__10668_ (
);

FILL SFILL3480x53050 (
);

FILL FILL_0__10248_ (
);

OAI21X1 _10533_ (
    .A(_1852_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .C(_1853_),
    .Y(_1823_[15])
);

OAI21X1 _10113_ (
    .A(_1633_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .C(_1634_),
    .Y(_1628_[3])
);

FILL SFILL68600x72050 (
);

FILL FILL_6__14447_ (
);

FILL FILL_6__14027_ (
);

FILL FILL_4__15481_ (
);

FILL FILL_4__15061_ (
);

FILL FILL_2__9641_ (
);

FILL FILL_3__14894_ (
);

FILL FILL_3__14474_ (
);

FILL FILL_2__9221_ (
);

FILL FILL_3__14054_ (
);

FILL FILL112120x48050 (
);

FILL FILL_4__9987_ (
);

FILL FILL_4__9147_ (
);

FILL FILL_2__13887_ (
);

FILL FILL_2__13467_ (
);

FILL FILL_0__14081_ (
);

FILL FILL_5__14801_ (
);

FILL FILL_6_CLKBUF1_insert162 (
);

FILL SFILL89800x9050 (
);

FILL FILL_3__7984_ (
);

FILL FILL_0__9887_ (
);

FILL FILL_3__7564_ (
);

FILL FILL_0__9467_ (
);

OAI21X1 _11738_ (
    .A(_2168_),
    .B(_2198_),
    .C(_2462__bF$buf3),
    .Y(_2835_)
);

AOI21X1 _11318_ (
    .A(_2408_),
    .B(_2422_),
    .C(_2436_),
    .Y(_2437_)
);

FILL FILL_6_CLKBUF1_insert168 (
);

FILL FILL_1__13821_ (
);

FILL SFILL28840x52050 (
);

FILL FILL_1__13401_ (
);

FILL FILL_4__16266_ (
);

FILL FILL_6__10367_ (
);

FILL FILL_3__15679_ (
);

FILL FILL_3__15259_ (
);

FILL FILL_1__16293_ (
);

FILL SFILL33800x35050 (
);

FILL FILL_5__8851_ (
);

FILL SFILL64200x26050 (
);

FILL FILL_3__10394_ (
);

FILL FILL_5__8011_ (
);

OAI21X1 _15991_ (
    .A(_6446_),
    .B(_5535__bF$buf4),
    .C(_6447_),
    .Y(_6448_)
);

NAND2X1 _15571_ (
    .A(_6038_),
    .B(_6032_),
    .Y(_6039_)
);

FILL FILL_0__15286_ (
);

NAND3X1 _15151_ (
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf3),
    .Y(_5629_)
);

FILL FILL_3__16200_ (
);

FILL FILL_1__8843_ (
);

FILL FILL_5__10301_ (
);

FILL FILL_1__8003_ (
);

FILL FILL_2__15613_ (
);

FILL FILL_3__8769_ (
);

FILL FILL_3__8349_ (
);

FILL FILL_1__14606_ (
);

NAND2X1 _7493_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_315_)
);

NAND2X1 _7073_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_96_)
);

FILL FILL_4__12186_ (
);

FILL FILL_5__9636_ (
);

FILL FILL_3__11599_ (
);

FILL FILL_5__9216_ (
);

FILL FILL_3__11179_ (
);

OAI21X1 _16356_ (
    .A(_6790_),
    .B(gnd),
    .C(_6791_),
    .Y(_6769_[11])
);

AOI21X1 _11491_ (
    .A(_2602_),
    .B(_2603_),
    .C(_2300_),
    .Y(_2604_)
);

FILL FILL_5__11926_ (
);

INVX2 _11071_ (
    .A(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2190_)
);

FILL FILL_3__12960_ (
);

FILL FILL_1__9628_ (
);

FILL FILL_5__11506_ (
);

FILL FILL_1__9208_ (
);

FILL FILL_3__12120_ (
);

FILL FILL_4__7633_ (
);

FILL FILL_4__10919_ (
);

FILL FILL_4__7213_ (
);

FILL FILL_2__11953_ (
);

FILL FILL_5__14398_ (
);

FILL FILL_2__11533_ (
);

FILL FILL_2__11113_ (
);

NAND2X1 _8698_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_915_)
);

FILL FILL_3_CLKBUF1_insert111 (
);

FILL FILL_3_CLKBUF1_insert112 (
);

DFFSR _8278_ (
    .Q(\datapath_1.regfile_1.regOut[11] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_653_[0])
);

FILL FILL_3_CLKBUF1_insert113 (
);

FILL FILL_3_CLKBUF1_insert114 (
);

FILL FILL_1__10946_ (
);

FILL FILL_3_CLKBUF1_insert115 (
);

FILL FILL_3_CLKBUF1_insert116 (
);

FILL FILL_1__10526_ (
);

FILL FILL_3_CLKBUF1_insert117 (
);

FILL FILL_1__10106_ (
);

FILL SFILL18840x50050 (
);

FILL FILL_3_CLKBUF1_insert118 (
);

FILL FILL_3_CLKBUF1_insert119 (
);

FILL FILL_0__7953_ (
);

FILL FILL_0__7113_ (
);

FILL FILL_6__8500_ (
);

FILL FILL_4__14752_ (
);

FILL FILL_4__14332_ (
);

NAND2X1 _12696_ (
    .A(memoryOutData[0]),
    .B(IRWrite_bF$buf2),
    .Y(_3554_)
);

NAND3X1 _12276_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3198__bF$buf2),
    .Y(_3246_)
);

FILL FILL_2__8912_ (
);

FILL FILL_3__13745_ (
);

FILL FILL_3__13325_ (
);

FILL FILL_4__8838_ (
);

FILL FILL_2__12738_ (
);

FILL FILL_0__13772_ (
);

FILL FILL_2__12318_ (
);

FILL FILL_0__13352_ (
);

FILL FILL_0__8738_ (
);

FILL FILL_5__16124_ (
);

FILL FILL_0__8318_ (
);

FILL FILL_1__9381_ (
);

FILL FILL_4__15957_ (
);

FILL FILL_4__15537_ (
);

FILL FILL_4__15117_ (
);

FILL FILL_2__16151_ (
);

FILL FILL_4__10672_ (
);

FILL FILL_4__10252_ (
);

FILL SFILL23320x26050 (
);

FILL FILL_1__15984_ (
);

FILL FILL_1__15564_ (
);

FILL FILL_1__15144_ (
);

FILL FILL_5__7702_ (
);

FILL FILL_0__14977_ (
);

INVX1 _14842_ (
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_5325_)
);

FILL FILL_0__14557_ (
);

FILL FILL_0__14137_ (
);

NAND3X1 _14422_ (
    .A(_4905_),
    .B(_4906_),
    .C(_4913_),
    .Y(_4914_)
);

INVX1 _14002_ (
    .A(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_4503_)
);

FILL FILL_5__12884_ (
);

FILL FILL_5__12464_ (
);

FILL FILL_5__12044_ (
);

FILL FILL_4__8591_ (
);

FILL FILL_4__11877_ (
);

FILL FILL_4__11457_ (
);

FILL SFILL48920x44050 (
);

FILL FILL_2__12491_ (
);

FILL FILL_4__11037_ (
);

FILL FILL_2__12071_ (
);

FILL FILL_6__8097_ (
);

FILL FILL_1__16349_ (
);

FILL FILL_5__8907_ (
);

FILL FILL_1__11484_ (
);

FILL FILL_1__11064_ (
);

NOR3X1 _15627_ (
    .A(_6088_),
    .B(_6090_),
    .C(_6092_),
    .Y(_6093_)
);

NOR3X1 _15207_ (
    .A(_5673_),
    .B(_5664_),
    .C(_5683_),
    .Y(_5684_)
);

FILL FILL_0__10897_ (
);

FILL FILL_0__8491_ (
);

OAI21X1 _10762_ (
    .A(_1964_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1965_),
    .Y(_1953_[6])
);

FILL FILL_2__8089_ (
);

FILL FILL_0__8071_ (
);

DFFSR _10342_ (
    .Q(\datapath_1.regfile_1.regOut[27] [16]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_1693_[16])
);

FILL FILL_0__10057_ (
);

FILL FILL_3__11811_ (
);

FILL FILL_4__15290_ (
);

FILL FILL_4__6904_ (
);

FILL SFILL13720x38050 (
);

FILL SFILL44120x29050 (
);

FILL FILL_2__9870_ (
);

FILL FILL_5__13669_ (
);

FILL FILL_2__10804_ (
);

FILL FILL_5__13249_ (
);

NAND2X1 _7969_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_551_)
);

FILL FILL_2__9030_ (
);

FILL FILL_3__14283_ (
);

FILL SFILL109560x18050 (
);

NAND2X1 _7549_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_332_)
);

DFFSR _7129_ (
    .Q(\datapath_1.regfile_1.regOut[2] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_68_[3])
);

FILL FILL_4__9796_ (
);

FILL FILL_4__9376_ (
);

FILL SFILL109400x7050 (
);

FILL FILL_2__13696_ (
);

FILL FILL_2__13276_ (
);

FILL FILL_5__14610_ (
);

NAND2X1 _8910_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1036_)
);

FILL FILL_1__12269_ (
);

FILL FILL_4__13603_ (
);

FILL FILL_3__7373_ (
);

FILL FILL_0__9276_ (
);

OAI21X1 _11967_ (
    .A(_3018_),
    .B(IorD_bF$buf7),
    .C(_3019_),
    .Y(_1_[26])
);

NAND3X1 _11547_ (
    .A(_2410_),
    .B(_2552_),
    .C(_2648_),
    .Y(_2657_)
);

FILL FILL_5_CLKBUF1_insert150 (
);

NOR2X1 _11127_ (
    .A(\datapath_1.alu_1.ALUInA [19]),
    .B(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2246_)
);

FILL FILL_5_CLKBUF1_insert151 (
);

FILL FILL_5_CLKBUF1_insert152 (
);

FILL FILL_1__13630_ (
);

FILL FILL_5__7299_ (
);

FILL FILL_5_CLKBUF1_insert153 (
);

FILL FILL_1__13210_ (
);

FILL FILL_4__16075_ (
);

FILL FILL_5_CLKBUF1_insert154 (
);

FILL FILL_5_CLKBUF1_insert155 (
);

FILL FILL_5_CLKBUF1_insert156 (
);

FILL FILL_5_CLKBUF1_insert157 (
);

FILL FILL_6__10176_ (
);

FILL FILL_5_CLKBUF1_insert158 (
);

FILL FILL_5_CLKBUF1_insert159 (
);

FILL FILL_0__12623_ (
);

FILL FILL_3__15488_ (
);

FILL FILL_0__12203_ (
);

FILL FILL_3__15068_ (
);

FILL FILL_6_BUFX2_insert940 (
);

FILL FILL_5__8660_ (
);

FILL FILL_5__8240_ (
);

AOI22X1 _15380_ (
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .B(_5785_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_5852_)
);

FILL FILL_6_BUFX2_insert945 (
);

FILL FILL_0__15095_ (
);

FILL FILL_5__15815_ (
);

FILL FILL_5__10950_ (
);

FILL FILL_1__8652_ (
);

FILL FILL_5__10530_ (
);

FILL FILL_1__8232_ (
);

FILL FILL_5__10110_ (
);

FILL FILL_4__14808_ (
);

FILL FILL_2__15842_ (
);

FILL FILL_3__8998_ (
);

FILL FILL_2__15422_ (
);

FILL FILL_3__8578_ (
);

FILL FILL_2__15002_ (
);

FILL FILL_1__14835_ (
);

FILL FILL_1__14415_ (
);

FILL FILL_0__13828_ (
);

FILL FILL_0__13408_ (
);

FILL SFILL38840x49050 (
);

FILL FILL_2__6995_ (
);

FILL FILL_5__9865_ (
);

FILL FILL_5__9025_ (
);

FILL SFILL99560x22050 (
);

AOI22X1 _16165_ (
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_6617_)
);

FILL SFILL3560x41050 (
);

FILL FILL_1__9857_ (
);

FILL FILL_5__11735_ (
);

FILL SFILL24200x63050 (
);

FILL FILL_5__11315_ (
);

FILL FILL_1__9017_ (
);

FILL FILL_4__7862_ (
);

FILL FILL_2__16207_ (
);

FILL FILL_4__7442_ (
);

FILL FILL_4__10308_ (
);

FILL FILL_2__11762_ (
);

FILL FILL_2__11342_ (
);

FILL FILL_6__7368_ (
);

INVX1 _8087_ (
    .A(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_609_)
);

FILL FILL112200x36050 (
);

FILL SFILL99480x29050 (
);

FILL FILL_1__10755_ (
);

FILL FILL_0__7762_ (
);

FILL FILL_0__7342_ (
);

FILL FILL_4__14981_ (
);

FILL FILL_4__14561_ (
);

FILL FILL_4__14141_ (
);

AOI22X1 _12085_ (
    .A(\datapath_1.ALUResult [24]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3110_)
);

FILL FILL_3__13974_ (
);

FILL FILL_2__8721_ (
);

FILL FILL_3__13554_ (
);

FILL FILL_3__13134_ (
);

FILL SFILL28920x40050 (
);

FILL FILL_4__8647_ (
);

FILL FILL_4__8227_ (
);

FILL FILL_5_BUFX2_insert960 (
);

FILL FILL_5_BUFX2_insert961 (
);

FILL FILL_2__12967_ (
);

FILL FILL_5_BUFX2_insert962 (
);

FILL FILL_5_BUFX2_insert963 (
);

FILL FILL_2__12127_ (
);

FILL FILL_0__13581_ (
);

FILL FILL_5_BUFX2_insert964 (
);

FILL FILL_0__13161_ (
);

FILL FILL_5_BUFX2_insert965 (
);

FILL FILL_5_BUFX2_insert966 (
);

FILL FILL_5_BUFX2_insert967 (
);

FILL FILL_5_BUFX2_insert968 (
);

FILL FILL_5_BUFX2_insert969 (
);

FILL FILL_0__8967_ (
);

FILL FILL_5__16353_ (
);

FILL FILL_0__8127_ (
);

NAND2X1 _10818_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_2003_)
);

FILL SFILL28840x47050 (
);

FILL FILL_1__12901_ (
);

FILL FILL_4__15766_ (
);

FILL FILL_4__15346_ (
);

FILL FILL_2__16380_ (
);

FILL FILL_4__10061_ (
);

FILL FILL_2__9926_ (
);

FILL FILL_2__9506_ (
);

FILL FILL_3__14759_ (
);

FILL FILL_1__15793_ (
);

FILL FILL_3__14339_ (
);

FILL FILL_1__15373_ (
);

FILL FILL_5__7931_ (
);

FILL FILL_0__14786_ (
);

FILL FILL_0__14366_ (
);

INVX1 _14651_ (
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_5138_)
);

INVX1 _14231_ (
    .A(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_4727_)
);

FILL FILL_3__15700_ (
);

FILL FILL_1__7503_ (
);

FILL FILL_6__13280_ (
);

FILL SFILL89480x27050 (
);

FILL FILL_3__7849_ (
);

FILL FILL_3__7429_ (
);

FILL FILL_5__12273_ (
);

NAND2X1 _6993_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_63_)
);

FILL FILL_4__11686_ (
);

FILL FILL_4__11266_ (
);

FILL FILL_1__16158_ (
);

FILL FILL_3__10679_ (
);

FILL FILL_5__8716_ (
);

FILL FILL_3__10259_ (
);

FILL FILL_1__11293_ (
);

NAND2X1 _15856_ (
    .A(_6315_),
    .B(_6313_),
    .Y(_6316_)
);

OAI22X1 _15436_ (
    .A(_5466__bF$buf4),
    .B(_4403_),
    .C(_4395_),
    .D(_5483__bF$buf2),
    .Y(_5907_)
);

INVX8 _15016_ (
    .A(_5495__bF$buf3),
    .Y(_5496_)
);

NOR2X1 _10991_ (
    .A(_2107_),
    .B(_2109_),
    .Y(_2110_)
);

NAND2X1 _10571_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1879_)
);

FILL FILL_0__10286_ (
);

NAND2X1 _10151_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1660_)
);

FILL FILL_3_BUFX2_insert1040 (
);

FILL FILL_1__8708_ (
);

FILL FILL_3_BUFX2_insert1041 (
);

FILL FILL_3_BUFX2_insert1042 (
);

FILL FILL_3__11620_ (
);

FILL FILL_3_BUFX2_insert1043 (
);

FILL FILL_3__11200_ (
);

FILL FILL_3_BUFX2_insert1044 (
);

FILL FILL_3_BUFX2_insert1045 (
);

FILL FILL_3_BUFX2_insert1046 (
);

FILL FILL_3_BUFX2_insert1047 (
);

FILL FILL_3_BUFX2_insert1048 (
);

FILL FILL_5__13898_ (
);

FILL SFILL103640x54050 (
);

FILL FILL_3_BUFX2_insert1049 (
);

FILL FILL_5__13478_ (
);

FILL SFILL18040x62050 (
);

DFFSR _7778_ (
    .Q(\datapath_1.regfile_1.regOut[7] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_393_[12])
);

FILL FILL_3__14092_ (
);

INVX1 _7358_ (
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_245_)
);

FILL SFILL18840x45050 (
);

FILL FILL_2__13085_ (
);

FILL FILL_1__12498_ (
);

FILL FILL_1__12078_ (
);

FILL FILL_4__13832_ (
);

FILL SFILL79880x39050 (
);

FILL FILL_4__13412_ (
);

FILL FILL_3__7182_ (
);

OAI21X1 _11776_ (
    .A(_2558_),
    .B(_2851_),
    .C(_2869_),
    .Y(_2870_)
);

FILL FILL_0__9085_ (
);

INVX1 _11356_ (
    .A(_2473_),
    .Y(\datapath_1.ALUResult [30])
);

FILL FILL_3__12825_ (
);

FILL FILL_3__12405_ (
);

FILL FILL_4_CLKBUF1_insert140 (
);

FILL FILL_4_CLKBUF1_insert141 (
);

FILL FILL_2__11818_ (
);

FILL FILL_4_CLKBUF1_insert142 (
);

FILL FILL_0__12852_ (
);

FILL FILL_0__12432_ (
);

FILL FILL_3__15297_ (
);

FILL FILL_4_CLKBUF1_insert143 (
);

FILL FILL_4_CLKBUF1_insert144 (
);

FILL FILL_0__12012_ (
);

FILL FILL_4_CLKBUF1_insert145 (
);

FILL FILL_4_CLKBUF1_insert146 (
);

FILL FILL_4_CLKBUF1_insert147 (
);

FILL SFILL38920x5050 (
);

FILL FILL_4_CLKBUF1_insert148 (
);

FILL FILL_4_CLKBUF1_insert149 (
);

FILL FILL_5__15624_ (
);

FILL FILL_5__15204_ (
);

FILL FILL_0__7818_ (
);

INVX1 _9924_ (
    .A(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_1549_)
);

INVX1 _9504_ (
    .A(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_1330_)
);

FILL FILL_1__8881_ (
);

FILL FILL_1__8461_ (
);

FILL FILL_4__14617_ (
);

FILL FILL_2__15651_ (
);

FILL FILL_2__15231_ (
);

FILL FILL_3__8387_ (
);

FILL FILL_1__14644_ (
);

FILL FILL_1__14224_ (
);

FILL FILL_0__13637_ (
);

INVX1 _13922_ (
    .A(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_4425_)
);

FILL FILL_0__13217_ (
);

NOR2X1 _13502_ (
    .A(_4009_),
    .B(_4012_),
    .Y(_4013_)
);

FILL SFILL69480x68050 (
);

FILL FILL_5__9674_ (
);

FILL FILL_5__9254_ (
);

FILL FILL_6__12971_ (
);

NAND2X1 _16394_ (
    .A(gnd),
    .B(gnd),
    .Y(_6817_)
);

FILL FILL_6__12131_ (
);

FILL FILL_5__16409_ (
);

FILL FILL_5__11964_ (
);

FILL FILL_5__11544_ (
);

FILL FILL_1__9666_ (
);

FILL FILL_1__9246_ (
);

FILL FILL_5__11124_ (
);

FILL SFILL69080x54050 (
);

FILL FILL_2__16016_ (
);

FILL FILL_4__7671_ (
);

FILL FILL_4__10957_ (
);

FILL FILL_4__7251_ (
);

FILL SFILL48920x39050 (
);

FILL FILL_2__11991_ (
);

FILL FILL_4__10537_ (
);

FILL FILL_2__11571_ (
);

FILL FILL_4__10117_ (
);

FILL FILL_2__11151_ (
);

FILL FILL_1__15849_ (
);

FILL FILL_1__15429_ (
);

FILL FILL_1__15009_ (
);

FILL FILL_1__10564_ (
);

FILL FILL_1__10144_ (
);

INVX1 _14707_ (
    .A(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_5193_)
);

FILL FILL_0__7991_ (
);

FILL FILL_2__7589_ (
);

BUFX2 BUFX2_insert780 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf4)
);

FILL FILL_0__7571_ (
);

FILL FILL_2__7169_ (
);

BUFX2 BUFX2_insert781 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf3)
);

BUFX2 BUFX2_insert782 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf2)
);

BUFX2 BUFX2_insert783 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf1)
);

FILL FILL_6__13756_ (
);

BUFX2 BUFX2_insert784 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf0)
);

FILL FILL_6__13336_ (
);

BUFX2 BUFX2_insert785 (
    .A(_3997_),
    .Y(_3997__bF$buf3)
);

FILL FILL_4__14790_ (
);

BUFX2 BUFX2_insert786 (
    .A(_3997_),
    .Y(_3997__bF$buf2)
);

FILL FILL_4__14370_ (
);

BUFX2 BUFX2_insert787 (
    .A(_3997_),
    .Y(_3997__bF$buf1)
);

BUFX2 BUFX2_insert788 (
    .A(_3997_),
    .Y(_3997__bF$buf0)
);

BUFX2 BUFX2_insert789 (
    .A(_5532_),
    .Y(_5532__bF$buf3)
);

FILL FILL_2__8950_ (
);

FILL FILL_5__12749_ (
);

FILL FILL_3__13783_ (
);

FILL FILL_5__12329_ (
);

FILL FILL_2__8530_ (
);

FILL FILL_3__13363_ (
);

FILL FILL_2__8110_ (
);

FILL FILL_4__8876_ (
);

FILL FILL_4__8456_ (
);

FILL FILL_2__12776_ (
);

FILL FILL_2__12356_ (
);

FILL FILL_0__13390_ (
);

FILL FILL_1__11769_ (
);

FILL FILL_1__11349_ (
);

FILL SFILL3640x74050 (
);

FILL FILL_3__6873_ (
);

FILL FILL_5__16162_ (
);

FILL FILL_0__8776_ (
);

FILL FILL_0__8356_ (
);

NAND2X1 _10627_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1896_)
);

DFFSR _10207_ (
    .Q(\datapath_1.regfile_1.regOut[26] [9]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_1628_[9])
);

FILL SFILL43880x81050 (
);

FILL FILL_4__15995_ (
);

FILL FILL_1__12710_ (
);

FILL FILL_4__15575_ (
);

FILL FILL_4__15155_ (
);

OAI21X1 _13099_ (
    .A(_3696_),
    .B(PCEn_bF$buf1),
    .C(_3697_),
    .Y(_3685_[6])
);

FILL FILL_4__10290_ (
);

FILL FILL_3__14988_ (
);

FILL FILL_2__9735_ (
);

FILL FILL_3__14568_ (
);

FILL FILL_0__11703_ (
);

FILL FILL_3__14148_ (
);

FILL FILL_1__15182_ (
);

FILL FILL_5__7740_ (
);

FILL FILL_5__7320_ (
);

FILL SFILL59080x52050 (
);

NOR2X1 _14880_ (
    .A(_5362_),
    .B(_5352_),
    .Y(_5363_)
);

FILL FILL_0__14595_ (
);

FILL FILL_0__14175_ (
);

NAND3X1 _14460_ (
    .A(_4949_),
    .B(_4950_),
    .C(_4948_),
    .Y(_4951_)
);

NOR2X1 _14040_ (
    .A(_4539_),
    .B(_3960_),
    .Y(_4540_)
);

FILL SFILL38920x37050 (
);

FILL FILL_1__7732_ (
);

FILL FILL_1__7312_ (
);

FILL FILL_2__14922_ (
);

FILL FILL_2__14502_ (
);

FILL FILL_3__7238_ (
);

FILL FILL_5__12082_ (
);

FILL FILL_1__13915_ (
);

FILL FILL_4__11495_ (
);

FILL FILL_4__11075_ (
);

FILL FILL_0__12908_ (
);

FILL FILL_1__16387_ (
);

FILL FILL_5__8525_ (
);

FILL FILL_3__10488_ (
);

FILL FILL_3__10068_ (
);

FILL FILL_5__8105_ (
);

FILL SFILL59000x50050 (
);

OAI22X1 _15665_ (
    .A(_4687_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf1),
    .D(_6129_),
    .Y(_6130_)
);

NOR3X1 _15245_ (
    .A(_5494_),
    .B(_5517_),
    .C(_5697_),
    .Y(_5721_)
);

FILL SFILL3560x36050 (
);

NAND2X1 _10380_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1772_)
);

FILL FILL_5__10815_ (
);

FILL FILL_1__8517_ (
);

FILL FILL_2__15707_ (
);

FILL FILL_4__6942_ (
);

FILL FILL_0__16321_ (
);

FILL FILL_2__10422_ (
);

FILL FILL_5__13287_ (
);

FILL SFILL9240x57050 (
);

FILL FILL_6__6868_ (
);

FILL FILL_2__10002_ (
);

INVX1 _7587_ (
    .A(\datapath_1.regfile_1.regOut[6] [15]),
    .Y(_357_)
);

INVX1 _7167_ (
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_138_)
);

FILL FILL_3__9804_ (
);

FILL FILL_0__6842_ (
);

FILL FILL_4__13641_ (
);

FILL FILL_4__13221_ (
);

INVX2 _11585_ (
    .A(_2263_),
    .Y(_2692_)
);

FILL SFILL49080x50050 (
);

OAI21X1 _11165_ (
    .A(_2275_),
    .B(_2262_),
    .C(_2283_),
    .Y(_2284_)
);

FILL FILL_2__7801_ (
);

FILL FILL_3__12634_ (
);

FILL FILL_3__12214_ (
);

FILL SFILL28920x35050 (
);

FILL FILL_4__7727_ (
);

FILL FILL_4__7307_ (
);

FILL FILL_2__11627_ (
);

FILL FILL_0__12661_ (
);

FILL FILL_2__11207_ (
);

FILL FILL_0__12241_ (
);

FILL FILL_2__14099_ (
);

FILL FILL_5__15853_ (
);

FILL FILL_5__15433_ (
);

FILL FILL_0__7627_ (
);

FILL FILL_5__15013_ (
);

FILL FILL_0__7207_ (
);

INVX1 _9733_ (
    .A(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_1442_)
);

DFFSR _9313_ (
    .Q(\datapath_1.regfile_1.regOut[19] [11]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_1173_[11])
);

FILL FILL_1__8270_ (
);

FILL FILL_4__14846_ (
);

FILL FILL_4__14426_ (
);

FILL FILL_2__15880_ (
);

FILL FILL_4__14006_ (
);

FILL FILL_2__15460_ (
);

FILL FILL_2__15040_ (
);

FILL FILL_3__8196_ (
);

FILL FILL_3__13839_ (
);

FILL FILL_1__14873_ (
);

FILL FILL_3__13419_ (
);

FILL FILL_1__14453_ (
);

FILL FILL_1__14033_ (
);

FILL FILL_0__13866_ (
);

FILL FILL_0__13446_ (
);

INVX1 _13731_ (
    .A(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_4238_)
);

INVX1 _13311_ (
    .A(_3793_),
    .Y(_3844_)
);

FILL FILL_0__13026_ (
);

FILL FILL_5__9483_ (
);

FILL FILL_5__16218_ (
);

FILL FILL_3__6929_ (
);

FILL FILL_1__9895_ (
);

FILL FILL_5__11773_ (
);

FILL FILL_1__9475_ (
);

FILL FILL_5__11353_ (
);

FILL FILL_2__16245_ (
);

FILL FILL_4__7480_ (
);

FILL SFILL63960x73050 (
);

FILL FILL_4__10766_ (
);

FILL FILL_4__7060_ (
);

FILL SFILL94360x64050 (
);

FILL FILL_2__11380_ (
);

FILL SFILL103720x42050 (
);

FILL FILL_1__15658_ (
);

FILL FILL_1__15238_ (
);

FILL FILL_1__10793_ (
);

FILL FILL_1__10373_ (
);

INVX1 _14936_ (
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_5417_)
);

INVX1 _14516_ (
    .A(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_5006_)
);

FILL SFILL98680x72050 (
);

FILL FILL_0__7380_ (
);

FILL SFILL79160x44050 (
);

FILL FILL_3__10700_ (
);

FILL FILL_5__12978_ (
);

FILL FILL_3__13592_ (
);

FILL FILL_5__12138_ (
);

BUFX2 _6858_ (
    .A(_1_[20]),
    .Y(memoryAddress[20])
);

FILL FILL_3__13172_ (
);

FILL SFILL18680x5050 (
);

FILL FILL_4__8265_ (
);

FILL FILL_2__12585_ (
);

FILL FILL_2__12165_ (
);

FILL SFILL13800x50 (
);

FILL FILL_1__11998_ (
);

FILL FILL_1__11578_ (
);

FILL FILL_1__11158_ (
);

FILL FILL_4__12912_ (
);

FILL FILL_5__16391_ (
);

FILL FILL_0__8585_ (
);

DFFSR _10856_ (
    .Q(\datapath_1.regfile_1.regOut[31] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1953_[18])
);

INVX1 _10436_ (
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_1809_)
);

INVX1 _10016_ (
    .A(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_1590_)
);

FILL FILL_3__11905_ (
);

FILL FILL_4__15384_ (
);

FILL SFILL8760x81050 (
);

FILL FILL_0__11932_ (
);

FILL FILL_3__14797_ (
);

FILL FILL_2__9544_ (
);

FILL FILL_2__9124_ (
);

FILL FILL_3__14377_ (
);

FILL FILL_0__11512_ (
);

FILL SFILL114600x81050 (
);

FILL FILL_5__14704_ (
);

FILL SFILL53960x71050 (
);

FILL SFILL84360x62050 (
);

FILL FILL_1__7961_ (
);

FILL FILL_1__7121_ (
);

FILL FILL_2__14731_ (
);

FILL FILL_3__7887_ (
);

FILL FILL_2__14311_ (
);

FILL FILL_3__7467_ (
);

FILL FILL_3__7047_ (
);

FILL FILL_1__13724_ (
);

FILL FILL_1__13304_ (
);

FILL FILL_4__16169_ (
);

FILL FILL_0__12717_ (
);

FILL FILL_1__16196_ (
);

FILL FILL_5__8754_ (
);

FILL FILL_5__8334_ (
);

FILL FILL_3__10297_ (
);

NOR2X1 _15894_ (
    .A(_4968_),
    .B(_5534__bF$buf2),
    .Y(_6353_)
);

FILL FILL_0__15189_ (
);

FILL FILL_6__11211_ (
);

NAND2X1 _15474_ (
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .B(_5570__bF$buf0),
    .Y(_5944_)
);

FILL FILL_5__15909_ (
);

NAND3X1 _15054_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5477_),
    .C(_5461_),
    .Y(_5534_)
);

FILL FILL_3__16103_ (
);

FILL FILL_5__10624_ (
);

FILL FILL_1__8746_ (
);

FILL FILL_1__8326_ (
);

FILL FILL_2__15936_ (
);

FILL FILL_2__15516_ (
);

FILL FILL_0__16130_ (
);

FILL FILL_2__10651_ (
);

FILL FILL_2__10231_ (
);

FILL FILL_5__13096_ (
);

FILL FILL_1__14929_ (
);

DFFSR _7396_ (
    .Q(\datapath_1.regfile_1.regOut[4] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_198_[14])
);

FILL FILL_1__14509_ (
);

FILL FILL_4__12089_ (
);

FILL FILL_3__9613_ (
);

FILL FILL_5__9539_ (
);

FILL SFILL114520x43050 (
);

FILL FILL_5__9119_ (
);

FILL FILL_6__12836_ (
);

FILL FILL_4__13870_ (
);

FILL FILL_4__13450_ (
);

NOR2X1 _16259_ (
    .A(_6701_),
    .B(_6708_),
    .Y(_6709_)
);

FILL FILL_4__13030_ (
);

INVX1 _11394_ (
    .A(_2203_),
    .Y(_2511_)
);

FILL FILL_5__11829_ (
);

FILL FILL_2__7610_ (
);

FILL FILL_3__12863_ (
);

FILL FILL_5__11409_ (
);

FILL FILL_3__12443_ (
);

FILL FILL_3__12023_ (
);

FILL FILL_4__7956_ (
);

FILL FILL_4__7116_ (
);

FILL FILL_2__11856_ (
);

FILL FILL_0__12890_ (
);

FILL FILL_2__11436_ (
);

FILL FILL_0__12470_ (
);

FILL FILL_2__11016_ (
);

FILL FILL_0__12050_ (
);

FILL FILL_1__10429_ (
);

FILL SFILL38200x42050 (
);

FILL FILL_1__10009_ (
);

FILL SFILL3640x69050 (
);

FILL FILL_5__15662_ (
);

FILL FILL_5__15242_ (
);

FILL FILL_0__7856_ (
);

FILL FILL_0__7436_ (
);

DFFSR _9962_ (
    .Q(\datapath_1.regfile_1.regOut[24] [20]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_1498_[20])
);

OAI21X1 _9542_ (
    .A(_1354_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1355_),
    .Y(_1303_[26])
);

OAI21X1 _9122_ (
    .A(_1135_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1136_),
    .Y(_1108_[14])
);

FILL FILL_4__14655_ (
);

FILL FILL_4__14235_ (
);

OAI21X1 _12599_ (
    .A(_3444_),
    .B(vdd),
    .C(_3445_),
    .Y(_3425_[10])
);

NAND2X1 _12179_ (
    .A(ALUSrcA_bF$buf6),
    .B(\datapath_1.a [21]),
    .Y(_3173_)
);

FILL SFILL3560x7050 (
);

FILL FILL_3__13648_ (
);

FILL FILL_3__13228_ (
);

FILL FILL_1__14682_ (
);

FILL FILL_1__14262_ (
);

FILL FILL_0_BUFX2_insert420 (
);

FILL FILL_0_BUFX2_insert421 (
);

FILL FILL_0_BUFX2_insert422 (
);

FILL SFILL59080x47050 (
);

FILL FILL112280x80050 (
);

FILL FILL_0_BUFX2_insert423 (
);

FILL FILL_0__13675_ (
);

FILL FILL_0_BUFX2_insert424 (
);

NOR2X1 _13960_ (
    .A(_4461_),
    .B(_4458_),
    .Y(_4462_)
);

FILL FILL_0__13255_ (
);

FILL FILL_0_BUFX2_insert425 (
);

NOR2X1 _13540_ (
    .A(_4049_),
    .B(_4046_),
    .Y(_4050_)
);

OAI21X1 _13120_ (
    .A(_3710_),
    .B(PCEn_bF$buf3),
    .C(_3711_),
    .Y(_3685_[13])
);

FILL FILL_0_BUFX2_insert426 (
);

FILL FILL_0_BUFX2_insert427 (
);

FILL FILL_0_BUFX2_insert428 (
);

FILL FILL_0_BUFX2_insert429 (
);

FILL FILL_5__9292_ (
);

FILL FILL_5__16027_ (
);

FILL SFILL3640x24050 (
);

FILL FILL_5__11582_ (
);

FILL FILL_1__9284_ (
);

FILL FILL_5__11162_ (
);

FILL SFILL104520x41050 (
);

FILL FILL_2__16054_ (
);

FILL SFILL43880x31050 (
);

FILL FILL_4__10995_ (
);

FILL FILL_4__10575_ (
);

FILL FILL_4__10155_ (
);

FILL FILL_1__15887_ (
);

FILL FILL_1__15467_ (
);

FILL FILL_1__15047_ (
);

FILL FILL_5__7605_ (
);

FILL SFILL59000x45050 (
);

FILL FILL_1__10182_ (
);

AOI21X1 _14745_ (
    .A(\datapath_1.regfile_1.regOut[11] [27]),
    .B(_3950__bF$buf2),
    .C(_5229_),
    .Y(_5230_)
);

INVX1 _14325_ (
    .A(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_4819_)
);

FILL SFILL104440x48050 (
);

FILL FILL_0__15821_ (
);

FILL FILL_0__15401_ (
);

FILL FILL_5__12787_ (
);

FILL FILL_5__12367_ (
);

FILL FILL_4__8494_ (
);

FILL SFILL33880x74050 (
);

FILL FILL_4__8074_ (
);

FILL FILL_2__12394_ (
);

FILL FILL_1__11387_ (
);

FILL FILL_4__12721_ (
);

FILL FILL_4__12301_ (
);

FILL FILL_0__8394_ (
);

FILL SFILL33480x60050 (
);

INVX1 _10665_ (
    .A(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_1921_)
);

INVX1 _10245_ (
    .A(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_1702_)
);

FILL FILL_6__14999_ (
);

FILL FILL_3__11714_ (
);

FILL FILL_4__15193_ (
);

FILL FILL_2__10707_ (
);

FILL FILL_2__9773_ (
);

FILL FILL_2__9353_ (
);

FILL FILL_0__11741_ (
);

FILL FILL_3__14186_ (
);

FILL FILL_0__11321_ (
);

FILL FILL_6__15940_ (
);

FILL FILL_4__9279_ (
);

FILL FILL_2__13599_ (
);

FILL SFILL28520x16050 (
);

FILL FILL_5__14933_ (
);

FILL FILL_5__14513_ (
);

DFFSR _8813_ (
    .Q(\datapath_1.regfile_1.regOut[15] [23]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_913_[23])
);

FILL FILL_1__7350_ (
);

FILL FILL_4__13926_ (
);

FILL FILL_2__14960_ (
);

FILL FILL_4__13506_ (
);

FILL FILL_2__14540_ (
);

FILL SFILL18600x52050 (
);

FILL FILL_3__7696_ (
);

FILL FILL_0__9599_ (
);

FILL FILL_2__14120_ (
);

FILL SFILL49000x43050 (
);

FILL FILL_1__13953_ (
);

FILL FILL_1__13533_ (
);

FILL FILL_4__16398_ (
);

FILL FILL_1__13113_ (
);

FILL SFILL94440x52050 (
);

DFFSR _12811_ (
    .Q(\datapath_1.PCJump [22]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3490_[20])
);

FILL FILL_0__12526_ (
);

FILL FILL_0__12106_ (
);

FILL FILL_5__8983_ (
);

FILL FILL_5__8143_ (
);

FILL FILL_6__11860_ (
);

OAI22X1 _15283_ (
    .A(_5485__bF$buf2),
    .B(_4230_),
    .C(_5483__bF$buf1),
    .D(_4206_),
    .Y(_5758_)
);

FILL FILL_5__15718_ (
);

FILL FILL_3__16332_ (
);

FILL FILL_1__8975_ (
);

FILL FILL_5__10433_ (
);

FILL FILL_1__8135_ (
);

FILL FILL_5__10013_ (
);

FILL FILL_2__15745_ (
);

FILL FILL_2__15325_ (
);

FILL FILL_4__6980_ (
);

FILL FILL_2__10880_ (
);

FILL FILL_2__10040_ (
);

FILL FILL_1__14738_ (
);

FILL FILL_1__14318_ (
);

FILL FILL_3__9422_ (
);

FILL FILL_3__9002_ (
);

FILL FILL_2__6898_ (
);

FILL FILL_0__6880_ (
);

FILL FILL_5__9768_ (
);

FILL FILL_5__9348_ (
);

NAND2X1 _16068_ (
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .B(_5570__bF$buf1),
    .Y(_6523_)
);

FILL SFILL23800x70050 (
);

FILL FILL_5__11638_ (
);

FILL FILL_5__11218_ (
);

FILL FILL_3__12252_ (
);

FILL FILL_4__7765_ (
);

FILL FILL_4__7345_ (
);

FILL FILL_2__11665_ (
);

FILL FILL_2__11245_ (
);

FILL SFILL39000x41050 (
);

FILL SFILL94360x14050 (
);

FILL FILL_1__10658_ (
);

FILL FILL_1__10238_ (
);

FILL FILL_5__15891_ (
);

FILL FILL_5__15471_ (
);

FILL FILL_5__15051_ (
);

FILL FILL_0__7245_ (
);

OAI21X1 _9771_ (
    .A(_1466_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1467_),
    .Y(_1433_[17])
);

FILL SFILL84440x50050 (
);

OAI21X1 _9351_ (
    .A(_1247_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1248_),
    .Y(_1238_[5])
);

FILL FILL_4__14884_ (
);

FILL FILL_4__14464_ (
);

FILL FILL_4__14044_ (
);

FILL FILL_3__13877_ (
);

FILL FILL_2__8624_ (
);

FILL FILL_2__8204_ (
);

FILL FILL_3__13457_ (
);

FILL FILL_1__14491_ (
);

FILL FILL_3__13037_ (
);

FILL FILL_1__14071_ (
);

FILL FILL_0__13484_ (
);

FILL SFILL114600x76050 (
);

FILL SFILL53960x66050 (
);

FILL SFILL84360x57050 (
);

FILL FILL_4__9911_ (
);

FILL FILL_2__13811_ (
);

FILL FILL_3__6967_ (
);

FILL FILL_5__16256_ (
);

FILL FILL_5__11391_ (
);

FILL FILL_1__9093_ (
);

FILL FILL_4__15669_ (
);

FILL FILL_4__15249_ (
);

FILL FILL_2__16283_ (
);

FILL FILL_4__10384_ (
);

FILL FILL_0__9811_ (
);

FILL SFILL8760x31050 (
);

FILL FILL_2__9409_ (
);

FILL FILL_1__15696_ (
);

FILL FILL_1__15276_ (
);

FILL FILL_5__7834_ (
);

FILL FILL_5__7414_ (
);

OAI22X1 _14974_ (
    .A(_3941_),
    .B(_5454_),
    .C(_3902__bF$buf2),
    .D(_5453_),
    .Y(_5455_)
);

FILL FILL_0__14689_ (
);

INVX1 _14554_ (
    .A(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_5043_)
);

FILL FILL_0__14269_ (
);

AOI22X1 _14134_ (
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .B(_4225_),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_4632_)
);

FILL FILL_3__15603_ (
);

FILL SFILL114600x31050 (
);

FILL FILL_1__7826_ (
);

FILL SFILL53960x21050 (
);

FILL SFILL84360x12050 (
);

FILL FILL_0__15630_ (
);

FILL FILL_0__15210_ (
);

FILL FILL_5__12596_ (
);

FILL FILL_5__12176_ (
);

BUFX2 _6896_ (
    .A(_2_[26]),
    .Y(memoryWriteData[26])
);

FILL FILL_4__11589_ (
);

FILL FILL_4__11169_ (
);

FILL FILL_5__8619_ (
);

FILL FILL_1__11196_ (
);

NAND3X1 _15759_ (
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf4),
    .Y(_6222_)
);

NAND2X1 _15339_ (
    .A(\datapath_1.regfile_1.regOut[20] [7]),
    .B(_5785_),
    .Y(_5812_)
);

FILL FILL_4__12530_ (
);

FILL FILL_4__12110_ (
);

NOR3X1 _10894_ (
    .A(\aluControl_1.inst [3]),
    .B(_2039_),
    .C(_2024_),
    .Y(_2040_)
);

FILL FILL_0__10189_ (
);

DFFSR _10474_ (
    .Q(\datapath_1.regfile_1.regOut[28] [20]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_1758_[20])
);

FILL FILL_5__10909_ (
);

OAI21X1 _10054_ (
    .A(_1614_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1615_),
    .Y(_1563_[26])
);

FILL FILL_3__11943_ (
);

FILL SFILL43960x64050 (
);

FILL FILL_3__11523_ (
);

FILL FILL_3__11103_ (
);

FILL FILL_0__16415_ (
);

FILL FILL_2__10936_ (
);

FILL FILL_0__11970_ (
);

FILL FILL_2__10516_ (
);

FILL FILL_2__9162_ (
);

FILL FILL_0__11550_ (
);

FILL FILL_0__11130_ (
);

FILL FILL_4__9088_ (
);

FILL FILL_5__14742_ (
);

FILL FILL_0__6936_ (
);

FILL FILL_5__14322_ (
);

OAI21X1 _8622_ (
    .A(_883_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_884_),
    .Y(_848_[18])
);

OAI21X1 _8202_ (
    .A(_664_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_665_),
    .Y(_653_[6])
);

FILL FILL_4__13735_ (
);

FILL FILL_4__13315_ (
);

FILL FILL_3__7085_ (
);

AOI21X1 _11679_ (
    .A(_2164_),
    .B(_2778_),
    .C(_2458_),
    .Y(_2780_)
);

NAND2X1 _11259_ (
    .A(_2164_),
    .B(_2165_),
    .Y(_2378_)
);

FILL FILL_3__12728_ (
);

FILL FILL_1__13762_ (
);

FILL FILL_3__12308_ (
);

FILL SFILL64840x60050 (
);

FILL FILL_1__13342_ (
);

FILL FILL112280x75050 (
);

FILL FILL_0__12755_ (
);

OAI21X1 _12620_ (
    .A(_3458_),
    .B(vdd),
    .C(_3459_),
    .Y(_3425_[17])
);

FILL FILL_0__12335_ (
);

NAND2X1 _12200_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.a [28]),
    .Y(_3187_)
);

FILL FILL_6__16114_ (
);

FILL FILL_5__8372_ (
);

FILL FILL_5__15947_ (
);

INVX4 _15092_ (
    .A(_5545__bF$buf2),
    .Y(_5571_)
);

FILL FILL_5__15527_ (
);

FILL FILL_5__15107_ (
);

FILL FILL_3__16141_ (
);

DFFSR _9827_ (
    .Q(\datapath_1.regfile_1.regOut[23] [13]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_1433_[13])
);

FILL SFILL3640x19050 (
);

NAND2X1 _9407_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1286_)
);

FILL FILL_5__10662_ (
);

FILL FILL_1__8784_ (
);

FILL FILL_5__10242_ (
);

FILL FILL_1__8364_ (
);

FILL FILL_2__15974_ (
);

FILL SFILL104520x36050 (
);

FILL FILL_2__15554_ (
);

FILL SFILL43880x26050 (
);

FILL FILL_2__15134_ (
);

FILL FILL_1__14967_ (
);

FILL FILL_1__14547_ (
);

FILL FILL_1__14127_ (
);

FILL FILL_3__9651_ (
);

FILL FILL_3__9231_ (
);

NOR2X1 _13825_ (
    .A(_4326_),
    .B(_4329_),
    .Y(_4330_)
);

AND2X2 _13405_ (
    .A(_3892_),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .Y(_3917_)
);

FILL FILL112280x30050 (
);

FILL FILL_5__9997_ (
);

FILL FILL_5__9157_ (
);

FILL FILL_6__12454_ (
);

FILL FILL_6__12034_ (
);

NOR3X1 _16297_ (
    .A(_5515__bF$buf0),
    .B(_5428_),
    .C(_5521__bF$buf2),
    .Y(_6746_)
);

FILL FILL_0__14901_ (
);

FILL FILL_5__11867_ (
);

FILL FILL_1__9989_ (
);

FILL FILL_5__11447_ (
);

FILL FILL_1__9149_ (
);

FILL FILL_3__12481_ (
);

FILL FILL_5__11027_ (
);

FILL FILL_3__12061_ (
);

FILL FILL_2__16339_ (
);

FILL FILL_4__7994_ (
);

FILL SFILL33880x69050 (
);

FILL FILL_4__7574_ (
);

FILL FILL_2__11894_ (
);

FILL FILL_2__11474_ (
);

FILL FILL_2__11054_ (
);

FILL FILL_1__10887_ (
);

FILL FILL_1__10047_ (
);

FILL FILL_4__11801_ (
);

FILL FILL_5__15280_ (
);

FILL FILL_0__7474_ (
);

FILL FILL_0__7054_ (
);

DFFSR _9580_ (
    .Q(\datapath_1.regfile_1.regOut[21] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1303_[22])
);

NAND2X1 _9160_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1162_)
);

FILL FILL_6__13659_ (
);

FILL FILL_6__13239_ (
);

FILL FILL_4__14693_ (
);

FILL FILL_4__14273_ (
);

FILL FILL_2__8853_ (
);

FILL FILL_3__13686_ (
);

FILL FILL_0__10821_ (
);

FILL FILL_2__8013_ (
);

FILL FILL_3__13266_ (
);

FILL FILL_0__10401_ (
);

FILL FILL_6__14600_ (
);

FILL FILL_0_BUFX2_insert800 (
);

FILL FILL_4__8779_ (
);

FILL FILL_4__8359_ (
);

FILL FILL_0_BUFX2_insert801 (
);

FILL FILL_0_BUFX2_insert802 (
);

FILL FILL_0_BUFX2_insert803 (
);

FILL FILL_2__12259_ (
);

FILL FILL_0_BUFX2_insert804 (
);

FILL FILL_0__13293_ (
);

FILL FILL_0_BUFX2_insert805 (
);

FILL SFILL33880x24050 (
);

FILL FILL_0_BUFX2_insert806 (
);

FILL FILL_0_BUFX2_insert807 (
);

FILL FILL_0_BUFX2_insert808 (
);

FILL FILL_0_BUFX2_insert809 (
);

FILL FILL_1__6850_ (
);

FILL FILL_4__9720_ (
);

FILL FILL_4__9300_ (
);

FILL FILL_2__13620_ (
);

FILL SFILL49000x38050 (
);

FILL FILL_5__16065_ (
);

FILL FILL_0__8259_ (
);

FILL FILL_4__15898_ (
);

FILL FILL_1__12613_ (
);

FILL FILL_4__15478_ (
);

FILL FILL_4__15058_ (
);

FILL FILL_2__16092_ (
);

FILL SFILL94440x47050 (
);

FILL FILL_4__10193_ (
);

FILL FILL_2__9638_ (
);

FILL FILL_0__9620_ (
);

FILL FILL_2__9218_ (
);

FILL FILL_0__11606_ (
);

FILL FILL_1__15085_ (
);

FILL FILL_5__7223_ (
);

FILL FILL_0__14498_ (
);

AOI22X1 _14783_ (
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .B(_4090_),
    .C(_3948_),
    .D(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_5268_)
);

INVX1 _14363_ (
    .A(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_4856_)
);

FILL FILL_0__14078_ (
);

FILL FILL_3__15832_ (
);

FILL FILL_3__15412_ (
);

FILL FILL_1__7635_ (
);

FILL FILL_1__7215_ (
);

FILL FILL_2__14825_ (
);

FILL FILL_2__14405_ (
);

FILL FILL_1__13818_ (
);

FILL FILL_4__11398_ (
);

FILL FILL_3__8502_ (
);

FILL FILL_5__8848_ (
);

FILL FILL_5__8008_ (
);

NOR2X1 _15988_ (
    .A(_6443_),
    .B(_6444_),
    .Y(_6445_)
);

NOR3X1 _15568_ (
    .A(_6034_),
    .B(_5459__bF$buf0),
    .C(_6035_),
    .Y(_6036_)
);

INVX1 _15148_ (
    .A(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_5626_)
);

OAI21X1 _10283_ (
    .A(_1726_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1727_),
    .Y(_1693_[17])
);

FILL SFILL23880x22050 (
);

FILL FILL_3__11752_ (
);

FILL FILL_3__11332_ (
);

FILL FILL_4__6845_ (
);

FILL FILL_0__16224_ (
);

FILL FILL111800x38050 (
);

FILL FILL_2__10745_ (
);

FILL FILL_2__9391_ (
);

FILL FILL_2__10325_ (
);

FILL SFILL109720x81050 (
);

FILL FILL_5__14971_ (
);

FILL FILL_5__14551_ (
);

FILL FILL_5__14131_ (
);

OAI21X1 _8851_ (
    .A(_995_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_996_),
    .Y(_978_[9])
);

DFFSR _8431_ (
    .Q(\datapath_1.regfile_1.regOut[12] [25]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_718_[25])
);

NAND2X1 _8011_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_579_)
);

FILL FILL_4__13964_ (
);

FILL FILL_4__13544_ (
);

FILL FILL_4__13124_ (
);

NAND3X1 _11488_ (
    .A(_2599_),
    .B(_2595_),
    .C(_2601_),
    .Y(\datapath_1.ALUResult [26])
);

NOR2X1 _11068_ (
    .A(_2180_),
    .B(_2186_),
    .Y(_2187_)
);

FILL SFILL23800x20050 (
);

FILL FILL_2__7704_ (
);

FILL FILL_3__12957_ (
);

FILL FILL_1__13991_ (
);

FILL FILL_3__12117_ (
);

FILL FILL_1__13571_ (
);

FILL FILL_1__13151_ (
);

FILL FILL_0__12984_ (
);

FILL FILL_0__12144_ (
);

FILL SFILL74200x1050 (
);

FILL FILL_5__15756_ (
);

FILL FILL_5__15336_ (
);

FILL FILL_3__16370_ (
);

NAND2X1 _9636_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1398_)
);

NAND2X1 _9216_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1179_)
);

FILL FILL_5__10891_ (
);

FILL FILL_1__8593_ (
);

FILL FILL_5__10051_ (
);

FILL FILL_4__14749_ (
);

FILL FILL_2__15783_ (
);

FILL FILL_4__14329_ (
);

FILL FILL_2__15363_ (
);

FILL FILL_3__8099_ (
);

FILL SFILL8760x26050 (
);

FILL FILL_2__8909_ (
);

FILL SFILL13800x63050 (
);

FILL FILL_1__14776_ (
);

FILL FILL_1__14356_ (
);

FILL FILL_5__6914_ (
);

FILL FILL_3__9880_ (
);

FILL FILL_0__13769_ (
);

FILL FILL_0__13349_ (
);

NOR2X1 _13634_ (
    .A(_4139_),
    .B(_4142_),
    .Y(_4143_)
);

FILL FILL_3__9040_ (
);

INVX1 _13214_ (
    .A(\datapath_1.a3 [3]),
    .Y(_3757_)
);

FILL FILL_5__9386_ (
);

FILL SFILL114600x26050 (
);

FILL SFILL53960x16050 (
);

FILL FILL_1__6906_ (
);

FILL FILL_0__14710_ (
);

FILL FILL_1__9798_ (
);

FILL FILL_5__11676_ (
);

FILL FILL_1__9378_ (
);

FILL FILL_5__11256_ (
);

FILL FILL_3__12290_ (
);

FILL FILL_2__16148_ (
);

FILL FILL_4__10669_ (
);

FILL FILL_4__10249_ (
);

FILL FILL_2__11283_ (
);

FILL FILL_2_BUFX2_insert330 (
);

FILL FILL_1__10696_ (
);

FILL FILL_1__10276_ (
);

FILL FILL_2_BUFX2_insert331 (
);

FILL FILL_2_BUFX2_insert332 (
);

INVX1 _14839_ (
    .A(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_5322_)
);

FILL FILL_2_BUFX2_insert333 (
);

FILL FILL_2_BUFX2_insert334 (
);

INVX1 _14419_ (
    .A(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_4911_)
);

FILL FILL_4__11610_ (
);

FILL FILL_2_BUFX2_insert335 (
);

FILL FILL_2_BUFX2_insert336 (
);

FILL FILL_2_BUFX2_insert337 (
);

FILL FILL_2_BUFX2_insert338 (
);

FILL FILL_2_BUFX2_insert339 (
);

FILL SFILL43960x59050 (
);

FILL FILL_4__14082_ (
);

FILL FILL_0__15915_ (
);

FILL FILL_2__8242_ (
);

FILL FILL_3__13495_ (
);

FILL FILL_0__10630_ (
);

FILL FILL_4__8588_ (
);

FILL FILL112360x63050 (
);

FILL FILL_2__12488_ (
);

FILL FILL_2__12068_ (
);

FILL FILL_5__13822_ (
);

FILL FILL_5__13402_ (
);

FILL FILL_2_BUFX2_insert1050 (
);

FILL FILL_2_BUFX2_insert1051 (
);

FILL FILL_2_BUFX2_insert1052 (
);

OAI21X1 _7702_ (
    .A(_412_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .C(_413_),
    .Y(_393_[10])
);

FILL FILL_2_BUFX2_insert1053 (
);

FILL FILL_2_BUFX2_insert1054 (
);

FILL FILL_2_BUFX2_insert1055 (
);

FILL FILL_2_BUFX2_insert1056 (
);

FILL FILL_2_BUFX2_insert1057 (
);

FILL SFILL64040x72050 (
);

FILL FILL_2_BUFX2_insert1058 (
);

FILL FILL_5__16294_ (
);

FILL FILL_0__8488_ (
);

FILL FILL_2_BUFX2_insert1059 (
);

FILL FILL_6__9875_ (
);

FILL FILL_0__8068_ (
);

OAI21X1 _10759_ (
    .A(_1962_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .C(_1963_),
    .Y(_1953_[5])
);

DFFSR _10339_ (
    .Q(\datapath_1.regfile_1.regOut[27] [13]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_1693_[13])
);

FILL FILL_3__11808_ (
);

FILL FILL_1__12842_ (
);

FILL FILL_1__12422_ (
);

FILL FILL_4__15287_ (
);

FILL FILL_1__12002_ (
);

FILL FILL_2__9867_ (
);

FILL FILL_0__11835_ (
);

FILL SFILL68360x80050 (
);

INVX1 _11700_ (
    .A(_2799_),
    .Y(\datapath_1.ALUResult [12])
);

FILL FILL_0__11415_ (
);

FILL FILL_2__9027_ (
);

FILL FILL_5__7872_ (
);

FILL FILL_5__7452_ (
);

FILL FILL_5__7032_ (
);

INVX1 _14592_ (
    .A(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_5081_)
);

INVX1 _14172_ (
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_4669_)
);

FILL FILL_5__14607_ (
);

FILL FILL_3__15641_ (
);

NAND2X1 _8907_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1034_)
);

FILL FILL_3__15221_ (
);

FILL FILL_1__7864_ (
);

FILL FILL_1__7444_ (
);

FILL FILL_2__14634_ (
);

FILL FILL_2__14214_ (
);

FILL FILL_1__13627_ (
);

FILL FILL_1__13207_ (
);

FILL FILL_1_BUFX2_insert350 (
);

FILL FILL_3__8731_ (
);

FILL FILL_1_BUFX2_insert351 (
);

FILL FILL_3__8311_ (
);

NAND2X1 _12905_ (
    .A(vdd),
    .B(\datapath_1.rd1 [27]),
    .Y(_3609_)
);

FILL FILL_1_BUFX2_insert352 (
);

FILL FILL_1_BUFX2_insert353 (
);

FILL FILL112280x25050 (
);

FILL FILL_1_BUFX2_insert354 (
);

FILL FILL_1__16099_ (
);

FILL FILL_1_BUFX2_insert355 (
);

FILL FILL_1_BUFX2_insert356 (
);

FILL FILL_5__8657_ (
);

FILL FILL_1_BUFX2_insert357 (
);

FILL FILL_5__8237_ (
);

FILL FILL_1_BUFX2_insert358 (
);

FILL FILL_1_BUFX2_insert359 (
);

INVX1 _15797_ (
    .A(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_6259_)
);

INVX1 _15377_ (
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_5849_)
);

FILL FILL_3__16006_ (
);

FILL FILL_5__10947_ (
);

DFFSR _10092_ (
    .Q(\datapath_1.regfile_1.regOut[25] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1563_[22])
);

FILL FILL_3__11981_ (
);

FILL FILL_1__8649_ (
);

FILL FILL_5__10527_ (
);

FILL FILL_1__8229_ (
);

FILL FILL_3__11561_ (
);

FILL FILL_5__10107_ (
);

FILL FILL_3__11141_ (
);

FILL FILL_2__15839_ (
);

FILL FILL_2__15419_ (
);

FILL FILL_0__16033_ (
);

FILL FILL_2__10974_ (
);

FILL FILL_2__10554_ (
);

FILL FILL_2__10134_ (
);

NAND2X1 _7299_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_206_)
);

FILL FILL_3__9936_ (
);

FILL FILL_3__9516_ (
);

FILL FILL_5__14780_ (
);

FILL FILL_0__6974_ (
);

FILL FILL_5__14360_ (
);

NAND2X1 _8660_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_910_)
);

NAND2X1 _8240_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_691_)
);

FILL FILL_4__13773_ (
);

FILL FILL_4__13353_ (
);

NAND2X1 _11297_ (
    .A(_2263_),
    .B(_2264_),
    .Y(_2416_)
);

FILL FILL_2__7933_ (
);

FILL FILL_3__12766_ (
);

FILL FILL_3__12346_ (
);

FILL FILL_1__13380_ (
);

FILL FILL_4__7859_ (
);

FILL FILL_4__7439_ (
);

FILL FILL_2__11759_ (
);

FILL FILL_2__11339_ (
);

FILL SFILL33880x19050 (
);

FILL FILL_0__12373_ (
);

FILL FILL_5__15985_ (
);

FILL FILL_2__12700_ (
);

FILL FILL_5__15565_ (
);

FILL FILL_0__7759_ (
);

FILL FILL_5__15145_ (
);

NAND2X1 _9865_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1510_)
);

FILL FILL_0__7339_ (
);

DFFSR _9445_ (
    .Q(\datapath_1.regfile_1.regOut[20] [15]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_1238_[15])
);

INVX1 _9025_ (
    .A(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_1092_)
);

FILL FILL_5__10280_ (
);

FILL FILL_4__14978_ (
);

FILL FILL_4__14558_ (
);

FILL FILL_4__14138_ (
);

FILL FILL_2__15592_ (
);

FILL FILL_2__15172_ (
);

FILL FILL_2__8718_ (
);

FILL FILL_0__8700_ (
);

FILL FILL_1__14585_ (
);

FILL FILL_1__14165_ (
);

FILL FILL_0__13998_ (
);

NOR2X1 _13863_ (
    .A(_4356_),
    .B(_4366_),
    .Y(_4367_)
);

FILL FILL_0__13578_ (
);

NAND3X1 _13443_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3883_),
    .C(_3888_),
    .Y(_3955_)
);

FILL FILL_0__13158_ (
);

INVX1 _13023_ (
    .A(_2_[24]),
    .Y(_3667_)
);

FILL FILL_3__14912_ (
);

FILL FILL_2__13905_ (
);

FILL FILL_5__11485_ (
);

FILL FILL_5__11065_ (
);

FILL FILL_2__16377_ (
);

FILL FILL_4__10898_ (
);

FILL FILL_4__7192_ (
);

FILL FILL_4__10058_ (
);

FILL FILL_0__9905_ (
);

FILL FILL_2__11092_ (
);

FILL FILL_5__7928_ (
);

FILL FILL_5__7508_ (
);

FILL SFILL79400x4050 (
);

INVX1 _14648_ (
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_5135_)
);

INVX1 _14228_ (
    .A(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_4724_)
);

FILL FILL_0__7092_ (
);

FILL FILL_1__16311_ (
);

FILL SFILL23880x17050 (
);

FILL FILL_3__10832_ (
);

FILL FILL_3__10412_ (
);

FILL FILL_0__15724_ (
);

FILL FILL_0__15304_ (
);

FILL FILL_2__8891_ (
);

FILL FILL_2__8471_ (
);

FILL FILL_4__8397_ (
);

FILL FILL_2__12297_ (
);

FILL SFILL8440x45050 (
);

FILL FILL_5__13631_ (
);

FILL FILL_5__13211_ (
);

OAI21X1 _7931_ (
    .A(_524_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_525_),
    .Y(_523_[1])
);

DFFSR _7511_ (
    .Q(\datapath_1.regfile_1.regOut[5] [1]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_263_[1])
);

FILL FILL_4__12624_ (
);

FILL FILL_4__12204_ (
);

FILL FILL_6__9684_ (
);

NOR2X1 _10988_ (
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2107_)
);

NAND2X1 _10568_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1877_)
);

FILL SFILL23800x15050 (
);

NAND2X1 _10148_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1658_)
);

FILL FILL_3__11617_ (
);

FILL FILL_1__12651_ (
);

FILL FILL_1__12231_ (
);

FILL FILL_4__15096_ (
);

FILL FILL_2__9676_ (
);

FILL FILL_2__9256_ (
);

FILL FILL_0__11644_ (
);

FILL FILL_0__11224_ (
);

FILL FILL_3__14089_ (
);

FILL SFILL104360x2050 (
);

FILL FILL_6__15843_ (
);

FILL FILL_5__7681_ (
);

FILL FILL_5__14836_ (
);

FILL FILL_3__15870_ (
);

FILL FILL_5__14416_ (
);

FILL FILL_3__15450_ (
);

NAND2X1 _8716_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_927_)
);

FILL FILL_3__15030_ (
);

FILL FILL_1__7673_ (
);

FILL FILL_1__7253_ (
);

FILL FILL_4__13829_ (
);

FILL FILL_2__14863_ (
);

FILL FILL_4__13409_ (
);

FILL FILL_2__14443_ (
);

FILL FILL_2__14023_ (
);

FILL FILL_3__7599_ (
);

FILL FILL_3__7179_ (
);

FILL FILL_1__13856_ (
);

FILL FILL_1__13436_ (
);

FILL FILL_1__13016_ (
);

FILL FILL_3__8960_ (
);

FILL FILL_0__12849_ (
);

NAND2X1 _12714_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[6]),
    .Y(_3502_)
);

FILL FILL_0__12429_ (
);

FILL FILL_3__8120_ (
);

FILL FILL_0__12009_ (
);

FILL FILL_5__8886_ (
);

FILL FILL_5__8466_ (
);

FILL FILL_1_BUFX2_insert20 (
);

FILL FILL_1_BUFX2_insert21 (
);

FILL FILL_6__11763_ (
);

FILL FILL_1_BUFX2_insert22 (
);

FILL FILL_1_BUFX2_insert23 (
);

INVX1 _15186_ (
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_5663_)
);

FILL FILL_1_BUFX2_insert24 (
);

FILL FILL_1_BUFX2_insert25 (
);

FILL FILL_1_BUFX2_insert26 (
);

FILL FILL_3__16235_ (
);

FILL FILL_1_BUFX2_insert27 (
);

FILL FILL_1_BUFX2_insert28 (
);

FILL FILL_1_BUFX2_insert29 (
);

FILL FILL_5__10756_ (
);

FILL FILL_1__8878_ (
);

FILL FILL_1__8458_ (
);

FILL FILL_3__11790_ (
);

FILL FILL_3__11370_ (
);

FILL FILL_2__15648_ (
);

FILL FILL_2__15228_ (
);

FILL FILL_4__6883_ (
);

FILL FILL_0__16262_ (
);

FILL FILL_2__10783_ (
);

FILL FILL_2__10363_ (
);

FILL SFILL13800x13050 (
);

FILL FILL_3__9745_ (
);

INVX1 _13919_ (
    .A(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_4422_)
);

FILL SFILL49720x9050 (
);

FILL FILL_4__13582_ (
);

FILL FILL_4__13162_ (
);

FILL FILL_2__7742_ (
);

FILL FILL_3__12995_ (
);

FILL FILL_3__12575_ (
);

FILL FILL_2__7322_ (
);

FILL FILL_3__12155_ (
);

FILL FILL_4__7248_ (
);

FILL FILL112360x58050 (
);

FILL FILL_2__11988_ (
);

FILL FILL_2__11568_ (
);

FILL FILL_2__11148_ (
);

FILL FILL_0__12182_ (
);

FILL FILL_5__12902_ (
);

FILL SFILL49000x2050 (
);

FILL SFILL64040x67050 (
);

FILL FILL_5__15794_ (
);

FILL FILL_5__15374_ (
);

FILL FILL_0__7988_ (
);

FILL FILL_0__7568_ (
);

INVX1 _9674_ (
    .A(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_1423_)
);

INVX1 _9254_ (
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_1204_)
);

FILL FILL_1__11922_ (
);

FILL FILL_4__14787_ (
);

FILL FILL_4__14367_ (
);

FILL FILL_1__11502_ (
);

FILL SFILL24360x40050 (
);

FILL FILL_2__8527_ (
);

FILL FILL_0__10915_ (
);

FILL FILL_2__8107_ (
);

FILL FILL_1__14394_ (
);

FILL FILL_5__6952_ (
);

OAI22X1 _13672_ (
    .A(_4178_),
    .B(_3944__bF$buf3),
    .C(_3959_),
    .D(_4179_),
    .Y(_4180_)
);

FILL FILL_0__13387_ (
);

NOR2X1 _13252_ (
    .A(_3794_),
    .B(_3792_),
    .Y(_3795_)
);

FILL FILL112360x13050 (
);

FILL FILL_3__14721_ (
);

FILL FILL_3__14301_ (
);

FILL FILL_1__6944_ (
);

FILL FILL_2__13714_ (
);

FILL FILL_5__16159_ (
);

FILL FILL_5__11294_ (
);

FILL FILL_1__12707_ (
);

FILL FILL_2__16186_ (
);

FILL FILL_4__10287_ (
);

FILL FILL_3__7811_ (
);

FILL SFILL89240x71050 (
);

FILL FILL_1__15599_ (
);

FILL FILL_1__15179_ (
);

FILL FILL_5__7737_ (
);

FILL FILL_2_BUFX2_insert710 (
);

FILL FILL_5__7317_ (
);

FILL FILL_2_BUFX2_insert711 (
);

FILL FILL_2_BUFX2_insert712 (
);

AOI22X1 _14877_ (
    .A(_3950__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [29]),
    .C(\datapath_1.regfile_1.regOut[31] [29]),
    .D(_3995__bF$buf1),
    .Y(_5360_)
);

FILL FILL_2_BUFX2_insert713 (
);

NOR2X1 _14457_ (
    .A(_4944_),
    .B(_4947_),
    .Y(_4948_)
);

FILL FILL_2_BUFX2_insert714 (
);

FILL FILL_2_BUFX2_insert715 (
);

AOI22X1 _14037_ (
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .B(_4005__bF$buf1),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_4537_)
);

FILL FILL_3__15926_ (
);

FILL FILL_2_BUFX2_insert716 (
);

FILL FILL_3__15506_ (
);

FILL FILL_2_BUFX2_insert717 (
);

FILL FILL_2_BUFX2_insert718 (
);

FILL FILL_2_BUFX2_insert719 (
);

FILL FILL_1__16120_ (
);

FILL FILL_1__7729_ (
);

FILL FILL_1__7309_ (
);

FILL FILL_3__10641_ (
);

FILL FILL_2__14919_ (
);

FILL FILL_0__15953_ (
);

FILL FILL_0__15533_ (
);

FILL FILL_0__15113_ (
);

FILL FILL_5__12499_ (
);

FILL SFILL54040x65050 (
);

FILL FILL_5__12079_ (
);

FILL FILL_5__13860_ (
);

FILL FILL_5__13440_ (
);

FILL FILL_5__13020_ (
);

NAND2X1 _7740_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_439_)
);

NAND2X1 _7320_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_220_)
);

FILL FILL_1__11099_ (
);

FILL FILL_6__11819_ (
);

FILL FILL_4__12853_ (
);

FILL FILL_4__12433_ (
);

FILL FILL_4__12013_ (
);

NAND2X1 _10797_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1989_)
);

FILL FILL_6__9493_ (
);

NAND2X1 _10377_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1770_)
);

FILL FILL_3__11846_ (
);

FILL FILL_1__12880_ (
);

FILL FILL_3__11426_ (
);

FILL FILL_1__12460_ (
);

FILL FILL_3__11006_ (
);

FILL FILL_1__12040_ (
);

FILL FILL_4__6939_ (
);

FILL FILL_0__16318_ (
);

FILL FILL_2__9485_ (
);

FILL FILL_0__11873_ (
);

FILL FILL_2__10419_ (
);

FILL FILL_0__11453_ (
);

FILL FILL_0__11033_ (
);

FILL FILL_5__7490_ (
);

FILL FILL_5__7070_ (
);

FILL FILL_5__14645_ (
);

FILL FILL_5__14225_ (
);

FILL FILL_0__6839_ (
);

DFFSR _8945_ (
    .Q(\datapath_1.regfile_1.regOut[16] [27]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_978_[27])
);

INVX1 _8525_ (
    .A(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_840_)
);

INVX1 _8105_ (
    .A(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_621_)
);

FILL FILL_1__7482_ (
);

FILL FILL_1__7062_ (
);

FILL FILL_4__13638_ (
);

FILL FILL_4__13218_ (
);

FILL FILL_2__14672_ (
);

FILL FILL_2__14252_ (
);

FILL FILL_1__13665_ (
);

FILL FILL_1__13245_ (
);

FILL FILL_1_BUFX2_insert730 (
);

FILL FILL_1_BUFX2_insert731 (
);

FILL SFILL59160x4050 (
);

FILL FILL_0__12658_ (
);

DFFSR _12943_ (
    .Q(\datapath_1.a [24]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3555_[24])
);

FILL FILL_1_BUFX2_insert732 (
);

INVX1 _12523_ (
    .A(ALUOut[28]),
    .Y(_3415_)
);

FILL FILL_1_BUFX2_insert733 (
);

FILL FILL_0__12238_ (
);

NAND3X1 _12103_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[29]),
    .C(_3032__bF$buf0),
    .Y(_3123_)
);

FILL FILL_1_BUFX2_insert734 (
);

FILL FILL_1_BUFX2_insert735 (
);

FILL FILL_5__8695_ (
);

FILL FILL_1_BUFX2_insert736 (
);

FILL SFILL79160x76050 (
);

FILL SFILL59080x9050 (
);

FILL FILL_6__16017_ (
);

FILL FILL_1_BUFX2_insert737 (
);

FILL FILL_5__8275_ (
);

FILL SFILL44040x63050 (
);

FILL FILL_1_BUFX2_insert738 (
);

FILL FILL_1_BUFX2_insert739 (
);

FILL FILL_3__16044_ (
);

FILL FILL_5__10565_ (
);

FILL FILL_1__8267_ (
);

FILL FILL_5__10145_ (
);

FILL FILL_2__15877_ (
);

FILL FILL_2__15457_ (
);

FILL FILL_2__15037_ (
);

FILL FILL_0__16071_ (
);

FILL FILL_2__10172_ (
);

FILL FILL_3__9974_ (
);

FILL FILL_3__9554_ (
);

FILL FILL_3__9134_ (
);

INVX1 _13728_ (
    .A(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_4235_)
);

NAND2X1 _13308_ (
    .A(_3841_),
    .B(_3839_),
    .Y(_3842_)
);

FILL FILL_1__15811_ (
);

FILL SFILL109400x50050 (
);

FILL FILL_6__12357_ (
);

FILL FILL_4__13391_ (
);

FILL FILL_0__14804_ (
);

FILL FILL_2__7971_ (
);

FILL FILL_2__7551_ (
);

BUFX2 BUFX2_insert400 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf1 )
);

BUFX2 BUFX2_insert401 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf0 )
);

FILL FILL_3__12384_ (
);

BUFX2 BUFX2_insert402 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf7)
);

FILL SFILL88840x36050 (
);

BUFX2 BUFX2_insert403 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf6)
);

BUFX2 BUFX2_insert404 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf5)
);

FILL FILL_4__7477_ (
);

BUFX2 BUFX2_insert405 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf4)
);

BUFX2 BUFX2_insert406 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf3)
);

FILL FILL_4__7057_ (
);

BUFX2 BUFX2_insert407 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf2)
);

FILL FILL_2__11797_ (
);

BUFX2 BUFX2_insert408 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf1)
);

FILL FILL_2__11377_ (
);

BUFX2 BUFX2_insert409 (
    .A(MemToReg),
    .Y(MemToReg_bF$buf0)
);

FILL FILL_5__12711_ (
);

FILL SFILL114680x70050 (
);

FILL FILL_4__11704_ (
);

FILL FILL_5__15183_ (
);

FILL FILL_6__8764_ (
);

FILL FILL_0__7377_ (
);

INVX1 _9483_ (
    .A(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_1316_)
);

DFFSR _9063_ (
    .Q(\datapath_1.regfile_1.regOut[17] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_1043_[17])
);

FILL FILL_4__14596_ (
);

FILL FILL_1__11731_ (
);

FILL FILL_4__14176_ (
);

FILL FILL_1__11311_ (
);

FILL SFILL69160x74050 (
);

FILL FILL_2__8756_ (
);

FILL FILL_2__8336_ (
);

FILL FILL_3__13589_ (
);

FILL FILL_0__10304_ (
);

FILL FILL_3__13169_ (
);

FILL FILL_6__14503_ (
);

FILL SFILL74120x57050 (
);

INVX1 _13481_ (
    .A(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_3992_)
);

DFFSR _13061_ (
    .Q(_2_[14]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3620_[14])
);

FILL FILL_5__13916_ (
);

FILL FILL_3__14950_ (
);

FILL FILL_3__14530_ (
);

FILL FILL_3__14110_ (
);

FILL FILL_4_BUFX2_insert240 (
);

FILL FILL_4__9623_ (
);

FILL FILL_4_BUFX2_insert241 (
);

FILL FILL_4_BUFX2_insert242 (
);

FILL FILL_4__12909_ (
);

FILL FILL_4_BUFX2_insert243 (
);

FILL FILL_2__13943_ (
);

FILL FILL_5__16388_ (
);

FILL FILL_4_BUFX2_insert244 (
);

FILL FILL_2__13523_ (
);

FILL FILL_4_BUFX2_insert245 (
);

FILL FILL_2__13103_ (
);

FILL FILL_6__9549_ (
);

FILL FILL_4_BUFX2_insert246 (
);

FILL FILL_4_BUFX2_insert247 (
);

FILL FILL_4_BUFX2_insert248 (
);

FILL FILL_4_BUFX2_insert249 (
);

FILL FILL_1__12516_ (
);

FILL FILL_0__11929_ (
);

FILL FILL_3__7620_ (
);

FILL FILL_0__9523_ (
);

FILL FILL_0__9103_ (
);

FILL FILL_3__7200_ (
);

FILL FILL_0__11509_ (
);

FILL FILL_5__7966_ (
);

FILL FILL_5__7546_ (
);

FILL FILL_4__16322_ (
);

OAI22X1 _14686_ (
    .A(_3982__bF$buf2),
    .B(_5171_),
    .C(_3971__bF$buf2),
    .D(_5172_),
    .Y(_5173_)
);

INVX1 _14266_ (
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_4761_)
);

FILL SFILL74120x12050 (
);

FILL FILL_3__15735_ (
);

FILL FILL_3__15315_ (
);

FILL FILL_1__7958_ (
);

FILL FILL_3__10870_ (
);

FILL FILL_1__7118_ (
);

FILL FILL_3__10450_ (
);

FILL SFILL28840x6050 (
);

FILL FILL_3__10030_ (
);

FILL FILL_2__14728_ (
);

FILL FILL_2__14308_ (
);

FILL FILL_0__15762_ (
);

FILL SFILL99320x61050 (
);

FILL FILL_0__15342_ (
);

FILL FILL_3__8825_ (
);

FILL SFILL8760x2050 (
);

FILL FILL_3__8405_ (
);

FILL SFILL8680x7050 (
);

FILL SFILL68840x77050 (
);

FILL FILL_4__12662_ (
);

FILL FILL_4__12242_ (
);

FILL SFILL64120x55050 (
);

INVX1 _10186_ (
    .A(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_1683_)
);

FILL SFILL33960x50 (
);

FILL FILL_3__11655_ (
);

FILL FILL_3__11235_ (
);

FILL FILL_0__16127_ (
);

NAND2X1 _16412_ (
    .A(gnd),
    .B(gnd),
    .Y(_6829_)
);

FILL FILL_2__10648_ (
);

FILL FILL_2__9294_ (
);

FILL FILL_0__11682_ (
);

FILL FILL_0__11262_ (
);

FILL FILL_3_BUFX2_insert260 (
);

FILL FILL_3_BUFX2_insert261 (
);

FILL FILL_5__14874_ (
);

FILL FILL_3_BUFX2_insert262 (
);

FILL FILL_5__14454_ (
);

FILL FILL_3_BUFX2_insert263 (
);

FILL FILL_5__14034_ (
);

FILL FILL_3_BUFX2_insert264 (
);

FILL FILL_3_BUFX2_insert265 (
);

INVX1 _8754_ (
    .A(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_952_)
);

INVX1 _8334_ (
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_733_)
);

FILL FILL_3_BUFX2_insert266 (
);

FILL FILL_3_BUFX2_insert267 (
);

FILL FILL_1__7291_ (
);

FILL FILL_3_BUFX2_insert268 (
);

FILL FILL_4__13867_ (
);

FILL FILL_3_BUFX2_insert269 (
);

FILL FILL_4__13447_ (
);

FILL FILL_2__14481_ (
);

FILL FILL_4__13027_ (
);

FILL FILL_2__14061_ (
);

FILL FILL_2__7607_ (
);

FILL SFILL64120x10050 (
);

FILL FILL_1__13894_ (
);

FILL FILL_1__13474_ (
);

FILL FILL_0__12887_ (
);

INVX1 _12752_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_3527_)
);

FILL FILL_0__12467_ (
);

FILL FILL_0__12047_ (
);

NAND3X1 _12332_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf0),
    .Y(_3288_)
);

FILL FILL_3__13801_ (
);

FILL FILL_5__8084_ (
);

FILL FILL_5__15659_ (
);

FILL FILL_5__15239_ (
);

DFFSR _9959_ (
    .Q(\datapath_1.regfile_1.regOut[24] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_1498_[17])
);

FILL FILL_3__16273_ (
);

OAI21X1 _9539_ (
    .A(_1352_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1353_),
    .Y(_1303_[25])
);

FILL SFILL64040x17050 (
);

FILL FILL_5__10794_ (
);

OAI21X1 _9119_ (
    .A(_1133_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1134_),
    .Y(_1108_[13])
);

FILL FILL_1__8496_ (
);

FILL FILL_5__10374_ (
);

FILL FILL_1__8076_ (
);

FILL FILL_2__15686_ (
);

FILL FILL_2__15266_ (
);

FILL SFILL14360x78050 (
);

FILL SFILL89240x66050 (
);

FILL SFILL54120x53050 (
);

FILL FILL_1__14679_ (
);

FILL FILL_1__14259_ (
);

FILL FILL_0_BUFX2_insert390 (
);

FILL FILL_0_BUFX2_insert391 (
);

FILL FILL_0_BUFX2_insert392 (
);

FILL FILL_3__9783_ (
);

FILL FILL_0_BUFX2_insert393 (
);

FILL FILL_0_BUFX2_insert394 (
);

INVX1 _13957_ (
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_4459_)
);

FILL FILL_3__9363_ (
);

FILL FILL_0_BUFX2_insert395 (
);

INVX1 _13537_ (
    .A(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_4047_)
);

FILL FILL_0_BUFX2_insert396 (
);

OAI21X1 _13117_ (
    .A(_3708_),
    .B(PCEn_bF$buf2),
    .C(_3709_),
    .Y(_3685_[12])
);

FILL FILL_0_BUFX2_insert397 (
);

FILL FILL_0_BUFX2_insert398 (
);

FILL FILL_1__15620_ (
);

FILL FILL_5__9289_ (
);

FILL FILL_0_BUFX2_insert399 (
);

FILL FILL_1__15200_ (
);

FILL FILL_0__14613_ (
);

FILL FILL_5__11999_ (
);

FILL FILL_5__11579_ (
);

FILL FILL_2__7360_ (
);

FILL FILL_5__11159_ (
);

FILL FILL_3__12193_ (
);

FILL FILL_4__7286_ (
);

FILL FILL_2__11186_ (
);

FILL FILL_5__12520_ (
);

FILL FILL_5__12100_ (
);

FILL SFILL89240x21050 (
);

FILL FILL_1__10179_ (
);

FILL FILL_4__11933_ (
);

FILL FILL_4__11513_ (
);

FILL FILL_2_BUFX2_insert70 (
);

FILL FILL_6__8573_ (
);

FILL FILL_0__7186_ (
);

FILL FILL_1__16405_ (
);

OAI21X1 _9292_ (
    .A(_1228_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .C(_1229_),
    .Y(_1173_[28])
);

FILL FILL_2_BUFX2_insert71 (
);

FILL FILL_2_BUFX2_insert72 (
);

FILL FILL_2_BUFX2_insert73 (
);

FILL FILL_3__10926_ (
);

FILL FILL_2_BUFX2_insert74 (
);

FILL FILL_1__11960_ (
);

FILL FILL_3__10506_ (
);

FILL SFILL18680x41050 (
);

FILL FILL_2_BUFX2_insert75 (
);

FILL FILL_1__11540_ (
);

FILL FILL_2_BUFX2_insert76 (
);

FILL FILL_1__11120_ (
);

FILL FILL_2_BUFX2_insert77 (
);

FILL FILL_0__15818_ (
);

FILL FILL_2_BUFX2_insert78 (
);

FILL FILL_2_BUFX2_insert79 (
);

FILL FILL_2__8985_ (
);

FILL FILL_0__10953_ (
);

FILL FILL_0__10533_ (
);

FILL FILL_3__13398_ (
);

FILL FILL_2__8145_ (
);

FILL FILL_0__10113_ (
);

FILL FILL_5__6990_ (
);

FILL SFILL54040x15050 (
);

AND2X2 _13290_ (
    .A(_3827_),
    .B(_3817_),
    .Y(_3828_)
);

FILL FILL_5__13725_ (
);

FILL FILL_5__13305_ (
);

INVX1 _7605_ (
    .A(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_369_)
);

FILL FILL_1__6982_ (
);

FILL FILL_4__9852_ (
);

FILL FILL_4__12718_ (
);

FILL FILL_4__9012_ (
);

FILL FILL_2__13752_ (
);

FILL FILL_2__13332_ (
);

FILL FILL_5__16197_ (
);

FILL FILL_1__12745_ (
);

FILL FILL_1__12325_ (
);

FILL FILL_0__9752_ (
);

FILL FILL_0__11738_ (
);

FILL FILL_0__11318_ (
);

NAND2X1 _11603_ (
    .A(_2462__bF$buf1),
    .B(_2694_),
    .Y(_2709_)
);

FILL SFILL44040x58050 (
);

FILL FILL_5__7355_ (
);

FILL FILL_4__16131_ (
);

INVX1 _14495_ (
    .A(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_4986_)
);

AOI21X1 _14075_ (
    .A(_4574_),
    .B(_4548_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [12])
);

FILL FILL_3__15964_ (
);

FILL FILL_3__15544_ (
);

FILL FILL_3__15124_ (
);

FILL FILL_1__7347_ (
);

FILL FILL_2__14957_ (
);

FILL FILL_0__15991_ (
);

FILL FILL_2__14537_ (
);

FILL FILL_0__15571_ (
);

FILL FILL_2__14117_ (
);

FILL FILL_0__15151_ (
);

FILL FILL_3__8634_ (
);

DFFSR _12808_ (
    .Q(\datapath_1.PCJump [19]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3490_[17])
);

FILL FILL_3__8214_ (
);

FILL SFILL8520x28050 (
);

FILL SFILL109400x45050 (
);

FILL FILL_4__12891_ (
);

FILL FILL_4__12471_ (
);

FILL SFILL44040x13050 (
);

FILL FILL_4__12051_ (
);

FILL FILL_3__16329_ (
);

FILL FILL_3__11884_ (
);

FILL FILL_5__9921_ (
);

FILL FILL_3__11464_ (
);

FILL FILL_5__9501_ (
);

FILL FILL_3__11044_ (
);

FILL FILL_4__6977_ (
);

FILL SFILL69240x62050 (
);

FILL FILL_0__16356_ (
);

NOR3X1 _16221_ (
    .A(_5515__bF$buf1),
    .B(_5337_),
    .C(_5521__bF$buf0),
    .Y(_6672_)
);

FILL FILL_2__10877_ (
);

FILL FILL_2__10037_ (
);

FILL FILL_0__11491_ (
);

FILL FILL_0__11071_ (
);

FILL FILL_1__9913_ (
);

FILL FILL_6__15690_ (
);

FILL FILL_6__15270_ (
);

FILL FILL_3__9419_ (
);

FILL FILL_5__14683_ (
);

FILL FILL_5__14263_ (
);

FILL FILL_0__6877_ (
);

FILL FILL_6__7844_ (
);

INVX1 _8983_ (
    .A(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_1064_)
);

DFFSR _8563_ (
    .Q(\datapath_1.regfile_1.regOut[13] [29]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_783_[29])
);

OAI21X1 _8143_ (
    .A(_645_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .C(_646_),
    .Y(_588_[29])
);

FILL FILL_1__10811_ (
);

FILL FILL_4__13676_ (
);

FILL FILL_4__13256_ (
);

FILL FILL_2__14290_ (
);

FILL FILL_2__7836_ (
);

FILL FILL_2__7416_ (
);

FILL FILL_3__12249_ (
);

FILL FILL_1__13283_ (
);

FILL FILL_0__12696_ (
);

INVX1 _12981_ (
    .A(_2_[10]),
    .Y(_3639_)
);

DFFSR _12561_ (
    .Q(ALUOut[26]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3360_[26])
);

FILL FILL_0__12276_ (
);

OAI21X1 _12141_ (
    .A(_3146_),
    .B(ALUSrcA_bF$buf7),
    .C(_3147_),
    .Y(\datapath_1.alu_1.ALUInA [8])
);

FILL FILL_3__13610_ (
);

FILL FILL_4__8703_ (
);

FILL FILL_6__11190_ (
);

FILL FILL_5__15888_ (
);

FILL FILL_2__12603_ (
);

FILL FILL_5__15468_ (
);

FILL FILL_5__15048_ (
);

OAI21X1 _9768_ (
    .A(_1464_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .C(_1465_),
    .Y(_1433_[16])
);

FILL FILL_6__8629_ (
);

FILL FILL_3__16082_ (
);

OAI21X1 _9348_ (
    .A(_1245_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1246_),
    .Y(_1238_[4])
);

FILL FILL_5__10183_ (
);

FILL FILL_2__15495_ (
);

FILL FILL_2__15075_ (
);

FILL SFILL69160x24050 (
);

FILL FILL_0__8603_ (
);

FILL FILL_1__14488_ (
);

FILL FILL_1__14068_ (
);

FILL FILL_4__15822_ (
);

FILL FILL_4__15402_ (
);

FILL FILL_3__9592_ (
);

INVX1 _13766_ (
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_4272_)
);

FILL FILL_3__9172_ (
);

INVX1 _13346_ (
    .A(_3843_),
    .Y(_3865_)
);

FILL FILL_3__14815_ (
);

FILL FILL_5__9098_ (
);

FILL FILL_4__9908_ (
);

FILL FILL_2__13808_ (
);

FILL SFILL99320x56050 (
);

FILL FILL_0__14842_ (
);

FILL FILL_0__14422_ (
);

FILL FILL_0__14002_ (
);

FILL FILL_5__11388_ (
);

FILL FILL_4__7095_ (
);

FILL SFILL28760x76050 (
);

FILL FILL_0__9808_ (
);

FILL SFILL59160x67050 (
);

FILL FILL_6__10708_ (
);

FILL FILL_4__11742_ (
);

FILL FILL_4__11322_ (
);

FILL FILL_1__16214_ (
);

FILL FILL_3__10315_ (
);

OAI22X1 _15912_ (
    .A(_5466__bF$buf3),
    .B(_4952_),
    .C(_4955_),
    .D(_5483__bF$buf4),
    .Y(_6371_)
);

FILL FILL_0__15627_ (
);

FILL FILL_0__15207_ (
);

FILL FILL_2__8374_ (
);

FILL FILL_0__10762_ (
);

FILL SFILL99320x11050 (
);

FILL FILL_5__13954_ (
);

FILL FILL_5__13534_ (
);

FILL FILL_5__13114_ (
);

FILL SFILL28760x31050 (
);

INVX1 _7834_ (
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_481_)
);

FILL SFILL59160x22050 (
);

INVX1 _7414_ (
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_326_)
);

FILL FILL_4_BUFX2_insert620 (
);

FILL FILL_4__9661_ (
);

FILL FILL_4_BUFX2_insert621 (
);

FILL FILL_4_BUFX2_insert622 (
);

FILL FILL_4__9241_ (
);

FILL FILL_4_BUFX2_insert623 (
);

FILL FILL_4__12527_ (
);

FILL FILL_2__13981_ (
);

FILL FILL_4_BUFX2_insert624 (
);

FILL FILL_4__12107_ (
);

FILL FILL_2__13561_ (
);

FILL FILL_4_BUFX2_insert625 (
);

FILL FILL_2__13141_ (
);

FILL FILL_4_BUFX2_insert626 (
);

FILL FILL_6__9167_ (
);

FILL FILL_4_BUFX2_insert627 (
);

FILL SFILL99240x18050 (
);

FILL FILL_4_BUFX2_insert628 (
);

FILL FILL_4_BUFX2_insert629 (
);

FILL FILL_1__12974_ (
);

FILL FILL_1__12134_ (
);

FILL FILL_0__9981_ (
);

FILL FILL_2__9999_ (
);

FILL FILL_0__11967_ (
);

FILL FILL_0__9141_ (
);

AOI22X1 _11832_ (
    .A(_2478_),
    .B(_2920_),
    .C(_2357_),
    .D(_2341__bF$buf2),
    .Y(_2921_)
);

FILL FILL_2__9159_ (
);

FILL FILL_0__11547_ (
);

FILL SFILL89320x54050 (
);

INVX1 _11412_ (
    .A(_2316_),
    .Y(_2529_)
);

FILL FILL_0__11127_ (
);

FILL FILL_6__15746_ (
);

FILL FILL_6__15326_ (
);

FILL FILL_5__7584_ (
);

FILL FILL_5__7164_ (
);

FILL FILL_4__16360_ (
);

FILL FILL_6__10041_ (
);

FILL FILL_5__14739_ (
);

FILL FILL_5__14319_ (
);

FILL FILL_3__15773_ (
);

FILL FILL_3__15353_ (
);

FILL SFILL18760x74050 (
);

OAI21X1 _8619_ (
    .A(_881_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .C(_882_),
    .Y(_848_[17])
);

FILL FILL_1__7996_ (
);

FILL FILL_1__7576_ (
);

FILL FILL_2__14766_ (
);

FILL FILL_2__14346_ (
);

FILL FILL_0__15380_ (
);

FILL FILL_1__13759_ (
);

FILL FILL_1__13339_ (
);

FILL FILL_3__8863_ (
);

FILL FILL_3__8443_ (
);

OAI21X1 _12617_ (
    .A(_3456_),
    .B(vdd),
    .C(_3457_),
    .Y(_3425_[16])
);

FILL FILL_5__8789_ (
);

FILL FILL_1__14700_ (
);

FILL FILL_4_BUFX2_insert1000 (
);

FILL FILL_5__8369_ (
);

FILL FILL_4_BUFX2_insert1001 (
);

FILL FILL_4_BUFX2_insert1002 (
);

FILL FILL_4_BUFX2_insert1003 (
);

FILL FILL_6__11666_ (
);

FILL FILL_4_BUFX2_insert1004 (
);

FILL FILL_6__11246_ (
);

FILL FILL_4_BUFX2_insert1005 (
);

FILL FILL_4__12280_ (
);

NAND2X1 _15089_ (
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .B(_5567_),
    .Y(_5568_)
);

FILL FILL_4_BUFX2_insert1006 (
);

FILL FILL_4_BUFX2_insert1007 (
);

FILL FILL_4_BUFX2_insert1008 (
);

FILL FILL_3__16138_ (
);

FILL FILL_4_BUFX2_insert1009 (
);

FILL FILL_5__10659_ (
);

FILL FILL_2__6860_ (
);

FILL FILL_5__10239_ (
);

FILL FILL_5__9730_ (
);

FILL FILL_3__11693_ (
);

FILL FILL_3__11273_ (
);

AOI21X1 _16450_ (
    .A(Branch),
    .B(ALUZero),
    .C(PCWrite),
    .Y(_6835_)
);

FILL FILL_0__16165_ (
);

OAI21X1 _16030_ (
    .A(_6484_),
    .B(_5535__bF$buf2),
    .C(_6485_),
    .Y(_6486_)
);

FILL FILL_2__10686_ (
);

FILL FILL_2__10266_ (
);

FILL FILL_1__9722_ (
);

FILL FILL_5__11600_ (
);

FILL FILL_3__9648_ (
);

FILL FILL_3_BUFX2_insert640 (
);

FILL FILL_3__9228_ (
);

FILL FILL_3_BUFX2_insert641 (
);

FILL FILL_3_BUFX2_insert642 (
);

FILL FILL_5__14492_ (
);

FILL FILL_3_BUFX2_insert643 (
);

FILL FILL_3_BUFX2_insert644 (
);

FILL FILL_5__14072_ (
);

FILL FILL_1__15905_ (
);

FILL FILL_3_BUFX2_insert645 (
);

DFFSR _8792_ (
    .Q(\datapath_1.regfile_1.regOut[15] [2]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_913_[2])
);

FILL FILL_3_BUFX2_insert646 (
);

OAI21X1 _8372_ (
    .A(_757_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_758_),
    .Y(_718_[20])
);

FILL FILL_3_BUFX2_insert647 (
);

FILL SFILL79320x52050 (
);

FILL FILL_3_BUFX2_insert648 (
);

FILL SFILL18680x36050 (
);

FILL FILL_3_BUFX2_insert649 (
);

FILL FILL_4__13485_ (
);

FILL FILL_1__10620_ (
);

FILL FILL_3__12898_ (
);

FILL FILL_2__7225_ (
);

FILL FILL_3__12478_ (
);

FILL FILL111960x65050 (
);

FILL FILL_3__12058_ (
);

FILL FILL_1__13092_ (
);

FILL FILL_6__13812_ (
);

OAI21X1 _12790_ (
    .A(_3551_),
    .B(IRWrite_bF$buf4),
    .C(_3552_),
    .Y(_3490_[31])
);

FILL FILL_0__12085_ (
);

INVX1 _12370_ (
    .A(ALUOut[9]),
    .Y(_3312_)
);

FILL FILL_4__8512_ (
);

FILL FILL_5__15697_ (
);

FILL FILL_2__12832_ (
);

FILL FILL_2__12412_ (
);

FILL FILL_5__15277_ (
);

OAI21X1 _9997_ (
    .A(_1576_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1577_),
    .Y(_1563_[7])
);

DFFSR _9577_ (
    .Q(\datapath_1.regfile_1.regOut[21] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1303_[19])
);

NAND2X1 _9157_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1160_)
);

FILL FILL_1__11825_ (
);

FILL FILL_1__11405_ (
);

FILL FILL_0__8832_ (
);

FILL FILL_0__10818_ (
);

FILL FILL_1__14297_ (
);

FILL FILL_5__6855_ (
);

FILL FILL_0_BUFX2_insert770 (
);

FILL FILL_4__15631_ (
);

FILL FILL_0_BUFX2_insert771 (
);

FILL FILL_4__15211_ (
);

FILL FILL_0_BUFX2_insert772 (
);

FILL FILL111960x20050 (
);

FILL FILL_0_BUFX2_insert773 (
);

FILL FILL_0_BUFX2_insert774 (
);

OAI22X1 _13995_ (
    .A(_4494_),
    .B(_3893__bF$buf1),
    .C(_3944__bF$buf3),
    .D(_4495_),
    .Y(_4496_)
);

INVX1 _13575_ (
    .A(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_4085_)
);

FILL FILL_0_BUFX2_insert775 (
);

FILL FILL_0_BUFX2_insert776 (
);

NAND2X1 _13155_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [25]),
    .Y(_3735_)
);

FILL FILL_0_BUFX2_insert777 (
);

FILL FILL_3__14624_ (
);

FILL FILL_0_BUFX2_insert778 (
);

FILL FILL_3__14204_ (
);

FILL FILL_0_BUFX2_insert779 (
);

FILL FILL_1__6847_ (
);

FILL SFILL79240x14050 (
);

FILL FILL_2__13617_ (
);

FILL FILL_0__14651_ (
);

FILL FILL_0__14231_ (
);

FILL FILL_5__11197_ (
);

FILL FILL_2__16089_ (
);

FILL FILL111880x27050 (
);

FILL FILL_3__7714_ (
);

FILL FILL_0__9617_ (
);

FILL FILL_4__16416_ (
);

FILL FILL_4__11971_ (
);

FILL FILL_6__10517_ (
);

FILL FILL_4__11551_ (
);

FILL FILL_4__11131_ (
);

FILL FILL_3__15829_ (
);

FILL FILL_3__15409_ (
);

FILL FILL_6__8191_ (
);

FILL FILL_1__16023_ (
);

FILL FILL_3__10964_ (
);

FILL FILL_3__10544_ (
);

FILL FILL_3__10124_ (
);

FILL SFILL53640x72050 (
);

FILL SFILL69240x57050 (
);

FILL FILL_0__15856_ (
);

OAI22X1 _15721_ (
    .A(_5504__bF$buf1),
    .B(_4724_),
    .C(_5527__bF$buf1),
    .D(_4715_),
    .Y(_6185_)
);

FILL FILL_0__15436_ (
);

OAI22X1 _15301_ (
    .A(_5774_),
    .B(_5544__bF$buf2),
    .C(_5569_),
    .D(_4289_),
    .Y(_5775_)
);

FILL FILL_0__15016_ (
);

FILL FILL_0__10991_ (
);

FILL FILL_0__10571_ (
);

FILL FILL_2__8183_ (
);

FILL FILL_0__10151_ (
);

FILL FILL_5__13763_ (
);

FILL FILL_5__13343_ (
);

FILL FILL_6__6924_ (
);

DFFSR _7643_ (
    .Q(\datapath_1.regfile_1.regOut[6] [5]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_328_[5])
);

OAI21X1 _7223_ (
    .A(_174_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_175_),
    .Y(_133_[21])
);

FILL FILL_4__9890_ (
);

FILL FILL_4__9470_ (
);

FILL FILL_4__12756_ (
);

FILL FILL_2__13790_ (
);

FILL FILL_4__12336_ (
);

FILL FILL_2__13370_ (
);

FILL FILL_2__6916_ (
);

FILL FILL_3__11749_ (
);

FILL FILL_1__12783_ (
);

FILL FILL_3__11329_ (
);

FILL FILL_1__12363_ (
);

FILL FILL_0__9790_ (
);

FILL FILL_0__9370_ (
);

FILL FILL_2__9388_ (
);

FILL FILL_0__11776_ (
);

FILL SFILL104360x82050 (
);

FILL SFILL69240x12050 (
);

FILL FILL_0__11356_ (
);

AOI21X1 _11641_ (
    .A(_2209_),
    .B(_2743_),
    .C(_2162_),
    .Y(_2744_)
);

NOR2X1 _11221_ (
    .A(ALUControl[1]),
    .B(ALUControl[0]),
    .Y(_2340_)
);

FILL FILL_5__14968_ (
);

FILL FILL_5__14548_ (
);

FILL FILL_5__14128_ (
);

FILL FILL_3__15582_ (
);

OAI21X1 _8848_ (
    .A(_993_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_994_),
    .Y(_978_[8])
);

FILL FILL_3__15162_ (
);

DFFSR _8428_ (
    .Q(\datapath_1.regfile_1.regOut[12] [22]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_718_[22])
);

NAND2X1 _8008_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_577_)
);

FILL FILL_2__14995_ (
);

FILL FILL_2__14575_ (
);

FILL FILL_2__14155_ (
);

FILL SFILL69160x19050 (
);

FILL FILL_1__13988_ (
);

FILL FILL_1__13568_ (
);

FILL FILL_1__13148_ (
);

FILL FILL_4__14902_ (
);

FILL FILL_3__8252_ (
);

OAI21X1 _12846_ (
    .A(_3568_),
    .B(vdd),
    .C(_3569_),
    .Y(_3555_[7])
);

OAI21X1 _12426_ (
    .A(_3348_),
    .B(MemToReg_bF$buf4),
    .C(_3349_),
    .Y(\datapath_1.mux_wd3.dout [27])
);

NAND3X1 _12006_ (
    .A(_3048_),
    .B(_3049_),
    .C(_3050_),
    .Y(\datapath_1.mux_pcsrc.dout [4])
);

FILL FILL_5__8598_ (
);

FILL FILL_0__13922_ (
);

FILL FILL_3__16367_ (
);

FILL FILL_0__13502_ (
);

FILL FILL_5__10888_ (
);

FILL FILL_5__10048_ (
);

FILL FILL_3__11082_ (
);

FILL FILL_0__16394_ (
);

FILL FILL_2__10495_ (
);

FILL FILL_1__9531_ (
);

FILL FILL_1__9111_ (
);

FILL FILL_2__16301_ (
);

FILL FILL_3__9877_ (
);

FILL FILL_3__9037_ (
);

FILL FILL_4__10822_ (
);

FILL FILL_4__10402_ (
);

FILL FILL_1__15714_ (
);

DFFSR _8181_ (
    .Q(\datapath_1.regfile_1.regOut[10] [31]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_588_[31])
);

FILL FILL_4__13294_ (
);

FILL FILL_0__14707_ (
);

FILL FILL_2__7874_ (
);

FILL FILL_2_CLKBUF1_insert1074 (
);

FILL FILL_2__7454_ (
);

FILL FILL_3__12287_ (
);

FILL FILL_2_CLKBUF1_insert1075 (
);

FILL FILL_2__7034_ (
);

FILL FILL_2_CLKBUF1_insert1076 (
);

FILL FILL_2_CLKBUF1_insert1077 (
);

FILL FILL_2_CLKBUF1_insert1078 (
);

FILL FILL_2_CLKBUF1_insert1079 (
);

FILL SFILL89400x42050 (
);

FILL FILL_5__12614_ (
);

FILL SFILL28760x26050 (
);

FILL SFILL43560x32050 (
);

INVX1 _6914_ (
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_10_)
);

FILL FILL_4__8741_ (
);

FILL FILL_4__8321_ (
);

FILL FILL_4__11607_ (
);

FILL FILL_2__12641_ (
);

FILL FILL_5__15086_ (
);

FILL FILL_2__12221_ (
);

FILL FILL_6__8247_ (
);

NAND2X1 _9386_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1272_)
);

FILL FILL_4__14499_ (
);

FILL FILL_1__11634_ (
);

FILL FILL_1__11214_ (
);

FILL FILL_4__14079_ (
);

FILL FILL_2__8659_ (
);

FILL FILL_0__8641_ (
);

FILL SFILL89320x49050 (
);

NAND2X1 _10912_ (
    .A(_2046_),
    .B(_2052_),
    .Y(_2057_)
);

FILL FILL_0__10627_ (
);

FILL FILL_2__8239_ (
);

FILL FILL_0__8221_ (
);

FILL FILL_6_BUFX2_insert24 (
);

FILL FILL_4__15860_ (
);

FILL FILL_6__14406_ (
);

FILL FILL_4__15440_ (
);

FILL FILL_6_BUFX2_insert29 (
);

FILL FILL_4__15020_ (
);

FILL FILL_0__13099_ (
);

INVX1 _13384_ (
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_3896_)
);

FILL FILL_5__13819_ (
);

FILL FILL_2__9600_ (
);

FILL FILL_3__14853_ (
);

FILL FILL_3__14433_ (
);

FILL FILL_3__14013_ (
);

FILL FILL_4__9526_ (
);

FILL FILL_4__9106_ (
);

FILL FILL_2__13846_ (
);

FILL FILL_0__14880_ (
);

FILL FILL_2__13426_ (
);

FILL FILL_0__14460_ (
);

FILL FILL_2__13006_ (
);

FILL FILL_0__14040_ (
);

FILL FILL_1__12839_ (
);

FILL FILL_1__12419_ (
);

FILL FILL_0__9846_ (
);

FILL FILL_3__7943_ (
);

FILL FILL_0__9426_ (
);

FILL FILL_3__7103_ (
);

FILL FILL_0__9006_ (
);

FILL FILL_5__7869_ (
);

FILL FILL_5__7449_ (
);

FILL FILL_4__16225_ (
);

INVX1 _14589_ (
    .A(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_5078_)
);

FILL FILL_4__11780_ (
);

NAND2X1 _14169_ (
    .A(_4659_),
    .B(_4666_),
    .Y(_4667_)
);

FILL FILL_4__11360_ (
);

FILL FILL_3__15638_ (
);

FILL FILL_3__15218_ (
);

FILL FILL_1__16252_ (
);

FILL FILL_3__10773_ (
);

FILL SFILL79400x40050 (
);

FILL SFILL18760x24050 (
);

FILL FILL_0__15665_ (
);

NAND3X1 _15950_ (
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf1),
    .Y(_6408_)
);

FILL FILL_0__15245_ (
);

OAI22X1 _15530_ (
    .A(_5534__bF$buf0),
    .B(_4503_),
    .C(_5998_),
    .D(_5549__bF$buf3),
    .Y(_5999_)
);

OAI22X1 _15110_ (
    .A(_5472__bF$buf2),
    .B(_4010_),
    .C(_3992_),
    .D(_5527__bF$buf3),
    .Y(_5589_)
);

FILL FILL_0__10380_ (
);

FILL FILL_3__8728_ (
);

FILL FILL_5__13992_ (
);

FILL FILL_5__13572_ (
);

FILL FILL_5__13152_ (
);

OAI21X1 _7872_ (
    .A(_505_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .C(_506_),
    .Y(_458_[24])
);

OAI21X1 _7452_ (
    .A(_286_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_287_),
    .Y(_263_[12])
);

FILL SFILL79320x47050 (
);

OAI21X1 _7032_ (
    .A(_131_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_132_),
    .Y(_68_[0])
);

FILL FILL_4__12985_ (
);

FILL FILL_4__12145_ (
);

DFFSR _10089_ (
    .Q(\datapath_1.regfile_1.regOut[25] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1563_[19])
);

FILL FILL_3__11978_ (
);

FILL FILL_3__11558_ (
);

FILL FILL_1__12592_ (
);

FILL FILL_3__11138_ (
);

FILL FILL_1__12172_ (
);

INVX1 _16315_ (
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_6764_)
);

NAND3X1 _11870_ (
    .A(_2473_),
    .B(_2955_),
    .C(_2956_),
    .Y(_2957_)
);

FILL FILL_0__11585_ (
);

FILL FILL_0__11165_ (
);

INVX1 _11450_ (
    .A(_2420_),
    .Y(_2566_)
);

INVX1 _11030_ (
    .A(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2149_)
);

FILL FILL_2__11912_ (
);

FILL FILL_5__14777_ (
);

FILL FILL_5__14357_ (
);

FILL FILL_3__15391_ (
);

NAND2X1 _8657_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_908_)
);

NAND2X1 _8237_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_689_)
);

FILL FILL_1__7194_ (
);

FILL FILL_1__10905_ (
);

FILL FILL_2__14384_ (
);

FILL SFILL114440x72050 (
);

FILL SFILL94440x9050 (
);

FILL FILL_1__13797_ (
);

FILL FILL_1__13377_ (
);

FILL FILL_4__14711_ (
);

FILL FILL_3__8481_ (
);

NAND2X1 _12655_ (
    .A(vdd),
    .B(memoryOutData[29]),
    .Y(_3483_)
);

FILL FILL_3__8061_ (
);

NAND3X1 _12235_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3215_)
);

FILL FILL_3__13704_ (
);

FILL FILL_0__13731_ (
);

FILL SFILL105000x4050 (
);

FILL FILL_0__13311_ (
);

FILL FILL_3__16176_ (
);

FILL FILL_5__10697_ (
);

FILL FILL_5__10277_ (
);

FILL FILL_1__8399_ (
);

FILL FILL_2__15589_ (
);

FILL FILL_2__15169_ (
);

FILL SFILL69320x45050 (
);

FILL FILL_1__9760_ (
);

FILL FILL_1__9340_ (
);

FILL FILL_4__15916_ (
);

FILL FILL_2__16110_ (
);

FILL FILL_3__9266_ (
);

FILL SFILL29160x56050 (
);

FILL FILL_4__10631_ (
);

FILL FILL_3__14909_ (
);

FILL FILL_1__15943_ (
);

FILL FILL_1__15523_ (
);

FILL FILL_1__15103_ (
);

FILL FILL_0__14936_ (
);

NAND3X1 _14801_ (
    .A(_5276_),
    .B(_5277_),
    .C(_5284_),
    .Y(_5285_)
);

FILL FILL_0__14516_ (
);

FILL FILL_2__7683_ (
);

FILL FILL_3__12096_ (
);

FILL FILL_4__7189_ (
);

FILL FILL_2__11089_ (
);

FILL FILL_5__12843_ (
);

FILL FILL_5__12423_ (
);

FILL FILL_5__12003_ (
);

FILL FILL_4__8970_ (
);

FILL FILL_4__11836_ (
);

FILL FILL_4__8130_ (
);

FILL FILL_2__12870_ (
);

FILL FILL_4__11416_ (
);

FILL FILL_2__12450_ (
);

FILL FILL_2__12030_ (
);

FILL FILL_0__7089_ (
);

DFFSR _9195_ (
    .Q(\datapath_1.regfile_1.regOut[18] [21]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1108_[21])
);

FILL FILL_6__8056_ (
);

FILL FILL_1__16308_ (
);

FILL FILL_3__10829_ (
);

FILL FILL_3__10409_ (
);

FILL FILL_1__11863_ (
);

FILL FILL_1__11443_ (
);

FILL FILL_1__11023_ (
);

FILL FILL_0__8870_ (
);

FILL FILL_2__8888_ (
);

FILL FILL_0__8450_ (
);

FILL FILL_2__8468_ (
);

DFFSR _10721_ (
    .Q(\datapath_1.regfile_1.regOut[30] [11]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1888_[11])
);

FILL FILL_0__10436_ (
);

OAI21X1 _10301_ (
    .A(_1738_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1739_),
    .Y(_1693_[23])
);

FILL FILL_0__10016_ (
);

FILL FILL_5__6893_ (
);

DFFSR _13193_ (
    .Q(\datapath_1.mux_iord.din0 [18]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3685_[18])
);

FILL FILL_5__13628_ (
);

FILL FILL_5__13208_ (
);

FILL FILL_3__14662_ (
);

FILL FILL_3__14242_ (
);

OAI21X1 _7928_ (
    .A(_586_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .C(_587_),
    .Y(_523_[0])
);

NAND2X1 _7508_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_325_)
);

FILL FILL_1__6885_ (
);

FILL FILL_4__9755_ (
);

FILL FILL_4__9335_ (
);

FILL FILL_2__13655_ (
);

FILL SFILL99400x39050 (
);

FILL FILL_2__13235_ (
);

FILL FILL_1__12648_ (
);

FILL SFILL3400x58050 (
);

FILL FILL_1__12228_ (
);

FILL FILL_0__9655_ (
);

FILL FILL_3__7752_ (
);

FILL FILL112440x83050 (
);

FILL FILL_3__7332_ (
);

INVX1 _11926_ (
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_2992_)
);

FILL FILL_0__9235_ (
);

NAND2X1 _11506_ (
    .A(_2462__bF$buf1),
    .B(_2612_),
    .Y(_2618_)
);

FILL FILL_5__7678_ (
);

FILL SFILL104360x32050 (
);

FILL FILL_4__16034_ (
);

FILL SFILL64440x8050 (
);

FILL FILL_6__10135_ (
);

AOI22X1 _14398_ (
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .B(_3885_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_4891_)
);

FILL FILL_3__15867_ (
);

FILL FILL_3__15447_ (
);

FILL FILL_3__15027_ (
);

FILL FILL_1__16061_ (
);

FILL SFILL3800x27050 (
);

FILL FILL_3__10162_ (
);

FILL FILL_6_BUFX2_insert531 (
);

FILL SFILL64120x2050 (
);

FILL FILL_0__15894_ (
);

FILL FILL_0__15474_ (
);

FILL FILL_0__15054_ (
);

FILL FILL_6_BUFX2_insert536 (
);

FILL SFILL64040x7050 (
);

FILL FILL_1__8611_ (
);

FILL FILL_2__15801_ (
);

FILL FILL_3__8957_ (
);

FILL FILL_3__8117_ (
);

FILL FILL_5__13381_ (
);

OAI21X1 _7681_ (
    .A(_398_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .C(_399_),
    .Y(_393_[3])
);

DFFSR _7261_ (
    .Q(\datapath_1.regfile_1.regOut[3] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_133_[7])
);

FILL FILL_4__12374_ (
);

FILL FILL_2__6954_ (
);

FILL FILL_3__11787_ (
);

FILL FILL_5__9404_ (
);

FILL FILL_3__11367_ (
);

FILL FILL_0__16259_ (
);

AOI21X1 _16124_ (
    .A(_6577_),
    .B(_6556_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [26])
);

FILL FILL_0__11394_ (
);

FILL SFILL89400x37050 (
);

FILL FILL_6__15173_ (
);

FILL FILL_4__7821_ (
);

FILL FILL_5__14586_ (
);

FILL FILL_2__11721_ (
);

FILL FILL_5__14166_ (
);

FILL FILL_2__11301_ (
);

NAND2X1 _8886_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1020_)
);

NAND2X1 _8466_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_801_)
);

FILL FILL_6__7327_ (
);

FILL SFILL33640x63050 (
);

DFFSR _8046_ (
    .Q(\datapath_1.regfile_1.regOut[9] [24]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_523_[24])
);

FILL FILL_4__13999_ (
);

FILL FILL_4__13579_ (
);

FILL FILL_4__13159_ (
);

FILL FILL_2__14193_ (
);

FILL FILL_2__7739_ (
);

FILL FILL_0__7721_ (
);

FILL FILL_2__7319_ (
);

FILL FILL_0__7301_ (
);

FILL FILL_4__14940_ (
);

FILL FILL_4__14520_ (
);

FILL FILL_4__14100_ (
);

FILL FILL_0__12599_ (
);

NAND2X1 _12884_ (
    .A(vdd),
    .B(\datapath_1.rd1 [20]),
    .Y(_3595_)
);

FILL FILL_0__12179_ (
);

NAND2X1 _12464_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [8]),
    .Y(_3376_)
);

NAND3X1 _12044_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [14]),
    .C(_3034__bF$buf3),
    .Y(_3079_)
);

FILL FILL_3__13933_ (
);

FILL FILL_3__13513_ (
);

FILL FILL_4__8606_ (
);

FILL SFILL94280x43050 (
);

FILL FILL_5_BUFX2_insert550 (
);

FILL FILL_6__11093_ (
);

FILL FILL_5_BUFX2_insert551 (
);

FILL FILL_2__12506_ (
);

FILL FILL_5_BUFX2_insert552 (
);

FILL FILL_0__13960_ (
);

FILL FILL_5_BUFX2_insert553 (
);

FILL FILL_0__13540_ (
);

FILL FILL_0__13120_ (
);

FILL FILL_5_BUFX2_insert554 (
);

FILL FILL_5_BUFX2_insert555 (
);

FILL FILL_5_BUFX2_insert556 (
);

FILL FILL_5_BUFX2_insert557 (
);

FILL FILL_5_BUFX2_insert558 (
);

FILL FILL_1__11919_ (
);

FILL FILL_5_BUFX2_insert559 (
);

FILL FILL_2__15398_ (
);

FILL FILL_5__16312_ (
);

FILL SFILL79800x49050 (
);

FILL FILL_0__8506_ (
);

FILL SFILL33960x39050 (
);

FILL FILL_5__6949_ (
);

FILL FILL_4__15725_ (
);

FILL FILL_4__15305_ (
);

FILL FILL_3__9495_ (
);

FILL FILL_1_BUFX2_insert1084 (
);

OAI22X1 _13669_ (
    .A(_4176_),
    .B(_3941_),
    .C(_3960_),
    .D(_4175_),
    .Y(_4177_)
);

NOR2X1 _13249_ (
    .A(_3765_),
    .B(_3791_),
    .Y(_3792_)
);

FILL FILL_1_BUFX2_insert1085 (
);

FILL FILL_4__10440_ (
);

FILL FILL_4__10020_ (
);

FILL FILL_1_BUFX2_insert1086 (
);

FILL FILL_1_BUFX2_insert1087 (
);

FILL FILL_3__14718_ (
);

FILL FILL_1_BUFX2_insert1088 (
);

FILL FILL_1__15752_ (
);

FILL FILL_1_BUFX2_insert1089 (
);

FILL FILL_1__15332_ (
);

FILL SFILL94200x41050 (
);

FILL SFILL18760x19050 (
);

FILL FILL_0__14745_ (
);

INVX1 _14610_ (
    .A(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_5098_)
);

FILL FILL_0__14325_ (
);

FILL FILL_2__7492_ (
);

FILL FILL_2__7072_ (
);

FILL SFILL79000x21050 (
);

FILL FILL_3__7808_ (
);

FILL FILL_5__12652_ (
);

FILL FILL_5__12232_ (
);

OAI21X1 _6952_ (
    .A(_34_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .C(_35_),
    .Y(_3_[16])
);

FILL FILL_2_BUFX2_insert680 (
);

FILL SFILL8680x60050 (
);

FILL FILL_2_BUFX2_insert681 (
);

FILL FILL_2_BUFX2_insert682 (
);

FILL SFILL34040x6050 (
);

FILL FILL_2_BUFX2_insert683 (
);

FILL FILL_2_BUFX2_insert684 (
);

FILL FILL_4__11645_ (
);

FILL SFILL74280x4050 (
);

FILL FILL_2_BUFX2_insert685 (
);

FILL FILL_4__11225_ (
);

FILL FILL_2_BUFX2_insert686 (
);

FILL FILL_2_BUFX2_insert687 (
);

FILL FILL_2_BUFX2_insert688 (
);

FILL SFILL4280x59050 (
);

FILL FILL_2_BUFX2_insert689 (
);

FILL FILL_1__16117_ (
);

FILL FILL_3__10638_ (
);

FILL FILL_1__11672_ (
);

FILL FILL_1__11252_ (
);

FILL SFILL33400x3050 (
);

OAI22X1 _15815_ (
    .A(_5569_),
    .B(_6275_),
    .C(_5523_),
    .D(_4884_),
    .Y(_6276_)
);

FILL SFILL84280x41050 (
);

FILL FILL_2__8697_ (
);

NAND3X1 _10950_ (
    .A(_2071_),
    .B(_2063_),
    .C(_2082_),
    .Y(_2083_)
);

FILL FILL_0__10665_ (
);

FILL FILL_2__8277_ (
);

OAI21X1 _10530_ (
    .A(_1850_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1851_),
    .Y(_1823_[14])
);

FILL FILL_0__10245_ (
);

OAI21X1 _10110_ (
    .A(_1631_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .C(_1632_),
    .Y(_1628_[2])
);

FILL SFILL23160x54050 (
);

FILL FILL_5__13857_ (
);

FILL FILL_5__13437_ (
);

FILL FILL_3__14891_ (
);

FILL FILL_3__14471_ (
);

FILL FILL_5__13017_ (
);

FILL FILL_3__14051_ (
);

NAND2X1 _7737_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_437_)
);

NAND2X1 _7317_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_218_)
);

FILL FILL_4__9984_ (
);

FILL FILL_4__9144_ (
);

FILL FILL_2__13884_ (
);

FILL SFILL114440x67050 (
);

FILL FILL_2__13464_ (
);

FILL FILL_2__13044_ (
);

FILL SFILL109080x70050 (
);

FILL FILL_1__12877_ (
);

FILL FILL_1__12457_ (
);

FILL FILL_1__12037_ (
);

FILL FILL_6_CLKBUF1_insert132 (
);

FILL FILL_0__9884_ (
);

FILL FILL_3__7981_ (
);

FILL FILL_3__7561_ (
);

FILL FILL_0__9464_ (
);

FILL FILL_0__9044_ (
);

OAI21X1 _11735_ (
    .A(_2386_),
    .B(_2347__bF$buf3),
    .C(_2831_),
    .Y(_2832_)
);

FILL FILL_6_CLKBUF1_insert137 (
);

AOI21X1 _11315_ (
    .A(_2219_),
    .B(_2433_),
    .C(_2223_),
    .Y(_2434_)
);

FILL FILL_6__15649_ (
);

FILL FILL_5__7487_ (
);

FILL FILL_6__15229_ (
);

FILL FILL_4__16263_ (
);

FILL FILL_5__7067_ (
);

FILL FILL_3__15676_ (
);

FILL FILL_3__15256_ (
);

FILL FILL_1__16290_ (
);

FILL FILL_1__7479_ (
);

FILL FILL_3__10391_ (
);

FILL FILL_1__7059_ (
);

FILL FILL_2__14669_ (
);

FILL FILL_2__14249_ (
);

FILL FILL_0__15283_ (
);

FILL SFILL114440x22050 (
);

FILL FILL_1__8840_ (
);

FILL FILL_1__8000_ (
);

FILL FILL_2__15610_ (
);

FILL FILL_3__8766_ (
);

FILL FILL_3__8346_ (
);

FILL FILL_1__14603_ (
);

NAND2X1 _7490_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_313_)
);

NAND2X1 _7070_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_94_)
);

FILL FILL_6__11569_ (
);

FILL FILL_6__11149_ (
);

FILL FILL_4__12183_ (
);

FILL SFILL114360x29050 (
);

FILL FILL_5__9633_ (
);

FILL FILL_3__11596_ (
);

FILL FILL_5__9213_ (
);

FILL FILL_3__11176_ (
);

FILL FILL_6__12510_ (
);

FILL FILL_0__16068_ (
);

OAI21X1 _16353_ (
    .A(_6788_),
    .B(gnd),
    .C(_6789_),
    .Y(_6769_[10])
);

FILL FILL_2__10169_ (
);

FILL FILL_5__11923_ (
);

FILL FILL_1__9625_ (
);

FILL FILL_5__11503_ (
);

FILL FILL_4__7630_ (
);

FILL FILL_4__10916_ (
);

FILL FILL_4__7210_ (
);

FILL FILL_2__11950_ (
);

FILL FILL_5__14395_ (
);

FILL FILL_2__11530_ (
);

FILL FILL_2__11110_ (
);

NAND2X1 _8695_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .Y(_977_)
);

FILL FILL_1__15808_ (
);

FILL SFILL64280x82050 (
);

INVX1 _8275_ (
    .A(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_714_)
);

FILL FILL_1__10943_ (
);

FILL FILL_4__13388_ (
);

FILL FILL_1__10523_ (
);

FILL FILL_1__10103_ (
);

FILL FILL_0__7950_ (
);

FILL FILL_2__7968_ (
);

BUFX2 BUFX2_insert370 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf5 )
);

FILL FILL_2__7548_ (
);

FILL FILL_0__7110_ (
);

BUFX2 BUFX2_insert371 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf4 )
);

BUFX2 BUFX2_insert372 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf3 )
);

BUFX2 BUFX2_insert373 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf2 )
);

BUFX2 BUFX2_insert374 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf1 )
);

FILL FILL_6__13715_ (
);

BUFX2 BUFX2_insert375 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf0 )
);

BUFX2 BUFX2_insert376 (
    .A(_3196_),
    .Y(_3196__bF$buf4)
);

BUFX2 BUFX2_insert377 (
    .A(_3196_),
    .Y(_3196__bF$buf3)
);

BUFX2 BUFX2_insert378 (
    .A(_3196_),
    .Y(_3196__bF$buf2)
);

DFFSR _12693_ (
    .Q(\datapath_1.Data [30]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[30])
);

BUFX2 BUFX2_insert379 (
    .A(_3196_),
    .Y(_3196__bF$buf1)
);

AOI22X1 _12273_ (
    .A(_2_[14]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [14]),
    .Y(_3244_)
);

FILL FILL_5__12708_ (
);

FILL FILL_3__13742_ (
);

FILL FILL_3__13322_ (
);

FILL FILL_4__8835_ (
);

FILL FILL_2__12735_ (
);

FILL FILL_2__12315_ (
);

FILL FILL_1__11728_ (
);

FILL FILL_1__11308_ (
);

FILL FILL112440x78050 (
);

FILL FILL_5__16121_ (
);

FILL FILL_0__8735_ (
);

FILL FILL_0__8315_ (
);

FILL SFILL104360x27050 (
);

FILL FILL_4__15954_ (
);

FILL FILL_4__15534_ (
);

FILL FILL_4__15114_ (
);

AOI22X1 _13898_ (
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .B(_4225_),
    .C(_3885_),
    .D(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_4401_)
);

INVX1 _13478_ (
    .A(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_3989_)
);

DFFSR _13058_ (
    .Q(_2_[11]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3620_[11])
);

FILL FILL_3__14947_ (
);

FILL FILL_1__15981_ (
);

FILL FILL_3__14527_ (
);

FILL FILL_1__15561_ (
);

FILL FILL_3__14107_ (
);

FILL FILL_1__15141_ (
);

FILL FILL112040x64050 (
);

FILL FILL_0__14974_ (
);

FILL FILL_0__14554_ (
);

FILL FILL_0__14134_ (
);

FILL SFILL79320x50 (
);

FILL FILL_3__7617_ (
);

FILL FILL_5__12881_ (
);

FILL FILL_5__12461_ (
);

FILL FILL_5__12041_ (
);

FILL FILL112440x33050 (
);

FILL FILL_4__16319_ (
);

FILL FILL_4__11874_ (
);

FILL FILL_4__11454_ (
);

FILL FILL_4__11034_ (
);

FILL FILL_1__16346_ (
);

FILL FILL_5__8904_ (
);

FILL FILL_3__10447_ (
);

FILL FILL_3__10027_ (
);

FILL FILL_1__11481_ (
);

FILL FILL_1__11061_ (
);

FILL FILL_0__15759_ (
);

FILL FILL_0__15339_ (
);

NOR2X1 _15624_ (
    .A(_6089_),
    .B(_5539__bF$buf3),
    .Y(_6090_)
);

OAI22X1 _15204_ (
    .A(_5472__bF$buf1),
    .B(_4116_),
    .C(_4097_),
    .D(_5483__bF$buf3),
    .Y(_5681_)
);

FILL FILL_0__10894_ (
);

FILL FILL_2__8086_ (
);

FILL FILL_0__10054_ (
);

FILL FILL_4__6901_ (
);

FILL FILL_5__13666_ (
);

FILL FILL_2__10801_ (
);

FILL FILL_5__13246_ (
);

FILL FILL_3__14280_ (
);

NAND2X1 _7966_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_549_)
);

NAND2X1 _7546_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_330_)
);

DFFSR _7126_ (
    .Q(\datapath_1.regfile_1.regOut[2] [0]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_68_[0])
);

FILL FILL_4__9793_ (
);

FILL FILL_4__9373_ (
);

FILL FILL_4__12659_ (
);

FILL FILL_4__12239_ (
);

FILL FILL_2__13693_ (
);

FILL FILL_2__13273_ (
);

FILL FILL_1__12266_ (
);

FILL FILL_4__13600_ (
);

NAND2X1 _16409_ (
    .A(gnd),
    .B(gnd),
    .Y(_6827_)
);

FILL FILL_3__7370_ (
);

FILL FILL_0__9273_ (
);

OAI21X1 _11964_ (
    .A(_3016_),
    .B(IorD_bF$buf6),
    .C(_3017_),
    .Y(_1_[25])
);

FILL FILL_0__11679_ (
);

FILL FILL_0__11259_ (
);

AOI22X1 _11544_ (
    .A(_2219_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf0),
    .D(_2217_),
    .Y(_2654_)
);

FILL FILL_5_CLKBUF1_insert120 (
);

INVX1 _11124_ (
    .A(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2243_)
);

FILL FILL_5_CLKBUF1_insert121 (
);

FILL FILL_5_CLKBUF1_insert122 (
);

FILL FILL_5__7296_ (
);

FILL FILL_5_CLKBUF1_insert123 (
);

FILL FILL_5_CLKBUF1_insert124 (
);

FILL FILL_4__16072_ (
);

FILL FILL_5_CLKBUF1_insert125 (
);

FILL SFILL94280x38050 (
);

FILL FILL_5_CLKBUF1_insert126 (
);

FILL FILL_5_CLKBUF1_insert127 (
);

FILL FILL_5_CLKBUF1_insert128 (
);

FILL FILL_5_CLKBUF1_insert129 (
);

FILL FILL_0__12620_ (
);

FILL FILL_3__15485_ (
);

FILL FILL_3__15065_ (
);

FILL FILL_0__12200_ (
);

FILL FILL_1__7288_ (
);

FILL FILL_2__14898_ (
);

FILL FILL_2__14478_ (
);

FILL SFILL115240x21050 (
);

FILL FILL_2__14058_ (
);

FILL FILL_6_BUFX2_insert914 (
);

FILL FILL_0__15092_ (
);

FILL FILL_5__15812_ (
);

FILL SFILL58840x62050 (
);

FILL FILL_4__14805_ (
);

FILL FILL_3__8995_ (
);

FILL FILL_3__8575_ (
);

INVX1 _12749_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_3525_)
);

AOI22X1 _12329_ (
    .A(_2_[28]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3286_)
);

FILL FILL_1__14832_ (
);

FILL FILL_1__14412_ (
);

FILL FILL_0__13825_ (
);

FILL FILL_0__13405_ (
);

FILL FILL_2__6992_ (
);

FILL FILL_5__9862_ (
);

FILL FILL_5__9022_ (
);

FILL SFILL23640x56050 (
);

FILL FILL_0__16297_ (
);

NAND2X1 _16162_ (
    .A(_6614_),
    .B(_6609_),
    .Y(_6615_)
);

FILL SFILL79000x16050 (
);

FILL FILL_2__10398_ (
);

FILL FILL_5__11732_ (
);

FILL FILL_1__9854_ (
);

FILL FILL_5__11312_ (
);

FILL FILL_1__9014_ (
);

FILL SFILL8680x55050 (
);

FILL FILL_2__16204_ (
);

FILL FILL_4__10305_ (
);

FILL FILL_1__15617_ (
);

INVX1 _8084_ (
    .A(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_607_)
);

FILL FILL_1__10752_ (
);

FILL FILL_2__7357_ (
);

FILL SFILL69080x50 (
);

FILL SFILL53400x74050 (
);

FILL SFILL109480x79050 (
);

NAND3X1 _12082_ (
    .A(_3105_),
    .B(_3106_),
    .C(_3107_),
    .Y(\datapath_1.mux_pcsrc.dout [23])
);

FILL FILL_5__12517_ (
);

FILL FILL_3__13971_ (
);

FILL FILL_3__13551_ (
);

FILL SFILL8600x53050 (
);

FILL FILL_3__13131_ (
);

FILL FILL_4__8644_ (
);

FILL FILL_4__8224_ (
);

FILL FILL_5_BUFX2_insert930 (
);

FILL FILL_2__12964_ (
);

FILL FILL_5_BUFX2_insert931 (
);

FILL SFILL8680x10050 (
);

FILL FILL_5_BUFX2_insert932 (
);

FILL FILL_2__12124_ (
);

FILL FILL_5_BUFX2_insert933 (
);

FILL FILL_5_BUFX2_insert934 (
);

FILL FILL_5_BUFX2_insert935 (
);

OAI21X1 _9289_ (
    .A(_1226_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .C(_1227_),
    .Y(_1173_[27])
);

FILL FILL_5_BUFX2_insert936 (
);

FILL FILL_5_BUFX2_insert937 (
);

FILL FILL_1__11957_ (
);

FILL FILL_5_BUFX2_insert938 (
);

FILL FILL_5_BUFX2_insert939 (
);

FILL FILL_1__11537_ (
);

FILL FILL_1__11117_ (
);

FILL SFILL84200x34050 (
);

FILL SFILL74280x79050 (
);

FILL FILL_0__8964_ (
);

FILL FILL_5__16350_ (
);

NAND2X1 _10815_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_2001_)
);

FILL FILL_0__8124_ (
);

FILL FILL_5__6987_ (
);

FILL FILL_4__15763_ (
);

FILL FILL_4__15343_ (
);

FILL SFILL13640x54050 (
);

NOR2X1 _13287_ (
    .A(_3781_),
    .B(_3825_),
    .Y(\datapath_1.regfile_1.regEn [5])
);

FILL FILL_2__9923_ (
);

FILL FILL_3__14756_ (
);

FILL FILL_2__9503_ (
);

FILL FILL_1__15790_ (
);

FILL FILL_3__14336_ (
);

FILL SFILL109480x34050 (
);

FILL FILL_1__15370_ (
);

FILL FILL_1__6979_ (
);

FILL FILL_4__9849_ (
);

FILL FILL_4__9429_ (
);

FILL FILL_4__9009_ (
);

FILL FILL_2__13749_ (
);

FILL FILL_2__13329_ (
);

FILL FILL_0__14783_ (
);

FILL FILL_0__14363_ (
);

FILL SFILL17960x62050 (
);

FILL SFILL114440x17050 (
);

FILL FILL_1__7500_ (
);

FILL FILL_3__7846_ (
);

FILL FILL_0__9749_ (
);

FILL FILL_3__7426_ (
);

FILL FILL_5__12270_ (
);

FILL SFILL74280x34050 (
);

NAND2X1 _6990_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_61_)
);

FILL FILL_4__16128_ (
);

FILL FILL_4__11683_ (
);

FILL FILL_4__11263_ (
);

FILL SFILL99480x83050 (
);

FILL FILL_1__16155_ (
);

FILL FILL_5__8713_ (
);

FILL FILL_3__10676_ (
);

FILL FILL_3__10256_ (
);

FILL FILL_1__11290_ (
);

FILL FILL_0__15988_ (
);

FILL FILL_0__15568_ (
);

AOI22X1 _15853_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [20]),
    .C(\datapath_1.regfile_1.regOut[22] [20]),
    .D(_5650_),
    .Y(_6313_)
);

NAND3X1 _15433_ (
    .A(_5898_),
    .B(_5899_),
    .C(_5903_),
    .Y(_5904_)
);

FILL FILL_0__15148_ (
);

OR2X2 _15013_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5493_)
);

FILL FILL_0__10283_ (
);

FILL FILL_3_BUFX2_insert1010 (
);

FILL FILL_1__8705_ (
);

FILL FILL_3_BUFX2_insert1011 (
);

FILL FILL_6__14482_ (
);

FILL FILL_3_BUFX2_insert1012 (
);

FILL FILL_3_BUFX2_insert1013 (
);

FILL FILL_3_BUFX2_insert1014 (
);

FILL FILL_3_BUFX2_insert1015 (
);

FILL FILL_3_BUFX2_insert1016 (
);

FILL FILL_3_BUFX2_insert1017 (
);

FILL FILL_3_BUFX2_insert1018 (
);

FILL FILL_5__13895_ (
);

FILL FILL_5__13475_ (
);

FILL FILL_3_BUFX2_insert1019 (
);

FILL SFILL74200x32050 (
);

FILL SFILL13560x16050 (
);

DFFSR _7775_ (
    .Q(\datapath_1.regfile_1.regOut[7] [9]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_393_[9])
);

FILL SFILL95160x30050 (
);

INVX1 _7355_ (
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_243_)
);

FILL FILL_4__12888_ (
);

FILL FILL_4__12468_ (
);

FILL FILL_4__12048_ (
);

FILL FILL_2__13082_ (
);

FILL FILL_5__9918_ (
);

FILL FILL_1__12495_ (
);

FILL FILL_1__12075_ (
);

NOR3X1 _16218_ (
    .A(_6664_),
    .B(_6668_),
    .C(_6665_),
    .Y(_6669_)
);

NOR2X1 _11773_ (
    .A(_2867_),
    .B(_2858_),
    .Y(_2868_)
);

FILL FILL_0__9082_ (
);

FILL FILL_0__11488_ (
);

OAI21X1 _11353_ (
    .A(_2456_),
    .B(_2117_),
    .C(_2470__bF$buf3),
    .Y(_2471_)
);

FILL FILL_0__11068_ (
);

FILL FILL_3__12402_ (
);

FILL SFILL104440x15050 (
);

FILL FILL_2__11815_ (
);

FILL FILL_4_CLKBUF1_insert111 (
);

FILL FILL_4_CLKBUF1_insert112 (
);

FILL FILL_3__15294_ (
);

FILL FILL_4_CLKBUF1_insert113 (
);

FILL FILL_4_CLKBUF1_insert114 (
);

FILL FILL_4_CLKBUF1_insert115 (
);

FILL FILL_4_CLKBUF1_insert116 (
);

FILL FILL112120x52050 (
);

FILL FILL_1__7097_ (
);

FILL FILL_4_CLKBUF1_insert117 (
);

FILL FILL_1__10808_ (
);

FILL FILL_4_CLKBUF1_insert118 (
);

FILL FILL_4_CLKBUF1_insert119 (
);

FILL FILL_2__14287_ (
);

FILL FILL_5__15621_ (
);

FILL FILL_5__15201_ (
);

FILL FILL_0__7815_ (
);

INVX1 _9921_ (
    .A(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_1547_)
);

INVX1 _9501_ (
    .A(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_1328_)
);

FILL FILL_4__14614_ (
);

FILL FILL_3__8384_ (
);

INVX1 _12978_ (
    .A(_2_[9]),
    .Y(_3637_)
);

DFFSR _12558_ (
    .Q(ALUOut[23]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3360_[23])
);

OAI21X1 _12138_ (
    .A(_3144_),
    .B(ALUSrcA_bF$buf7),
    .C(_3145_),
    .Y(\datapath_1.alu_1.ALUInA [7])
);

FILL FILL_3__13607_ (
);

FILL FILL_1__14641_ (
);

FILL FILL112040x59050 (
);

FILL FILL_1__14221_ (
);

FILL FILL_0__13634_ (
);

FILL FILL_0__13214_ (
);

FILL FILL_3__16079_ (
);

FILL FILL_5__9671_ (
);

FILL FILL_5__9251_ (
);

FILL SFILL64200x30050 (
);

NAND2X1 _16391_ (
    .A(gnd),
    .B(gnd),
    .Y(_6815_)
);

FILL FILL_5__16406_ (
);

FILL FILL_5__11961_ (
);

FILL FILL_1__9663_ (
);

FILL FILL_5__11541_ (
);

FILL FILL112440x28050 (
);

FILL FILL_1__9243_ (
);

FILL FILL_5__11121_ (
);

FILL FILL_4__15819_ (
);

FILL FILL_2__16013_ (
);

FILL FILL_4__10954_ (
);

FILL FILL_3__9169_ (
);

FILL FILL_4__10534_ (
);

FILL FILL_4__10114_ (
);

FILL FILL_1__15846_ (
);

FILL FILL_1__15426_ (
);

FILL FILL_1__15006_ (
);

FILL FILL_1__10981_ (
);

FILL FILL_1__10561_ (
);

FILL FILL_1__10141_ (
);

FILL FILL112040x14050 (
);

FILL FILL_0__14839_ (
);

INVX1 _14704_ (
    .A(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_5190_)
);

FILL FILL_0__14419_ (
);

FILL FILL_2__7586_ (
);

BUFX2 BUFX2_insert750 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf4 )
);

BUFX2 BUFX2_insert751 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf3 )
);

FILL FILL_2__7166_ (
);

BUFX2 BUFX2_insert752 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf2 )
);

BUFX2 BUFX2_insert753 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf1 )
);

BUFX2 BUFX2_insert754 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf0 )
);

BUFX2 BUFX2_insert755 (
    .A(_3198_),
    .Y(_3198__bF$buf4)
);

BUFX2 BUFX2_insert756 (
    .A(_3198_),
    .Y(_3198__bF$buf3)
);

BUFX2 BUFX2_insert757 (
    .A(_3198_),
    .Y(_3198__bF$buf2)
);

BUFX2 BUFX2_insert758 (
    .A(_3198_),
    .Y(_3198__bF$buf1)
);

BUFX2 BUFX2_insert759 (
    .A(_3198_),
    .Y(_3198__bF$buf0)
);

FILL FILL_5__12746_ (
);

FILL FILL_3__13780_ (
);

FILL FILL_5__12326_ (
);

FILL FILL_3__13360_ (
);

FILL FILL_4__8873_ (
);

FILL FILL_4__8453_ (
);

FILL FILL_4__11739_ (
);

FILL FILL_2__12773_ (
);

FILL FILL_4__11319_ (
);

FILL FILL_2__12353_ (
);

OAI21X1 _9098_ (
    .A(_1119_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .C(_1120_),
    .Y(_1108_[6])
);

FILL FILL_1__11766_ (
);

FILL FILL_1__11346_ (
);

NAND3X1 _15909_ (
    .A(_6362_),
    .B(_6363_),
    .C(_6367_),
    .Y(_6368_)
);

FILL FILL_0__8773_ (
);

FILL FILL_3__6870_ (
);

FILL FILL_0__8353_ (
);

FILL FILL_0__10759_ (
);

NAND2X1 _10624_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1894_)
);

DFFSR _10204_ (
    .Q(\datapath_1.regfile_1.regOut[26] [6]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_1628_[6])
);

FILL FILL_6__14958_ (
);

FILL FILL_4__15992_ (
);

FILL FILL_4__15572_ (
);

FILL FILL_4__15152_ (
);

OAI21X1 _13096_ (
    .A(_3694_),
    .B(PCEn_bF$buf3),
    .C(_3695_),
    .Y(_3685_[5])
);

FILL FILL_3__14985_ (
);

FILL FILL_2__9732_ (
);

FILL FILL_3__14565_ (
);

FILL FILL_0__11700_ (
);

FILL FILL_3__14145_ (
);

FILL FILL_4_BUFX2_insert590 (
);

FILL FILL_4_BUFX2_insert591 (
);

FILL FILL_4__9658_ (
);

FILL FILL_4_BUFX2_insert592 (
);

FILL FILL_4__9238_ (
);

FILL FILL_2__13978_ (
);

FILL FILL_4_BUFX2_insert593 (
);

FILL FILL_4_BUFX2_insert594 (
);

FILL FILL_2__13558_ (
);

FILL FILL_4_BUFX2_insert595 (
);

FILL FILL_0__14592_ (
);

FILL FILL_2__13138_ (
);

FILL FILL_0__14172_ (
);

FILL FILL_4_BUFX2_insert596 (
);

FILL FILL_4_BUFX2_insert597 (
);

FILL FILL_4_BUFX2_insert598 (
);

FILL FILL_4_BUFX2_insert599 (
);

FILL FILL_0__9978_ (
);

FILL FILL_0__9138_ (
);

NOR2X1 _11829_ (
    .A(_2913_),
    .B(_2918_),
    .Y(_2919_)
);

FILL FILL_3__7235_ (
);

AOI21X1 _11409_ (
    .A(_2238_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_)
);

FILL FILL_1__13912_ (
);

FILL FILL_4__16357_ (
);

FILL FILL_4__11492_ (
);

FILL FILL_4__11072_ (
);

FILL FILL_0__12905_ (
);

FILL FILL_1__16384_ (
);

FILL FILL_5__8522_ (
);

FILL FILL_5__8102_ (
);

FILL FILL_3__10065_ (
);

FILL FILL_0__15797_ (
);

FILL FILL_0__15377_ (
);

AOI22X1 _15662_ (
    .A(_5565__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [15]),
    .C(\datapath_1.regfile_1.regOut[5] [15]),
    .D(_5700_),
    .Y(_6127_)
);

NAND2X1 _15242_ (
    .A(_5475_),
    .B(_5460_),
    .Y(_5718_)
);

FILL FILL_5__10812_ (
);

FILL FILL_1__8514_ (
);

FILL FILL_2__15704_ (
);

FILL FILL_5__13284_ (
);

INVX1 _7584_ (
    .A(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_355_)
);

INVX1 _7164_ (
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_136_)
);

FILL FILL_4__12697_ (
);

FILL FILL_4__12277_ (
);

FILL FILL_3__9801_ (
);

FILL FILL_2__6857_ (
);

FILL FILL_5__9727_ (
);

DFFSR _16447_ (
    .Q(\datapath_1.regfile_1.regOut[0] [30]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_6769_[30])
);

NOR2X1 _16027_ (
    .A(_6482_),
    .B(_6480_),
    .Y(_6483_)
);

AOI21X1 _11582_ (
    .A(_2523_),
    .B(_2688_),
    .C(_2263_),
    .Y(_2689_)
);

FILL FILL_0__11297_ (
);

OAI21X1 _11162_ (
    .A(_2223_),
    .B(_2224_),
    .C(_2280_),
    .Y(_2281_)
);

FILL FILL_1__9719_ (
);

FILL SFILL8600x48050 (
);

FILL FILL_3__12631_ (
);

FILL FILL_6__15076_ (
);

FILL FILL_3__12211_ (
);

FILL FILL_4__7724_ (
);

FILL FILL_4__7304_ (
);

FILL SFILL13720x42050 (
);

FILL FILL_5__14489_ (
);

FILL FILL_2__11624_ (
);

FILL FILL_5__14069_ (
);

FILL FILL_2__11204_ (
);

OAI21X1 _8789_ (
    .A(_974_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .C(_975_),
    .Y(_913_[31])
);

OAI21X1 _8369_ (
    .A(_755_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .C(_756_),
    .Y(_718_[19])
);

FILL FILL_1__10617_ (
);

FILL SFILL53800x38050 (
);

FILL SFILL94760x7050 (
);

FILL FILL_2__14096_ (
);

FILL SFILL84200x29050 (
);

FILL FILL_5__15850_ (
);

FILL FILL_5__15430_ (
);

FILL FILL_5__15010_ (
);

FILL FILL_0__7624_ (
);

FILL FILL_0__7204_ (
);

INVX1 _9730_ (
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_1440_)
);

DFFSR _9310_ (
    .Q(\datapath_1.regfile_1.regOut[19] [8]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_1173_[8])
);

FILL FILL_1__13089_ (
);

FILL FILL_4__14843_ (
);

FILL FILL_4__14423_ (
);

FILL FILL_4__14003_ (
);

FILL SFILL13640x49050 (
);

OAI21X1 _12787_ (
    .A(_3549_),
    .B(IRWrite_bF$buf4),
    .C(_3550_),
    .Y(_3490_[30])
);

FILL FILL_3__8193_ (
);

INVX1 _12367_ (
    .A(ALUOut[8]),
    .Y(_3310_)
);

FILL FILL_3__13836_ (
);

FILL SFILL109480x29050 (
);

FILL FILL_1__14870_ (
);

FILL FILL_3__13416_ (
);

FILL FILL_1__14450_ (
);

FILL FILL_1__14030_ (
);

FILL FILL_4__8509_ (
);

FILL FILL_2__12829_ (
);

FILL FILL_0__13863_ (
);

FILL FILL_2__12409_ (
);

FILL FILL_0__13443_ (
);

FILL FILL_0__13023_ (
);

FILL FILL_5__9480_ (
);

FILL FILL_3__6926_ (
);

FILL FILL_5__16215_ (
);

FILL FILL_0__8829_ (
);

FILL FILL_1__9892_ (
);

FILL FILL_5__11770_ (
);

FILL SFILL74280x29050 (
);

FILL FILL_1__9472_ (
);

FILL FILL_5__11350_ (
);

FILL FILL_4__15628_ (
);

FILL FILL_4__15208_ (
);

FILL FILL_2__16242_ (
);

FILL FILL_3__9398_ (
);

FILL FILL_4__10763_ (
);

FILL SFILL99480x78050 (
);

FILL FILL_1__15655_ (
);

FILL FILL_1__15235_ (
);

FILL FILL_1__10790_ (
);

FILL FILL_1__10370_ (
);

INVX1 _14933_ (
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_5414_)
);

FILL FILL_0__14648_ (
);

FILL FILL_0__14228_ (
);

INVX1 _14513_ (
    .A(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_5003_)
);

FILL SFILL34120x31050 (
);

FILL FILL_5__12975_ (
);

FILL SFILL74200x27050 (
);

FILL FILL_5__12135_ (
);

BUFX2 _6855_ (
    .A(_1_[17]),
    .Y(memoryAddress[17])
);

FILL FILL_4__8262_ (
);

FILL FILL_4__11968_ (
);

FILL FILL_4__11548_ (
);

FILL FILL_2__12582_ (
);

FILL FILL_4__11128_ (
);

FILL FILL_2__12162_ (
);

FILL FILL_1__11995_ (
);

FILL SFILL109560x50 (
);

FILL FILL_1__11575_ (
);

FILL SFILL99480x33050 (
);

FILL FILL_1__11155_ (
);

OAI22X1 _15718_ (
    .A(_4718_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf1),
    .D(_4751_),
    .Y(_6182_)
);

FILL FILL_0__10988_ (
);

FILL FILL_0__8582_ (
);

DFFSR _10853_ (
    .Q(\datapath_1.regfile_1.regOut[31] [15]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_1953_[15])
);

FILL FILL_0__10568_ (
);

FILL FILL_0__10148_ (
);

INVX1 _10433_ (
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_1807_)
);

INVX1 _10013_ (
    .A(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_1588_)
);

FILL FILL_3__11902_ (
);

FILL FILL_4__15381_ (
);

FILL FILL_3__14794_ (
);

FILL FILL_2__9541_ (
);

FILL FILL_2__9121_ (
);

FILL FILL_3__14374_ (
);

FILL FILL_4__9887_ (
);

FILL FILL_4__9467_ (
);

FILL FILL_2__13787_ (
);

FILL FILL_2__13367_ (
);

FILL FILL_5__14701_ (
);

FILL SFILL24520x43050 (
);

FILL SFILL89800x8050 (
);

FILL FILL_0__9787_ (
);

FILL FILL_3__7884_ (
);

FILL FILL_3__7464_ (
);

FILL FILL_0__9367_ (
);

FILL FILL_3__7044_ (
);

NAND3X1 _11638_ (
    .A(_2739_),
    .B(_2741_),
    .C(_2735_),
    .Y(\datapath_1.ALUResult [16])
);

NAND2X1 _11218_ (
    .A(_2334_),
    .B(_2336_),
    .Y(_2337_)
);

FILL FILL_1__13721_ (
);

FILL SFILL28840x51050 (
);

FILL FILL_1__13301_ (
);

FILL FILL_4__16166_ (
);

FILL FILL_6__10687_ (
);

FILL FILL_3__15999_ (
);

FILL FILL_0__12714_ (
);

FILL FILL_3__15579_ (
);

FILL FILL_3__15159_ (
);

FILL SFILL89400x7050 (
);

FILL FILL_1__16193_ (
);

FILL SFILL33800x34050 (
);

FILL FILL_5__8751_ (
);

FILL SFILL64200x25050 (
);

FILL FILL_5__8331_ (
);

FILL FILL_3__10294_ (
);

AOI21X1 _15891_ (
    .A(_6326_),
    .B(_6350_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [20])
);

FILL FILL_0__15186_ (
);

NOR2X1 _15471_ (
    .A(_5940_),
    .B(_5939_),
    .Y(_5941_)
);

FILL FILL_5__15906_ (
);

NOR3X1 _15051_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .C(_5459__bF$buf1),
    .Y(_5531_)
);

FILL FILL_3__16100_ (
);

FILL FILL_1__8743_ (
);

FILL FILL_5__10621_ (
);

FILL FILL_1__8323_ (
);

FILL FILL_2__15933_ (
);

FILL FILL_2__15513_ (
);

FILL FILL_3__8249_ (
);

FILL FILL_5__13093_ (
);

FILL FILL_1__14926_ (
);

DFFSR _7393_ (
    .Q(\datapath_1.regfile_1.regOut[4] [11]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_198_[11])
);

FILL FILL_1__14506_ (
);

FILL FILL_4__12086_ (
);

FILL FILL_3__9610_ (
);

FILL FILL_0__13919_ (
);

FILL FILL_5__9536_ (
);

FILL FILL_3__11499_ (
);

FILL FILL_5__9116_ (
);

FILL FILL_3__11079_ (
);

FILL FILL_6__12413_ (
);

OAI22X1 _16256_ (
    .A(_5384_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf3),
    .D(_6705_),
    .Y(_6706_)
);

INVX1 _11391_ (
    .A(_2196_),
    .Y(_2508_)
);

FILL FILL_5__11826_ (
);

FILL FILL_3__12860_ (
);

FILL FILL_1__9528_ (
);

FILL FILL_5__11406_ (
);

FILL FILL_3__12440_ (
);

FILL FILL_1__9108_ (
);

FILL FILL_3__12020_ (
);

FILL FILL_4__7953_ (
);

FILL FILL_4__7113_ (
);

FILL FILL_4__10819_ (
);

FILL FILL_2__11853_ (
);

FILL FILL_5__14298_ (
);

FILL FILL_2__11433_ (
);

FILL FILL_2__11013_ (
);

OAI21X1 _8598_ (
    .A(_867_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .C(_868_),
    .Y(_848_[10])
);

DFFSR _8178_ (
    .Q(\datapath_1.regfile_1.regOut[10] [28]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_588_[28])
);

FILL FILL_1__10426_ (
);

FILL FILL_1__10006_ (
);

FILL FILL_0__7853_ (
);

FILL FILL_0__7433_ (
);

FILL FILL_6__13618_ (
);

FILL FILL_4__14652_ (
);

FILL FILL_4__14232_ (
);

FILL SFILL54200x23050 (
);

OAI21X1 _12596_ (
    .A(_3442_),
    .B(vdd),
    .C(_3443_),
    .Y(_3425_[9])
);

NAND2X1 _12176_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [20]),
    .Y(_3171_)
);

FILL FILL_3__13645_ (
);

FILL FILL_3__13225_ (
);

FILL FILL_4__8738_ (
);

FILL FILL_4__8318_ (
);

FILL FILL_2__12638_ (
);

FILL FILL_0__13672_ (
);

FILL FILL_2__12218_ (
);

FILL FILL_0__13252_ (
);

FILL SFILL23720x39050 (
);

FILL FILL_0__8638_ (
);

FILL FILL_5__16024_ (
);

INVX2 _10909_ (
    .A(_2054_),
    .Y(_2055_)
);

FILL FILL_0__8218_ (
);

FILL FILL_1__9281_ (
);

FILL FILL_4__15857_ (
);

FILL FILL_4__15437_ (
);

FILL FILL_4__15017_ (
);

FILL FILL_2__16051_ (
);

FILL FILL_4__10992_ (
);

FILL FILL_4__10572_ (
);

FILL FILL_4__10152_ (
);

FILL FILL_1__15884_ (
);

FILL FILL_1__15464_ (
);

FILL FILL_1__15044_ (
);

FILL FILL_5__7602_ (
);

FILL FILL_0__14877_ (
);

FILL FILL_0__14457_ (
);

AOI21X1 _14742_ (
    .A(_5201_),
    .B(_5227_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [26])
);

FILL FILL_0__14037_ (
);

NAND3X1 _14322_ (
    .A(_4807_),
    .B(_4808_),
    .C(_4815_),
    .Y(_4816_)
);

FILL FILL_5__12784_ (
);

FILL FILL_5__12364_ (
);

FILL FILL_4__8491_ (
);

FILL FILL_4__11777_ (
);

FILL FILL_4__8071_ (
);

FILL FILL_4__11357_ (
);

FILL SFILL48920x43050 (
);

FILL FILL_2__12391_ (
);

FILL SFILL13320x68050 (
);

FILL FILL_1__16249_ (
);

FILL FILL_1__11384_ (
);

INVX1 _15947_ (
    .A(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_6405_)
);

FILL SFILL99160x8050 (
);

OAI22X1 _15527_ (
    .A(_5518__bF$buf3),
    .B(_5995_),
    .C(_5503__bF$buf2),
    .D(_5994_),
    .Y(_5996_)
);

INVX1 _15107_ (
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_5586_)
);

FILL FILL_0__10797_ (
);

FILL FILL_0__8391_ (
);

INVX1 _10662_ (
    .A(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_1919_)
);

FILL FILL_0__10377_ (
);

INVX1 _10242_ (
    .A(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_1700_)
);

FILL FILL_3__11711_ (
);

FILL FILL_4__15190_ (
);

FILL SFILL13720x37050 (
);

FILL FILL_5__13989_ (
);

FILL FILL_2__9770_ (
);

FILL FILL_5__13569_ (
);

FILL FILL_2__10704_ (
);

FILL FILL_5__13149_ (
);

FILL FILL_2__9350_ (
);

OAI21X1 _7869_ (
    .A(_503_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .C(_504_),
    .Y(_458_[23])
);

FILL FILL_3__14183_ (
);

FILL SFILL109560x17050 (
);

OAI21X1 _7449_ (
    .A(_284_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_285_),
    .Y(_263_[11])
);

FILL FILL_4_BUFX2_insert970 (
);

DFFSR _7029_ (
    .Q(\datapath_1.regfile_1.regOut[1] [31]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_3_[31])
);

FILL FILL_4_BUFX2_insert971 (
);

FILL FILL_4__9276_ (
);

FILL FILL_4_BUFX2_insert972 (
);

FILL FILL_4_BUFX2_insert973 (
);

FILL SFILL109400x6050 (
);

FILL FILL_2__13596_ (
);

FILL FILL_4_BUFX2_insert974 (
);

FILL FILL_4_BUFX2_insert975 (
);

FILL FILL_4_BUFX2_insert976 (
);

FILL FILL_4_BUFX2_insert977 (
);

FILL FILL_5__14930_ (
);

FILL FILL_5__14510_ (
);

FILL FILL_4_BUFX2_insert978 (
);

FILL FILL_4_BUFX2_insert979 (
);

DFFSR _8810_ (
    .Q(\datapath_1.regfile_1.regOut[15] [20]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_913_[20])
);

FILL FILL_1__12589_ (
);

FILL FILL_1__12169_ (
);

FILL FILL_4__13923_ (
);

FILL FILL_4__13503_ (
);

FILL FILL_3__7693_ (
);

FILL FILL_0__9596_ (
);

NOR2X1 _11867_ (
    .A(\datapath_1.ALUResult [22]),
    .B(\datapath_1.ALUResult [19]),
    .Y(_2954_)
);

AOI21X1 _11447_ (
    .A(_2360_),
    .B(_2362_),
    .C(_2562_),
    .Y(_2563_)
);

OR2X2 _11027_ (
    .A(_2140_),
    .B(_2145_),
    .Y(_2146_)
);

FILL FILL_3__12916_ (
);

FILL FILL_1__13950_ (
);

FILL FILL_4__16395_ (
);

FILL FILL_1__13530_ (
);

FILL FILL_5__7199_ (
);

FILL FILL_1__13110_ (
);

FILL FILL_2__11909_ (
);

FILL FILL_3__15388_ (
);

FILL FILL_0__12523_ (
);

FILL FILL_0__12103_ (
);

FILL FILL_5__8980_ (
);

FILL FILL_5__8140_ (
);

NOR2X1 _15280_ (
    .A(_5753_),
    .B(_5754_),
    .Y(_5755_)
);

FILL FILL_5__15715_ (
);

FILL SFILL38920x41050 (
);

FILL FILL_1__8972_ (
);

FILL FILL_5__10430_ (
);

FILL FILL_5__10010_ (
);

FILL FILL_1__8132_ (
);

FILL FILL_4__14708_ (
);

FILL FILL_2__15742_ (
);

FILL FILL_2__15322_ (
);

FILL FILL_3__8898_ (
);

FILL FILL_3__8478_ (
);

FILL FILL_3__8058_ (
);

FILL FILL_1__14735_ (
);

FILL FILL_1__14315_ (
);

FILL FILL_0__13728_ (
);

FILL FILL_0__13308_ (
);

FILL SFILL38840x48050 (
);

FILL FILL_2__6895_ (
);

FILL FILL_5__9765_ (
);

FILL FILL_5__9345_ (
);

FILL FILL_0_BUFX2_insert1090 (
);

FILL FILL_0_BUFX2_insert1091 (
);

FILL FILL_0_BUFX2_insert1092 (
);

FILL FILL_0_BUFX2_insert1093 (
);

NOR2X1 _16065_ (
    .A(_6519_),
    .B(_6517_),
    .Y(_6520_)
);

FILL SFILL3560x40050 (
);

FILL FILL_5__11635_ (
);

FILL FILL_1__9757_ (
);

FILL FILL_5__11215_ (
);

FILL FILL_1__9337_ (
);

FILL FILL_3_BUFX2_insert990 (
);

FILL FILL_2__16107_ (
);

FILL FILL_4__7762_ (
);

FILL FILL_3_BUFX2_insert991 (
);

FILL FILL_4__7342_ (
);

FILL FILL_3_BUFX2_insert992 (
);

FILL FILL_4__10628_ (
);

FILL FILL_3_BUFX2_insert993 (
);

FILL FILL_2__11662_ (
);

FILL FILL_3_BUFX2_insert994 (
);

FILL FILL_2__11242_ (
);

FILL FILL_3_BUFX2_insert995 (
);

FILL FILL_3_BUFX2_insert996 (
);

FILL FILL_3_BUFX2_insert997 (
);

FILL FILL_3_BUFX2_insert998 (
);

FILL FILL_3_BUFX2_insert999 (
);

FILL SFILL99480x28050 (
);

FILL FILL_1__10655_ (
);

FILL FILL_1__10235_ (
);

FILL FILL_0__7242_ (
);

FILL FILL_4__14881_ (
);

FILL FILL_4__14461_ (
);

FILL FILL_4__14041_ (
);

FILL SFILL69240x2050 (
);

FILL FILL_3__13874_ (
);

FILL FILL_2__8621_ (
);

FILL FILL_2__8201_ (
);

FILL FILL_3__13454_ (
);

FILL FILL_3__13034_ (
);

FILL FILL_4__8967_ (
);

FILL FILL_4__8127_ (
);

FILL FILL_2__12867_ (
);

FILL FILL_2__12447_ (
);

FILL FILL_2__12027_ (
);

FILL FILL_0__13481_ (
);

FILL FILL_5__16253_ (
);

FILL FILL_0__8867_ (
);

FILL FILL_3__6964_ (
);

FILL FILL_0__8447_ (
);

DFFSR _10718_ (
    .Q(\datapath_1.regfile_1.regOut[30] [8]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_1888_[8])
);

FILL FILL_1__9090_ (
);

FILL SFILL28840x46050 (
);

FILL FILL_4__15666_ (
);

FILL FILL_4__15246_ (
);

FILL FILL_2__16280_ (
);

FILL FILL_4__10381_ (
);

FILL FILL_2__9406_ (
);

FILL FILL_3__14659_ (
);

FILL FILL_3__14239_ (
);

FILL FILL_1__15693_ (
);

FILL FILL_1__15273_ (
);

FILL SFILL33800x29050 (
);

FILL SFILL18920x82050 (
);

FILL FILL_5__7831_ (
);

OAI22X1 _14971_ (
    .A(_5451_),
    .B(_3931__bF$buf3),
    .C(_3966__bF$buf2),
    .D(_5450_),
    .Y(_5452_)
);

FILL FILL_0__14686_ (
);

INVX1 _14551_ (
    .A(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_5040_)
);

FILL FILL_0__14266_ (
);

INVX2 _14131_ (
    .A(_3936__bF$buf0),
    .Y(_4629_)
);

FILL FILL_3__15600_ (
);

FILL FILL_1__7823_ (
);

FILL FILL_3__7749_ (
);

FILL FILL_3__7329_ (
);

FILL FILL_5__12593_ (
);

FILL FILL_5__12173_ (
);

BUFX2 _6893_ (
    .A(_2_[23]),
    .Y(memoryWriteData[23])
);

FILL FILL_4__11586_ (
);

FILL FILL_4__11166_ (
);

FILL FILL_1__16058_ (
);

FILL FILL_3__10999_ (
);

FILL FILL_5__8616_ (
);

FILL FILL_3__10579_ (
);

FILL FILL_3__10159_ (
);

FILL FILL_1__11193_ (
);

OAI22X1 _15756_ (
    .A(_5489__bF$buf3),
    .B(_6218_),
    .C(_4771_),
    .D(_5504__bF$buf0),
    .Y(_6219_)
);

NAND3X1 _15336_ (
    .A(_5803_),
    .B(_5809_),
    .C(_5799_),
    .Y(_5810_)
);

INVX1 _10891_ (
    .A(_2019_),
    .Y(_2037_)
);

FILL FILL_0__10186_ (
);

DFFSR _10471_ (
    .Q(\datapath_1.regfile_1.regOut[28] [17]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_1758_[17])
);

FILL FILL_5__10906_ (
);

OAI21X1 _10051_ (
    .A(_1612_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1613_),
    .Y(_1563_[25])
);

FILL FILL_1__8608_ (
);

FILL FILL_3__11940_ (
);

FILL FILL_6__14385_ (
);

FILL FILL_3__11520_ (
);

FILL FILL_3__11100_ (
);

FILL FILL_0__16412_ (
);

FILL FILL_2__10933_ (
);

FILL FILL_5__13798_ (
);

FILL FILL_5__13378_ (
);

FILL FILL_2__10513_ (
);

OAI21X1 _7678_ (
    .A(_396_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .C(_397_),
    .Y(_393_[2])
);

DFFSR _7258_ (
    .Q(\datapath_1.regfile_1.regOut[3] [4]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_133_[4])
);

FILL FILL_4__9085_ (
);

FILL SFILL58120x57050 (
);

FILL FILL_0__6933_ (
);

FILL SFILL79080x55050 (
);

FILL FILL_1__12398_ (
);

FILL FILL_4__13732_ (
);

FILL SFILL54200x18050 (
);

FILL FILL_4__13312_ (
);

FILL FILL_3__7082_ (
);

NAND2X1 _11676_ (
    .A(_2165_),
    .B(_2757_),
    .Y(_2777_)
);

OAI21X1 _11256_ (
    .A(_2366_),
    .B(_2372_),
    .C(_2374_),
    .Y(_2375_)
);

FILL FILL_3__12725_ (
);

FILL FILL_3__12305_ (
);

FILL FILL_4__7818_ (
);

FILL FILL_2__11718_ (
);

FILL FILL_0__12752_ (
);

FILL FILL_3__15197_ (
);

FILL FILL_0__12332_ (
);

FILL SFILL38920x4050 (
);

FILL FILL_5__15944_ (
);

FILL SFILL38840x9050 (
);

FILL FILL_5__15524_ (
);

FILL FILL_0__7718_ (
);

FILL FILL_5__15104_ (
);

DFFSR _9824_ (
    .Q(\datapath_1.regfile_1.regOut[23] [10]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_1433_[10])
);

NAND2X1 _9404_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1284_)
);

FILL FILL_1__8781_ (
);

FILL FILL_1__8361_ (
);

FILL FILL_4__14937_ (
);

FILL SFILL79080x10050 (
);

FILL FILL_2__15971_ (
);

FILL FILL_4__14517_ (
);

FILL FILL_2__15551_ (
);

FILL FILL_2__15131_ (
);

FILL FILL_1__14964_ (
);

FILL FILL_1__14544_ (
);

FILL FILL_1__14124_ (
);

FILL FILL_0__13957_ (
);

INVX1 _13822_ (
    .A(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_4327_)
);

FILL FILL_0__13537_ (
);

INVX1 _13402_ (
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_3914_)
);

FILL FILL_0__13117_ (
);

FILL FILL_5__9994_ (
);

FILL SFILL109240x36050 (
);

FILL FILL_5__9154_ (
);

AOI22X1 _16294_ (
    .A(\datapath_1.regfile_1.regOut[31] [31]),
    .B(_5571_),
    .C(_5570__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_6743_)
);

FILL FILL_5__16309_ (
);

FILL FILL_1__9986_ (
);

FILL FILL_5__11864_ (
);

FILL FILL_5__11444_ (
);

FILL FILL_1__9146_ (
);

FILL FILL_5__11024_ (
);

FILL SFILL69080x53050 (
);

FILL FILL_4__7991_ (
);

FILL FILL_2__16336_ (
);

FILL FILL_4__7571_ (
);

FILL SFILL48920x38050 (
);

FILL FILL_4__10437_ (
);

FILL FILL_2__11891_ (
);

FILL FILL_4__10017_ (
);

FILL FILL_2__11471_ (
);

FILL FILL_2__11051_ (
);

FILL FILL_6__7497_ (
);

FILL FILL_1__15749_ (
);

FILL FILL_1__15329_ (
);

FILL FILL_1__10884_ (
);

FILL FILL_1__10044_ (
);

NAND3X1 _14607_ (
    .A(_5093_),
    .B(_5094_),
    .C(_5092_),
    .Y(_5095_)
);

FILL FILL_0__7891_ (
);

FILL FILL_0__7471_ (
);

FILL FILL_2__7489_ (
);

FILL FILL_0__7051_ (
);

FILL FILL_2__7069_ (
);

FILL FILL_4__14690_ (
);

FILL FILL_4__14270_ (
);

FILL FILL_5__12649_ (
);

FILL FILL_2__8850_ (
);

FILL FILL_3__13683_ (
);

FILL FILL_5__12229_ (
);

FILL FILL_3__13263_ (
);

OAI21X1 _6949_ (
    .A(_32_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .C(_33_),
    .Y(_3_[15])
);

FILL FILL_2__8010_ (
);

FILL FILL_4__8776_ (
);

FILL FILL_4__8356_ (
);

FILL FILL_2__12256_ (
);

FILL FILL_0__13290_ (
);

FILL FILL_1__11669_ (
);

FILL FILL_1__11249_ (
);

FILL SFILL3640x73050 (
);

FILL FILL_5__16062_ (
);

NOR2X1 _10947_ (
    .A(\control_1.op [0]),
    .B(\control_1.op [1]),
    .Y(_2080_)
);

FILL FILL_0__8256_ (
);

FILL FILL_6__9643_ (
);

OAI21X1 _10527_ (
    .A(_1848_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .C(_1849_),
    .Y(_1823_[13])
);

OAI21X1 _10107_ (
    .A(_1629_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .C(_1630_),
    .Y(_1628_[1])
);

FILL FILL_4__15895_ (
);

FILL FILL_1__12610_ (
);

FILL FILL_4__15475_ (
);

FILL FILL_4__15055_ (
);

FILL SFILL34600x28050 (
);

FILL FILL_4__10190_ (
);

FILL FILL_2__9635_ (
);

FILL FILL_3__14888_ (
);

FILL FILL_2__9215_ (
);

FILL FILL_3__14468_ (
);

FILL FILL_0__11603_ (
);

FILL FILL_3__14048_ (
);

FILL FILL_1__15082_ (
);

FILL FILL_6__15802_ (
);

FILL FILL_5__7220_ (
);

FILL SFILL59080x51050 (
);

FILL FILL_0__14495_ (
);

INVX1 _14780_ (
    .A(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_5265_)
);

FILL FILL_0__14075_ (
);

INVX1 _14360_ (
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_4853_)
);

FILL SFILL38920x36050 (
);

FILL FILL_1__7632_ (
);

FILL FILL_1__7212_ (
);

FILL SFILL99160x47050 (
);

FILL FILL_2__14822_ (
);

FILL FILL_2__14402_ (
);

FILL FILL_3__7978_ (
);

FILL FILL_3__7558_ (
);

FILL FILL_1__13815_ (
);

FILL FILL_4__11395_ (
);

FILL FILL_1__16287_ (
);

FILL FILL_5__8845_ (
);

FILL FILL_3__10388_ (
);

FILL FILL_5__8005_ (
);

NOR3X1 _15985_ (
    .A(_5515__bF$buf1),
    .B(_5051_),
    .C(_5521__bF$buf0),
    .Y(_6442_)
);

FILL FILL_6__11722_ (
);

NOR2X1 _15565_ (
    .A(_4566_),
    .B(_5539__bF$buf2),
    .Y(_6033_)
);

NOR3X1 _15145_ (
    .A(_5515__bF$buf2),
    .B(_4058_),
    .C(_5521__bF$buf1),
    .Y(_5623_)
);

OAI21X1 _10280_ (
    .A(_1724_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1725_),
    .Y(_1693_[16])
);

FILL FILL_1__8837_ (
);

FILL SFILL104440x52050 (
);

FILL FILL_2__15607_ (
);

FILL FILL_4__6842_ (
);

FILL FILL_0__16221_ (
);

FILL FILL_2__10742_ (
);

FILL FILL_2__10322_ (
);

NAND2X1 _7487_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_311_)
);

NAND2X1 _7067_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_92_)
);

FILL FILL_4__13961_ (
);

FILL FILL_4__13541_ (
);

FILL FILL_4__13121_ (
);

NOR2X1 _11485_ (
    .A(_2598_),
    .B(_2597_),
    .Y(_2599_)
);

NOR2X1 _11065_ (
    .A(_2182_),
    .B(_2183_),
    .Y(_2184_)
);

FILL FILL_3__12954_ (
);

FILL FILL_2__7701_ (
);

FILL FILL_3__12534_ (
);

FILL FILL_3__12114_ (
);

FILL SFILL28920x34050 (
);

FILL FILL_4__7627_ (
);

FILL FILL_4__7207_ (
);

FILL FILL_2__11947_ (
);

FILL FILL_0__12981_ (
);

FILL FILL_2__11527_ (
);

FILL FILL_2__11107_ (
);

FILL FILL_0__12141_ (
);

FILL SFILL28040x58050 (
);

FILL SFILL28520x20050 (
);

FILL FILL_5__15753_ (
);

FILL FILL_0__7947_ (
);

FILL FILL_5__15333_ (
);

NAND2X1 _9633_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1396_)
);

FILL FILL_0__7107_ (
);

NAND2X1 _9213_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1177_)
);

FILL FILL_1__8590_ (
);

FILL FILL_4__14746_ (
);

FILL FILL_2__15780_ (
);

FILL FILL_4__14326_ (
);

FILL FILL_2__15360_ (
);

FILL FILL_3__8096_ (
);

FILL FILL_2__8906_ (
);

FILL FILL_3__13739_ (
);

FILL FILL_3__13319_ (
);

FILL FILL_1__14773_ (
);

FILL FILL_1__14353_ (
);

FILL FILL_5__6911_ (
);

FILL FILL_0__13766_ (
);

FILL FILL_0__13346_ (
);

INVX1 _13631_ (
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_4140_)
);

INVX2 _13211_ (
    .A(_3753_),
    .Y(_3754_)
);

FILL FILL_5__9383_ (
);

FILL FILL_1__6903_ (
);

FILL SFILL90040x55050 (
);

FILL FILL_5__16118_ (
);

FILL FILL_1__9795_ (
);

FILL FILL_5__11673_ (
);

FILL FILL_5__11253_ (
);

FILL FILL_1__9375_ (
);

FILL FILL_2__16145_ (
);

FILL FILL_4__7380_ (
);

FILL SFILL63960x72050 (
);

FILL FILL_4__10666_ (
);

FILL SFILL94360x63050 (
);

FILL FILL_4__10246_ (
);

FILL FILL_2__11280_ (
);

FILL FILL_1__15978_ (
);

FILL FILL_1__15558_ (
);

FILL FILL_1__15138_ (
);

FILL FILL_2_BUFX2_insert300 (
);

FILL FILL_1__10693_ (
);

FILL FILL_2_BUFX2_insert301 (
);

FILL FILL_1__10273_ (
);

FILL FILL_2_BUFX2_insert302 (
);

FILL FILL_2_BUFX2_insert303 (
);

INVX1 _14836_ (
    .A(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_5319_)
);

FILL FILL_2_BUFX2_insert304 (
);

INVX1 _14416_ (
    .A(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_4908_)
);

FILL FILL_2_BUFX2_insert305 (
);

FILL FILL_2_BUFX2_insert306 (
);

FILL FILL_2__7298_ (
);

FILL FILL_2_BUFX2_insert307 (
);

FILL FILL_2_BUFX2_insert308 (
);

FILL FILL_2_BUFX2_insert309 (
);

FILL FILL_0__15912_ (
);

FILL FILL_5__12878_ (
);

FILL FILL_5__12458_ (
);

FILL FILL_5__12038_ (
);

FILL FILL_3__13492_ (
);

FILL FILL_4__8585_ (
);

FILL SFILL18680x4050 (
);

FILL FILL_2__12485_ (
);

FILL FILL_2__12065_ (
);

FILL FILL_2_BUFX2_insert1020 (
);

FILL FILL_2_BUFX2_insert1021 (
);

FILL FILL_2_BUFX2_insert1022 (
);

FILL FILL_1__11898_ (
);

FILL FILL_2_BUFX2_insert1023 (
);

FILL FILL_1__11478_ (
);

FILL FILL_2_BUFX2_insert1024 (
);

FILL FILL_1__11058_ (
);

FILL FILL_2_BUFX2_insert1025 (
);

FILL FILL_2_BUFX2_insert1026 (
);

FILL FILL_2_BUFX2_insert1027 (
);

FILL FILL_2_BUFX2_insert1028 (
);

FILL FILL_5__16291_ (
);

FILL FILL_2_BUFX2_insert1029 (
);

FILL FILL_0__8485_ (
);

FILL FILL_0__8065_ (
);

OAI21X1 _10756_ (
    .A(_1960_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .C(_1961_),
    .Y(_1953_[4])
);

FILL FILL_6__9032_ (
);

DFFSR _10336_ (
    .Q(\datapath_1.regfile_1.regOut[27] [10]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_1693_[10])
);

FILL FILL_3__11805_ (
);

FILL FILL_4__15284_ (
);

FILL SFILL8760x80050 (
);

FILL FILL_2__9864_ (
);

FILL FILL_3__14697_ (
);

FILL FILL_0__11832_ (
);

FILL FILL_3__14277_ (
);

FILL FILL_0__11412_ (
);

FILL FILL_2__9024_ (
);

FILL SFILL114600x80050 (
);

FILL FILL_5__14604_ (
);

FILL SFILL53960x70050 (
);

FILL SFILL84360x61050 (
);

NAND2X1 _8904_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1032_)
);

FILL FILL_1__7861_ (
);

FILL FILL_1__7441_ (
);

FILL FILL_2__14631_ (
);

FILL FILL_2__14211_ (
);

FILL FILL_3__7367_ (
);

FILL FILL_1__13624_ (
);

FILL FILL_4__16069_ (
);

FILL FILL_1_BUFX2_insert320 (
);

FILL FILL_1_BUFX2_insert321 (
);

FILL FILL_0__12617_ (
);

FILL FILL_1_BUFX2_insert322 (
);

NAND2X1 _12902_ (
    .A(vdd),
    .B(\datapath_1.rd1 [26]),
    .Y(_3607_)
);

FILL FILL_1_BUFX2_insert323 (
);

FILL FILL_1_BUFX2_insert324 (
);

FILL FILL_1__16096_ (
);

FILL FILL_1_BUFX2_insert325 (
);

FILL FILL_5__8654_ (
);

FILL FILL_1_BUFX2_insert326 (
);

FILL FILL_3__10197_ (
);

FILL FILL_5__8234_ (
);

FILL FILL_1_BUFX2_insert327 (
);

FILL FILL_1_BUFX2_insert328 (
);

FILL FILL_1_BUFX2_insert329 (
);

FILL FILL_6_BUFX2_insert884 (
);

NAND3X1 _15794_ (
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .B(_5471__bF$buf4),
    .C(_5531__bF$buf0),
    .Y(_6256_)
);

AOI22X1 _15374_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [8]),
    .C(\datapath_1.regfile_1.regOut[22] [8]),
    .D(_5650_),
    .Y(_5846_)
);

FILL FILL_0__15089_ (
);

FILL FILL_5__15809_ (
);

FILL FILL_3__16003_ (
);

FILL FILL_6_BUFX2_insert889 (
);

FILL FILL_5__10944_ (
);

FILL FILL_1__8646_ (
);

FILL FILL_5__10524_ (
);

FILL FILL_1__8226_ (
);

FILL FILL_5__10104_ (
);

FILL FILL_2__15836_ (
);

FILL FILL_2__15416_ (
);

FILL FILL_0__16450_ (
);

FILL FILL_0__16030_ (
);

FILL FILL_2__10971_ (
);

FILL FILL_2__10551_ (
);

FILL FILL_2__10131_ (
);

FILL FILL_1__14829_ (
);

NAND2X1 _7296_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_204_)
);

FILL FILL_1__14409_ (
);

FILL FILL_3__9933_ (
);

FILL FILL_3__9513_ (
);

FILL FILL_0__6971_ (
);

FILL FILL_2__6989_ (
);

FILL FILL_5__9859_ (
);

FILL SFILL114520x42050 (
);

FILL FILL_5__9019_ (
);

FILL FILL_4__13770_ (
);

FILL FILL_6__12316_ (
);

FILL FILL_4__13350_ (
);

INVX1 _16159_ (
    .A(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_6612_)
);

NAND2X1 _11294_ (
    .A(_2231_),
    .B(_2236_),
    .Y(_2413_)
);

FILL FILL_2__7930_ (
);

FILL FILL_5__11729_ (
);

FILL FILL_3__12763_ (
);

FILL FILL_5__11309_ (
);

FILL FILL_3__12343_ (
);

FILL FILL_4__7856_ (
);

FILL FILL_4__7436_ (
);

FILL FILL_2__11756_ (
);

FILL FILL_0__12790_ (
);

FILL FILL_2__11336_ (
);

FILL FILL_0__12370_ (
);

FILL FILL_1__10749_ (
);

FILL SFILL3640x68050 (
);

FILL FILL_5__15982_ (
);

FILL FILL_5__15562_ (
);

FILL FILL_0__7756_ (
);

FILL FILL_5__15142_ (
);

FILL FILL_0__7336_ (
);

NAND2X1 _9862_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1508_)
);

FILL FILL_6__8723_ (
);

DFFSR _9442_ (
    .Q(\datapath_1.regfile_1.regOut[20] [12]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_1238_[12])
);

INVX1 _9022_ (
    .A(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_1090_)
);

FILL SFILL43880x75050 (
);

FILL FILL_4__14975_ (
);

FILL FILL_4__14555_ (
);

FILL FILL_4__14135_ (
);

INVX1 _12499_ (
    .A(ALUOut[20]),
    .Y(_3399_)
);

NAND3X1 _12079_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[23]),
    .C(_3032__bF$buf4),
    .Y(_3105_)
);

FILL FILL_2__8715_ (
);

FILL FILL_3__13968_ (
);

FILL SFILL3560x6050 (
);

FILL FILL_3__13548_ (
);

FILL FILL_1__14582_ (
);

FILL FILL_3__13128_ (
);

FILL FILL_1__14162_ (
);

FILL FILL_0__13995_ (
);

OAI22X1 _13860_ (
    .A(_4363_),
    .B(_3936__bF$buf2),
    .C(_3954__bF$buf1),
    .D(_4362_),
    .Y(_4364_)
);

FILL FILL_0__13575_ (
);

INVX1 _13440_ (
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_3952_)
);

FILL FILL_0__13155_ (
);

INVX1 _13020_ (
    .A(_2_[23]),
    .Y(_3665_)
);

FILL FILL_2__13902_ (
);

FILL FILL_5__16347_ (
);

FILL FILL_6__9508_ (
);

FILL SFILL3640x23050 (
);

FILL FILL_5__11482_ (
);

FILL FILL_5__11062_ (
);

FILL FILL_2__16374_ (
);

FILL SFILL104520x40050 (
);

FILL SFILL43880x30050 (
);

FILL FILL_4__10895_ (
);

FILL FILL_0__9902_ (
);

FILL FILL_4__10055_ (
);

FILL FILL_1__15787_ (
);

FILL FILL_1__15367_ (
);

FILL FILL_5__7505_ (
);

NAND2X1 _14645_ (
    .A(_5125_),
    .B(_5132_),
    .Y(_5133_)
);

AOI22X1 _14225_ (
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .B(_3891__bF$buf3),
    .C(_4051__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_4721_)
);

FILL FILL_6__13694_ (
);

FILL SFILL104440x47050 (
);

FILL FILL_0__15721_ (
);

FILL FILL_0__15301_ (
);

FILL FILL_5__12267_ (
);

NAND2X1 _6987_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_59_)
);

FILL FILL_4__8394_ (
);

FILL SFILL33880x73050 (
);

FILL FILL_2__12294_ (
);

FILL FILL_1__11287_ (
);

FILL FILL_4__12621_ (
);

FILL FILL_4__12201_ (
);

DFFSR _10985_ (
    .Q(\control_1.reg_state.dout [1]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_2098_[1])
);

FILL SFILL49080x44050 (
);

NAND2X1 _10565_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1875_)
);

NAND2X1 _10145_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1656_)
);

FILL FILL_3__11614_ (
);

FILL FILL_4__15093_ (
);

FILL FILL_2__9673_ (
);

FILL FILL_2__9253_ (
);

FILL FILL_0__11641_ (
);

FILL FILL_0__11221_ (
);

FILL FILL_3__14086_ (
);

FILL FILL_4__9599_ (
);

FILL FILL_2__13499_ (
);

FILL FILL_2__13079_ (
);

FILL FILL_5__14833_ (
);

FILL FILL_5__14413_ (
);

NAND2X1 _8713_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_925_)
);

FILL FILL_1__7670_ (
);

FILL FILL_1__7250_ (
);

FILL FILL_4__13826_ (
);

FILL FILL_2__14860_ (
);

FILL FILL_4__13406_ (
);

FILL FILL_2__14440_ (
);

FILL FILL_2__14020_ (
);

FILL FILL_0__9499_ (
);

FILL FILL_3__7596_ (
);

FILL FILL_3__7176_ (
);

FILL FILL_0__9079_ (
);

FILL FILL_1__13853_ (
);

FILL FILL_1__13433_ (
);

FILL FILL_4__16298_ (
);

FILL FILL_1__13013_ (
);

FILL SFILL94440x51050 (
);

FILL FILL_0__12846_ (
);

NAND2X1 _12711_ (
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[5]),
    .Y(_3500_)
);

FILL FILL_0__12426_ (
);

FILL FILL_0__12006_ (
);

FILL FILL_5__8883_ (
);

FILL FILL_5__8463_ (
);

NOR2X1 _15183_ (
    .A(_5659_),
    .B(_5657_),
    .Y(_5660_)
);

FILL FILL_5__15618_ (
);

FILL FILL_3__16232_ (
);

INVX1 _9918_ (
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .Y(_1545_)
);

FILL FILL_5__10753_ (
);

FILL FILL_1__8875_ (
);

FILL FILL_1__8455_ (
);

FILL FILL_2__15645_ (
);

FILL FILL_2__15225_ (
);

FILL FILL_4__6880_ (
);

FILL SFILL94360x58050 (
);

FILL FILL_2__10780_ (
);

FILL FILL_2__10360_ (
);

FILL FILL_1__14638_ (
);

FILL FILL_1__14218_ (
);

FILL FILL_3__9742_ (
);

OAI22X1 _13916_ (
    .A(_3947__bF$buf0),
    .B(_4417_),
    .C(_3977__bF$buf0),
    .D(_4418_),
    .Y(_4419_)
);

FILL SFILL79160x38050 (
);

FILL FILL_5__9668_ (
);

FILL FILL_5__9248_ (
);

FILL FILL_6__12965_ (
);

NAND2X1 _16388_ (
    .A(gnd),
    .B(gnd),
    .Y(_6813_)
);

FILL SFILL39400x54050 (
);

FILL FILL_5__11958_ (
);

FILL FILL_3__12992_ (
);

FILL FILL_5__11538_ (
);

FILL FILL_3__12572_ (
);

FILL FILL_5__11118_ (
);

FILL FILL_3__12152_ (
);

FILL FILL_4__7245_ (
);

FILL FILL_2__11985_ (
);

FILL FILL_2__11565_ (
);

FILL FILL_2__11145_ (
);

FILL SFILL94360x13050 (
);

FILL FILL_1__10978_ (
);

FILL FILL_1__10558_ (
);

FILL FILL_1__10138_ (
);

FILL FILL_5__15791_ (
);

FILL FILL_5__15371_ (
);

FILL FILL_0__7985_ (
);

FILL FILL_0__7565_ (
);

INVX1 _9671_ (
    .A(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_1421_)
);

INVX1 _9251_ (
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_1202_)
);

FILL FILL_4__14784_ (
);

FILL FILL_4__14364_ (
);

FILL SFILL8760x75050 (
);

FILL FILL111720x49050 (
);

FILL FILL_0__10912_ (
);

FILL FILL_3__13777_ (
);

FILL FILL_2__8524_ (
);

FILL FILL_3__13357_ (
);

FILL FILL_2__8104_ (
);

FILL FILL_1__14391_ (
);

FILL FILL_0__13384_ (
);

FILL SFILL53960x65050 (
);

FILL SFILL29000x83050 (
);

FILL SFILL84360x56050 (
);

FILL FILL_1__6941_ (
);

FILL FILL_4__9811_ (
);

FILL FILL_2__13711_ (
);

FILL FILL_3__6867_ (
);

FILL FILL_5__16156_ (
);

FILL FILL_5__11291_ (
);

FILL FILL_4__15989_ (
);

FILL FILL_1__12704_ (
);

FILL FILL_4__15569_ (
);

FILL FILL_4__15149_ (
);

FILL FILL_2__16183_ (
);

FILL FILL_4__10284_ (
);

FILL FILL_2__9729_ (
);

FILL SFILL8760x30050 (
);

FILL FILL_1__15596_ (
);

FILL FILL_1__15176_ (
);

FILL FILL_5__7734_ (
);

FILL FILL_5__7314_ (
);

FILL FILL_0__14589_ (
);

INVX1 _14874_ (
    .A(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_5357_)
);

INVX1 _14454_ (
    .A(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_4945_)
);

FILL FILL_0__14169_ (
);

NOR2X1 _14034_ (
    .A(_4533_),
    .B(_3944__bF$buf0),
    .Y(_4534_)
);

FILL FILL_3__15923_ (
);

FILL FILL_3__15503_ (
);

FILL SFILL114600x30050 (
);

FILL FILL_1__7726_ (
);

FILL FILL_1__7306_ (
);

FILL SFILL84360x11050 (
);

FILL FILL_2__14916_ (
);

FILL FILL_0__15950_ (
);

FILL FILL_0__15530_ (
);

FILL FILL_0__15110_ (
);

FILL FILL_5__12496_ (
);

FILL FILL_5__12076_ (
);

FILL FILL_1__13909_ (
);

FILL FILL_4__11489_ (
);

FILL FILL_4__11069_ (
);

FILL SFILL114520x37050 (
);

FILL FILL_5__8519_ (
);

FILL FILL_1__11096_ (
);

AOI22X1 _15659_ (
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .B(_5693_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_6124_)
);

FILL FILL_4__12850_ (
);

FILL FILL_4__12430_ (
);

OAI22X1 _15239_ (
    .A(_5713_),
    .B(_5545__bF$buf2),
    .C(_5485__bF$buf3),
    .D(_5714_),
    .Y(_5715_)
);

FILL SFILL3720x56050 (
);

FILL FILL_4__12010_ (
);

NAND2X1 _10794_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1987_)
);

NAND2X1 _10374_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1768_)
);

FILL FILL_5__10809_ (
);

FILL FILL_3__11843_ (
);

FILL SFILL43960x63050 (
);

FILL FILL_6__14288_ (
);

FILL FILL_3__11423_ (
);

FILL SFILL74360x54050 (
);

FILL FILL_3__11003_ (
);

FILL FILL_4__6936_ (
);

FILL FILL_0__16315_ (
);

FILL FILL_2__10836_ (
);

FILL FILL_2__9482_ (
);

FILL FILL_0__11870_ (
);

FILL FILL_2__10416_ (
);

FILL FILL_0__11450_ (
);

FILL FILL_0__11030_ (
);

FILL FILL_5__14642_ (
);

FILL FILL_0__6836_ (
);

FILL FILL_5__14222_ (
);

DFFSR _8942_ (
    .Q(\datapath_1.regfile_1.regOut[16] [24]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_978_[24])
);

FILL FILL_6__7803_ (
);

INVX1 _8522_ (
    .A(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_838_)
);

INVX1 _8102_ (
    .A(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_619_)
);

FILL FILL_4__13635_ (
);

FILL FILL_4__13215_ (
);

NAND3X1 _11999_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[3]),
    .C(_3032__bF$buf0),
    .Y(_3045_)
);

NOR2X1 _11579_ (
    .A(_2686_),
    .B(_2680_),
    .Y(_2687_)
);

OAI21X1 _11159_ (
    .A(_2227_),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .C(_2277_),
    .Y(_2278_)
);

FILL SFILL3720x11050 (
);

FILL FILL_3__12628_ (
);

FILL FILL_1__13662_ (
);

FILL FILL_3__12208_ (
);

FILL FILL_1__13242_ (
);

FILL FILL112280x74050 (
);

FILL FILL_1_BUFX2_insert700 (
);

FILL FILL_1_BUFX2_insert701 (
);

FILL FILL_0__12655_ (
);

DFFSR _12940_ (
    .Q(\datapath_1.a [21]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3555_[21])
);

FILL FILL_1_BUFX2_insert702 (
);

FILL FILL_1_BUFX2_insert703 (
);

INVX1 _12520_ (
    .A(ALUOut[27]),
    .Y(_3413_)
);

FILL FILL_0__12235_ (
);

FILL FILL_1_BUFX2_insert704 (
);

NAND3X1 _12100_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [28]),
    .C(_3034__bF$buf2),
    .Y(_3121_)
);

FILL FILL_1_BUFX2_insert705 (
);

FILL FILL_1_BUFX2_insert706 (
);

FILL FILL_1_BUFX2_insert707 (
);

FILL FILL_5__8272_ (
);

FILL FILL_1_BUFX2_insert708 (
);

FILL FILL_1_BUFX2_insert709 (
);

FILL FILL_5__15847_ (
);

FILL FILL_5__15427_ (
);

FILL FILL_5__15007_ (
);

INVX1 _9727_ (
    .A(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_1438_)
);

FILL FILL_3__16041_ (
);

FILL SFILL3640x18050 (
);

FILL FILL_5__10982_ (
);

DFFSR _9307_ (
    .Q(\datapath_1.regfile_1.regOut[19] [5]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_1173_[5])
);

FILL FILL_5__10562_ (
);

FILL FILL_1__8264_ (
);

FILL FILL_5__10142_ (
);

FILL FILL_2__15874_ (
);

FILL SFILL104520x35050 (
);

FILL FILL_2__15454_ (
);

FILL FILL_2__15034_ (
);

FILL FILL_1__14867_ (
);

FILL FILL_1__14447_ (
);

FILL FILL_1__14027_ (
);

FILL SFILL59000x39050 (
);

FILL FILL_3__9551_ (
);

FILL FILL_3__9131_ (
);

OAI22X1 _13725_ (
    .A(_4231_),
    .B(_3949_),
    .C(_3881_),
    .D(_4230_),
    .Y(_4232_)
);

OAI21X1 _13305_ (
    .A(\datapath_1.a3 [0]),
    .B(_3791_),
    .C(_3839_),
    .Y(_3840_)
);

FILL FILL_5__9897_ (
);

FILL FILL_5__9477_ (
);

FILL FILL_6__12774_ (
);

INVX1 _16197_ (
    .A(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_6649_)
);

FILL FILL_0__14801_ (
);

FILL FILL_1__9889_ (
);

FILL FILL_5__11767_ (
);

FILL FILL_5__11347_ (
);

FILL FILL_1__9469_ (
);

FILL FILL_3__12381_ (
);

FILL FILL_2__16239_ (
);

FILL SFILL33880x68050 (
);

FILL FILL_4__7474_ (
);

FILL FILL_4__7054_ (
);

FILL FILL_2__11794_ (
);

FILL FILL_2__11374_ (
);

FILL FILL_1__10787_ (
);

FILL FILL_1__10367_ (
);

FILL FILL_4__11701_ (
);

FILL FILL_5__15180_ (
);

FILL FILL_0__7374_ (
);

INVX1 _9480_ (
    .A(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_1314_)
);

DFFSR _9060_ (
    .Q(\datapath_1.regfile_1.regOut[17] [14]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_1043_[14])
);

FILL FILL_4__14593_ (
);

FILL FILL_4__14173_ (
);

FILL FILL_2__8753_ (
);

FILL FILL_3__13586_ (
);

FILL FILL_2__8333_ (
);

FILL FILL_0__10301_ (
);

FILL FILL_3__13166_ (
);

FILL FILL_4__8259_ (
);

FILL FILL_2__12999_ (
);

FILL FILL_2__12579_ (
);

FILL FILL_2__12159_ (
);

FILL SFILL33880x23050 (
);

FILL FILL_5__13913_ (
);

FILL FILL_4__9620_ (
);

FILL FILL_4__12906_ (
);

FILL FILL_2__13940_ (
);

FILL FILL_0__8999_ (
);

FILL FILL_5__16385_ (
);

FILL FILL_2__13520_ (
);

FILL SFILL49000x37050 (
);

FILL SFILL104440x50 (
);

FILL FILL_0__8579_ (
);

FILL FILL_2__13100_ (
);

FILL FILL_6__9126_ (
);

FILL FILL_4__15798_ (
);

FILL FILL_4__15378_ (
);

FILL FILL_1__12513_ (
);

FILL SFILL94440x46050 (
);

FILL FILL_0__9940_ (
);

FILL FILL_0__11926_ (
);

FILL FILL_0__9520_ (
);

FILL FILL_2__9538_ (
);

FILL FILL_0__9100_ (
);

FILL FILL_0__11506_ (
);

FILL FILL_2__9118_ (
);

FILL FILL_6__15705_ (
);

FILL FILL_5__7963_ (
);

FILL FILL_5__7543_ (
);

FILL FILL_5__7123_ (
);

FILL FILL_0__14398_ (
);

OAI22X1 _14683_ (
    .A(_5169_),
    .B(_3949_),
    .C(_3978_),
    .D(_5168_),
    .Y(_5170_)
);

NAND3X1 _14263_ (
    .A(_4757_),
    .B(_4758_),
    .C(_4756_),
    .Y(_4759_)
);

FILL FILL_6__10000_ (
);

FILL SFILL23880x66050 (
);

FILL FILL_3__15732_ (
);

FILL FILL_3__15312_ (
);

FILL FILL_1__7955_ (
);

FILL FILL_1__7115_ (
);

FILL FILL_2__14725_ (
);

FILL FILL_2__14305_ (
);

FILL FILL_1__13718_ (
);

FILL FILL_4__11298_ (
);

FILL FILL_3__8822_ (
);

FILL FILL_3__8402_ (
);

FILL FILL_5__8748_ (
);

FILL FILL_5__8328_ (
);

NOR2X1 _15888_ (
    .A(_6344_),
    .B(_6347_),
    .Y(_6348_)
);

FILL FILL_6__11625_ (
);

FILL FILL_6__11205_ (
);

AOI22X1 _15468_ (
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [10]),
    .C(\datapath_1.regfile_1.regOut[5] [10]),
    .D(_5700_),
    .Y(_5938_)
);

FILL SFILL23800x64050 (
);

OAI22X1 _15048_ (
    .A(_5526__bF$buf3),
    .B(_3970_),
    .C(_3934_),
    .D(_5527__bF$buf4),
    .Y(_5528_)
);

INVX1 _10183_ (
    .A(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_1681_)
);

FILL FILL_5__10618_ (
);

FILL SFILL23880x21050 (
);

FILL FILL_3__11652_ (
);

FILL FILL_3__11232_ (
);

FILL FILL_0__16124_ (
);

FILL FILL_2__10645_ (
);

FILL FILL_2__9291_ (
);

FILL SFILL23400x50050 (
);

FILL FILL112360x3050 (
);

FILL FILL_3_BUFX2_insert230 (
);

FILL FILL_3__9607_ (
);

FILL FILL_3_BUFX2_insert231 (
);

FILL FILL_5__14871_ (
);

FILL FILL_3_BUFX2_insert232 (
);

FILL FILL_5__14451_ (
);

FILL FILL_3_BUFX2_insert233 (
);

FILL FILL_5__14031_ (
);

FILL FILL_3_BUFX2_insert234 (
);

INVX1 _8751_ (
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_950_)
);

FILL FILL_3_BUFX2_insert235 (
);

INVX1 _8331_ (
    .A(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_731_)
);

FILL FILL_3_BUFX2_insert236 (
);

FILL FILL_3_BUFX2_insert237 (
);

FILL FILL_3_BUFX2_insert238 (
);

FILL FILL_4__13864_ (
);

FILL FILL_3_BUFX2_insert239 (
);

FILL FILL_4__13444_ (
);

FILL FILL_4__13024_ (
);

NOR2X1 _11388_ (
    .A(_2504_),
    .B(_2193_),
    .Y(_2505_)
);

FILL FILL_3__12857_ (
);

FILL FILL_2__7604_ (
);

FILL FILL_3__12437_ (
);

FILL FILL_1__13891_ (
);

FILL FILL_3__12017_ (
);

FILL FILL_1__13471_ (
);

FILL FILL_0__12884_ (
);

FILL FILL_0__12464_ (
);

FILL FILL_0__12044_ (
);

FILL FILL_5__8081_ (
);

FILL FILL_5__15656_ (
);

FILL FILL_5__15236_ (
);

DFFSR _9956_ (
    .Q(\datapath_1.regfile_1.regOut[24] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_1498_[14])
);

FILL FILL_3__16270_ (
);

OAI21X1 _9536_ (
    .A(_1350_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1351_),
    .Y(_1303_[24])
);

FILL FILL_5__10791_ (
);

OAI21X1 _9116_ (
    .A(_1131_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .C(_1132_),
    .Y(_1108_[12])
);

FILL FILL_5__10371_ (
);

FILL FILL_1__8493_ (
);

FILL FILL_1__8073_ (
);

FILL FILL_4__14649_ (
);

FILL FILL_4__14229_ (
);

FILL FILL_2__15683_ (
);

FILL FILL_2__15263_ (
);

FILL SFILL8760x25050 (
);

FILL SFILL13800x62050 (
);

FILL FILL_1__14676_ (
);

FILL FILL_1__14256_ (
);

FILL FILL_0_BUFX2_insert360 (
);

FILL SFILL74040x73050 (
);

FILL FILL_0_BUFX2_insert361 (
);

FILL FILL_0_BUFX2_insert362 (
);

FILL FILL_3__9780_ (
);

FILL FILL_0_BUFX2_insert363 (
);

FILL FILL_3__9360_ (
);

FILL FILL_0__13669_ (
);

FILL FILL_0_BUFX2_insert364 (
);

INVX1 _13954_ (
    .A(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_4456_)
);

FILL FILL_0__13249_ (
);

FILL FILL_0_BUFX2_insert365 (
);

INVX1 _13534_ (
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_4044_)
);

OAI21X1 _13114_ (
    .A(_3706_),
    .B(PCEn_bF$buf2),
    .C(_3707_),
    .Y(_3685_[11])
);

FILL FILL_0_BUFX2_insert366 (
);

FILL FILL_0_BUFX2_insert367 (
);

FILL FILL_0_BUFX2_insert368 (
);

FILL FILL_0_BUFX2_insert369 (
);

FILL FILL_5__9286_ (
);

FILL SFILL114600x25050 (
);

FILL SFILL53960x15050 (
);

FILL FILL_6__12583_ (
);

FILL FILL_0__14610_ (
);

FILL FILL_5__11996_ (
);

FILL FILL_5__11576_ (
);

FILL FILL_1__9278_ (
);

FILL FILL_5__11156_ (
);

FILL FILL_3__12190_ (
);

FILL FILL_2__16048_ (
);

FILL FILL_4__10989_ (
);

FILL FILL_4__10569_ (
);

FILL FILL_4__10149_ (
);

FILL FILL_2__11183_ (
);

FILL FILL_1__10176_ (
);

FILL FILL_4__11930_ (
);

AOI22X1 _14739_ (
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .B(_4135_),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_5225_)
);

INVX1 _14319_ (
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_4813_)
);

FILL FILL_4__11510_ (
);

FILL FILL_0__7183_ (
);

FILL FILL_2_BUFX2_insert40 (
);

FILL FILL_2_BUFX2_insert41 (
);

FILL FILL_1__16402_ (
);

FILL FILL_2_BUFX2_insert42 (
);

FILL SFILL43960x58050 (
);

FILL FILL_3__10923_ (
);

FILL FILL_2_BUFX2_insert43 (
);

FILL FILL_2_BUFX2_insert44 (
);

FILL FILL_3__10503_ (
);

FILL FILL_2_BUFX2_insert45 (
);

FILL FILL_2_BUFX2_insert46 (
);

FILL FILL_0__15815_ (
);

FILL FILL_2_BUFX2_insert47 (
);

FILL FILL_2_BUFX2_insert48 (
);

FILL FILL_2_BUFX2_insert49 (
);

FILL FILL_2__8982_ (
);

FILL FILL_0__10950_ (
);

FILL FILL_2__8142_ (
);

FILL FILL_0__10530_ (
);

FILL FILL_3__13395_ (
);

FILL FILL_0__10110_ (
);

FILL FILL_4__8488_ (
);

FILL FILL_4__8068_ (
);

FILL FILL112360x62050 (
);

FILL FILL_2__12388_ (
);

FILL FILL_5__13722_ (
);

FILL FILL_5__13302_ (
);

FILL FILL_0_CLKBUF1_insert1080 (
);

FILL FILL_0_CLKBUF1_insert1081 (
);

FILL FILL_0_CLKBUF1_insert1082 (
);

INVX1 _7602_ (
    .A(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_367_)
);

FILL FILL_0_CLKBUF1_insert1083 (
);

FILL FILL_4__12715_ (
);

FILL SFILL64040x71050 (
);

FILL FILL_5__16194_ (
);

FILL FILL_0__8388_ (
);

INVX1 _10659_ (
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_1917_)
);

INVX1 _10239_ (
    .A(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_1698_)
);

FILL FILL_3__11708_ (
);

FILL FILL_1__12742_ (
);

FILL FILL_4__15187_ (
);

FILL FILL_1__12322_ (
);

FILL SFILL43960x13050 (
);

FILL FILL112280x69050 (
);

FILL FILL_2__9767_ (
);

FILL FILL_2__9347_ (
);

FILL FILL_0__11735_ (
);

NAND3X1 _11600_ (
    .A(_2696_),
    .B(_2699_),
    .C(_2706_),
    .Y(\datapath_1.ALUResult [19])
);

FILL FILL_0__11315_ (
);

FILL FILL_5__7352_ (
);

INVX1 _14492_ (
    .A(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_4983_)
);

NOR2X1 _14072_ (
    .A(_4568_),
    .B(_4571_),
    .Y(_4572_)
);

FILL FILL_5__14927_ (
);

FILL FILL_5__14507_ (
);

FILL FILL_3__15961_ (
);

FILL FILL_3__15541_ (
);

DFFSR _8807_ (
    .Q(\datapath_1.regfile_1.regOut[15] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_913_[17])
);

FILL FILL_3__15121_ (
);

FILL FILL_1__7764_ (
);

FILL FILL_1__7344_ (
);

FILL FILL_2__14954_ (
);

FILL FILL_2__14534_ (
);

FILL FILL_2__14114_ (
);

FILL FILL_1__13947_ (
);

FILL FILL_1__13527_ (
);

FILL FILL_1__13107_ (
);

FILL SFILL84360x2050 (
);

FILL FILL_3__8631_ (
);

DFFSR _12805_ (
    .Q(\datapath_1.PCJump [16]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[14])
);

FILL FILL_3__8211_ (
);

FILL FILL_5__8977_ (
);

FILL FILL_5__8137_ (
);

NAND3X1 _15697_ (
    .A(_6159_),
    .B(_6160_),
    .C(_6158_),
    .Y(_6161_)
);

NAND3X1 _15277_ (
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf1),
    .Y(_5752_)
);

FILL FILL_3__16326_ (
);

FILL FILL_1__8969_ (
);

FILL FILL_5__10427_ (
);

FILL FILL_3__11881_ (
);

FILL FILL_5__10007_ (
);

FILL FILL_3__11461_ (
);

FILL FILL_1__8129_ (
);

FILL FILL_3__11041_ (
);

FILL FILL_2__15739_ (
);

FILL FILL_4__6974_ (
);

FILL FILL_2__15319_ (
);

FILL FILL_0__16353_ (
);

FILL FILL_2__10874_ (
);

FILL FILL_2__10034_ (
);

FILL FILL_1__9910_ (
);

OAI21X1 _7199_ (
    .A(_158_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_159_),
    .Y(_133_[13])
);

FILL FILL_3__9416_ (
);

FILL FILL_5__14680_ (
);

FILL FILL_5__14260_ (
);

FILL FILL_0__6874_ (
);

INVX1 _8980_ (
    .A(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_1062_)
);

DFFSR _8560_ (
    .Q(\datapath_1.regfile_1.regOut[13] [26]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_783_[26])
);

FILL FILL_6__7421_ (
);

OAI21X1 _8140_ (
    .A(_643_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_644_),
    .Y(_588_[28])
);

FILL FILL_6__12639_ (
);

FILL FILL_4__13673_ (
);

FILL FILL_4__13253_ (
);

NOR2X1 _11197_ (
    .A(_2315_),
    .B(_2310_),
    .Y(_2316_)
);

FILL FILL_2__7833_ (
);

FILL FILL_3__12246_ (
);

FILL FILL_1__13280_ (
);

FILL FILL_4__7759_ (
);

FILL FILL_4__7339_ (
);

FILL FILL_2__11659_ (
);

FILL FILL_2__11239_ (
);

FILL SFILL33880x18050 (
);

FILL FILL_0__12273_ (
);

FILL FILL_4__8700_ (
);

FILL FILL_5__15885_ (
);

FILL FILL_2__12600_ (
);

FILL FILL_5__15465_ (
);

FILL FILL_5__15045_ (
);

OAI21X1 _9765_ (
    .A(_1462_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .C(_1463_),
    .Y(_1433_[15])
);

FILL FILL_0__7239_ (
);

FILL FILL_6__8206_ (
);

OAI21X1 _9345_ (
    .A(_1243_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .C(_1244_),
    .Y(_1238_[3])
);

FILL FILL_5__10180_ (
);

FILL FILL_4__14878_ (
);

FILL FILL_4__14458_ (
);

FILL FILL_4__14038_ (
);

FILL FILL_2__15492_ (
);

FILL FILL_2__15072_ (
);

FILL FILL_0__8600_ (
);

FILL FILL_2__8618_ (
);

FILL FILL_1__14485_ (
);

FILL FILL_1__14065_ (
);

FILL FILL_0__13898_ (
);

NOR2X1 _13763_ (
    .A(_4268_),
    .B(_3959_),
    .Y(_4269_)
);

FILL FILL_0__13478_ (
);

NOR2X1 _13343_ (
    .A(_3862_),
    .B(_3863_),
    .Y(_3864_)
);

FILL FILL_3__14812_ (
);

FILL FILL_5__9095_ (
);

FILL SFILL79160x80050 (
);

FILL FILL_4__9905_ (
);

FILL FILL_6__12392_ (
);

FILL FILL_2__13805_ (
);

FILL FILL_5__11385_ (
);

FILL FILL_1__9087_ (
);

FILL FILL_2__16277_ (
);

FILL FILL_4__10798_ (
);

FILL FILL_4__7092_ (
);

FILL FILL_4__10378_ (
);

FILL FILL_0__9805_ (
);

FILL FILL_5__7828_ (
);

AOI21X1 _14968_ (
    .A(\datapath_1.regfile_1.regOut[24] [31]),
    .B(_4079__bF$buf0),
    .C(_5448_),
    .Y(_5449_)
);

NOR2X1 _14548_ (
    .A(_5027_),
    .B(_5037_),
    .Y(_5038_)
);

OAI22X1 _14128_ (
    .A(_4625_),
    .B(_3972__bF$buf1),
    .C(_3920_),
    .D(_4624_),
    .Y(_4626_)
);

FILL SFILL84520x32050 (
);

FILL FILL_1__16211_ (
);

FILL SFILL23880x16050 (
);

FILL FILL_6__13597_ (
);

FILL FILL_3__10312_ (
);

FILL FILL_0__15624_ (
);

FILL SFILL53960x9050 (
);

FILL FILL_0__15204_ (
);

FILL FILL_2__8371_ (
);

FILL SFILL105000x53050 (
);

FILL FILL_2__12197_ (
);

FILL FILL_5__13951_ (
);

FILL FILL_5__13531_ (
);

FILL FILL_5__13111_ (
);

INVX1 _7831_ (
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_479_)
);

DFFSR _7411_ (
    .Q(\datapath_1.regfile_1.regOut[4] [29]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_198_[29])
);

FILL FILL_4__12524_ (
);

FILL FILL_4__12104_ (
);

AOI21X1 _10888_ (
    .A(_2027_),
    .B(_2033_),
    .C(_2026_),
    .Y(_2035_)
);

FILL FILL_0__8197_ (
);

DFFSR _10468_ (
    .Q(\datapath_1.regfile_1.regOut[28] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_1758_[14])
);

OAI21X1 _10048_ (
    .A(_1610_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .C(_1611_),
    .Y(_1563_[24])
);

FILL FILL_3__11937_ (
);

FILL FILL_1__12971_ (
);

FILL FILL_3__11517_ (
);

FILL FILL_1__12131_ (
);

FILL FILL_0__16409_ (
);

FILL FILL_2__9996_ (
);

FILL FILL_0__11964_ (
);

FILL FILL_2__9156_ (
);

FILL FILL_0__11544_ (
);

FILL FILL_0__11124_ (
);

FILL FILL_5__7581_ (
);

FILL FILL_5__7161_ (
);

FILL SFILL74120x61050 (
);

FILL FILL_5__14736_ (
);

FILL FILL_5__14316_ (
);

FILL FILL_3__15770_ (
);

FILL FILL_3__15350_ (
);

OAI21X1 _8616_ (
    .A(_879_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .C(_880_),
    .Y(_848_[16])
);

FILL FILL_1__7993_ (
);

FILL FILL_1__7573_ (
);

FILL FILL_4__13729_ (
);

FILL FILL_4__13309_ (
);

FILL FILL_2__14763_ (
);

FILL FILL_2__14343_ (
);

FILL FILL_3__7499_ (
);

FILL FILL_3__7079_ (
);

FILL SFILL13800x57050 (
);

FILL FILL_1__13756_ (
);

FILL FILL_1__13336_ (
);

FILL FILL_3__8860_ (
);

FILL FILL_0__12749_ (
);

FILL FILL_3__8440_ (
);

OAI21X1 _12614_ (
    .A(_3454_),
    .B(vdd),
    .C(_3455_),
    .Y(_3425_[15])
);

FILL FILL_3__8020_ (
);

FILL FILL_0__12329_ (
);

FILL FILL_5__8786_ (
);

FILL FILL_5__8366_ (
);

INVX8 _15086_ (
    .A(_5523_),
    .Y(_5565_)
);

FILL FILL_3__16135_ (
);

FILL FILL_5__10656_ (
);

FILL FILL_1__8778_ (
);

FILL FILL_1__8358_ (
);

FILL FILL_3__11690_ (
);

FILL FILL_5__10236_ (
);

FILL FILL_3__11270_ (
);

FILL FILL_2__15968_ (
);

FILL FILL_2__15548_ (
);

FILL FILL_2__15128_ (
);

FILL FILL_0__16162_ (
);

FILL FILL_2__10683_ (
);

FILL FILL_2__10263_ (
);

FILL SFILL13800x12050 (
);

FILL FILL_3_BUFX2_insert610 (
);

FILL FILL_3__9645_ (
);

INVX1 _13819_ (
    .A(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_4324_)
);

FILL FILL_3__9225_ (
);

FILL FILL_3_BUFX2_insert611 (
);

FILL FILL_3_BUFX2_insert612 (
);

FILL FILL_3_BUFX2_insert613 (
);

FILL FILL_3_BUFX2_insert614 (
);

FILL FILL_1__15902_ (
);

FILL FILL_3_BUFX2_insert615 (
);

FILL FILL_3_BUFX2_insert616 (
);

FILL FILL_3_BUFX2_insert617 (
);

FILL FILL_3_BUFX2_insert618 (
);

FILL FILL_3_BUFX2_insert619 (
);

FILL FILL_4__13482_ (
);

FILL FILL_3__12895_ (
);

FILL FILL_2__7222_ (
);

FILL FILL_3__12475_ (
);

FILL FILL_3__12055_ (
);

FILL FILL_4__7988_ (
);

FILL FILL_4__7568_ (
);

FILL FILL112360x57050 (
);

FILL FILL_2__11888_ (
);

FILL FILL_2__11468_ (
);

FILL FILL_2__11048_ (
);

FILL FILL_0__12082_ (
);

FILL SFILL49000x1050 (
);

FILL SFILL64040x66050 (
);

FILL FILL_5__15694_ (
);

FILL FILL_0__7888_ (
);

FILL FILL_5__15274_ (
);

OAI21X1 _9994_ (
    .A(_1574_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .C(_1575_),
    .Y(_1563_[6])
);

FILL FILL_0__7468_ (
);

DFFSR _9574_ (
    .Q(\datapath_1.regfile_1.regOut[21] [16]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_1303_[16])
);

FILL FILL_0__7048_ (
);

NAND2X1 _9154_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1158_)
);

FILL SFILL23640x2050 (
);

FILL FILL_1__11822_ (
);

FILL FILL_4__14687_ (
);

FILL FILL_4__14267_ (
);

FILL FILL_1__11402_ (
);

FILL FILL_2__8847_ (
);

FILL FILL_0__10815_ (
);

FILL FILL_2__8007_ (
);

FILL FILL_1__14294_ (
);

FILL FILL_5__6852_ (
);

FILL FILL_0_BUFX2_insert740 (
);

FILL FILL_0_BUFX2_insert741 (
);

FILL FILL_0_BUFX2_insert742 (
);

FILL FILL_0_BUFX2_insert743 (
);

OAI22X1 _13992_ (
    .A(_4492_),
    .B(_3936__bF$buf0),
    .C(_3955__bF$buf0),
    .D(_4491_),
    .Y(_4493_)
);

FILL FILL_0_BUFX2_insert744 (
);

FILL FILL_0__13287_ (
);

FILL FILL_0_BUFX2_insert745 (
);

INVX1 _13572_ (
    .A(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_4082_)
);

NAND2X1 _13152_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_pcsrc.dout [24]),
    .Y(_3733_)
);

FILL FILL_0_BUFX2_insert746 (
);

FILL FILL_0_BUFX2_insert747 (
);

FILL FILL112360x12050 (
);

FILL FILL_3__14621_ (
);

FILL FILL_0_BUFX2_insert748 (
);

FILL FILL_0_BUFX2_insert749 (
);

FILL FILL_3__14201_ (
);

FILL FILL_1__6844_ (
);

FILL FILL_2__13614_ (
);

FILL FILL_5__16059_ (
);

FILL SFILL64040x21050 (
);

FILL FILL_5__11194_ (
);

FILL FILL_1__12607_ (
);

FILL FILL_2__16086_ (
);

FILL FILL_4__10187_ (
);

FILL FILL_0__9614_ (
);

FILL FILL_3__7711_ (
);

FILL SFILL89240x70050 (
);

FILL FILL112280x19050 (
);

FILL FILL_1__15499_ (
);

FILL FILL_1__15079_ (
);

FILL FILL_5__7637_ (
);

FILL FILL_5__7217_ (
);

FILL FILL_4__16413_ (
);

INVX1 _14777_ (
    .A(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_5262_)
);

AOI21X1 _14357_ (
    .A(_4827_),
    .B(_4850_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [18])
);

FILL FILL_3__15826_ (
);

FILL FILL_3__15406_ (
);

FILL FILL_1__16020_ (
);

FILL FILL_3__10961_ (
);

FILL FILL_1__7629_ (
);

FILL FILL_3__10541_ (
);

FILL FILL_1__7209_ (
);

FILL FILL_3__10121_ (
);

FILL FILL_2__14819_ (
);

FILL FILL_0__15853_ (
);

FILL FILL_0__15433_ (
);

FILL FILL_0__15013_ (
);

FILL FILL_5__12399_ (
);

FILL SFILL54040x64050 (
);

FILL FILL_3__8916_ (
);

FILL FILL_5__13760_ (
);

FILL FILL_5__13340_ (
);

DFFSR _7640_ (
    .Q(\datapath_1.regfile_1.regOut[6] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_328_[2])
);

OAI21X1 _7220_ (
    .A(_172_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_173_),
    .Y(_133_[20])
);

FILL FILL_4__12753_ (
);

FILL FILL_4__12333_ (
);

OAI21X1 _10697_ (
    .A(_1941_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1942_),
    .Y(_1888_[27])
);

OAI21X1 _10277_ (
    .A(_1722_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1723_),
    .Y(_1693_[15])
);

FILL FILL_2__6913_ (
);

FILL FILL_3__11746_ (
);

FILL FILL_1__12780_ (
);

FILL FILL_3__11326_ (
);

FILL FILL_1__12360_ (
);

FILL FILL_4__6839_ (
);

FILL FILL_0__16218_ (
);

FILL FILL_2__10319_ (
);

FILL FILL_0__11773_ (
);

FILL FILL_2__9385_ (
);

FILL FILL_0__11353_ (
);

FILL FILL_6__15552_ (
);

FILL FILL_6__15132_ (
);

FILL FILL_5__14965_ (
);

FILL FILL_5__14545_ (
);

FILL FILL_5__14125_ (
);

OAI21X1 _8845_ (
    .A(_991_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_992_),
    .Y(_978_[7])
);

DFFSR _8425_ (
    .Q(\datapath_1.regfile_1.regOut[12] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_718_[19])
);

NAND2X1 _8005_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_575_)
);

FILL FILL_4__13958_ (
);

FILL FILL_2__14992_ (
);

FILL FILL_4__13538_ (
);

FILL FILL_2__14572_ (
);

FILL FILL_4__13118_ (
);

FILL FILL_2__14152_ (
);

FILL FILL_1__13985_ (
);

FILL FILL_1__13565_ (
);

FILL FILL_1__13145_ (
);

FILL SFILL58920x1050 (
);

FILL FILL_0__12978_ (
);

FILL SFILL59160x3050 (
);

OAI21X1 _12843_ (
    .A(_3566_),
    .B(vdd),
    .C(_3567_),
    .Y(_3555_[6])
);

FILL FILL_0__12138_ (
);

OAI21X1 _12423_ (
    .A(_3346_),
    .B(MemToReg_bF$buf6),
    .C(_3347_),
    .Y(\datapath_1.mux_wd3.dout [26])
);

NAND3X1 _12003_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[4]),
    .C(_3032__bF$buf2),
    .Y(_3048_)
);

FILL FILL_5__8595_ (
);

FILL SFILL79160x75050 (
);

FILL SFILL59080x8050 (
);

FILL SFILL44040x62050 (
);

FILL SFILL58280x34050 (
);

FILL FILL_6__11052_ (
);

FILL FILL_3__16364_ (
);

FILL FILL_5__10885_ (
);

FILL FILL_1__8587_ (
);

FILL FILL_5__10045_ (
);

FILL FILL_2__15777_ (
);

FILL FILL_2__15357_ (
);

FILL FILL_0__16391_ (
);

FILL FILL_2__10492_ (
);

FILL FILL_5__6908_ (
);

FILL FILL_3__9874_ (
);

INVX1 _13628_ (
    .A(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_4137_)
);

FILL FILL_3__9034_ (
);

FILL SFILL109480x9050 (
);

INVX2 _13208_ (
    .A(\datapath_1.a3 [0]),
    .Y(_3751_)
);

FILL FILL_1__15711_ (
);

FILL FILL_4__13291_ (
);

FILL FILL_0__14704_ (
);

FILL FILL_2__7871_ (
);

FILL FILL_2__7451_ (
);

FILL FILL_2__7031_ (
);

FILL FILL_3__12284_ (
);

FILL FILL_4__7377_ (
);

FILL FILL_2__11697_ (
);

FILL FILL_2__11277_ (
);

FILL SFILL8440x39050 (
);

FILL FILL_5__12611_ (
);

INVX1 _6911_ (
    .A(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_8_)
);

FILL FILL_2_BUFX2_insert270 (
);

FILL FILL_2_BUFX2_insert271 (
);

FILL FILL_2_BUFX2_insert272 (
);

FILL FILL_2_BUFX2_insert273 (
);

FILL FILL_2_BUFX2_insert274 (
);

FILL FILL_4__11604_ (
);

FILL FILL_2_BUFX2_insert275 (
);

FILL FILL_5__15083_ (
);

FILL FILL_0__7697_ (
);

FILL FILL_2_BUFX2_insert276 (
);

FILL FILL_2_BUFX2_insert277 (
);

NAND2X1 _9383_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1270_)
);

FILL FILL_2_BUFX2_insert278 (
);

FILL FILL_2_BUFX2_insert279 (
);

FILL FILL_4__14496_ (
);

FILL FILL_1__11631_ (
);

FILL FILL_1__11211_ (
);

FILL FILL_4__14076_ (
);

FILL SFILL69160x73050 (
);

FILL FILL_0__15909_ (
);

FILL FILL_2__8656_ (
);

FILL FILL_0__10624_ (
);

FILL FILL_2__8236_ (
);

FILL FILL_3__13489_ (
);

NAND3X1 _13381_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3892_),
    .C(_3880_),
    .Y(_3893_)
);

FILL FILL_0__13096_ (
);

FILL FILL_5__13816_ (
);

FILL FILL_3__14850_ (
);

FILL FILL_3__14430_ (
);

FILL FILL_3__14010_ (
);

FILL FILL_4__9523_ (
);

FILL FILL_4__9103_ (
);

FILL FILL_2__13843_ (
);

FILL FILL_2__13423_ (
);

FILL FILL_5__16288_ (
);

FILL SFILL109320x11050 (
);

FILL FILL_2__13003_ (
);

FILL FILL_1__12836_ (
);

FILL FILL_1__12416_ (
);

FILL FILL_3__7940_ (
);

FILL FILL_0__9423_ (
);

FILL FILL_0__11829_ (
);

FILL FILL_3__7100_ (
);

FILL FILL_0__9003_ (
);

FILL FILL_0__11409_ (
);

FILL FILL_5__7866_ (
);

FILL FILL_6__15608_ (
);

FILL FILL_5__7446_ (
);

FILL FILL_4__16222_ (
);

OAI22X1 _14586_ (
    .A(_3881_),
    .B(_5073_),
    .C(_3971__bF$buf1),
    .D(_5074_),
    .Y(_5075_)
);

INVX1 _14166_ (
    .A(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_4664_)
);

FILL SFILL74120x11050 (
);

FILL FILL_3__15635_ (
);

FILL FILL_3__15215_ (
);

FILL FILL_1__7858_ (
);

FILL FILL_1__7438_ (
);

FILL FILL_3__10770_ (
);

FILL SFILL28840x5050 (
);

FILL FILL_2__14628_ (
);

FILL FILL_0__15662_ (
);

FILL FILL_2__14208_ (
);

FILL SFILL99320x60050 (
);

FILL FILL_0__15242_ (
);

FILL FILL_1_BUFX2_insert290 (
);

FILL SFILL73960x50 (
);

FILL FILL_1_BUFX2_insert291 (
);

FILL FILL_3__8725_ (
);

FILL SFILL28760x80050 (
);

FILL SFILL74040x18050 (
);

FILL FILL_1_BUFX2_insert292 (
);

FILL FILL_1_BUFX2_insert293 (
);

FILL FILL_1_BUFX2_insert294 (
);

FILL FILL_1_BUFX2_insert295 (
);

FILL FILL_1_BUFX2_insert296 (
);

FILL SFILL8680x6050 (
);

FILL FILL_1_BUFX2_insert297 (
);

FILL FILL_1_BUFX2_insert298 (
);

FILL FILL_1_BUFX2_insert299 (
);

FILL FILL_4__12982_ (
);

FILL FILL_6__11528_ (
);

FILL FILL_6__11108_ (
);

FILL FILL_4__12142_ (
);

FILL SFILL64120x54050 (
);

DFFSR _10086_ (
    .Q(\datapath_1.regfile_1.regOut[25] [16]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_1563_[16])
);

FILL FILL_3__11975_ (
);

FILL FILL_3__11555_ (
);

FILL FILL_3__11135_ (
);

FILL FILL_0__16027_ (
);

NOR2X1 _16312_ (
    .A(_6760_),
    .B(_6758_),
    .Y(_6761_)
);

FILL FILL_2__10968_ (
);

FILL FILL_2__10548_ (
);

FILL FILL_2__10128_ (
);

FILL FILL_0__11582_ (
);

FILL FILL_0__11162_ (
);

FILL SFILL99640x36050 (
);

FILL FILL_5__14774_ (
);

FILL FILL_0__6968_ (
);

FILL FILL_5__14354_ (
);

NAND2X1 _8654_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_906_)
);

NAND2X1 _8234_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_687_)
);

FILL FILL_1__7191_ (
);

FILL FILL_1__10902_ (
);

FILL FILL_4__13767_ (
);

FILL FILL_4__13347_ (
);

FILL FILL_2__14381_ (
);

FILL FILL_2__7927_ (
);

FILL FILL_2__7507_ (
);

FILL FILL_1__13794_ (
);

FILL FILL_1__13374_ (
);

FILL FILL_0__12787_ (
);

NAND2X1 _12652_ (
    .A(vdd),
    .B(memoryOutData[28]),
    .Y(_3481_)
);

FILL FILL_0__12367_ (
);

NAND3X1 _12232_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\aluControl_1.inst [4]),
    .C(_3198__bF$buf2),
    .Y(_3213_)
);

FILL FILL_3__13701_ (
);

FILL SFILL89640x79050 (
);

FILL FILL_5__15979_ (
);

FILL FILL_5__15559_ (
);

FILL FILL_5__15139_ (
);

NAND2X1 _9859_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1506_)
);

FILL FILL_3__16173_ (
);

DFFSR _9439_ (
    .Q(\datapath_1.regfile_1.regOut[20] [9]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_1238_[9])
);

FILL SFILL64040x16050 (
);

INVX1 _9019_ (
    .A(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_1088_)
);

FILL FILL_5__10694_ (
);

FILL FILL_1__8396_ (
);

FILL FILL_5__10274_ (
);

FILL FILL_2__15586_ (
);

FILL FILL_2__15166_ (
);

FILL SFILL89240x65050 (
);

FILL FILL_1__14999_ (
);

FILL SFILL54120x52050 (
);

FILL FILL_1__14579_ (
);

FILL FILL_1__14159_ (
);

FILL FILL_4__15913_ (
);

FILL FILL_3__9683_ (
);

OAI22X1 _13857_ (
    .A(_4360_),
    .B(_3935__bF$buf3),
    .C(_3966__bF$buf3),
    .D(_4359_),
    .Y(_4361_)
);

FILL FILL_3__9263_ (
);

NAND3X1 _13437_ (
    .A(_3898_),
    .B(_3903_),
    .C(_3919_),
    .Y(_3949_)
);

INVX1 _13017_ (
    .A(_2_[22]),
    .Y(_3663_)
);

FILL FILL_3__14906_ (
);

FILL FILL_1__15940_ (
);

FILL FILL_1__15520_ (
);

FILL FILL_1__15100_ (
);

FILL FILL_0__14933_ (
);

FILL FILL_0__14513_ (
);

FILL FILL_5__11899_ (
);

FILL SFILL54040x59050 (
);

FILL FILL_2__7680_ (
);

FILL FILL_5__11479_ (
);

FILL FILL_5__11059_ (
);

FILL FILL_3__12093_ (
);

FILL FILL_4__7186_ (
);

FILL FILL_2__11086_ (
);

FILL FILL_5__12840_ (
);

FILL FILL_5__12420_ (
);

FILL FILL_5__12000_ (
);

FILL FILL_1__10499_ (
);

FILL FILL_4__11833_ (
);

FILL FILL_4__11413_ (
);

FILL FILL_6__8893_ (
);

FILL FILL_0__7086_ (
);

DFFSR _9192_ (
    .Q(\datapath_1.regfile_1.regOut[18] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_1108_[18])
);

FILL FILL_1__16305_ (
);

FILL FILL_3__10826_ (
);

FILL FILL_3__10406_ (
);

FILL FILL_1__11860_ (
);

FILL SFILL18680x40050 (
);

FILL FILL_1__11440_ (
);

FILL FILL_1__11020_ (
);

FILL SFILL38680x1050 (
);

FILL FILL_0__15718_ (
);

FILL FILL_2__8885_ (
);

FILL FILL_2__8465_ (
);

FILL FILL_3__13298_ (
);

FILL FILL_0__10433_ (
);

FILL FILL_0__10013_ (
);

FILL FILL_5__6890_ (
);

FILL SFILL54040x14050 (
);

DFFSR _13190_ (
    .Q(\datapath_1.mux_iord.din0 [15]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3685_[15])
);

FILL FILL_5__13625_ (
);

DFFSR _7925_ (
    .Q(\datapath_1.regfile_1.regOut[8] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_458_[31])
);

NAND2X1 _7505_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_323_)
);

FILL SFILL79240x63050 (
);

FILL FILL_1__6882_ (
);

FILL FILL_4__9752_ (
);

FILL FILL_4__12618_ (
);

FILL FILL_2__13652_ (
);

FILL FILL_2__13232_ (
);

FILL FILL_5__16097_ (
);

FILL FILL_6__9678_ (
);

FILL FILL111880x76050 (
);

FILL FILL_1__12645_ (
);

FILL FILL_1__12225_ (
);

FILL FILL_0__9652_ (
);

FILL FILL_0__9232_ (
);

INVX1 _11923_ (
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_2990_)
);

FILL FILL_0__11638_ (
);

FILL FILL_0__11218_ (
);

AOI21X1 _11503_ (
    .A(_2615_),
    .B(_2613_),
    .C(_2610_),
    .Y(_2616_)
);

FILL FILL_5__7675_ (
);

FILL FILL_4__16451_ (
);

FILL FILL_4__16031_ (
);

INVX1 _14395_ (
    .A(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_4888_)
);

FILL FILL_3__15864_ (
);

FILL FILL_3__15444_ (
);

FILL FILL_3__15024_ (
);

FILL FILL_1__7247_ (
);

FILL FILL_6_BUFX2_insert500 (
);

FILL FILL_2__14857_ (
);

FILL FILL_2__14437_ (
);

FILL FILL_0__15891_ (
);

FILL FILL_2__14017_ (
);

FILL FILL_0__15471_ (
);

FILL FILL_6_BUFX2_insert505 (
);

FILL FILL_0__15051_ (
);

FILL FILL111880x31050 (
);

FILL FILL_3__8954_ (
);

NAND2X1 _12708_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[4]),
    .Y(_3498_)
);

FILL FILL_3__8114_ (
);

FILL SFILL8520x27050 (
);

FILL FILL_4__12371_ (
);

FILL SFILL44040x12050 (
);

FILL FILL_3__16229_ (
);

FILL FILL_2__6951_ (
);

FILL FILL_3__11784_ (
);

FILL FILL_5__9401_ (
);

FILL FILL_3__11364_ (
);

FILL FILL_4__6877_ (
);

FILL SFILL69240x61050 (
);

FILL FILL_0__16256_ (
);

NOR2X1 _16121_ (
    .A(_6571_),
    .B(_6574_),
    .Y(_6575_)
);

FILL FILL_2__10777_ (
);

FILL SFILL48360x20050 (
);

FILL FILL_0__11391_ (
);

FILL FILL_1__9813_ (
);

FILL FILL_3__9739_ (
);

FILL FILL_5__14583_ (
);

FILL FILL_5__14163_ (
);

NAND2X1 _8883_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1018_)
);

NAND2X1 _8463_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_799_)
);

DFFSR _8043_ (
    .Q(\datapath_1.regfile_1.regOut[9] [21]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_523_[21])
);

FILL FILL_4__13996_ (
);

FILL FILL_4__13576_ (
);

FILL FILL_4__13156_ (
);

FILL FILL_2__14190_ (
);

FILL FILL_2__7736_ (
);

FILL FILL_3__12989_ (
);

FILL FILL_3__12569_ (
);

FILL FILL_2__7316_ (
);

FILL FILL_3__12149_ (
);

FILL FILL_0__12596_ (
);

NAND2X1 _12881_ (
    .A(vdd),
    .B(\datapath_1.rd1 [19]),
    .Y(_3593_)
);

NAND2X1 _12461_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [7]),
    .Y(_3374_)
);

FILL FILL_0__12176_ (
);

AOI22X1 _12041_ (
    .A(\datapath_1.ALUResult [13]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3077_)
);

FILL FILL_3__13930_ (
);

FILL FILL_6__16375_ (
);

FILL FILL_3__13510_ (
);

FILL FILL_4__8603_ (
);

FILL FILL_5_BUFX2_insert520 (
);

FILL FILL_5_BUFX2_insert521 (
);

FILL FILL_5__15788_ (
);

FILL FILL_5__15368_ (
);

FILL FILL_2__12503_ (
);

FILL FILL_5_BUFX2_insert522 (
);

FILL FILL_5_BUFX2_insert523 (
);

INVX1 _9668_ (
    .A(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_1419_)
);

FILL FILL_5_BUFX2_insert524 (
);

INVX1 _9248_ (
    .A(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_1200_)
);

FILL FILL_5_BUFX2_insert525 (
);

FILL FILL_5_BUFX2_insert526 (
);

FILL FILL_5_BUFX2_insert527 (
);

FILL FILL_1__11916_ (
);

FILL FILL_5_BUFX2_insert528 (
);

FILL FILL_5_BUFX2_insert529 (
);

FILL FILL_2__15395_ (
);

FILL FILL_0__10909_ (
);

FILL FILL_0__8503_ (
);

FILL FILL_1__14388_ (
);

FILL FILL_5__6946_ (
);

FILL FILL_4__15722_ (
);

FILL FILL_1_BUFX2_insert1050 (
);

FILL FILL_4__15302_ (
);

FILL FILL_1_BUFX2_insert1051 (
);

FILL FILL_1_BUFX2_insert1052 (
);

FILL FILL_1_BUFX2_insert1053 (
);

FILL FILL_3__9492_ (
);

FILL FILL_1_BUFX2_insert1054 (
);

AOI22X1 _13666_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [4]),
    .C(\datapath_1.regfile_1.regOut[31] [4]),
    .D(_3995__bF$buf1),
    .Y(_4174_)
);

NAND2X1 _13246_ (
    .A(\datapath_1.a3 [3]),
    .B(_3771_),
    .Y(_3789_)
);

FILL FILL_1_BUFX2_insert1055 (
);

FILL FILL_1_BUFX2_insert1056 (
);

FILL FILL_1_BUFX2_insert1057 (
);

FILL FILL_3__14715_ (
);

FILL FILL_1_BUFX2_insert1058 (
);

FILL FILL_1_BUFX2_insert1059 (
);

FILL FILL_1__6938_ (
);

FILL FILL_4__9808_ (
);

FILL FILL_6__12295_ (
);

FILL FILL_2__13708_ (
);

FILL SFILL99320x55050 (
);

FILL FILL_0__14742_ (
);

FILL FILL_0__14322_ (
);

FILL SFILL19080x70050 (
);

FILL FILL_5__11288_ (
);

FILL SFILL28760x75050 (
);

FILL FILL_3__7805_ (
);

FILL SFILL59160x66050 (
);

FILL FILL_2_BUFX2_insert650 (
);

FILL FILL_2_BUFX2_insert651 (
);

FILL FILL_2_BUFX2_insert652 (
);

FILL FILL_2_BUFX2_insert653 (
);

FILL SFILL83640x77050 (
);

FILL FILL_2_BUFX2_insert654 (
);

FILL FILL_4__11642_ (
);

FILL SFILL64120x49050 (
);

FILL FILL_2_BUFX2_insert655 (
);

FILL FILL_4__11222_ (
);

FILL FILL_2_BUFX2_insert656 (
);

FILL FILL_2_BUFX2_insert657 (
);

FILL FILL_2_BUFX2_insert658 (
);

FILL FILL_2_BUFX2_insert659 (
);

FILL FILL_1__16114_ (
);

FILL FILL_3__10635_ (
);

FILL FILL_0__15947_ (
);

FILL FILL_0__15527_ (
);

AOI21X1 _15812_ (
    .A(_6248_),
    .B(_6273_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [18])
);

FILL FILL_0__15107_ (
);

FILL FILL_2__8694_ (
);

FILL FILL_0__10662_ (
);

FILL FILL_2__8274_ (
);

FILL SFILL99320x10050 (
);

FILL FILL_0__10242_ (
);

FILL FILL_6__14861_ (
);

FILL FILL_6__14441_ (
);

FILL FILL_5__13854_ (
);

FILL FILL_5__13434_ (
);

FILL FILL_5__13014_ (
);

FILL SFILL28760x30050 (
);

NAND2X1 _7734_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_435_)
);

FILL SFILL59160x21050 (
);

NAND2X1 _7314_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_216_)
);

FILL FILL_4__9981_ (
);

FILL FILL_4__9141_ (
);

FILL FILL_4__12847_ (
);

FILL FILL_2__13881_ (
);

FILL FILL_4__12427_ (
);

FILL FILL_2__13461_ (
);

FILL FILL_4__12007_ (
);

FILL FILL_2__13041_ (
);

FILL FILL_1__12874_ (
);

FILL FILL_1__12454_ (
);

FILL FILL_1__12034_ (
);

FILL FILL_0__9881_ (
);

FILL FILL_2__9899_ (
);

FILL FILL_0__11867_ (
);

FILL FILL_2__9479_ (
);

FILL FILL_0__9041_ (
);

FILL FILL_0__11447_ (
);

NAND2X1 _11732_ (
    .A(_2385_),
    .B(_2481__bF$buf0),
    .Y(_2829_)
);

FILL FILL_0__11027_ (
);

OAI21X1 _11312_ (
    .A(_2430_),
    .B(_2230_),
    .C(_2429_),
    .Y(_2431_)
);

FILL FILL_5__7484_ (
);

FILL FILL_5__7064_ (
);

FILL FILL_4__16260_ (
);

FILL FILL_6__10781_ (
);

FILL FILL_5__14639_ (
);

FILL FILL_3__15673_ (
);

FILL FILL_5__14219_ (
);

DFFSR _8939_ (
    .Q(\datapath_1.regfile_1.regOut[16] [21]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_978_[21])
);

FILL FILL_3__15253_ (
);

FILL SFILL18760x73050 (
);

INVX1 _8519_ (
    .A(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_836_)
);

FILL FILL_1__7476_ (
);

FILL FILL_1__7056_ (
);

FILL FILL_2__14666_ (
);

FILL FILL_2__14246_ (
);

FILL FILL_0__15280_ (
);

FILL FILL_1__13659_ (
);

FILL FILL_1__13239_ (
);

FILL FILL_1_BUFX2_insert670 (
);

FILL FILL_3__8763_ (
);

FILL FILL_1_BUFX2_insert671 (
);

FILL FILL_1_BUFX2_insert672 (
);

FILL FILL_3__8343_ (
);

DFFSR _12937_ (
    .Q(\datapath_1.a [18]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3555_[18])
);

INVX1 _12517_ (
    .A(ALUOut[26]),
    .Y(_3411_)
);

FILL FILL_1_BUFX2_insert673 (
);

FILL FILL_1_BUFX2_insert674 (
);

FILL FILL_1_BUFX2_insert675 (
);

FILL FILL_1_BUFX2_insert676 (
);

FILL FILL_5__8269_ (
);

FILL FILL_1__14600_ (
);

FILL FILL_1_BUFX2_insert677 (
);

FILL FILL_1_BUFX2_insert678 (
);

FILL FILL_1_BUFX2_insert679 (
);

FILL FILL_4__12180_ (
);

FILL SFILL89640x29050 (
);

FILL FILL_3__16038_ (
);

FILL FILL_5__10979_ (
);

FILL FILL_5__10559_ (
);

FILL FILL_3__11593_ (
);

FILL FILL_5__10139_ (
);

FILL FILL_5__9630_ (
);

FILL FILL_3__11173_ (
);

FILL FILL_5__9210_ (
);

OAI21X1 _16350_ (
    .A(_6786_),
    .B(gnd),
    .C(_6787_),
    .Y(_6769_[9])
);

FILL FILL_0__16065_ (
);

FILL FILL_2__10166_ (
);

FILL FILL_5__11920_ (
);

FILL FILL_1__9622_ (
);

FILL FILL_5__11500_ (
);

FILL SFILL89240x15050 (
);

FILL FILL_3__9548_ (
);

FILL FILL_4__10913_ (
);

FILL FILL_3__9128_ (
);

FILL FILL_5__14392_ (
);

FILL FILL_6__7973_ (
);

FILL FILL_1__15805_ (
);

DFFSR _8692_ (
    .Q(\datapath_1.regfile_1.regOut[14] [30]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_848_[30])
);

INVX1 _8272_ (
    .A(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_712_)
);

FILL SFILL79320x51050 (
);

FILL SFILL18680x35050 (
);

FILL FILL_1__10940_ (
);

FILL FILL_4__13385_ (
);

FILL FILL_1__10520_ (
);

FILL FILL_2__7965_ (
);

BUFX2 BUFX2_insert340 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf1 )
);

FILL FILL_2__7545_ (
);

BUFX2 BUFX2_insert341 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf0 )
);

FILL FILL_3__12378_ (
);

FILL FILL_2__7125_ (
);

FILL FILL111960x64050 (
);

BUFX2 BUFX2_insert342 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf4 )
);

BUFX2 BUFX2_insert343 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf3 )
);

BUFX2 BUFX2_insert344 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf2 )
);

BUFX2 BUFX2_insert345 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf1 )
);

BUFX2 BUFX2_insert346 (
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf0 )
);

FILL SFILL103880x13050 (
);

BUFX2 BUFX2_insert347 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf4)
);

BUFX2 BUFX2_insert348 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf3)
);

DFFSR _12690_ (
    .Q(\datapath_1.Data [27]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[27])
);

BUFX2 BUFX2_insert349 (
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf2)
);

NAND3X1 _12270_ (
    .A(_3239_),
    .B(_3240_),
    .C(_3241_),
    .Y(\datapath_1.alu_1.ALUInB [13])
);

FILL FILL_5__12705_ (
);

FILL FILL_4__8832_ (
);

FILL FILL_2__12732_ (
);

FILL FILL_5__15597_ (
);

FILL FILL_5__15177_ (
);

FILL FILL_2__12312_ (
);

INVX1 _9897_ (
    .A(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_1531_)
);

INVX1 _9477_ (
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_1312_)
);

DFFSR _9057_ (
    .Q(\datapath_1.regfile_1.regOut[17] [11]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_1043_[11])
);

FILL FILL_1__11725_ (
);

FILL FILL_1__11305_ (
);

FILL FILL_0__8732_ (
);

FILL FILL_0__8312_ (
);

FILL FILL_1__14197_ (
);

FILL FILL_6__14917_ (
);

FILL FILL_4__15951_ (
);

FILL FILL_4__15531_ (
);

FILL FILL_4__15111_ (
);

AOI22X1 _13895_ (
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .B(_4246_),
    .C(_4115_),
    .D(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_4398_)
);

NOR2X1 _13475_ (
    .A(_3986_),
    .B(_3963_),
    .Y(_3987_)
);

DFFSR _13055_ (
    .Q(_2_[8]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_3620_[8])
);

FILL FILL_3__14944_ (
);

FILL FILL_3__14524_ (
);

FILL FILL_3__14104_ (
);

FILL FILL_4__9617_ (
);

FILL FILL_2__13937_ (
);

FILL SFILL114360x83050 (
);

FILL FILL_0__14971_ (
);

FILL FILL_2__13517_ (
);

FILL FILL_0__14551_ (
);

FILL FILL_0__14131_ (
);

FILL FILL_5__11097_ (
);

FILL FILL_0__9937_ (
);

FILL FILL_3__7614_ (
);

FILL FILL_0__9517_ (
);

FILL FILL_4__16316_ (
);

FILL SFILL109400x39050 (
);

FILL FILL_6__10837_ (
);

FILL FILL_4__11871_ (
);

FILL FILL_4__11451_ (
);

FILL FILL_4__11031_ (
);

FILL FILL_3__15729_ (
);

FILL FILL_3__15309_ (
);

FILL FILL_1__16343_ (
);

FILL FILL_5__8901_ (
);

FILL FILL_3__10444_ (
);

FILL FILL_3__10024_ (
);

FILL SFILL69240x56050 (
);

FILL FILL_0__15756_ (
);

FILL FILL_0__15336_ (
);

INVX1 _15621_ (
    .A(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_6087_)
);

NOR2X1 _15201_ (
    .A(_5674_),
    .B(_5677_),
    .Y(_5678_)
);

FILL SFILL109000x25050 (
);

FILL FILL_0__10891_ (
);

FILL FILL_2__8083_ (
);

FILL FILL_0__10051_ (
);

FILL FILL_5__13663_ (
);

FILL FILL_5__13243_ (
);

NAND2X1 _7963_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_547_)
);

NAND2X1 _7543_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .Y(_392_)
);

INVX1 _7123_ (
    .A(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_129_)
);

FILL FILL_4__9790_ (
);

FILL FILL_4__9370_ (
);

FILL FILL_4__12656_ (
);

FILL FILL_4__12236_ (
);

FILL FILL_2__13690_ (
);

FILL FILL_2__13270_ (
);

FILL FILL_6__9296_ (
);

FILL FILL_3__11649_ (
);

FILL FILL_3__11229_ (
);

FILL FILL_1__12263_ (
);

NAND2X1 _16406_ (
    .A(gnd),
    .B(gnd),
    .Y(_6825_)
);

FILL FILL_0__9270_ (
);

OAI21X1 _11961_ (
    .A(_3014_),
    .B(IorD_bF$buf2),
    .C(_3015_),
    .Y(_1_[24])
);

FILL FILL_2__9288_ (
);

FILL FILL_0__11676_ (
);

FILL SFILL104360x81050 (
);

FILL SFILL69240x11050 (
);

FILL FILL_0__11256_ (
);

NAND3X1 _11541_ (
    .A(_2639_),
    .B(_2642_),
    .C(_2651_),
    .Y(\datapath_1.ALUResult [23])
);

NAND2X1 _11121_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2240_)
);

FILL FILL_6__15035_ (
);

FILL FILL_5__7293_ (
);

FILL FILL_6__10170_ (
);

FILL FILL_5__14868_ (
);

FILL FILL_5__14448_ (
);

FILL FILL_5__14028_ (
);

FILL FILL_3__15482_ (
);

FILL FILL_3__15062_ (
);

INVX1 _8748_ (
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_948_)
);

INVX1 _8328_ (
    .A(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_729_)
);

FILL FILL_2__14895_ (
);

FILL FILL_2__14475_ (
);

FILL FILL_2__14055_ (
);

FILL SFILL38760x27050 (
);

FILL SFILL69160x18050 (
);

FILL FILL_1__13888_ (
);

FILL FILL_1__13468_ (
);

FILL FILL_4__14802_ (
);

FILL FILL_3__8992_ (
);

FILL FILL_3__8572_ (
);

INVX1 _12746_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_3523_)
);

NAND3X1 _12326_ (
    .A(_3281_),
    .B(_3282_),
    .C(_3283_),
    .Y(\datapath_1.alu_1.ALUInB [27])
);

FILL FILL_5__8498_ (
);

FILL FILL_5__8078_ (
);

FILL FILL_0__13822_ (
);

FILL FILL_0__13402_ (
);

FILL FILL_3__16267_ (
);

FILL FILL_5__10788_ (
);

FILL FILL_5__10368_ (
);

FILL FILL_0__16294_ (
);

FILL FILL_2__10395_ (
);

FILL SFILL24040x48050 (
);

FILL FILL_1__9851_ (
);

FILL SFILL104280x43050 (
);

FILL FILL_1__9011_ (
);

FILL FILL_2__16201_ (
);

FILL FILL_3__9777_ (
);

FILL FILL_3__9357_ (
);

FILL FILL_4__10302_ (
);

FILL FILL_1__15614_ (
);

INVX1 _8081_ (
    .A(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_605_)
);

FILL FILL_0__14607_ (
);

FILL FILL_2__7354_ (
);

FILL FILL_3__12187_ (
);

FILL FILL_6__13521_ (
);

FILL FILL_5__12514_ (
);

FILL SFILL59160x16050 (
);

FILL FILL_4__8641_ (
);

FILL FILL_5_BUFX2_insert900 (
);

FILL FILL_4__11927_ (
);

FILL FILL_4__8221_ (
);

FILL FILL_2__12961_ (
);

FILL FILL_5_BUFX2_insert901 (
);

FILL FILL_4__11507_ (
);

FILL FILL_5_BUFX2_insert902 (
);

FILL FILL_5_BUFX2_insert903 (
);

FILL FILL_2__12121_ (
);

FILL FILL_5_BUFX2_insert904 (
);

FILL FILL_5_BUFX2_insert905 (
);

OAI21X1 _9286_ (
    .A(_1224_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1225_),
    .Y(_1173_[26])
);

FILL FILL_5_BUFX2_insert906 (
);

FILL FILL_5_BUFX2_insert907 (
);

FILL FILL_5_BUFX2_insert908 (
);

FILL FILL_1__11954_ (
);

FILL FILL_5_BUFX2_insert909 (
);

FILL FILL_4__14399_ (
);

FILL FILL_1__11534_ (
);

FILL FILL_1__11114_ (
);

FILL FILL_0__8961_ (
);

FILL FILL_2__8979_ (
);

FILL FILL_0__10947_ (
);

FILL SFILL89320x48050 (
);

FILL SFILL89800x10050 (
);

NAND2X1 _10812_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1999_)
);

FILL FILL_0__8121_ (
);

FILL FILL_2__8139_ (
);

FILL FILL_0__10527_ (
);

FILL FILL_0__10107_ (
);

FILL FILL_5__6984_ (
);

FILL FILL_4__15760_ (
);

FILL FILL_4__15340_ (
);

OAI21X1 _13284_ (
    .A(_3822_),
    .B(_3811_),
    .C(_3750_),
    .Y(_3823_)
);

FILL FILL_2__9920_ (
);

FILL FILL_5__13719_ (
);

FILL FILL_2__9500_ (
);

FILL FILL_3__14753_ (
);

FILL FILL_3__14333_ (
);

FILL SFILL49160x59050 (
);

FILL FILL_1__6976_ (
);

FILL FILL_4__9846_ (
);

FILL FILL_4__9426_ (
);

FILL FILL_4__9006_ (
);

FILL FILL_2__13746_ (
);

FILL FILL_2__13326_ (
);

FILL FILL_0__14780_ (
);

FILL FILL_0__14360_ (
);

FILL FILL_1__12739_ (
);

FILL FILL_1__12319_ (
);

FILL SFILL79000x70050 (
);

FILL FILL_3__7843_ (
);

FILL FILL_0__9746_ (
);

FILL FILL_3__7423_ (
);

FILL SFILL33960x43050 (
);

FILL FILL_5__7349_ (
);

FILL FILL_4__16125_ (
);

FILL FILL_6__10646_ (
);

OAI22X1 _14489_ (
    .A(_4979_),
    .B(_3935__bF$buf4),
    .C(_3924__bF$buf0),
    .D(_4978_),
    .Y(_4980_)
);

FILL FILL_4__11680_ (
);

INVX1 _14069_ (
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_4569_)
);

FILL FILL_4__11260_ (
);

FILL FILL_3__15958_ (
);

FILL FILL_3__15538_ (
);

FILL FILL_3__15118_ (
);

FILL FILL_1__16152_ (
);

FILL FILL_3__10673_ (
);

FILL FILL_5__8710_ (
);

FILL FILL_3__10253_ (
);

FILL SFILL18760x23050 (
);

FILL FILL_0__15985_ (
);

FILL FILL_0__15565_ (
);

NAND2X1 _15850_ (
    .A(_6304_),
    .B(_6310_),
    .Y(_6311_)
);

FILL FILL_0__15145_ (
);

INVX1 _15430_ (
    .A(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_5901_)
);

INVX8 _15010_ (
    .A(_5489__bF$buf0),
    .Y(_5490_)
);

FILL FILL_0__10280_ (
);

FILL FILL_1__8702_ (
);

FILL FILL_3__8628_ (
);

FILL FILL_3__8208_ (
);

FILL FILL_5__13892_ (
);

FILL FILL_5__13472_ (
);

DFFSR _7772_ (
    .Q(\datapath_1.regfile_1.regOut[7] [6]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_393_[6])
);

INVX1 _7352_ (
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_241_)
);

FILL SFILL79320x46050 (
);

FILL FILL_4__12885_ (
);

FILL FILL_4__12465_ (
);

FILL FILL_4__12045_ (
);

FILL FILL_5__9915_ (
);

FILL FILL_3__11878_ (
);

FILL FILL111960x59050 (
);

FILL FILL_3__11458_ (
);

FILL FILL_1__12492_ (
);

FILL FILL_3__11038_ (
);

FILL FILL_1__12072_ (
);

INVX1 _16215_ (
    .A(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_6666_)
);

FILL FILL_2__9097_ (
);

AOI21X1 _11770_ (
    .A(_2364_),
    .B(_2864_),
    .C(_2458_),
    .Y(_2865_)
);

FILL FILL_0__11485_ (
);

NOR2X1 _11350_ (
    .A(_2467_),
    .B(_2466_),
    .Y(_2468_)
);

FILL FILL_0__11065_ (
);

FILL FILL_1__9907_ (
);

FILL FILL_2__11812_ (
);

FILL FILL_5__14677_ (
);

FILL FILL_5__14257_ (
);

INVX1 _8977_ (
    .A(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_1060_)
);

FILL FILL_3__15291_ (
);

DFFSR _8557_ (
    .Q(\datapath_1.regfile_1.regOut[13] [23]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_783_[23])
);

OAI21X1 _8137_ (
    .A(_641_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_642_),
    .Y(_588_[27])
);

FILL FILL_1__7094_ (
);

FILL FILL_1__10805_ (
);

FILL FILL_2__14284_ (
);

FILL SFILL114440x71050 (
);

FILL FILL_0__7812_ (
);

FILL SFILL94440x8050 (
);

FILL FILL_1__13697_ (
);

FILL FILL_1__13277_ (
);

FILL FILL_4__14611_ (
);

FILL FILL111960x14050 (
);

FILL FILL_3__8381_ (
);

INVX1 _12975_ (
    .A(_2_[8]),
    .Y(_3635_)
);

DFFSR _12555_ (
    .Q(ALUOut[20]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3360_[20])
);

OAI21X1 _12135_ (
    .A(_3142_),
    .B(ALUSrcA_bF$buf4),
    .C(_3143_),
    .Y(\datapath_1.alu_1.ALUInA [6])
);

FILL FILL_3__13604_ (
);

FILL FILL_0__13631_ (
);

FILL FILL_0__13211_ (
);

FILL FILL_3__16076_ (
);

FILL FILL_5__10177_ (
);

FILL FILL_2__15489_ (
);

FILL FILL_2__15069_ (
);

FILL FILL_5__16403_ (
);

FILL FILL_1__9660_ (
);

FILL FILL_1__9240_ (
);

FILL FILL_4__15816_ (
);

FILL FILL_2__16010_ (
);

FILL FILL_4__10951_ (
);

FILL FILL_3__9166_ (
);

FILL FILL_4__10531_ (
);

FILL FILL_4__10111_ (
);

FILL FILL_3__14809_ (
);

FILL FILL_6__7591_ (
);

FILL FILL_1__15843_ (
);

FILL FILL_1__15423_ (
);

FILL FILL_1__15003_ (
);

FILL FILL_0__14836_ (
);

NOR2X1 _14701_ (
    .A(_5183_),
    .B(_5186_),
    .Y(_5187_)
);

FILL FILL_0__14416_ (
);

BUFX2 BUFX2_insert720 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf7 )
);

FILL FILL_2__7583_ (
);

BUFX2 BUFX2_insert721 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf6 )
);

FILL FILL_2__7163_ (
);

BUFX2 BUFX2_insert722 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf5 )
);

BUFX2 BUFX2_insert723 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf4 )
);

BUFX2 BUFX2_insert724 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf3 )
);

BUFX2 BUFX2_insert725 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf2 )
);

BUFX2 BUFX2_insert726 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf1 )
);

FILL FILL_4__7089_ (
);

BUFX2 BUFX2_insert727 (
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf0 )
);

BUFX2 BUFX2_insert728 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf4 )
);

BUFX2 BUFX2_insert729 (
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf3 )
);

FILL FILL_5__12743_ (
);

FILL FILL_5__12323_ (
);

FILL FILL_4__8870_ (
);

FILL FILL_4__8450_ (
);

FILL FILL_4__11736_ (
);

FILL FILL_2__12770_ (
);

FILL FILL_4__11316_ (
);

FILL FILL_2__12350_ (
);

FILL FILL_6__8376_ (
);

FILL FILL_1__16208_ (
);

OAI21X1 _9095_ (
    .A(_1117_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .C(_1118_),
    .Y(_1108_[5])
);

FILL FILL_3__10309_ (
);

FILL FILL_1__11763_ (
);

FILL FILL_1__11343_ (
);

INVX1 _15906_ (
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_6365_)
);

FILL FILL_2__8788_ (
);

FILL FILL_0__8770_ (
);

FILL SFILL104360x76050 (
);

FILL FILL_0__10756_ (
);

FILL FILL_2__8368_ (
);

FILL FILL_0__8350_ (
);

NAND2X1 _10621_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1892_)
);

DFFSR _10201_ (
    .Q(\datapath_1.regfile_1.regOut[26] [3]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_1628_[3])
);

OAI21X1 _13093_ (
    .A(_3692_),
    .B(PCEn_bF$buf1),
    .C(_3693_),
    .Y(_3685_[4])
);

FILL FILL_5__13948_ (
);

FILL FILL_3__14982_ (
);

FILL FILL_5__13528_ (
);

FILL FILL_3__14562_ (
);

FILL FILL_5__13108_ (
);

FILL FILL_3__14142_ (
);

INVX1 _7828_ (
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_477_)
);

DFFSR _7408_ (
    .Q(\datapath_1.regfile_1.regOut[4] [26]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_198_[26])
);

FILL FILL_4_BUFX2_insert560 (
);

FILL FILL_4__9655_ (
);

FILL FILL_4_BUFX2_insert561 (
);

FILL FILL_4_BUFX2_insert562 (
);

FILL FILL_4__9235_ (
);

FILL FILL_4_BUFX2_insert563 (
);

FILL FILL_2__13975_ (
);

FILL FILL_4_BUFX2_insert564 (
);

FILL FILL_2__13555_ (
);

FILL SFILL99400x38050 (
);

FILL FILL_4_BUFX2_insert565 (
);

FILL FILL_2__13135_ (
);

FILL FILL_4_BUFX2_insert566 (
);

FILL FILL_4_BUFX2_insert567 (
);

FILL FILL_4_BUFX2_insert568 (
);

FILL FILL_4_BUFX2_insert569 (
);

FILL FILL_1__12968_ (
);

FILL FILL_1__12128_ (
);

FILL FILL_0__9975_ (
);

FILL FILL_0__9555_ (
);

FILL FILL112440x82050 (
);

FILL FILL_3__7232_ (
);

FILL FILL_0__9135_ (
);

AOI21X1 _11826_ (
    .A(_2353_),
    .B(_2359_),
    .C(_2458_),
    .Y(_2916_)
);

INVX2 _11406_ (
    .A(_2269_),
    .Y(_2523_)
);

FILL FILL_5__7998_ (
);

FILL FILL_5__7578_ (
);

FILL SFILL104360x31050 (
);

FILL FILL_4__16354_ (
);

FILL FILL_5__7158_ (
);

NAND3X1 _14298_ (
    .A(_4784_),
    .B(_4785_),
    .C(_4792_),
    .Y(_4793_)
);

FILL FILL_0__12902_ (
);

FILL FILL_3__15767_ (
);

FILL FILL_3__15347_ (
);

FILL FILL_1__16381_ (
);

FILL FILL_3__10062_ (
);

FILL SFILL64120x1050 (
);

FILL FILL_0__15794_ (
);

FILL FILL_0__15374_ (
);

FILL FILL_1__8511_ (
);

FILL FILL_2__15701_ (
);

FILL FILL_3__8857_ (
);

FILL FILL_3__8017_ (
);

FILL FILL_5__13281_ (
);

INVX1 _7581_ (
    .A(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_353_)
);

INVX1 _7161_ (
    .A(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_134_)
);

FILL FILL_4__12274_ (
);

FILL FILL_2__6854_ (
);

FILL FILL_3__11687_ (
);

FILL FILL_5__9724_ (
);

FILL FILL_3__11267_ (
);

FILL FILL_0__16159_ (
);

DFFSR _16444_ (
    .Q(\datapath_1.regfile_1.regOut[0] [27]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_6769_[27])
);

OAI22X1 _16024_ (
    .A(_6479_),
    .B(_5501_),
    .C(_5524__bF$buf3),
    .D(_5127_),
    .Y(_6480_)
);

FILL FILL_0__11294_ (
);

FILL FILL_3_BUFX2_insert580 (
);

FILL FILL_4__7721_ (
);

FILL SFILL113800x4050 (
);

FILL FILL_3_BUFX2_insert581 (
);

FILL FILL_4__7301_ (
);

FILL FILL_3_BUFX2_insert582 (
);

FILL FILL_3_BUFX2_insert583 (
);

FILL FILL_5__14486_ (
);

FILL FILL_2__11621_ (
);

FILL FILL_3_BUFX2_insert584 (
);

FILL FILL_5__14066_ (
);

FILL FILL_2__11201_ (
);

FILL FILL_3_BUFX2_insert585 (
);

OAI21X1 _8786_ (
    .A(_972_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_973_),
    .Y(_913_[30])
);

FILL FILL_3_BUFX2_insert586 (
);

OAI21X1 _8366_ (
    .A(_753_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_754_),
    .Y(_718_[18])
);

FILL FILL_3_BUFX2_insert587 (
);

FILL FILL_3_BUFX2_insert588 (
);

FILL FILL_3_BUFX2_insert589 (
);

FILL FILL_4__13899_ (
);

FILL FILL_1__10614_ (
);

FILL FILL_4__13479_ (
);

FILL FILL_2__14093_ (
);

FILL SFILL73720x58050 (
);

FILL FILL_0__7621_ (
);

FILL FILL_0__7201_ (
);

FILL FILL_2__7219_ (
);

FILL FILL_1__13086_ (
);

FILL FILL_4__14840_ (
);

FILL FILL_4__14420_ (
);

FILL FILL_4__14000_ (
);

OAI21X1 _12784_ (
    .A(_3547_),
    .B(IRWrite_bF$buf4),
    .C(_3548_),
    .Y(_3490_[29])
);

FILL FILL_0__12499_ (
);

FILL FILL_3__8190_ (
);

INVX1 _12364_ (
    .A(ALUOut[7]),
    .Y(_3308_)
);

FILL FILL_0__12079_ (
);

FILL FILL_3__13833_ (
);

FILL FILL_3__13413_ (
);

FILL FILL_6__16278_ (
);

FILL FILL_4__8506_ (
);

FILL FILL_2__12826_ (
);

FILL FILL_2__12406_ (
);

FILL FILL_0__13860_ (
);

FILL FILL_0__13440_ (
);

FILL FILL_0__13020_ (
);

FILL FILL_1__11819_ (
);

FILL FILL_2__15298_ (
);

FILL FILL_3__6923_ (
);

FILL FILL_5__16212_ (
);

FILL FILL_0__8826_ (
);

FILL SFILL33960x38050 (
);

FILL FILL_5__6849_ (
);

FILL FILL_4__15625_ (
);

FILL FILL_4__15205_ (
);

AOI22X1 _13989_ (
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .B(_3942__bF$buf2),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_4490_)
);

FILL FILL_3__9395_ (
);

FILL FILL_4__10760_ (
);

INVX8 _13569_ (
    .A(_3920_),
    .Y(_4079_)
);

NAND2X1 _13149_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [23]),
    .Y(_3731_)
);

FILL FILL_3__14618_ (
);

FILL FILL_1__15652_ (
);

FILL FILL_1__15232_ (
);

FILL SFILL94200x40050 (
);

FILL SFILL18760x18050 (
);

FILL FILL_6__12198_ (
);

FILL FILL_0__14645_ (
);

AOI22X1 _14930_ (
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .B(_4225_),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_5411_)
);

FILL FILL_0__14225_ (
);

AOI21X1 _14510_ (
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .B(_4079__bF$buf3),
    .C(_4999_),
    .Y(_5000_)
);

FILL FILL_3__7708_ (
);

FILL FILL_5__12972_ (
);

FILL FILL_5__12132_ (
);

BUFX2 _6852_ (
    .A(_1_[14]),
    .Y(memoryAddress[14])
);

FILL FILL_4__11965_ (
);

FILL SFILL33720x8050 (
);

FILL FILL_4__11545_ (
);

FILL FILL_4__11125_ (
);

FILL FILL_1__16017_ (
);

FILL FILL_3__10958_ (
);

FILL FILL_1__11992_ (
);

FILL FILL_3__10538_ (
);

FILL SFILL84200x83050 (
);

FILL FILL_1__11572_ (
);

FILL FILL_3__10118_ (
);

FILL FILL_1__11152_ (
);

NOR3X1 _15715_ (
    .A(_4728_),
    .B(\datapath_1.PCJump_27_bF$buf3 ),
    .C(_5519_),
    .Y(_6179_)
);

FILL SFILL84280x40050 (
);

FILL FILL_2__8597_ (
);

DFFSR _10850_ (
    .Q(\datapath_1.regfile_1.regOut[31] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_1953_[12])
);

FILL FILL_0__10565_ (
);

INVX1 _10430_ (
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_1805_)
);

FILL FILL_0__10145_ (
);

INVX1 _10010_ (
    .A(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_1586_)
);

FILL FILL_6__14764_ (
);

FILL FILL_6__14344_ (
);

FILL SFILL110120x58050 (
);

FILL SFILL109480x83050 (
);

FILL FILL_5__13757_ (
);

FILL FILL_5__13337_ (
);

FILL FILL_3__14791_ (
);

FILL FILL_3__14371_ (
);

OAI21X1 _7637_ (
    .A(_389_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_390_),
    .Y(_328_[31])
);

OAI21X1 _7217_ (
    .A(_170_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_171_),
    .Y(_133_[19])
);

FILL FILL_4__9884_ (
);

FILL FILL_4__9464_ (
);

FILL FILL_4__9044_ (
);

FILL FILL_2__13784_ (
);

FILL SFILL114440x66050 (
);

FILL FILL_2__13364_ (
);

FILL FILL_1__12777_ (
);

FILL FILL_1__12357_ (
);

FILL FILL_0__9784_ (
);

FILL FILL_3__7881_ (
);

FILL FILL_3__7461_ (
);

FILL FILL_0__9364_ (
);

FILL FILL_3__7041_ (
);

NOR2X1 _11635_ (
    .A(_2736_),
    .B(_2738_),
    .Y(_2739_)
);

NOR2X1 _11215_ (
    .A(ALUControl[0]),
    .B(_2333_),
    .Y(_2334_)
);

FILL FILL_4__16163_ (
);

FILL FILL_6__10264_ (
);

FILL FILL_3__15996_ (
);

FILL FILL_0__12711_ (
);

FILL FILL_3__15576_ (
);

FILL FILL_3__15156_ (
);

FILL FILL_1__16190_ (
);

FILL FILL_1__7799_ (
);

FILL FILL_1__7379_ (
);

FILL FILL_3__10291_ (
);

FILL FILL_2__14989_ (
);

FILL FILL_2__14569_ (
);

FILL FILL_2__14149_ (
);

FILL FILL_0__15183_ (
);

FILL FILL_5__15903_ (
);

FILL FILL_1__8740_ (
);

FILL FILL_1__8320_ (
);

FILL FILL_2__15930_ (
);

FILL FILL_2__15510_ (
);

FILL SFILL74200x81050 (
);

FILL FILL_3__8246_ (
);

FILL FILL_5__13090_ (
);

FILL FILL_1__14923_ (
);

DFFSR _7390_ (
    .Q(\datapath_1.regfile_1.regOut[4] [8]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_198_[8])
);

FILL FILL_1__14503_ (
);

FILL FILL_4__12083_ (
);

FILL FILL_0__13916_ (
);

FILL SFILL114360x28050 (
);

FILL FILL_5__9533_ (
);

FILL FILL_3__11496_ (
);

FILL FILL_5__9113_ (
);

FILL FILL_3__11076_ (
);

FILL FILL_0__16388_ (
);

AOI22X1 _16253_ (
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [30]),
    .C(\datapath_1.regfile_1.regOut[5] [30]),
    .D(_5700_),
    .Y(_6703_)
);

FILL FILL_2__10489_ (
);

FILL FILL_2__10069_ (
);

FILL FILL_5__11823_ (
);

FILL FILL_1__9525_ (
);

FILL FILL_5__11403_ (
);

FILL FILL_1__9105_ (
);

FILL FILL_4__7950_ (
);

FILL FILL_4__10816_ (
);

FILL FILL_4__7110_ (
);

FILL FILL_2__11850_ (
);

FILL FILL_5__14295_ (
);

FILL FILL_2__11430_ (
);

FILL FILL_2__11010_ (
);

FILL FILL_1__15708_ (
);

FILL FILL_6__7456_ (
);

OAI21X1 _8595_ (
    .A(_865_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .C(_866_),
    .Y(_848_[9])
);

DFFSR _8175_ (
    .Q(\datapath_1.regfile_1.regOut[10] [25]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_588_[25])
);

FILL FILL_1__10423_ (
);

FILL FILL_4__13288_ (
);

FILL FILL_1__10003_ (
);

FILL FILL_2__7868_ (
);

FILL FILL_0__7850_ (
);

FILL FILL_2__7448_ (
);

FILL FILL_0__7430_ (
);

OAI21X1 _12593_ (
    .A(_3440_),
    .B(vdd),
    .C(_3441_),
    .Y(_3425_[8])
);

NAND2X1 _12173_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [19]),
    .Y(_3169_)
);

FILL FILL_5__12608_ (
);

FILL FILL_3__13642_ (
);

FILL FILL_3__13222_ (
);

INVX1 _6908_ (
    .A(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_6_)
);

FILL FILL_4__8735_ (
);

FILL FILL_4__8315_ (
);

FILL FILL_2__12635_ (
);

FILL FILL_2__12215_ (
);

FILL FILL_1__11628_ (
);

FILL FILL_1__11208_ (
);

FILL FILL112440x77050 (
);

FILL FILL_0__8635_ (
);

FILL FILL_5__16021_ (
);

NAND2X1 _10906_ (
    .A(\control_1.reg_state.dout [2]),
    .B(_2052_),
    .Y(_2053_)
);

FILL FILL_6__9602_ (
);

FILL FILL_0__8215_ (
);

FILL SFILL104360x26050 (
);

FILL FILL_4__15854_ (
);

FILL FILL_4__15434_ (
);

FILL FILL_4__15014_ (
);

NOR2X1 _13798_ (
    .A(_4302_),
    .B(_3949_),
    .Y(_4303_)
);

NAND2X1 _13378_ (
    .A(_3889_),
    .B(_3888_),
    .Y(_3890_)
);

FILL FILL_3__14847_ (
);

FILL FILL_1__15881_ (
);

FILL FILL_3__14427_ (
);

FILL FILL_3__14007_ (
);

FILL FILL_1__15461_ (
);

FILL FILL_1__15041_ (
);

FILL FILL112040x63050 (
);

FILL FILL_0__14874_ (
);

FILL FILL_0__14454_ (
);

FILL FILL_0__14034_ (
);

FILL FILL_3__7937_ (
);

FILL FILL_5__12781_ (
);

FILL FILL_5__12361_ (
);

FILL FILL112440x32050 (
);

FILL FILL_4__16219_ (
);

FILL FILL_4__11774_ (
);

FILL FILL_4__11354_ (
);

FILL FILL_1__16246_ (
);

FILL FILL_3__10767_ (
);

FILL FILL_1__11381_ (
);

FILL FILL_0__15659_ (
);

NOR3X1 _15944_ (
    .A(_5515__bF$buf3),
    .B(_5003_),
    .C(_5521__bF$buf3),
    .Y(_6402_)
);

FILL FILL_0__15239_ (
);

OAI22X1 _15524_ (
    .A(_5466__bF$buf4),
    .B(_4517_),
    .C(_4500_),
    .D(_5526__bF$buf0),
    .Y(_5993_)
);

NOR3X1 _15104_ (
    .A(_5515__bF$buf2),
    .B(_4007_),
    .C(_5521__bF$buf1),
    .Y(_5583_)
);

FILL FILL_0__10794_ (
);

FILL FILL_0__10374_ (
);

FILL FILL_5__13986_ (
);

FILL FILL_2__10701_ (
);

FILL FILL_5__13566_ (
);

FILL FILL_5__13146_ (
);

FILL FILL_3__14180_ (
);

OAI21X1 _7866_ (
    .A(_501_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .C(_502_),
    .Y(_458_[22])
);

OAI21X1 _7446_ (
    .A(_282_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .C(_283_),
    .Y(_263_[10])
);

DFFSR _7026_ (
    .Q(\datapath_1.regfile_1.regOut[1] [28]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_3_[28])
);

FILL FILL_4_BUFX2_insert940 (
);

FILL FILL_4_BUFX2_insert941 (
);

FILL FILL_4__9273_ (
);

FILL FILL_4_BUFX2_insert942 (
);

FILL FILL_4__12979_ (
);

FILL FILL_4_BUFX2_insert943 (
);

FILL FILL_2__13593_ (
);

FILL FILL_4__12139_ (
);

FILL FILL_4_BUFX2_insert944 (
);

FILL FILL_4_BUFX2_insert945 (
);

FILL FILL_2__13173_ (
);

FILL FILL_4_BUFX2_insert946 (
);

FILL FILL_4_BUFX2_insert947 (
);

FILL FILL_4_BUFX2_insert948 (
);

FILL FILL_4_BUFX2_insert949 (
);

FILL SFILL39320x78050 (
);

FILL FILL_1__12586_ (
);

FILL FILL_1__12166_ (
);

FILL FILL_4__13920_ (
);

OAI22X1 _16309_ (
    .A(_5466__bF$buf1),
    .B(_5450_),
    .C(_5429_),
    .D(_5526__bF$buf4),
    .Y(_6758_)
);

FILL FILL_4__13500_ (
);

FILL FILL_3__7690_ (
);

FILL FILL_0__11999_ (
);

FILL FILL_0__9593_ (
);

NOR2X1 _11864_ (
    .A(\datapath_1.ALUResult [29]),
    .B(\datapath_1.ALUResult [15]),
    .Y(_2951_)
);

FILL FILL_0__9173_ (
);

FILL FILL_0__11579_ (
);

XNOR2X1 _11444_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2560_)
);

FILL FILL_0__11159_ (
);

AND2X2 _11024_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2143_)
);

FILL FILL_3__12913_ (
);

FILL FILL_5__7196_ (
);

FILL FILL_4__16392_ (
);

FILL SFILL94280x37050 (
);

FILL FILL_2__11906_ (
);

FILL FILL_3__15385_ (
);

FILL FILL_0__12520_ (
);

FILL FILL_0__12100_ (
);

FILL FILL_1__7188_ (
);

FILL FILL_2__14798_ (
);

FILL FILL_2__14378_ (
);

FILL FILL_5__15712_ (
);

FILL FILL_4__14705_ (
);

FILL FILL_3__8895_ (
);

FILL FILL_3__8475_ (
);

NAND2X1 _12649_ (
    .A(vdd),
    .B(memoryOutData[27]),
    .Y(_3479_)
);

FILL FILL_3__8055_ (
);

AOI22X1 _12229_ (
    .A(_2_[3]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf0),
    .D(\aluControl_1.inst [1]),
    .Y(_3211_)
);

FILL FILL_1__14732_ (
);

FILL FILL_1__14312_ (
);

FILL FILL_0__13725_ (
);

FILL FILL_0__13305_ (
);

FILL FILL_2__6892_ (
);

FILL FILL_5__9762_ (
);

FILL FILL_5__9342_ (
);

FILL FILL_0_BUFX2_insert1060 (
);

FILL FILL_0_BUFX2_insert1061 (
);

FILL FILL_0_BUFX2_insert1062 (
);

FILL FILL_0__16197_ (
);

FILL FILL_0_BUFX2_insert1063 (
);

FILL FILL_0_BUFX2_insert1064 (
);

OAI22X1 _16062_ (
    .A(_5526__bF$buf1),
    .B(_5172_),
    .C(_5151_),
    .D(_5527__bF$buf2),
    .Y(_6517_)
);

FILL SFILL79000x15050 (
);

FILL FILL_0_BUFX2_insert1065 (
);

FILL FILL_2__10298_ (
);

FILL FILL_0_BUFX2_insert1066 (
);

FILL FILL_0_BUFX2_insert1067 (
);

FILL FILL_0_BUFX2_insert1068 (
);

FILL FILL_1__9754_ (
);

FILL FILL_0_BUFX2_insert1069 (
);

FILL FILL_5__11632_ (
);

FILL FILL_1__9334_ (
);

FILL FILL_5__11212_ (
);

FILL SFILL8680x54050 (
);

FILL FILL_2__16104_ (
);

FILL FILL_3_BUFX2_insert960 (
);

FILL FILL_3_BUFX2_insert961 (
);

FILL FILL_4__10625_ (
);

FILL FILL_3_BUFX2_insert962 (
);

FILL SFILL109560x71050 (
);

FILL FILL_3_BUFX2_insert963 (
);

FILL FILL_3_BUFX2_insert964 (
);

FILL FILL_3_BUFX2_insert965 (
);

FILL FILL_1__15937_ (
);

FILL FILL_3_BUFX2_insert966 (
);

FILL FILL_1__15517_ (
);

FILL FILL_3_BUFX2_insert967 (
);

FILL FILL_3_BUFX2_insert968 (
);

FILL SFILL84200x78050 (
);

FILL FILL_3_BUFX2_insert969 (
);

FILL FILL_1__10652_ (
);

FILL FILL_4__13097_ (
);

FILL FILL_1__10232_ (
);

FILL FILL_2__7677_ (
);

FILL SFILL109480x78050 (
);

FILL FILL_5__12837_ (
);

FILL FILL_3__13871_ (
);

FILL FILL_5__12417_ (
);

FILL FILL_3__13451_ (
);

FILL SFILL8600x52050 (
);

FILL FILL_3__13031_ (
);

FILL FILL_4__8964_ (
);

FILL FILL_4__8124_ (
);

FILL FILL_2__12864_ (
);

FILL FILL_2__12444_ (
);

FILL FILL_2__12024_ (
);

DFFSR _9189_ (
    .Q(\datapath_1.regfile_1.regOut[18] [15]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_1108_[15])
);

FILL FILL_1__11857_ (
);

FILL FILL_1__11437_ (
);

FILL FILL_1__11017_ (
);

FILL SFILL84200x33050 (
);

FILL FILL_0__8864_ (
);

FILL FILL_3__6961_ (
);

FILL FILL_5__16250_ (
);

FILL FILL_0__8444_ (
);

DFFSR _10715_ (
    .Q(\datapath_1.regfile_1.regOut[30] [5]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_1888_[5])
);

FILL FILL_5__6887_ (
);

FILL FILL_4__15663_ (
);

FILL FILL_4__15243_ (
);

DFFSR _13187_ (
    .Q(\datapath_1.mux_iord.din0 [12]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3685_[12])
);

FILL SFILL88520x41050 (
);

FILL FILL_2__9403_ (
);

FILL FILL_3__14656_ (
);

FILL FILL_1__15690_ (
);

FILL FILL_3__14236_ (
);

FILL FILL_1__15270_ (
);

FILL FILL_1__6879_ (
);

FILL FILL_4__9749_ (
);

FILL FILL_2__13649_ (
);

FILL FILL_2__13229_ (
);

FILL FILL_0__14683_ (
);

FILL FILL_0__14263_ (
);

FILL SFILL114440x16050 (
);

FILL FILL_1__7820_ (
);

FILL FILL_0__9649_ (
);

FILL FILL_3__7746_ (
);

FILL FILL_0__9229_ (
);

FILL FILL_3__7326_ (
);

FILL FILL_5__12590_ (
);

FILL FILL_5__12170_ (
);

FILL SFILL74280x33050 (
);

BUFX2 _6890_ (
    .A(_2_[20]),
    .Y(memoryWriteData[20])
);

FILL FILL_4__16028_ (
);

FILL FILL_4__11583_ (
);

FILL FILL_4__11163_ (
);

FILL SFILL99480x82050 (
);

FILL FILL_1__16055_ (
);

FILL FILL_3__10996_ (
);

FILL FILL_5__8613_ (
);

FILL FILL_3__10576_ (
);

FILL FILL_3__10156_ (
);

FILL FILL_1__11190_ (
);

FILL FILL_0__15888_ (
);

FILL FILL_6_BUFX2_insert474 (
);

NOR2X1 _15753_ (
    .A(_6215_),
    .B(_6213_),
    .Y(_6216_)
);

FILL FILL_0__15468_ (
);

INVX1 _15333_ (
    .A(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_5807_)
);

FILL FILL_0__15048_ (
);

FILL FILL_0__10183_ (
);

FILL FILL_5__10903_ (
);

FILL FILL_1__8605_ (
);

FILL FILL_2__10930_ (
);

FILL FILL_5__13795_ (
);

FILL FILL_2__10510_ (
);

FILL FILL_5__13375_ (
);

OAI21X1 _7675_ (
    .A(_394_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .C(_395_),
    .Y(_393_[1])
);

DFFSR _7255_ (
    .Q(\datapath_1.regfile_1.regOut[3] [1]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_133_[1])
);

FILL FILL_4__12788_ (
);

FILL FILL_4__9082_ (
);

FILL FILL_4__12368_ (
);

FILL FILL_2__6948_ (
);

FILL FILL_0__6930_ (
);

FILL FILL_1__12395_ (
);

INVX1 _16118_ (
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_6572_)
);

FILL SFILL43720x47050 (
);

FILL FILL_0__11388_ (
);

OAI21X1 _11673_ (
    .A(_2773_),
    .B(_2774_),
    .C(_2772_),
    .Y(_2775_)
);

AOI21X1 _11253_ (
    .A(_2143_),
    .B(_2371_),
    .C(_2141_),
    .Y(_2372_)
);

FILL FILL_3__12722_ (
);

FILL FILL_6__15587_ (
);

FILL FILL_3__12302_ (
);

FILL SFILL104440x14050 (
);

FILL FILL_4__7815_ (
);

FILL FILL_2__11715_ (
);

FILL SFILL64200x74050 (
);

FILL FILL_3__15194_ (
);

FILL FILL112120x51050 (
);

FILL FILL_1__10708_ (
);

FILL FILL_2__14187_ (
);

FILL FILL_5__15941_ (
);

FILL FILL_5__15521_ (
);

FILL FILL_0__7715_ (
);

FILL FILL_5__15101_ (
);

DFFSR _9821_ (
    .Q(\datapath_1.regfile_1.regOut[23] [7]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_1433_[7])
);

NAND2X1 _9401_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1282_)
);

FILL FILL_4__14934_ (
);

FILL FILL_4__14514_ (
);

NAND2X1 _12878_ (
    .A(vdd),
    .B(\datapath_1.rd1 [18]),
    .Y(_3591_)
);

NAND2X1 _12458_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [6]),
    .Y(_3372_)
);

NAND3X1 _12038_ (
    .A(_3072_),
    .B(_3073_),
    .C(_3074_),
    .Y(\datapath_1.mux_pcsrc.dout [12])
);

FILL FILL_3__13927_ (
);

FILL FILL_1__14961_ (
);

FILL FILL_3__13507_ (
);

FILL FILL_1__14541_ (
);

FILL FILL112040x58050 (
);

FILL FILL_1__14121_ (
);

FILL FILL_5_BUFX2_insert490 (
);

FILL FILL_5_BUFX2_insert491 (
);

FILL FILL_5_BUFX2_insert492 (
);

FILL FILL_0__13954_ (
);

FILL FILL_5_BUFX2_insert493 (
);

FILL FILL_3__16399_ (
);

FILL FILL_0__13534_ (
);

FILL FILL_0__13114_ (
);

FILL FILL_5_BUFX2_insert494 (
);

FILL FILL_5_BUFX2_insert495 (
);

FILL FILL_5_BUFX2_insert496 (
);

FILL FILL_5__9991_ (
);

FILL FILL_5_BUFX2_insert497 (
);

FILL FILL_5__9151_ (
);

FILL FILL_5_BUFX2_insert498 (
);

FILL FILL_5_BUFX2_insert499 (
);

OAI22X1 _16291_ (
    .A(_5414_),
    .B(_5539__bF$buf0),
    .C(_5469__bF$buf2),
    .D(_5453_),
    .Y(_6740_)
);

FILL FILL_5__16306_ (
);

FILL FILL_1__9983_ (
);

FILL FILL_5__11861_ (
);

FILL FILL_5__11441_ (
);

FILL FILL112440x27050 (
);

FILL FILL_1__9143_ (
);

FILL FILL_5__11021_ (
);

FILL FILL_4__15719_ (
);

FILL FILL_2__16333_ (
);

FILL FILL_3__9489_ (
);

FILL FILL_4__10434_ (
);

FILL FILL_4__10014_ (
);

FILL FILL_1__15746_ (
);

FILL FILL_1__15326_ (
);

FILL FILL_6__7074_ (
);

FILL FILL_1__10881_ (
);

FILL FILL_1__10041_ (
);

FILL FILL112040x13050 (
);

FILL FILL_0__14739_ (
);

NOR2X1 _14604_ (
    .A(_5091_),
    .B(_5088_),
    .Y(_5092_)
);

FILL FILL_0__14319_ (
);

FILL FILL_2__7486_ (
);

FILL FILL_2__7066_ (
);

FILL FILL_5__12646_ (
);

FILL FILL_3__13680_ (
);

FILL FILL_5__12226_ (
);

FILL FILL_3__13260_ (
);

OAI21X1 _6946_ (
    .A(_30_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .C(_31_),
    .Y(_3_[14])
);

FILL FILL_4__8773_ (
);

FILL SFILL58520x80050 (
);

FILL FILL_4__8353_ (
);

FILL FILL_4__11639_ (
);

FILL FILL_4__11219_ (
);

FILL FILL_2__12253_ (
);

FILL FILL_1__11666_ (
);

FILL FILL_1__11246_ (
);

NOR2X1 _15809_ (
    .A(_6267_),
    .B(_6270_),
    .Y(_6271_)
);

FILL FILL_0__10659_ (
);

AOI21X1 _10944_ (
    .A(_2055_),
    .B(_2059_),
    .C(IRWrite_bF$buf2),
    .Y(_2078_)
);

FILL FILL_0__8253_ (
);

FILL FILL_0__10239_ (
);

OAI21X1 _10524_ (
    .A(_1846_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1847_),
    .Y(_1823_[12])
);

OAI21X1 _10104_ (
    .A(_1691_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1692_),
    .Y(_1628_[0])
);

FILL FILL_4__15892_ (
);

FILL FILL_4__15472_ (
);

FILL FILL_4__15052_ (
);

FILL FILL_2__9632_ (
);

FILL FILL_3__14885_ (
);

FILL FILL_3__14465_ (
);

FILL FILL_2__9212_ (
);

FILL FILL_0__11600_ (
);

FILL FILL_3__14045_ (
);

FILL FILL_4__9978_ (
);

FILL FILL_4__9138_ (
);

FILL FILL_2__13878_ (
);

FILL FILL_2__13458_ (
);

FILL FILL_0__14492_ (
);

FILL FILL_2__13038_ (
);

FILL FILL_0__14072_ (
);

FILL FILL_3__7975_ (
);

FILL FILL_0__9878_ (
);

FILL FILL_3__7555_ (
);

FILL FILL_0__9038_ (
);

OAI21X1 _11729_ (
    .A(_2197_),
    .B(_2388_),
    .C(_2825_),
    .Y(_2826_)
);

INVX1 _11309_ (
    .A(_2427_),
    .Y(_2428_)
);

FILL FILL_1__13812_ (
);

FILL FILL_4__16257_ (
);

FILL FILL_4__11392_ (
);

FILL FILL_1__16284_ (
);

FILL FILL_5__8842_ (
);

FILL FILL_3__10385_ (
);

FILL FILL_5__8002_ (
);

NOR2X1 _15982_ (
    .A(_6438_),
    .B(_6437_),
    .Y(_6439_)
);

FILL FILL_0__15697_ (
);

OAI22X1 _15562_ (
    .A(_4525_),
    .B(_5545__bF$buf1),
    .C(_5548__bF$buf2),
    .D(_6029_),
    .Y(_6030_)
);

FILL FILL_0__15277_ (
);

NOR2X1 _15142_ (
    .A(_5619_),
    .B(_5617_),
    .Y(_5620_)
);

FILL FILL_1__8834_ (
);

FILL SFILL8680x49050 (
);

FILL FILL_6__14191_ (
);

FILL FILL_2__15604_ (
);

FILL SFILL88600x74050 (
);

FILL SFILL27960x58050 (
);

NAND2X1 _7484_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_309_)
);

NAND2X1 _7064_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_90_)
);

FILL FILL_4__12597_ (
);

FILL FILL_4__12177_ (
);

FILL FILL_5__9627_ (
);

FILL FILL_5__9207_ (
);

OAI21X1 _16347_ (
    .A(_6784_),
    .B(gnd),
    .C(_6785_),
    .Y(_6769_[8])
);

NAND2X1 _11482_ (
    .A(_2285_),
    .B(_2341__bF$buf2),
    .Y(_2596_)
);

FILL FILL_0__11197_ (
);

FILL FILL_5__11917_ (
);

XNOR2X1 _11062_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2181_)
);

FILL FILL_3__12951_ (
);

FILL FILL_1__9619_ (
);

FILL SFILL8600x47050 (
);

FILL FILL_3__12531_ (
);

FILL FILL_3__12111_ (
);

FILL FILL_4__7624_ (
);

FILL FILL_4__7204_ (
);

FILL FILL_2__11944_ (
);

FILL SFILL13240x79050 (
);

FILL FILL_5__14389_ (
);

FILL FILL_2__11524_ (
);

FILL FILL_2__11104_ (
);

DFFSR _8689_ (
    .Q(\datapath_1.regfile_1.regOut[14] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_848_[27])
);

INVX1 _8269_ (
    .A(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_710_)
);

FILL FILL_1__10937_ (
);

FILL FILL_1__10517_ (
);

FILL SFILL84200x28050 (
);

FILL FILL_5__15750_ (
);

FILL FILL_0__7944_ (
);

FILL FILL_5__15330_ (
);

FILL FILL_0__7104_ (
);

NAND2X1 _9630_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1394_)
);

FILL SFILL48440x40050 (
);

NAND2X1 _9210_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1175_)
);

FILL FILL_4__14743_ (
);

FILL FILL_4__14323_ (
);

DFFSR _12687_ (
    .Q(\datapath_1.Data [24]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_3425_[24])
);

FILL FILL_3__8093_ (
);

NAND3X1 _12267_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3239_)
);

FILL FILL_2__8903_ (
);

FILL FILL_3__13736_ (
);

FILL FILL_3__13316_ (
);

FILL FILL_1__14770_ (
);

FILL FILL_1__14350_ (
);

FILL FILL_4__8829_ (
);

FILL FILL_2__12729_ (
);

FILL FILL_0__13763_ (
);

FILL FILL_2__12309_ (
);

FILL FILL_0__13343_ (
);

FILL FILL_5__9380_ (
);

FILL FILL_1__6900_ (
);

FILL FILL_0__8729_ (
);

FILL FILL_5__16115_ (
);

FILL FILL_1__9792_ (
);

FILL FILL_5__11670_ (
);

FILL SFILL74280x28050 (
);

FILL FILL_1__9372_ (
);

FILL FILL_5__11250_ (
);

FILL FILL_4__15948_ (
);

FILL FILL_4__15528_ (
);

FILL FILL_4__15108_ (
);

FILL FILL_2__16142_ (
);

FILL FILL_3__9298_ (
);

FILL FILL_4__10663_ (
);

FILL FILL_4__10243_ (
);

FILL FILL_1__15975_ (
);

FILL FILL_1__15555_ (
);

FILL FILL_1__15135_ (
);

FILL FILL_1__10690_ (
);

FILL FILL_1__10270_ (
);

FILL FILL_0__14968_ (
);

NOR2X1 _14833_ (
    .A(_5316_),
    .B(_5306_),
    .Y(_5317_)
);

FILL FILL_0__14548_ (
);

FILL FILL_0__14128_ (
);

AOI22X1 _14413_ (
    .A(_3950__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [20]),
    .C(\datapath_1.regfile_1.regOut[27] [20]),
    .D(_4129_),
    .Y(_4905_)
);

FILL FILL_2__7295_ (
);

FILL FILL_6__13042_ (
);

FILL FILL_5__12875_ (
);

FILL SFILL74200x26050 (
);

FILL FILL_5__12455_ (
);

FILL FILL_5__12035_ (
);

FILL FILL_4__8582_ (
);

FILL FILL_4__11868_ (
);

FILL FILL_4__11448_ (
);

FILL FILL_2__12482_ (
);

FILL FILL_4__11028_ (
);

FILL FILL_2__12062_ (
);

FILL FILL_1__11895_ (
);

FILL FILL_1__11475_ (
);

FILL SFILL99480x32050 (
);

FILL FILL_1__11055_ (
);

NAND3X1 _15618_ (
    .A(_6082_),
    .B(_6083_),
    .C(_6081_),
    .Y(_6084_)
);

FILL FILL_0__8482_ (
);

FILL FILL_0__10888_ (
);

OAI21X1 _10753_ (
    .A(_1958_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .C(_1959_),
    .Y(_1953_[3])
);

FILL FILL_0__8062_ (
);

FILL SFILL3480x51050 (
);

DFFSR _10333_ (
    .Q(\datapath_1.regfile_1.regOut[27] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_1693_[7])
);

FILL FILL_0__10048_ (
);

FILL FILL_3__11802_ (
);

FILL FILL_6__14667_ (
);

FILL FILL_6__14247_ (
);

FILL FILL_4__15281_ (
);

FILL SFILL33800x78050 (
);

FILL FILL_2__9861_ (
);

FILL SFILL64200x69050 (
);

FILL FILL_3__14694_ (
);

FILL FILL_2__9021_ (
);

FILL FILL_3__14274_ (
);

FILL FILL112120x46050 (
);

FILL FILL_4__9787_ (
);

FILL FILL_4__9367_ (
);

FILL FILL_2__13687_ (
);

FILL FILL_2__13267_ (
);

FILL FILL_5__14601_ (
);

NAND2X1 _8901_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1030_)
);

OAI21X1 _11958_ (
    .A(_3012_),
    .B(IorD_bF$buf5),
    .C(_3013_),
    .Y(_1_[23])
);

FILL FILL_3__7364_ (
);

FILL FILL_0__9267_ (
);

AOI21X1 _11538_ (
    .A(_2552_),
    .B(_2648_),
    .C(_2410_),
    .Y(_2649_)
);

NOR2X1 _11118_ (
    .A(_2231_),
    .B(_2236_),
    .Y(_2237_)
);

FILL FILL_1__13621_ (
);

FILL FILL_4__16066_ (
);

FILL FILL_3__15899_ (
);

FILL FILL_0__12614_ (
);

FILL FILL_3__15479_ (
);

FILL FILL_3__15059_ (
);

FILL SFILL89400x6050 (
);

FILL FILL_1__16093_ (
);

FILL SFILL33800x33050 (
);

FILL FILL_5__8651_ (
);

FILL SFILL64200x24050 (
);

FILL FILL_5__8231_ (
);

FILL FILL_3__10194_ (
);

FILL FILL_6_BUFX2_insert853 (
);

INVX1 _15791_ (
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_6253_)
);

NAND3X1 _15371_ (
    .A(_5840_),
    .B(_5843_),
    .C(_5835_),
    .Y(_5844_)
);

FILL FILL_0__15086_ (
);

FILL FILL_5__15806_ (
);

FILL FILL_6_BUFX2_insert858 (
);

FILL FILL_3__16000_ (
);

FILL FILL_5__10941_ (
);

FILL FILL_5__10521_ (
);

FILL FILL_1__8643_ (
);

FILL FILL_1__8223_ (
);

FILL FILL_2__15833_ (
);

FILL FILL_2__15413_ (
);

FILL FILL_3__8989_ (
);

FILL FILL_3__8569_ (
);

FILL FILL_3__8149_ (
);

FILL FILL_1__14826_ (
);

NAND2X1 _7293_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_202_)
);

FILL FILL_1__14406_ (
);

FILL FILL_3__9930_ (
);

FILL FILL_0__13819_ (
);

FILL FILL_3__9510_ (
);

FILL FILL_2__6986_ (
);

FILL FILL_5__9856_ (
);

FILL FILL_3__11399_ (
);

FILL FILL_5__9016_ (
);

FILL FILL_6__12733_ (
);

NOR2X1 _16156_ (
    .A(_6607_),
    .B(_6608_),
    .Y(_6609_)
);

NAND2X1 _11291_ (
    .A(_2218_),
    .B(_2409_),
    .Y(_2410_)
);

FILL FILL_1__9848_ (
);

FILL FILL_5__11726_ (
);

FILL FILL_3__12760_ (
);

FILL FILL_1__9428_ (
);

FILL FILL_5__11306_ (
);

FILL FILL_1__9008_ (
);

FILL FILL_3__12340_ (
);

FILL FILL_4__7853_ (
);

FILL FILL_4__7433_ (
);

FILL FILL_2__11753_ (
);

FILL FILL_5__14198_ (
);

FILL FILL_2__11333_ (
);

INVX1 _8498_ (
    .A(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_822_)
);

INVX1 _8078_ (
    .A(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_603_)
);

FILL FILL_1__10746_ (
);

FILL FILL_0__7753_ (
);

FILL FILL_0__7333_ (
);

FILL FILL_4__14972_ (
);

FILL FILL_4__14552_ (
);

FILL FILL_4__14132_ (
);

INVX1 _12496_ (
    .A(ALUOut[19]),
    .Y(_3397_)
);

NAND3X1 _12076_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump_22_bF$buf3 ),
    .C(_3034__bF$buf2),
    .Y(_3103_)
);

FILL FILL_2__8712_ (
);

FILL FILL_3__13965_ (
);

FILL FILL_3__13545_ (
);

FILL FILL_3__13125_ (
);

FILL FILL_4__8638_ (
);

FILL FILL_4__8218_ (
);

FILL FILL_5_BUFX2_insert870 (
);

FILL FILL_5_BUFX2_insert871 (
);

FILL FILL_2__12958_ (
);

FILL FILL_0__13992_ (
);

FILL FILL_5_BUFX2_insert872 (
);

FILL FILL_2__12118_ (
);

FILL FILL_5_BUFX2_insert873 (
);

FILL FILL_0__13572_ (
);

FILL FILL_0__13152_ (
);

FILL FILL_5_BUFX2_insert874 (
);

FILL FILL_5_BUFX2_insert875 (
);

FILL FILL_5_BUFX2_insert876 (
);

FILL FILL_5_BUFX2_insert877 (
);

FILL FILL_5_BUFX2_insert878 (
);

FILL FILL_5_BUFX2_insert879 (
);

FILL SFILL23720x38050 (
);

FILL FILL_5__16344_ (
);

FILL FILL_0__8958_ (
);

FILL FILL_0__8118_ (
);

NAND2X1 _10809_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1997_)
);

FILL FILL_4__15757_ (
);

FILL FILL_4__15337_ (
);

FILL FILL_2__16371_ (
);

FILL FILL_4__10892_ (
);

FILL FILL_2__9917_ (
);

FILL FILL_4__10052_ (
);

FILL FILL_1__15784_ (
);

FILL FILL_1__15364_ (
);

FILL SFILL59800x6050 (
);

FILL FILL_5__7502_ (
);

FILL FILL_0__14777_ (
);

INVX1 _14642_ (
    .A(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_5130_)
);

FILL FILL_0__14357_ (
);

INVX1 _14222_ (
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_4718_)
);

FILL FILL_5__12264_ (
);

NAND2X1 _6984_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_57_)
);

FILL FILL_4__8391_ (
);

FILL FILL_4__11677_ (
);

FILL FILL_4__11257_ (
);

FILL FILL_2__12291_ (
);

FILL FILL_1__16149_ (
);

FILL FILL_5__8707_ (
);

FILL FILL_1__11284_ (
);

INVX1 _15847_ (
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_6308_)
);

AOI22X1 _15427_ (
    .A(\datapath_1.regfile_1.regOut[1] [9]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_5898_)
);

AOI22X1 _15007_ (
    .A(_5486_),
    .B(\datapath_1.regfile_1.regOut[29] [0]),
    .C(\datapath_1.regfile_1.regOut[26] [0]),
    .D(_5484_),
    .Y(_5487_)
);

NAND2X1 _10982_ (
    .A(vdd),
    .B(\control_1.next [3]),
    .Y(_2106_)
);

FILL FILL_0__10697_ (
);

FILL FILL_0__10277_ (
);

NAND2X1 _10562_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1873_)
);

NAND2X1 _10142_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1654_)
);

FILL FILL_3__11611_ (
);

FILL FILL_4__15090_ (
);

FILL SFILL48840x49050 (
);

FILL FILL_5__13889_ (
);

FILL FILL_5__13469_ (
);

FILL FILL_2__9670_ (
);

FILL FILL_2__9250_ (
);

DFFSR _7769_ (
    .Q(\datapath_1.regfile_1.regOut[7] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_393_[3])
);

FILL FILL_3__14083_ (
);

FILL SFILL109560x16050 (
);

INVX1 _7349_ (
    .A(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_239_)
);

FILL FILL_4__9596_ (
);

FILL SFILL109400x5050 (
);

FILL FILL_2__13496_ (
);

FILL FILL_5__14830_ (
);

FILL FILL_5__14410_ (
);

FILL SFILL48440x35050 (
);

NAND2X1 _8710_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_923_)
);

FILL FILL_1__12489_ (
);

FILL FILL_1__12069_ (
);

FILL FILL_4__13823_ (
);

FILL FILL_4__13403_ (
);

FILL FILL_0__9496_ (
);

FILL FILL_3__7593_ (
);

INVX1 _11767_ (
    .A(_2372_),
    .Y(_2862_)
);

FILL FILL_3__7173_ (
);

NAND2X1 _11347_ (
    .A(_2115_),
    .B(_2341__bF$buf2),
    .Y(_2465_)
);

FILL FILL_1__13850_ (
);

FILL FILL_5__7099_ (
);

FILL FILL_1__13430_ (
);

FILL FILL_4__16295_ (
);

FILL FILL_1__13010_ (
);

FILL FILL_2__11809_ (
);

FILL FILL_0__12843_ (
);

FILL FILL_0__12423_ (
);

FILL FILL_3__15288_ (
);

FILL FILL_0__12003_ (
);

FILL FILL_5__8880_ (
);

FILL FILL_5__8460_ (
);

OAI22X1 _15180_ (
    .A(_4122_),
    .B(_5503__bF$buf0),
    .C(_5463__bF$buf3),
    .D(_5656_),
    .Y(_5657_)
);

FILL FILL_5__15615_ (
);

FILL FILL_0__7809_ (
);

INVX1 _9915_ (
    .A(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_1543_)
);

FILL FILL_1__8872_ (
);

FILL FILL_5__10750_ (
);

FILL FILL_1__8452_ (
);

FILL FILL_4__14608_ (
);

FILL FILL_2__15642_ (
);

FILL FILL_2__15222_ (
);

FILL FILL_3__8378_ (
);

FILL FILL_1__14635_ (
);

FILL FILL_1__14215_ (
);

FILL FILL_0__13628_ (
);

OAI22X1 _13913_ (
    .A(_4414_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf0),
    .D(_4415_),
    .Y(_4416_)
);

FILL FILL_0__13208_ (
);

FILL SFILL38840x47050 (
);

FILL FILL_5__9665_ (
);

FILL FILL_5__9245_ (
);

NAND2X1 _16385_ (
    .A(gnd),
    .B(gnd),
    .Y(_6811_)
);

FILL SFILL28920x83050 (
);

FILL FILL_5__11955_ (
);

FILL FILL_1__9657_ (
);

FILL FILL_5__11535_ (
);

FILL FILL_1__9237_ (
);

FILL FILL_5__11115_ (
);

FILL FILL_2__16007_ (
);

FILL FILL_4__10948_ (
);

FILL FILL_4__7242_ (
);

FILL FILL_4__10528_ (
);

FILL FILL_2__11982_ (
);

FILL FILL_2__11562_ (
);

FILL FILL_4__10108_ (
);

FILL FILL_2__11142_ (
);

FILL FILL112200x34050 (
);

FILL FILL_1__10975_ (
);

FILL SFILL99480x27050 (
);

FILL FILL_1__10555_ (
);

FILL FILL_1__10135_ (
);

FILL FILL_0__7982_ (
);

FILL FILL_0__7562_ (
);

BUFX2 BUFX2_insert690 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf6 )
);

FILL SFILL3480x46050 (
);

BUFX2 BUFX2_insert691 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf5 )
);

BUFX2 BUFX2_insert692 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf4 )
);

BUFX2 BUFX2_insert693 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf3 )
);

BUFX2 BUFX2_insert694 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf2 )
);

BUFX2 BUFX2_insert695 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf1 )
);

FILL FILL_4__14781_ (
);

BUFX2 BUFX2_insert696 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf0 )
);

FILL FILL_4__14361_ (
);

BUFX2 BUFX2_insert697 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf4 )
);

BUFX2 BUFX2_insert698 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf3 )
);

FILL SFILL69240x1050 (
);

BUFX2 BUFX2_insert699 (
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf2 )
);

FILL FILL_3__13774_ (
);

FILL FILL_2__8521_ (
);

FILL FILL_3__13354_ (
);

FILL FILL_2__8101_ (
);

FILL FILL_4__8867_ (
);

FILL FILL_4__8447_ (
);

FILL FILL_2__12767_ (
);

FILL FILL_2__12347_ (
);

FILL FILL_0__13381_ (
);

FILL FILL_0__8767_ (
);

FILL FILL_3__6864_ (
);

FILL FILL_5__16153_ (
);

FILL FILL_0__8347_ (
);

NAND2X1 _10618_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1890_)
);

FILL FILL_4__15986_ (
);

FILL FILL_1__12701_ (
);

FILL FILL_4__15566_ (
);

FILL FILL_4__15146_ (
);

FILL FILL_2__16180_ (
);

FILL FILL_4__10281_ (
);

FILL FILL_3__14979_ (
);

FILL FILL_2__9726_ (
);

FILL FILL_3__14559_ (
);

FILL FILL_3__14139_ (
);

FILL FILL_1__15593_ (
);

FILL FILL_1__15173_ (
);

FILL SFILL64200x19050 (
);

FILL FILL_5__7731_ (
);

FILL FILL_5__7311_ (
);

INVX1 _14871_ (
    .A(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_5354_)
);

FILL FILL_0__14586_ (
);

INVX1 _14451_ (
    .A(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_4942_)
);

FILL FILL_0__14166_ (
);

NOR2X1 _14031_ (
    .A(_4530_),
    .B(_4527_),
    .Y(_4531_)
);

FILL FILL_3__15920_ (
);

FILL FILL_3__15500_ (
);

FILL FILL_1__7723_ (
);

FILL FILL_1__7303_ (
);

FILL FILL_2__14913_ (
);

FILL FILL_3__7229_ (
);

FILL FILL_5__12493_ (
);

FILL FILL_5__12073_ (
);

FILL FILL_1__13906_ (
);

FILL FILL_4__11486_ (
);

FILL FILL_4__11066_ (
);

FILL FILL_1__16378_ (
);

FILL FILL_3__10899_ (
);

FILL FILL_5__8516_ (
);

FILL FILL_3__10059_ (
);

FILL FILL_1__11093_ (
);

NOR3X1 _15656_ (
    .A(_6120_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6121_)
);

OAI22X1 _15236_ (
    .A(_5480__bF$buf3),
    .B(_5711_),
    .C(_4187_),
    .D(_5569_),
    .Y(_5712_)
);

NAND2X1 _10791_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1985_)
);

NAND2X1 _10371_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1766_)
);

FILL FILL_5__10806_ (
);

FILL FILL_1__8508_ (
);

FILL FILL_3__11840_ (
);

FILL FILL_3__11420_ (
);

FILL FILL_3__11000_ (
);

FILL FILL_4__6933_ (
);

FILL SFILL63880x83050 (
);

FILL SFILL79480x68050 (
);

FILL FILL_0__16312_ (
);

FILL FILL_2__10833_ (
);

FILL FILL_5__13698_ (
);

FILL FILL_5__13278_ (
);

FILL FILL_2__10413_ (
);

INVX1 _7998_ (
    .A(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_570_)
);

INVX1 _7578_ (
    .A(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_351_)
);

INVX1 _7158_ (
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .Y(_196_)
);

FILL SFILL18840x43050 (
);

FILL FILL_1__12298_ (
);

FILL FILL_4__13632_ (
);

FILL FILL_4__13212_ (
);

NAND3X1 _11996_ (
    .A(PCSource_1_bF$buf2),
    .B(\aluControl_1.inst [0]),
    .C(_3034__bF$buf4),
    .Y(_3043_)
);

AND2X2 _11576_ (
    .A(_2659_),
    .B(_2670_),
    .Y(_2684_)
);

AND2X2 _11156_ (
    .A(_2270_),
    .B(_2274_),
    .Y(_2275_)
);

FILL FILL_3__12625_ (
);

FILL FILL_3__12205_ (
);

FILL FILL_4__7718_ (
);

FILL FILL_2__11618_ (
);

FILL FILL_0__12652_ (
);

FILL FILL_3__15097_ (
);

FILL FILL_0__12232_ (
);

FILL FILL_5__15844_ (
);

FILL SFILL38840x8050 (
);

FILL FILL_5__15424_ (
);

FILL FILL_5__15004_ (
);

FILL FILL_0__7618_ (
);

INVX1 _9724_ (
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_1436_)
);

DFFSR _9304_ (
    .Q(\datapath_1.regfile_1.regOut[19] [2]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_1173_[2])
);

FILL FILL_1__8261_ (
);

FILL FILL_4__14837_ (
);

FILL FILL_4__14417_ (
);

FILL FILL_2__15871_ (
);

FILL FILL_2__15451_ (
);

FILL FILL_2__15031_ (
);

FILL FILL_3__8187_ (
);

FILL FILL_1__14864_ (
);

FILL FILL_1__14444_ (
);

FILL FILL_1__14024_ (
);

FILL FILL_0__13857_ (
);

FILL FILL_0__13437_ (
);

OAI22X1 _13722_ (
    .A(_4227_),
    .B(_3910_),
    .C(_3978_),
    .D(_4228_),
    .Y(_4229_)
);

OAI21X1 _13302_ (
    .A(_3752_),
    .B(_3764_),
    .C(_3754_),
    .Y(_3837_)
);

FILL FILL_0__13017_ (
);

FILL FILL_5__9894_ (
);

FILL FILL_5__9474_ (
);

FILL FILL_6__12351_ (
);

OAI21X1 _16194_ (
    .A(_5527__bF$buf1),
    .B(_5282_),
    .C(_6645_),
    .Y(_6646_)
);

FILL FILL_5__16209_ (
);

FILL FILL_5__11764_ (
);

FILL FILL_1__9886_ (
);

FILL FILL_1__9466_ (
);

FILL FILL_5__11344_ (
);

FILL SFILL69080x52050 (
);

FILL FILL_2__16236_ (
);

FILL FILL_4__7891_ (
);

FILL FILL_4__7471_ (
);

FILL FILL_4__7051_ (
);

FILL FILL_4__10757_ (
);

FILL SFILL48920x37050 (
);

FILL FILL_2__11791_ (
);

FILL FILL_2__11371_ (
);

FILL FILL_1__15649_ (
);

FILL FILL_1__15229_ (
);

FILL FILL_1__10784_ (
);

FILL FILL_1__10364_ (
);

NAND3X1 _14927_ (
    .A(_5407_),
    .B(_5408_),
    .C(_5406_),
    .Y(_5409_)
);

NOR2X1 _14507_ (
    .A(_4993_),
    .B(_4996_),
    .Y(_4997_)
);

FILL FILL_0__7371_ (
);

FILL FILL_6__13976_ (
);

FILL SFILL69480x21050 (
);

FILL FILL_6__13556_ (
);

FILL FILL_4__14590_ (
);

FILL FILL_6__13136_ (
);

FILL FILL_4__14170_ (
);

FILL FILL_5__12969_ (
);

FILL FILL_2__8750_ (
);

FILL FILL_2__8330_ (
);

FILL FILL_5__12129_ (
);

FILL FILL_3__13583_ (
);

FILL FILL_3__13163_ (
);

BUFX2 _6849_ (
    .A(_1_[11]),
    .Y(memoryAddress[11])
);

FILL FILL_4__8256_ (
);

FILL FILL_2__12996_ (
);

FILL FILL_2__12576_ (
);

FILL FILL_2__12156_ (
);

FILL FILL_5__13910_ (
);

FILL FILL_1__11989_ (
);

FILL FILL_1__11569_ (
);

FILL FILL_1__11149_ (
);

FILL FILL_4__12903_ (
);

FILL FILL_5__16382_ (
);

FILL FILL_0__8996_ (
);

FILL FILL_0__8576_ (
);

DFFSR _10847_ (
    .Q(\datapath_1.regfile_1.regOut[31] [9]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_1953_[9])
);

INVX1 _10427_ (
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_1803_)
);

INVX1 _10007_ (
    .A(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_1584_)
);

FILL FILL_4__15795_ (
);

FILL FILL_4__15375_ (
);

FILL FILL_1__12510_ (
);

FILL FILL_2__9535_ (
);

FILL FILL_0__11923_ (
);

FILL FILL_3__14788_ (
);

FILL FILL_2__9115_ (
);

FILL FILL_3__14368_ (
);

FILL FILL_0__11503_ (
);

FILL FILL_5__7960_ (
);

FILL FILL_5__7120_ (
);

FILL SFILL3560x79050 (
);

FILL SFILL59080x50050 (
);

FILL FILL_0__14395_ (
);

NAND3X1 _14680_ (
    .A(_5156_),
    .B(_5159_),
    .C(_5166_),
    .Y(_5167_)
);

NOR2X1 _14260_ (
    .A(_4752_),
    .B(_4755_),
    .Y(_4756_)
);

FILL SFILL38920x35050 (
);

FILL SFILL34200x13050 (
);

FILL FILL_1__7952_ (
);

FILL FILL_1__7112_ (
);

FILL FILL_2__14722_ (
);

FILL FILL_3__7878_ (
);

FILL FILL_2__14302_ (
);

FILL FILL_3__7458_ (
);

FILL FILL_3__7038_ (
);

FILL FILL_1__13715_ (
);

FILL FILL_4__11295_ (
);

FILL FILL_0__12708_ (
);

FILL FILL_1__16187_ (
);

FILL FILL_5__8745_ (
);

FILL FILL_3__10288_ (
);

FILL FILL_5__8325_ (
);

FILL SFILL99560x15050 (
);

INVX1 _15885_ (
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_6345_)
);

NOR2X1 _15465_ (
    .A(_5933_),
    .B(_5934_),
    .Y(_5935_)
);

OAI22X1 _15045_ (
    .A(_5523_),
    .B(_3908_),
    .C(_3976_),
    .D(_5524__bF$buf0),
    .Y(_5525_)
);

FILL SFILL28920x78050 (
);

FILL SFILL3560x34050 (
);

INVX1 _10180_ (
    .A(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_1679_)
);

FILL FILL_1__8737_ (
);

FILL FILL_5__10615_ (
);

FILL FILL_1__8317_ (
);

FILL FILL_6__14094_ (
);

FILL FILL_2__15927_ (
);

FILL SFILL104440x51050 (
);

FILL FILL_2__15507_ (
);

FILL FILL_0__16121_ (
);

FILL FILL_2__10642_ (
);

FILL FILL_5__13087_ (
);

DFFSR _7387_ (
    .Q(\datapath_1.regfile_1.regOut[4] [5]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_198_[5])
);

FILL FILL112200x29050 (
);

FILL FILL_3__9604_ (
);

FILL FILL_4__13861_ (
);

FILL FILL_4__13441_ (
);

FILL FILL_4__13021_ (
);

AOI21X1 _11385_ (
    .A(_2497_),
    .B(_2499_),
    .C(_2501_),
    .Y(_2502_)
);

FILL FILL_2__7601_ (
);

FILL FILL_3__12854_ (
);

FILL FILL_3__12434_ (
);

FILL FILL_3__12014_ (
);

FILL SFILL28920x33050 (
);

FILL FILL_4__7947_ (
);

FILL FILL_4__7107_ (
);

FILL FILL_2__11847_ (
);

FILL FILL_0__12881_ (
);

FILL FILL_2__11427_ (
);

FILL FILL_0__12461_ (
);

FILL FILL_2__11007_ (
);

FILL FILL_0__12041_ (
);

FILL FILL_5__15653_ (
);

FILL FILL_0__7847_ (
);

FILL FILL_5__15233_ (
);

FILL FILL_0__7427_ (
);

DFFSR _9953_ (
    .Q(\datapath_1.regfile_1.regOut[24] [11]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1498_[11])
);

OAI21X1 _9533_ (
    .A(_1348_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1349_),
    .Y(_1303_[23])
);

OAI21X1 _9113_ (
    .A(_1129_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1130_),
    .Y(_1108_[11])
);

FILL FILL_1__8490_ (
);

FILL FILL_1__8070_ (
);

FILL FILL_4__14646_ (
);

FILL FILL_2__15680_ (
);

FILL FILL_4__14226_ (
);

FILL FILL_2__15260_ (
);

FILL FILL_3__13639_ (
);

FILL FILL_3__13219_ (
);

FILL FILL_1__14673_ (
);

FILL FILL_1__14253_ (
);

FILL FILL_0_BUFX2_insert330 (
);

FILL FILL_0_BUFX2_insert331 (
);

FILL FILL_0_BUFX2_insert332 (
);

FILL FILL_0_BUFX2_insert333 (
);

FILL FILL_0__13666_ (
);

FILL FILL_0_BUFX2_insert334 (
);

AOI22X1 _13951_ (
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .B(_4225_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_4453_)
);

FILL FILL_0__13246_ (
);

FILL FILL_0_BUFX2_insert335 (
);

NAND3X1 _13531_ (
    .A(_4039_),
    .B(_4041_),
    .C(_4037_),
    .Y(_4042_)
);

OAI21X1 _13111_ (
    .A(_3704_),
    .B(PCEn_bF$buf2),
    .C(_3705_),
    .Y(_3685_[10])
);

FILL FILL_0_BUFX2_insert336 (
);

FILL FILL_0_BUFX2_insert337 (
);

FILL FILL_0_BUFX2_insert338 (
);

FILL FILL_0_BUFX2_insert339 (
);

FILL FILL_5__9283_ (
);

FILL FILL_5__16018_ (
);

FILL FILL_5__11993_ (
);

FILL FILL_5__11573_ (
);

FILL SFILL28040x12050 (
);

FILL FILL_1__9275_ (
);

FILL FILL_5__11153_ (
);

FILL FILL_2__16045_ (
);

FILL SFILL63960x71050 (
);

FILL FILL_4__10566_ (
);

FILL SFILL94360x62050 (
);

FILL FILL_4__10146_ (
);

FILL FILL_2__11180_ (
);

FILL FILL_1__15878_ (
);

FILL FILL_1__15458_ (
);

FILL FILL_1__15038_ (
);

FILL FILL_1__10173_ (
);

FILL SFILL18920x31050 (
);

OAI22X1 _14736_ (
    .A(_5221_),
    .B(_3941_),
    .C(_3966__bF$buf0),
    .D(_5220_),
    .Y(_5222_)
);

INVX1 _14316_ (
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_4810_)
);

FILL SFILL58200x44050 (
);

FILL FILL_0__7180_ (
);

FILL FILL_2_BUFX2_insert10 (
);

FILL FILL_2__7198_ (
);

FILL FILL_2_BUFX2_insert11 (
);

FILL FILL_2_BUFX2_insert12 (
);

FILL FILL_3__10920_ (
);

FILL FILL_2_BUFX2_insert13 (
);

FILL FILL_3__10500_ (
);

FILL FILL_2_BUFX2_insert14 (
);

FILL FILL_2_BUFX2_insert15 (
);

FILL FILL_2_BUFX2_insert16 (
);

FILL FILL_2_BUFX2_insert17 (
);

FILL FILL_0__15812_ (
);

FILL SFILL94760x31050 (
);

FILL FILL_2_BUFX2_insert18 (
);

FILL FILL_2_BUFX2_insert19 (
);

FILL FILL_5__12778_ (
);

FILL FILL_5__12358_ (
);

FILL FILL_3__13392_ (
);

FILL FILL_4__8485_ (
);

FILL SFILL18680x3050 (
);

FILL FILL_4__8065_ (
);

FILL SFILL18840x38050 (
);

FILL FILL_2__12385_ (
);

FILL FILL_1__11798_ (
);

FILL FILL_1__11378_ (
);

FILL FILL_4__12712_ (
);

FILL FILL_5__16191_ (
);

FILL FILL_6__9772_ (
);

FILL FILL_0__8385_ (
);

INVX1 _10656_ (
    .A(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_1915_)
);

INVX1 _10236_ (
    .A(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_1696_)
);

FILL FILL_3__11705_ (
);

FILL FILL_4__15184_ (
);

FILL FILL_2__9764_ (
);

FILL FILL_2__9344_ (
);

FILL FILL_3__14597_ (
);

FILL FILL_0__11732_ (
);

FILL FILL_3__14177_ (
);

FILL FILL_0__11312_ (
);

FILL FILL_6__15511_ (
);

FILL FILL_5__14924_ (
);

FILL FILL_5__14504_ (
);

DFFSR _8804_ (
    .Q(\datapath_1.regfile_1.regOut[15] [14]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_913_[14])
);

FILL FILL_1__7761_ (
);

FILL FILL_1__7341_ (
);

FILL FILL_4__13917_ (
);

FILL FILL_2__14951_ (
);

FILL FILL_2__14531_ (
);

FILL FILL_3__7687_ (
);

FILL FILL_2__14111_ (
);

FILL FILL_1__13944_ (
);

FILL FILL_4__16389_ (
);

FILL FILL_1__13524_ (
);

FILL FILL_1__13104_ (
);

DFFSR _12802_ (
    .Q(\datapath_1.PCJump [13]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3490_[11])
);

FILL FILL_0__12517_ (
);

FILL SFILL53880x76050 (
);

FILL FILL_5__8974_ (
);

FILL FILL_5__8134_ (
);

NOR2X1 _15694_ (
    .A(_6156_),
    .B(_6157_),
    .Y(_6158_)
);

FILL FILL_6__11431_ (
);

FILL FILL_6__11011_ (
);

NOR2X1 _15274_ (
    .A(_5748_),
    .B(_5740_),
    .Y(_5749_)
);

FILL FILL_5__15709_ (
);

FILL FILL_3__16323_ (
);

FILL FILL_1__8966_ (
);

FILL FILL_5__10424_ (
);

FILL FILL_1__8126_ (
);

FILL FILL_5__10004_ (
);

FILL SFILL69080x47050 (
);

FILL FILL_2__15736_ (
);

FILL FILL_4__6971_ (
);

FILL FILL_2__15316_ (
);

FILL FILL_0__16350_ (
);

FILL FILL_2__10871_ (
);

FILL FILL_2__10451_ (
);

FILL FILL_2__10031_ (
);

FILL FILL_1__14729_ (
);

OAI21X1 _7196_ (
    .A(_156_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .C(_157_),
    .Y(_133_[12])
);

FILL FILL_1__14309_ (
);

FILL FILL_3__9413_ (
);

FILL FILL_2__6889_ (
);

FILL FILL_0__6871_ (
);

FILL FILL_5__9759_ (
);

FILL FILL_5__9339_ (
);

FILL SFILL114520x41050 (
);

FILL FILL_4__13670_ (
);

FILL FILL_4__13250_ (
);

NAND3X1 _16059_ (
    .A(_6502_),
    .B(_6513_),
    .C(_6508_),
    .Y(_6514_)
);

FILL SFILL3720x60050 (
);

NOR2X1 _11194_ (
    .A(\datapath_1.alu_1.ALUInB [26]),
    .B(_2312_),
    .Y(_2313_)
);

FILL FILL_5__11629_ (
);

FILL FILL_2__7830_ (
);

FILL FILL_5__11209_ (
);

FILL FILL_3__12243_ (
);

FILL FILL_4__7756_ (
);

FILL FILL_4__7336_ (
);

FILL FILL_2__11656_ (
);

FILL FILL_2__11236_ (
);

FILL FILL_0__12270_ (
);

FILL FILL_1__10649_ (
);

FILL FILL_5__15882_ (
);

FILL FILL_5__15462_ (
);

FILL FILL_5__15042_ (
);

OAI21X1 _9762_ (
    .A(_1460_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1461_),
    .Y(_1433_[14])
);

FILL FILL_0__7236_ (
);

OAI21X1 _9342_ (
    .A(_1241_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1242_),
    .Y(_1238_[2])
);

FILL SFILL43880x74050 (
);

FILL FILL_4__14875_ (
);

FILL FILL_4__14455_ (
);

FILL FILL_4__14035_ (
);

OAI21X1 _12399_ (
    .A(_3330_),
    .B(MemToReg_bF$buf6),
    .C(_3331_),
    .Y(\datapath_1.mux_wd3.dout [18])
);

FILL FILL_3__13868_ (
);

FILL FILL_2__8615_ (
);

FILL SFILL3560x5050 (
);

FILL FILL_3__13448_ (
);

FILL FILL_1__14482_ (
);

FILL FILL_3__13028_ (
);

FILL FILL_1__14062_ (
);

FILL SFILL59080x45050 (
);

FILL FILL_0__13895_ (
);

NAND3X1 _13760_ (
    .A(_4257_),
    .B(_4258_),
    .C(_4265_),
    .Y(_4266_)
);

FILL FILL_0__13475_ (
);

NOR2X1 _13340_ (
    .A(_3797_),
    .B(_3861_),
    .Y(\datapath_1.regfile_1.regEn [22])
);

FILL SFILL104920x53050 (
);

FILL FILL_5__9092_ (
);

FILL FILL_4__9902_ (
);

FILL FILL_2__13802_ (
);

FILL FILL_3__6958_ (
);

FILL FILL_5__16247_ (
);

FILL SFILL3640x22050 (
);

FILL FILL_5__11382_ (
);

FILL FILL_1__9084_ (
);

FILL FILL_2__16274_ (
);

FILL FILL_4__10795_ (
);

FILL FILL_4__10375_ (
);

FILL FILL_0__9802_ (
);

FILL FILL_1__15687_ (
);

FILL FILL_1__15267_ (
);

FILL FILL_5__7825_ (
);

AOI22X1 _14965_ (
    .A(\datapath_1.regfile_1.regOut[11] [31]),
    .B(_3950__bF$buf2),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_5446_)
);

OAI22X1 _14545_ (
    .A(_5034_),
    .B(_3971__bF$buf0),
    .C(_3924__bF$buf0),
    .D(_5033_),
    .Y(_5035_)
);

OAI22X1 _14125_ (
    .A(_4621_),
    .B(_3944__bF$buf3),
    .C(_3966__bF$buf0),
    .D(_4622_),
    .Y(_4623_)
);

FILL SFILL3560x29050 (
);

FILL FILL_1__7817_ (
);

FILL FILL_0__15621_ (
);

FILL FILL_0__15201_ (
);

FILL FILL_5__12587_ (
);

FILL FILL_5__12167_ (
);

BUFX2 _6887_ (
    .A(_2_[17]),
    .Y(memoryWriteData[17])
);

FILL SFILL33880x72050 (
);

FILL SFILL108760x54050 (
);

FILL FILL_2__12194_ (
);

FILL FILL_1__11187_ (
);

FILL FILL_4__12521_ (
);

FILL FILL_4__12101_ (
);

FILL SFILL28120x45050 (
);

FILL FILL_0__8194_ (
);

OR2X2 _10885_ (
    .A(\aluControl_1.inst [3]),
    .B(\aluControl_1.inst [2]),
    .Y(_2032_)
);

FILL SFILL49080x43050 (
);

DFFSR _10465_ (
    .Q(\datapath_1.regfile_1.regOut[28] [11]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_1758_[11])
);

OAI21X1 _10045_ (
    .A(_1608_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .C(_1609_),
    .Y(_1563_[23])
);

FILL FILL_3__11934_ (
);

FILL FILL_3__11514_ (
);

FILL SFILL28920x28050 (
);

FILL FILL_0__16406_ (
);

FILL SFILL89160x39050 (
);

FILL FILL_2__10927_ (
);

FILL FILL_2__9993_ (
);

FILL FILL_2__10507_ (
);

FILL FILL_0__11961_ (
);

FILL FILL_2__9153_ (
);

FILL FILL_0__11541_ (
);

FILL FILL_0__11121_ (
);

FILL FILL_4__9499_ (
);

FILL FILL_4__9079_ (
);

FILL FILL_2__13399_ (
);

FILL FILL_5__14733_ (
);

FILL FILL_0__6927_ (
);

FILL FILL_5__14313_ (
);

OAI21X1 _8613_ (
    .A(_877_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_878_),
    .Y(_848_[15])
);

FILL FILL_1__7990_ (
);

FILL FILL_1__7570_ (
);

FILL FILL_4__13726_ (
);

FILL FILL_4__13306_ (
);

FILL FILL_2__14760_ (
);

FILL FILL_2__14340_ (
);

FILL FILL_0__9399_ (
);

FILL FILL_3__7496_ (
);

FILL SFILL49000x41050 (
);

FILL FILL_3__7076_ (
);

FILL FILL_3__12719_ (
);

FILL FILL_1__13753_ (
);

FILL FILL_1__13333_ (
);

FILL FILL_4__16198_ (
);

FILL SFILL94440x50050 (
);

FILL FILL_0__12746_ (
);

OAI21X1 _12611_ (
    .A(_3452_),
    .B(vdd),
    .C(_3453_),
    .Y(_3425_[14])
);

FILL FILL_0__12326_ (
);

FILL FILL_5__8783_ (
);

FILL FILL_5__8363_ (
);

INVX2 _15083_ (
    .A(_5466__bF$buf2),
    .Y(_5562_)
);

FILL FILL_5__15938_ (
);

FILL FILL_5__15518_ (
);

FILL SFILL23880x70050 (
);

DFFSR _9818_ (
    .Q(\datapath_1.regfile_1.regOut[23] [4]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1433_[4])
);

FILL FILL_3__16132_ (
);

FILL FILL_1__8775_ (
);

FILL FILL_5__10653_ (
);

FILL FILL_1__8355_ (
);

FILL FILL_5__10233_ (
);

FILL FILL_2__15965_ (
);

FILL FILL_2__15545_ (
);

FILL FILL_2__15125_ (
);

FILL FILL_2__10680_ (
);

FILL FILL_2__10260_ (
);

FILL FILL_1__14958_ (
);

FILL FILL_1__14538_ (
);

FILL FILL_1__14118_ (
);

FILL SFILL18920x26050 (
);

FILL FILL_3__9642_ (
);

NOR2X1 _13816_ (
    .A(_4320_),
    .B(_4310_),
    .Y(_4321_)
);

FILL FILL_3__9222_ (
);

FILL FILL_5__9988_ (
);

FILL SFILL79160x37050 (
);

FILL FILL_5__9148_ (
);

NAND2X1 _16288_ (
    .A(\datapath_1.regfile_1.regOut[13] [31]),
    .B(_5576_),
    .Y(_6737_)
);

FILL SFILL39400x53050 (
);

FILL FILL_5__11858_ (
);

FILL FILL_3__12892_ (
);

FILL FILL_5__11438_ (
);

FILL FILL_3__12472_ (
);

FILL FILL_5__11018_ (
);

FILL FILL_3__12052_ (
);

FILL FILL_4__7985_ (
);

FILL FILL_4__7565_ (
);

FILL FILL_2__11885_ (
);

FILL FILL_2__11465_ (
);

FILL FILL_2__11045_ (
);

FILL SFILL94360x12050 (
);

FILL FILL_1__10878_ (
);

FILL FILL_1__10038_ (
);

FILL FILL_5__15691_ (
);

FILL FILL_0__7885_ (
);

FILL FILL_5__15271_ (
);

FILL FILL_0__7465_ (
);

OAI21X1 _9991_ (
    .A(_1572_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1573_),
    .Y(_1563_[5])
);

FILL FILL_6__8852_ (
);

FILL FILL_0__7045_ (
);

DFFSR _9571_ (
    .Q(\datapath_1.regfile_1.regOut[21] [13]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_1303_[13])
);

NAND2X1 _9151_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1156_)
);

FILL FILL_4__14684_ (
);

FILL FILL_4__14264_ (
);

FILL SFILL8760x74050 (
);

FILL FILL_2__8844_ (
);

FILL FILL_0__10812_ (
);

FILL FILL_3__13677_ (
);

FILL FILL_3__13257_ (
);

FILL FILL_2__8004_ (
);

FILL FILL_1__14291_ (
);

FILL FILL_0_BUFX2_insert710 (
);

FILL FILL_0_BUFX2_insert711 (
);

FILL FILL_0_BUFX2_insert712 (
);

FILL FILL_0_BUFX2_insert713 (
);

FILL FILL_0_BUFX2_insert714 (
);

FILL FILL_0__13284_ (
);

FILL FILL_0_BUFX2_insert715 (
);

FILL FILL_0_BUFX2_insert716 (
);

FILL SFILL53960x64050 (
);

FILL FILL_0_BUFX2_insert717 (
);

FILL SFILL84360x55050 (
);

FILL FILL_0_BUFX2_insert718 (
);

FILL FILL_0_BUFX2_insert719 (
);

FILL FILL_1__6841_ (
);

FILL FILL_2__13611_ (
);

FILL FILL_5__16056_ (
);

FILL FILL_6__9637_ (
);

FILL FILL_5__11191_ (
);

FILL FILL_4__15889_ (
);

FILL FILL_1__12604_ (
);

FILL FILL_4__15469_ (
);

FILL FILL_4__15049_ (
);

FILL FILL_2__16083_ (
);

FILL FILL_4__10184_ (
);

FILL FILL_0__9611_ (
);

FILL FILL_2__9629_ (
);

FILL FILL_2__9209_ (
);

FILL FILL_1__15496_ (
);

FILL FILL_1__15076_ (
);

FILL FILL_5__7634_ (
);

FILL FILL_4__16410_ (
);

FILL FILL_5__7214_ (
);

FILL FILL_0__14489_ (
);

AOI22X1 _14774_ (
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .B(_4005__bF$buf1),
    .C(_3995__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_5259_)
);

FILL FILL_0__14069_ (
);

AOI22X1 _14354_ (
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .B(_3894_),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_4848_)
);

FILL FILL_3__15823_ (
);

FILL FILL_3__15403_ (
);

FILL FILL_1__7626_ (
);

FILL FILL_1__7206_ (
);

FILL FILL_2__14816_ (
);

FILL FILL_0__15850_ (
);

FILL FILL_0__15430_ (
);

FILL FILL_0__15010_ (
);

FILL FILL_5__12396_ (
);

FILL FILL_1__13809_ (
);

FILL FILL_4__11389_ (
);

FILL FILL_3__8913_ (
);

FILL FILL_5__8839_ (
);

FILL SFILL114520x36050 (
);

INVX1 _15979_ (
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_6436_)
);

FILL FILL_4__12750_ (
);

NOR2X1 _15559_ (
    .A(_6025_),
    .B(_6026_),
    .Y(_6027_)
);

FILL FILL_4__12330_ (
);

OAI22X1 _15139_ (
    .A(_5569_),
    .B(_4047_),
    .C(_5483__bF$buf1),
    .D(_4082_),
    .Y(_5617_)
);

OAI21X1 _10694_ (
    .A(_1939_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .C(_1940_),
    .Y(_1888_[26])
);

OAI21X1 _10274_ (
    .A(_1720_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .C(_1721_),
    .Y(_1693_[14])
);

FILL FILL_5__10709_ (
);

FILL FILL_2__6910_ (
);

FILL FILL_3__11743_ (
);

FILL SFILL43960x62050 (
);

FILL FILL_3__11323_ (
);

FILL FILL_4__6836_ (
);

FILL FILL_0__16215_ (
);

FILL FILL_2__10316_ (
);

FILL FILL_2__9382_ (
);

FILL FILL_0__11770_ (
);

FILL FILL_0__11350_ (
);

FILL FILL_5__14962_ (
);

FILL FILL_5__14542_ (
);

FILL FILL_5__14122_ (
);

OAI21X1 _8842_ (
    .A(_989_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_990_),
    .Y(_978_[6])
);

DFFSR _8422_ (
    .Q(\datapath_1.regfile_1.regOut[12] [16]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_718_[16])
);

FILL SFILL43880x69050 (
);

NAND2X1 _8002_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_573_)
);

FILL FILL_4__13955_ (
);

FILL FILL_4__13535_ (
);

FILL FILL_4__13115_ (
);

INVX1 _11899_ (
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_2974_)
);

NAND3X1 _11479_ (
    .A(_2581_),
    .B(_2585_),
    .C(_2593_),
    .Y(\datapath_1.ALUResult [27])
);

AND2X2 _11059_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2178_)
);

FILL SFILL3720x10050 (
);

FILL FILL_3__12528_ (
);

FILL FILL_1__13982_ (
);

FILL FILL_3__12108_ (
);

FILL FILL_1__13562_ (
);

FILL FILL_1__13142_ (
);

FILL FILL112280x73050 (
);

FILL FILL_0__12975_ (
);

OAI21X1 _12840_ (
    .A(_3564_),
    .B(vdd),
    .C(_3565_),
    .Y(_3555_[5])
);

OAI21X1 _12420_ (
    .A(_3344_),
    .B(MemToReg_bF$buf0),
    .C(_3345_),
    .Y(\datapath_1.mux_wd3.dout [25])
);

FILL FILL_0__12135_ (
);

NAND3X1 _12000_ (
    .A(PCSource_1_bF$buf0),
    .B(\aluControl_1.inst [1]),
    .C(_3034__bF$buf0),
    .Y(_3046_)
);

FILL FILL_5__8592_ (
);

FILL FILL_6__16334_ (
);

FILL FILL_5_BUFX2_insert110 (
);

FILL FILL_5__15747_ (
);

FILL FILL_5__15327_ (
);

FILL FILL_6__8908_ (
);

FILL FILL_3__16361_ (
);

NAND2X1 _9627_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1392_)
);

FILL SFILL3640x17050 (
);

NAND2X1 _9207_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .Y(_1237_)
);

FILL FILL_5__10882_ (
);

FILL FILL_1__8584_ (
);

FILL FILL_5__10042_ (
);

FILL FILL_2__15774_ (
);

FILL SFILL104520x34050 (
);

FILL FILL_2__15354_ (
);

FILL SFILL43880x24050 (
);

FILL FILL_1__14767_ (
);

FILL FILL_1__14347_ (
);

FILL FILL_5__6905_ (
);

FILL FILL_3__9871_ (
);

AOI21X1 _13625_ (
    .A(\datapath_1.regfile_1.regOut[23] [3]),
    .B(_4038__bF$buf3),
    .C(_4133_),
    .Y(_4134_)
);

FILL FILL_3__9031_ (
);

DFFSR _13205_ (
    .Q(\datapath_1.PCJump [30]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[30])
);

FILL FILL_5__9797_ (
);

FILL FILL_5__9377_ (
);

FILL FILL_6__12254_ (
);

AOI22X1 _16097_ (
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .C(\datapath_1.regfile_1.regOut[5] [26]),
    .D(_5700_),
    .Y(_6551_)
);

FILL FILL_0__14701_ (
);

FILL FILL_1__9789_ (
);

FILL FILL_5__11667_ (
);

FILL FILL_1__9369_ (
);

FILL FILL_5__11247_ (
);

FILL FILL_3__12281_ (
);

FILL SFILL94520x83050 (
);

FILL FILL_2__16139_ (
);

FILL FILL_4__7374_ (
);

FILL FILL_2__11694_ (
);

FILL FILL_2__11274_ (
);

FILL FILL_1__10687_ (
);

FILL FILL_2_BUFX2_insert240 (
);

FILL FILL_2_BUFX2_insert241 (
);

FILL FILL_1__10267_ (
);

FILL FILL_2_BUFX2_insert242 (
);

FILL FILL_2_BUFX2_insert243 (
);

FILL FILL_2_BUFX2_insert244 (
);

FILL FILL_4__11601_ (
);

FILL FILL_2_BUFX2_insert245 (
);

FILL FILL_0__7694_ (
);

FILL FILL_2_BUFX2_insert246 (
);

FILL FILL_5__15080_ (
);

FILL SFILL49080x38050 (
);

FILL FILL_2_BUFX2_insert247 (
);

NAND2X1 _9380_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1268_)
);

FILL FILL_2_BUFX2_insert248 (
);

FILL FILL_2_BUFX2_insert249 (
);

FILL FILL_6__13879_ (
);

FILL FILL_6__13459_ (
);

FILL FILL_4__14493_ (
);

FILL FILL_4__14073_ (
);

FILL FILL_0__15906_ (
);

FILL FILL_2__8653_ (
);

FILL FILL_3__13486_ (
);

FILL FILL_2__8233_ (
);

FILL FILL_0__10621_ (
);

FILL FILL_4__8999_ (
);

FILL FILL_6__14820_ (
);

FILL FILL_4__8579_ (
);

FILL FILL_6__14400_ (
);

FILL FILL_2__12899_ (
);

FILL FILL_2__12479_ (
);

FILL FILL_2__12059_ (
);

FILL FILL_0__13093_ (
);

FILL FILL_5__13813_ (
);

FILL FILL_4__9940_ (
);

FILL FILL_4__9520_ (
);

FILL FILL_4__9100_ (
);

FILL FILL_2__13840_ (
);

FILL FILL_2__13420_ (
);

FILL FILL_3__6996_ (
);

FILL FILL_5__16285_ (
);

FILL FILL_0__8899_ (
);

FILL SFILL49000x36050 (
);

FILL FILL_2__13000_ (
);

FILL FILL_0__8479_ (
);

FILL FILL_0__8059_ (
);

FILL FILL_4__15698_ (
);

FILL FILL_1__12833_ (
);

FILL FILL_1__12413_ (
);

FILL FILL_4__15278_ (
);

FILL FILL_2__9858_ (
);

FILL FILL_0__9420_ (
);

FILL FILL_0__11826_ (
);

FILL FILL_0__9000_ (
);

FILL FILL_2__9018_ (
);

FILL FILL_0__11406_ (
);

FILL FILL_5__7863_ (
);

FILL FILL_5__7443_ (
);

OAI22X1 _14583_ (
    .A(_5070_),
    .B(_3893__bF$buf2),
    .C(_3944__bF$buf2),
    .D(_5071_),
    .Y(_5072_)
);

FILL FILL_0__14298_ (
);

FILL FILL_6__10320_ (
);

INVX1 _14163_ (
    .A(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_4661_)
);

FILL FILL_3__15632_ (
);

FILL FILL_3__15212_ (
);

FILL FILL_1__7855_ (
);

FILL FILL_1__7435_ (
);

FILL FILL_2__14625_ (
);

FILL FILL_2__14205_ (
);

FILL FILL_1__13618_ (
);

FILL FILL_4__11198_ (
);

FILL FILL_1_BUFX2_insert260 (
);

FILL FILL_1_BUFX2_insert261 (
);

FILL FILL_3__8722_ (
);

FILL FILL_1_BUFX2_insert262 (
);

FILL FILL_1_BUFX2_insert263 (
);

FILL FILL_1_BUFX2_insert264 (
);

FILL FILL_1_BUFX2_insert265 (
);

FILL FILL_1_BUFX2_insert266 (
);

FILL FILL_5__8648_ (
);

FILL FILL_5__8228_ (
);

FILL FILL_1_BUFX2_insert267 (
);

FILL FILL_1_BUFX2_insert268 (
);

FILL FILL_1_BUFX2_insert269 (
);

NOR3X1 _15788_ (
    .A(_5515__bF$buf0),
    .B(_6249_),
    .C(_5521__bF$buf2),
    .Y(_6250_)
);

OAI22X1 _15368_ (
    .A(_4304_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf2),
    .D(_4302_),
    .Y(_5841_)
);

FILL FILL_5__10938_ (
);

DFFSR _10083_ (
    .Q(\datapath_1.regfile_1.regOut[25] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_1563_[13])
);

FILL FILL_3__11972_ (
);

FILL FILL_5__10518_ (
);

FILL SFILL23880x20050 (
);

FILL FILL_3__11552_ (
);

FILL FILL_3__11132_ (
);

FILL FILL_0__16024_ (
);

FILL FILL_2__10965_ (
);

FILL FILL_2__10545_ (
);

FILL FILL_2__10125_ (
);

FILL SFILL63960x16050 (
);

FILL SFILL39000x34050 (
);

FILL FILL112360x2050 (
);

FILL FILL_3__9927_ (
);

FILL FILL_3__9507_ (
);

FILL FILL_5__14771_ (
);

FILL FILL_0__6965_ (
);

FILL FILL_5__14351_ (
);

FILL FILL112280x7050 (
);

FILL FILL_6__7932_ (
);

NAND2X1 _8651_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_904_)
);

NAND2X1 _8231_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_685_)
);

FILL FILL_4__13764_ (
);

FILL SFILL8760x69050 (
);

FILL FILL_4__13344_ (
);

AOI21X1 _11288_ (
    .A(_2379_),
    .B(_2395_),
    .C(_2406_),
    .Y(_2407_)
);

FILL FILL_3__12757_ (
);

FILL FILL_2__7504_ (
);

FILL FILL_1__13791_ (
);

FILL FILL_3__12337_ (
);

FILL FILL_1__13371_ (
);

FILL FILL_0__12784_ (
);

FILL FILL_0__12364_ (
);

FILL SFILL53960x59050 (
);

FILL FILL_5__15976_ (
);

FILL FILL_5__15556_ (
);

FILL FILL_5__15136_ (
);

NAND2X1 _9856_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1504_)
);

FILL FILL_3__16170_ (
);

DFFSR _9436_ (
    .Q(\datapath_1.regfile_1.regOut[20] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1238_[6])
);

INVX1 _9016_ (
    .A(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_1086_)
);

FILL FILL_5__10691_ (
);

FILL FILL_1__8393_ (
);

FILL FILL_5__10271_ (
);

FILL SFILL114200x55050 (
);

FILL FILL_4__14969_ (
);

FILL FILL_4__14549_ (
);

FILL FILL_4__14129_ (
);

FILL FILL_2__15583_ (
);

FILL FILL_2__15163_ (
);

FILL FILL_2__8709_ (
);

FILL SFILL13800x61050 (
);

FILL FILL_1__14996_ (
);

FILL FILL_1__14576_ (
);

FILL FILL_1__14156_ (
);

FILL FILL_4__15910_ (
);

FILL FILL_0__13989_ (
);

FILL FILL_3__9680_ (
);

AOI22X1 _13854_ (
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .B(_4246_),
    .C(_3998__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_4358_)
);

FILL FILL_0__13569_ (
);

FILL FILL_3__9260_ (
);

FILL FILL_0__13149_ (
);

AOI21X1 _13434_ (
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .B(_3942__bF$buf0),
    .C(_3945_),
    .Y(_3946_)
);

INVX1 _13014_ (
    .A(_2_[21]),
    .Y(_3661_)
);

FILL FILL_3__14903_ (
);

FILL SFILL114600x24050 (
);

FILL SFILL53960x14050 (
);

FILL FILL_0__14930_ (
);

FILL FILL_0__14510_ (
);

FILL FILL_5__11896_ (
);

FILL FILL_5__11476_ (
);

FILL FILL_1__9598_ (
);

FILL FILL_5__11056_ (
);

FILL FILL_3__12090_ (
);

FILL FILL_2__16368_ (
);

FILL FILL_4__7183_ (
);

FILL FILL_4__10889_ (
);

FILL FILL_4__10049_ (
);

FILL FILL_2__11083_ (
);

FILL FILL_1__10496_ (
);

INVX1 _14639_ (
    .A(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_5127_)
);

FILL FILL_4__11830_ (
);

INVX1 _14219_ (
    .A(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_4715_)
);

FILL FILL_4__11410_ (
);

FILL FILL_0__7083_ (
);

FILL FILL_6__8470_ (
);

FILL FILL_1__16302_ (
);

FILL FILL_3__10823_ (
);

FILL FILL_3__10403_ (
);

FILL FILL_0__15715_ (
);

FILL FILL_2__8882_ (
);

FILL FILL_2__8462_ (
);

FILL FILL_3__13295_ (
);

FILL FILL_0__10430_ (
);

FILL FILL_0__10010_ (
);

FILL FILL_4__8388_ (
);

FILL FILL112360x61050 (
);

FILL FILL_2__12288_ (
);

FILL FILL_5__13622_ (
);

DFFSR _7922_ (
    .Q(\datapath_1.regfile_1.regOut[8] [28]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_458_[28])
);

NAND2X1 _7502_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_321_)
);

FILL FILL_4__12615_ (
);

FILL SFILL64040x70050 (
);

FILL FILL_5__16094_ (
);

NAND2X1 _10979_ (
    .A(vdd),
    .B(\control_1.next [2]),
    .Y(_2104_)
);

NAND2X1 _10559_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1871_)
);

FILL FILL_6__9255_ (
);

NAND2X1 _10139_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1652_)
);

FILL FILL_3__11608_ (
);

FILL FILL_1__12642_ (
);

FILL FILL_1__12222_ (
);

FILL FILL_4__15087_ (
);

FILL SFILL43960x12050 (
);

FILL FILL112280x68050 (
);

FILL FILL_2__9667_ (
);

INVX1 _11920_ (
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_2988_)
);

FILL FILL_0__11635_ (
);

FILL FILL_2__9247_ (
);

FILL FILL_0__11215_ (
);

NAND3X1 _11500_ (
    .A(_2296_),
    .B(_2305_),
    .C(_2612_),
    .Y(_2613_)
);

FILL FILL_5__7672_ (
);

FILL FILL_5__7252_ (
);

INVX1 _14392_ (
    .A(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_4885_)
);

FILL FILL_5__14827_ (
);

FILL FILL_5__14407_ (
);

FILL FILL_3__15861_ (
);

FILL FILL_3__15441_ (
);

NAND2X1 _8707_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_921_)
);

FILL FILL_3__15021_ (
);

FILL FILL_1__7244_ (
);

FILL FILL_2__14854_ (
);

FILL SFILL43880x19050 (
);

FILL FILL_2__14434_ (
);

FILL FILL_2__14014_ (
);

FILL FILL_1__13847_ (
);

FILL FILL_1__13427_ (
);

FILL FILL_1__13007_ (
);

FILL FILL_3__8951_ (
);

FILL FILL_3__8531_ (
);

NAND2X1 _12705_ (
    .A(IRWrite_bF$buf1),
    .B(memoryOutData[3]),
    .Y(_3496_)
);

FILL FILL_3__8111_ (
);

FILL SFILL84280x6050 (
);

FILL FILL_5__8877_ (
);

FILL FILL_5__8457_ (
);

NOR2X1 _15597_ (
    .A(_6062_),
    .B(_6063_),
    .Y(_6064_)
);

NAND2X1 _15177_ (
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .B(_5494_),
    .Y(_5654_)
);

FILL FILL_3__16226_ (
);

FILL FILL_1__8869_ (
);

FILL FILL_5__10747_ (
);

FILL FILL_1__8449_ (
);

FILL FILL_3__11781_ (
);

FILL FILL_3__11361_ (
);

FILL FILL_2__15639_ (
);

FILL FILL_2__15219_ (
);

FILL FILL_4__6874_ (
);

FILL SFILL83560x8050 (
);

FILL FILL_0__16253_ (
);

FILL FILL_2__10774_ (
);

INVX1 _7099_ (
    .A(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_113_)
);

FILL FILL_1__9810_ (
);

FILL FILL_3__9736_ (
);

FILL FILL_5__14580_ (
);

FILL FILL_5__14160_ (
);

NAND2X1 _8880_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1016_)
);

NAND2X1 _8460_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_797_)
);

DFFSR _8040_ (
    .Q(\datapath_1.regfile_1.regOut[9] [18]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_523_[18])
);

FILL FILL_4__13993_ (
);

FILL FILL_4__13573_ (
);

FILL FILL_4__13153_ (
);

AOI21X1 _11097_ (
    .A(_2187_),
    .B(_2205_),
    .C(_2215_),
    .Y(_2216_)
);

FILL FILL_2__7733_ (
);

FILL FILL_3__12986_ (
);

FILL FILL_2__7313_ (
);

FILL FILL_3__12146_ (
);

FILL FILL_4__7239_ (
);

FILL FILL_2__11979_ (
);

FILL FILL_2__11559_ (
);

FILL FILL_0__12593_ (
);

FILL FILL_2__11139_ (
);

FILL SFILL33880x17050 (
);

FILL FILL_0__12173_ (
);

FILL FILL_4__8600_ (
);

FILL FILL_5__15785_ (
);

FILL FILL_5__15365_ (
);

FILL FILL_2__12500_ (
);

FILL FILL_0__7979_ (
);

FILL FILL_0__7559_ (
);

FILL FILL_6__8526_ (
);

INVX1 _9665_ (
    .A(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_1417_)
);

INVX1 _9245_ (
    .A(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_1198_)
);

FILL FILL_1__11913_ (
);

FILL FILL_4__14778_ (
);

FILL FILL_4__14358_ (
);

FILL FILL_2__15392_ (
);

FILL FILL_0__10906_ (
);

FILL FILL_2__8518_ (
);

FILL FILL_0__8500_ (
);

FILL FILL_1__14385_ (
);

FILL FILL_5__6943_ (
);

FILL FILL_1_BUFX2_insert1020 (
);

FILL FILL_1_BUFX2_insert1021 (
);

FILL FILL_1_BUFX2_insert1022 (
);

FILL FILL_0__13798_ (
);

FILL FILL_1_BUFX2_insert1023 (
);

NAND2X1 _13663_ (
    .A(_4170_),
    .B(_4163_),
    .Y(_4171_)
);

FILL FILL_0__13378_ (
);

FILL FILL_1_BUFX2_insert1024 (
);

NAND2X1 _13243_ (
    .A(_3750_),
    .B(_3754_),
    .Y(_3786_)
);

FILL FILL_1_BUFX2_insert1025 (
);

FILL FILL_1_BUFX2_insert1026 (
);

FILL FILL_3__14712_ (
);

FILL FILL_1_BUFX2_insert1027 (
);

FILL FILL_1_BUFX2_insert1028 (
);

FILL FILL_1_BUFX2_insert1029 (
);

FILL FILL_1__6935_ (
);

FILL FILL_4__9805_ (
);

FILL FILL_2__13705_ (
);

FILL FILL_5__11285_ (
);

FILL FILL_2__16177_ (
);

FILL FILL_4__10698_ (
);

FILL SFILL79720x8050 (
);

FILL FILL_4__10278_ (
);

FILL FILL_3__7802_ (
);

FILL FILL_5__7728_ (
);

FILL FILL_5__7308_ (
);

FILL FILL_2_BUFX2_insert620 (
);

FILL FILL_2_BUFX2_insert621 (
);

FILL FILL_2_BUFX2_insert622 (
);

AOI22X1 _14868_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [29]),
    .C(\datapath_1.regfile_1.regOut[18] [29]),
    .D(_4135_),
    .Y(_5351_)
);

FILL FILL_2_BUFX2_insert623 (
);

FILL SFILL23800x58050 (
);

FILL FILL_2_BUFX2_insert624 (
);

NAND3X1 _14448_ (
    .A(_4938_),
    .B(_4939_),
    .C(_4937_),
    .Y(_4940_)
);

FILL FILL_2_BUFX2_insert625 (
);

INVX1 _14028_ (
    .A(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_4528_)
);

FILL FILL_3__15917_ (
);

FILL FILL_2_BUFX2_insert626 (
);

FILL FILL_2_BUFX2_insert627 (
);

FILL FILL_2_BUFX2_insert628 (
);

FILL SFILL79320x7050 (
);

FILL FILL_1__16111_ (
);

FILL FILL_2_BUFX2_insert629 (
);

FILL SFILL23880x15050 (
);

FILL FILL_3__10632_ (
);

FILL FILL_0__15944_ (
);

FILL SFILL54280x5050 (
);

FILL FILL_0__15524_ (
);

FILL SFILL53960x8050 (
);

FILL FILL_0__15104_ (
);

FILL FILL_2__8271_ (
);

FILL SFILL39000x29050 (
);

FILL FILL_4__8197_ (
);

FILL FILL_2__12097_ (
);

FILL FILL_5__13851_ (
);

FILL FILL_5__13431_ (
);

FILL SFILL84440x38050 (
);

FILL FILL_5__13011_ (
);

FILL SFILL53560x7050 (
);

NAND2X1 _7731_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_433_)
);

NAND2X1 _7311_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_214_)
);

FILL FILL_4__12844_ (
);

FILL FILL_4__12424_ (
);

FILL FILL_4__12004_ (
);

NAND2X1 _10788_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1983_)
);

FILL FILL_0__8097_ (
);

NAND2X1 _10368_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1764_)
);

FILL SFILL23800x13050 (
);

FILL FILL_3__11837_ (
);

FILL SFILL104680x6050 (
);

FILL FILL_1__12871_ (
);

FILL FILL_3__11417_ (
);

FILL FILL_1__12451_ (
);

FILL FILL_1__12031_ (
);

FILL FILL_0__16309_ (
);

FILL FILL_2__9896_ (
);

FILL FILL_2__9476_ (
);

FILL FILL_0__11864_ (
);

FILL FILL_0__11444_ (
);

FILL FILL_0__11024_ (
);

FILL FILL_5__7481_ (
);

FILL FILL_5__7061_ (
);

FILL SFILL74120x60050 (
);

FILL FILL_5__14636_ (
);

FILL FILL_3__15670_ (
);

FILL FILL_5__14216_ (
);

FILL FILL_3__15250_ (
);

DFFSR _8936_ (
    .Q(\datapath_1.regfile_1.regOut[16] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_978_[18])
);

INVX1 _8516_ (
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_834_)
);

FILL FILL_1__7893_ (
);

FILL FILL_1__7473_ (
);

FILL FILL_1__7053_ (
);

FILL FILL_4__13629_ (
);

FILL FILL_4__13209_ (
);

FILL FILL_2__14663_ (
);

FILL FILL_2__14243_ (
);

FILL SFILL13800x56050 (
);

FILL FILL_3_BUFX2_insert80 (
);

FILL FILL_1__13656_ (
);

FILL FILL_3_BUFX2_insert81 (
);

FILL FILL_1__13236_ (
);

FILL FILL_3_BUFX2_insert82 (
);

FILL FILL_3_BUFX2_insert83 (
);

FILL SFILL74040x67050 (
);

FILL FILL_3_BUFX2_insert84 (
);

FILL FILL_3_BUFX2_insert85 (
);

FILL FILL_3_BUFX2_insert86 (
);

FILL FILL_1_BUFX2_insert640 (
);

FILL FILL_3_BUFX2_insert87 (
);

FILL FILL_3__8760_ (
);

FILL FILL_1_BUFX2_insert641 (
);

FILL FILL_0__12649_ (
);

FILL FILL_3_BUFX2_insert88 (
);

DFFSR _12934_ (
    .Q(\datapath_1.a [15]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_3555_[15])
);

FILL FILL_1_BUFX2_insert642 (
);

FILL FILL_3__8340_ (
);

FILL FILL_3_BUFX2_insert89 (
);

INVX1 _12514_ (
    .A(ALUOut[25]),
    .Y(_3409_)
);

FILL FILL_1_BUFX2_insert643 (
);

FILL FILL_0__12229_ (
);

FILL FILL_1_BUFX2_insert644 (
);

FILL FILL_1_BUFX2_insert645 (
);

FILL FILL_1_BUFX2_insert646 (
);

FILL FILL_5__8266_ (
);

FILL FILL_1_BUFX2_insert647 (
);

FILL FILL_1_BUFX2_insert648 (
);

FILL FILL_6__11983_ (
);

FILL FILL_1_BUFX2_insert649 (
);

FILL FILL_3__16035_ (
);

FILL FILL_5__10976_ (
);

FILL FILL_5__10556_ (
);

FILL FILL_5__10136_ (
);

FILL FILL_3__11590_ (
);

FILL FILL_1__8258_ (
);

FILL FILL_3__11170_ (
);

FILL FILL_2__15868_ (
);

FILL FILL_2__15448_ (
);

FILL FILL_2__15028_ (
);

FILL FILL_0__16062_ (
);

FILL FILL_2__10163_ (
);

FILL SFILL13800x11050 (
);

FILL FILL_3__9545_ (
);

FILL FILL_4__10910_ (
);

FILL FILL_3__9125_ (
);

AOI22X1 _13719_ (
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .B(_3942__bF$buf0),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_4226_)
);

FILL FILL_1__15802_ (
);

FILL FILL_6__7550_ (
);

FILL FILL_6__12768_ (
);

FILL FILL_4__13382_ (
);

FILL SFILL99240x71050 (
);

FILL FILL_2__7962_ (
);

FILL FILL_2__7542_ (
);

BUFX2 BUFX2_insert310 (
    .A(_2341_),
    .Y(_2341__bF$buf2)
);

FILL FILL_3__12375_ (
);

FILL FILL_2__7122_ (
);

BUFX2 BUFX2_insert311 (
    .A(_2341_),
    .Y(_2341__bF$buf1)
);

BUFX2 BUFX2_insert312 (
    .A(_2341_),
    .Y(_2341__bF$buf0)
);

BUFX2 BUFX2_insert313 (
    .A(_3966_),
    .Y(_3966__bF$buf3)
);

BUFX2 BUFX2_insert314 (
    .A(_3966_),
    .Y(_3966__bF$buf2)
);

FILL FILL_4__7888_ (
);

FILL FILL_4__7468_ (
);

BUFX2 BUFX2_insert315 (
    .A(_3966_),
    .Y(_3966__bF$buf1)
);

FILL FILL_4__7048_ (
);

BUFX2 BUFX2_insert316 (
    .A(_3966_),
    .Y(_3966__bF$buf0)
);

FILL FILL112360x56050 (
);

BUFX2 BUFX2_insert317 (
    .A(_5480_),
    .Y(_5480__bF$buf3)
);

FILL FILL_2__11788_ (
);

BUFX2 BUFX2_insert318 (
    .A(_5480_),
    .Y(_5480__bF$buf2)
);

FILL FILL_2__11368_ (
);

BUFX2 BUFX2_insert319 (
    .A(_5480_),
    .Y(_5480__bF$buf1)
);

FILL FILL_5__12702_ (
);

FILL FILL_6__16181_ (
);

FILL SFILL64040x65050 (
);

FILL FILL_5__15594_ (
);

FILL FILL_5__15174_ (
);

INVX1 _9894_ (
    .A(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_1529_)
);

FILL FILL_0__7368_ (
);

INVX1 _9474_ (
    .A(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_1310_)
);

FILL FILL_6__8335_ (
);

DFFSR _9054_ (
    .Q(\datapath_1.regfile_1.regOut[17] [8]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_1043_[8])
);

FILL SFILL23640x1050 (
);

FILL FILL_4__14587_ (
);

FILL FILL_1__11722_ (
);

FILL FILL_4__14167_ (
);

FILL FILL_1__11302_ (
);

FILL SFILL104600x17050 (
);

FILL FILL_2__8747_ (
);

FILL FILL_2__8327_ (
);

FILL FILL_1__14194_ (
);

INVX1 _13892_ (
    .A(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_4395_)
);

FILL SFILL108920x25050 (
);

OAI22X1 _13472_ (
    .A(_3981_),
    .B(_3982__bF$buf0),
    .C(_3983__bF$buf3),
    .D(_3980_),
    .Y(_3984_)
);

DFFSR _13052_ (
    .Q(_2_[5]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3620_[5])
);

FILL FILL_5__13907_ (
);

FILL FILL_3__14941_ (
);

FILL FILL112360x11050 (
);

FILL FILL_3__14521_ (
);

FILL FILL_3__14101_ (
);

FILL FILL_4__9614_ (
);

FILL FILL_2__13934_ (
);

FILL FILL_5__16379_ (
);

FILL FILL_2__13514_ (
);

FILL SFILL64040x20050 (
);

FILL FILL_5__11094_ (
);

FILL FILL_1__12507_ (
);

FILL FILL_0__9934_ (
);

FILL FILL_3__7611_ (
);

FILL FILL_0__9514_ (
);

FILL FILL112280x18050 (
);

FILL FILL_1__15399_ (
);

FILL FILL_5__7957_ (
);

FILL FILL_5__7117_ (
);

FILL FILL_4__16313_ (
);

INVX1 _14677_ (
    .A(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_5164_)
);

INVX1 _14257_ (
    .A(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_4753_)
);

FILL FILL_3__15726_ (
);

FILL FILL_3__15306_ (
);

FILL FILL_1__16340_ (
);

FILL FILL_1__7949_ (
);

FILL FILL_1__7109_ (
);

FILL FILL_3__10441_ (
);

FILL FILL_3__10021_ (
);

FILL FILL_2__14719_ (
);

FILL FILL_0__15753_ (
);

FILL FILL_0__15333_ (
);

FILL FILL_5__12299_ (
);

FILL SFILL54040x63050 (
);

FILL FILL_2__8080_ (
);

FILL FILL_5__13660_ (
);

FILL FILL_5__13240_ (
);

NAND2X1 _7960_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_545_)
);

DFFSR _7540_ (
    .Q(\datapath_1.regfile_1.regOut[5] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_263_[30])
);

INVX1 _7120_ (
    .A(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_127_)
);

FILL FILL_4__12653_ (
);

FILL FILL_4__12233_ (
);

DFFSR _10597_ (
    .Q(\datapath_1.regfile_1.regOut[29] [15]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_1823_[15])
);

INVX1 _10177_ (
    .A(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_1677_)
);

FILL FILL_3__11646_ (
);

FILL FILL_3__11226_ (
);

FILL FILL_1__12260_ (
);

FILL FILL_0__16118_ (
);

NAND2X1 _16403_ (
    .A(gnd),
    .B(gnd),
    .Y(_6823_)
);

FILL FILL_2__10639_ (
);

FILL FILL_2__9285_ (
);

FILL FILL_0__11673_ (
);

FILL FILL_0__11253_ (
);

FILL FILL_5__7290_ (
);

FILL FILL_5__14865_ (
);

FILL FILL_5__14445_ (
);

FILL FILL_5__14025_ (
);

FILL FILL_6__7606_ (
);

INVX1 _8745_ (
    .A(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_946_)
);

INVX1 _8325_ (
    .A(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_727_)
);

FILL FILL_4__13858_ (
);

FILL FILL_4__13438_ (
);

FILL FILL_2__14892_ (
);

FILL FILL_2__14472_ (
);

FILL FILL_4__13018_ (
);

FILL FILL_2__14052_ (
);

FILL FILL_1__13885_ (
);

FILL FILL_1__13465_ (
);

FILL FILL_1__13045_ (
);

FILL SFILL8520x76050 (
);

FILL FILL_0__12878_ (
);

FILL SFILL59160x2050 (
);

INVX1 _12743_ (
    .A(\datapath_1.PCJump [18]),
    .Y(_3521_)
);

FILL FILL_0__12458_ (
);

FILL FILL_0__12038_ (
);

NAND3X1 _12323_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3281_)
);

FILL FILL_6__16237_ (
);

FILL FILL_5__8495_ (
);

FILL SFILL79160x74050 (
);

FILL SFILL59080x7050 (
);

FILL FILL_5__8075_ (
);

FILL SFILL44040x61050 (
);

FILL FILL_3__16264_ (
);

FILL FILL_5__10785_ (
);

FILL FILL_1__8487_ (
);

FILL FILL_5__10365_ (
);

FILL FILL_1__8067_ (
);

FILL FILL_2__15677_ (
);

FILL FILL_2__15257_ (
);

FILL FILL_0__16291_ (
);

FILL FILL_2__10392_ (
);

FILL FILL_3__9774_ (
);

FILL FILL_3__9354_ (
);

OAI22X1 _13948_ (
    .A(_4449_),
    .B(_3972__bF$buf3),
    .C(_3920_),
    .D(_4448_),
    .Y(_4450_)
);

AOI22X1 _13528_ (
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .B(_3894_),
    .C(_4038__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_4039_)
);

OAI21X1 _13108_ (
    .A(_3702_),
    .B(PCEn_bF$buf2),
    .C(_3703_),
    .Y(_3685_[9])
);

FILL FILL_1__15611_ (
);

FILL FILL_6__12157_ (
);

FILL FILL_0__14604_ (
);

FILL FILL_2__7351_ (
);

FILL FILL_3__12184_ (
);

FILL FILL_4__7697_ (
);

FILL FILL_2__11597_ (
);

FILL FILL_2__11177_ (
);

FILL SFILL8440x38050 (
);

FILL FILL_5__12511_ (
);

FILL FILL_4__11924_ (
);

FILL FILL_4__11504_ (
);

FILL FILL_0__7597_ (
);

FILL FILL_0__7177_ (
);

OAI21X1 _9283_ (
    .A(_1222_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1223_),
    .Y(_1173_[25])
);

FILL FILL_3__10917_ (
);

FILL FILL_1__11951_ (
);

FILL FILL_4__14396_ (
);

FILL FILL_1__11531_ (
);

FILL SFILL38760x81050 (
);

FILL FILL_1__11111_ (
);

FILL FILL_0__15809_ (
);

FILL FILL_2__8976_ (
);

FILL FILL_0__10944_ (
);

FILL FILL_3__13389_ (
);

FILL FILL_0__10524_ (
);

FILL FILL_2__8136_ (
);

FILL FILL_0__10104_ (
);

FILL SFILL78840x77050 (
);

FILL FILL_6__14723_ (
);

FILL FILL_5__6981_ (
);

FILL FILL_6__14303_ (
);

FILL SFILL74120x55050 (
);

OAI21X1 _13281_ (
    .A(_3773_),
    .B(_3759_),
    .C(_3774_),
    .Y(_3820_)
);

FILL FILL_5__13716_ (
);

FILL FILL_3__14750_ (
);

FILL FILL_3__14330_ (
);

FILL FILL_1__6973_ (
);

FILL FILL_4__9423_ (
);

FILL FILL_4__12709_ (
);

FILL FILL_4__9003_ (
);

FILL FILL_2__13743_ (
);

FILL FILL_2__13323_ (
);

FILL FILL_5__16188_ (
);

FILL FILL_3__6899_ (
);

FILL FILL_1__12736_ (
);

FILL FILL_1__12316_ (
);

FILL FILL_0__9743_ (
);

FILL FILL_3__7840_ (
);

FILL FILL_3__7420_ (
);

FILL FILL_0__11729_ (
);

FILL FILL_0__11309_ (
);

FILL FILL_5__7346_ (
);

FILL FILL_4__16122_ (
);

OAI22X1 _14486_ (
    .A(_4975_),
    .B(_3902__bF$buf0),
    .C(_3971__bF$buf1),
    .D(_4976_),
    .Y(_4977_)
);

INVX1 _14066_ (
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_4566_)
);

FILL SFILL74120x10050 (
);

FILL FILL_3__15955_ (
);

FILL FILL_3__15535_ (
);

FILL FILL_3__15115_ (
);

FILL FILL_1__7758_ (
);

FILL FILL_3__10670_ (
);

FILL FILL_1__7338_ (
);

FILL FILL_3__10250_ (
);

FILL SFILL28840x4050 (
);

FILL FILL_2__14948_ (
);

FILL FILL_0__15982_ (
);

FILL FILL_2__14528_ (
);

FILL FILL_0__15562_ (
);

FILL FILL_2__14108_ (
);

FILL FILL_0__15142_ (
);

FILL SFILL28760x9050 (
);

FILL FILL_3__8625_ (
);

FILL FILL_3__8205_ (
);

FILL SFILL59160x70050 (
);

FILL SFILL8680x5050 (
);

FILL FILL_4__12882_ (
);

FILL FILL_4__12462_ (
);

FILL FILL_4__12042_ (
);

FILL SFILL64120x53050 (
);

FILL FILL_3__11875_ (
);

FILL FILL_5__9912_ (
);

FILL FILL_3__11455_ (
);

FILL FILL_3__11035_ (
);

FILL FILL_4__6968_ (
);

FILL FILL_0__16347_ (
);

AOI22X1 _16212_ (
    .A(_5971_),
    .B(\datapath_1.regfile_1.regOut[14] [29]),
    .C(\datapath_1.regfile_1.regOut[22] [29]),
    .D(_5650_),
    .Y(_6663_)
);

FILL FILL_2__10448_ (
);

FILL FILL_2__10028_ (
);

FILL FILL_0__11482_ (
);

FILL FILL_2__9094_ (
);

FILL FILL_0__11062_ (
);

FILL FILL_1__9904_ (
);

FILL FILL_5__14674_ (
);

FILL FILL_5__14254_ (
);

FILL FILL_0__6868_ (
);

INVX1 _8974_ (
    .A(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_1058_)
);

FILL FILL_6__7415_ (
);

DFFSR _8554_ (
    .Q(\datapath_1.regfile_1.regOut[13] [20]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_783_[20])
);

OAI21X1 _8134_ (
    .A(_639_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_640_),
    .Y(_588_[26])
);

FILL FILL_1__7091_ (
);

FILL FILL_4__13667_ (
);

FILL FILL_1__10802_ (
);

FILL FILL_4__13247_ (
);

FILL FILL_2__14281_ (
);

FILL FILL_2__7827_ (
);

FILL FILL_1__13694_ (
);

FILL FILL_1__13274_ (
);

INVX1 _12972_ (
    .A(_2_[7]),
    .Y(_3633_)
);

DFFSR _12552_ (
    .Q(ALUOut[17]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3360_[17])
);

FILL FILL_0__12267_ (
);

OAI21X1 _12132_ (
    .A(_3140_),
    .B(ALUSrcA_bF$buf0),
    .C(_3141_),
    .Y(\datapath_1.alu_1.ALUInA [5])
);

FILL SFILL28680x41050 (
);

FILL FILL_3__13601_ (
);

FILL FILL_5__15879_ (
);

FILL FILL_5__15459_ (
);

FILL FILL_5__15039_ (
);

FILL FILL_3__16073_ (
);

OAI21X1 _9759_ (
    .A(_1458_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .C(_1459_),
    .Y(_1433_[13])
);

OAI21X1 _9339_ (
    .A(_1239_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1240_),
    .Y(_1238_[1])
);

FILL SFILL64040x15050 (
);

FILL FILL_5__10174_ (
);

FILL FILL_2__15486_ (
);

FILL FILL_2__15066_ (
);

FILL FILL_5__16400_ (
);

FILL SFILL89240x64050 (
);

FILL FILL_1__14899_ (
);

FILL SFILL54120x51050 (
);

FILL FILL_1__14479_ (
);

FILL FILL_1__14059_ (
);

FILL FILL_4__15813_ (
);

FILL FILL_3__9163_ (
);

INVX1 _13757_ (
    .A(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_4263_)
);

NAND3X1 _13337_ (
    .A(_3799_),
    .B(_3856_),
    .C(_3859_),
    .Y(_3860_)
);

FILL FILL_3__14806_ (
);

FILL FILL_1__15840_ (
);

FILL FILL_5__9089_ (
);

FILL FILL_1__15420_ (
);

FILL FILL_1__15000_ (
);

FILL FILL_0__14833_ (
);

FILL FILL_0__14413_ (
);

FILL SFILL89640x33050 (
);

FILL FILL_5__11799_ (
);

FILL SFILL54040x58050 (
);

FILL FILL_2__7580_ (
);

FILL FILL_5__11379_ (
);

FILL FILL_2__7160_ (
);

FILL FILL_4__7086_ (
);

FILL FILL_5__12740_ (
);

FILL FILL_5__12320_ (
);

FILL FILL_1__10399_ (
);

FILL FILL_4__11733_ (
);

FILL FILL_4__11313_ (
);

OAI21X1 _9092_ (
    .A(_1115_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1116_),
    .Y(_1108_[4])
);

FILL FILL_1__16205_ (
);

FILL FILL_1__11760_ (
);

FILL FILL_3__10306_ (
);

FILL FILL_1__11340_ (
);

AOI22X1 _15903_ (
    .A(\datapath_1.regfile_1.regOut[1] [21]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_6362_)
);

FILL FILL_0__15618_ (
);

FILL FILL_2__8785_ (
);

FILL FILL_0__10753_ (
);

FILL FILL_2__8365_ (
);

FILL SFILL54040x13050 (
);

OAI21X1 _13090_ (
    .A(_3690_),
    .B(PCEn_bF$buf6),
    .C(_3691_),
    .Y(_3685_[3])
);

FILL FILL_5__13945_ (
);

FILL FILL_5__13525_ (
);

FILL FILL_5__13105_ (
);

INVX1 _7825_ (
    .A(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_475_)
);

DFFSR _7405_ (
    .Q(\datapath_1.regfile_1.regOut[4] [23]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_198_[23])
);

FILL SFILL79240x62050 (
);

FILL FILL_4_BUFX2_insert530 (
);

FILL FILL_4__9652_ (
);

FILL FILL_4_BUFX2_insert531 (
);

FILL FILL_4__9232_ (
);

FILL FILL_4_BUFX2_insert532 (
);

FILL FILL_4__12518_ (
);

FILL FILL_4_BUFX2_insert533 (
);

FILL FILL_2__13972_ (
);

FILL FILL_4_BUFX2_insert534 (
);

FILL FILL_2__13552_ (
);

FILL FILL_4_BUFX2_insert535 (
);

FILL FILL_2__13132_ (
);

FILL FILL_4_BUFX2_insert536 (
);

FILL FILL_4_BUFX2_insert537 (
);

FILL FILL_4_BUFX2_insert538 (
);

FILL FILL_4_BUFX2_insert539 (
);

FILL FILL111880x75050 (
);

FILL FILL_1__12965_ (
);

FILL FILL_1__12125_ (
);

FILL FILL_0__11958_ (
);

FILL FILL_0__9552_ (
);

FILL FILL_0__9132_ (
);

AOI21X1 _11823_ (
    .A(_2911_),
    .B(_2541_),
    .C(_2912_),
    .Y(_2913_)
);

FILL FILL_0__11538_ (
);

FILL FILL_0__11118_ (
);

NAND2X1 _11403_ (
    .A(_2265_),
    .B(_2519_),
    .Y(_2520_)
);

FILL FILL_5__7995_ (
);

FILL FILL_5__7575_ (
);

FILL SFILL44040x56050 (
);

FILL FILL_4__16351_ (
);

INVX1 _14295_ (
    .A(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_4790_)
);

FILL FILL_3__15764_ (
);

FILL FILL_3__15344_ (
);

FILL FILL_1__7987_ (
);

FILL FILL_1__7567_ (
);

FILL FILL_2__14757_ (
);

FILL FILL_0__15791_ (
);

FILL FILL_2__14337_ (
);

FILL FILL_0__15371_ (
);

FILL FILL_3__8854_ (
);

FILL FILL_3__8014_ (
);

OAI21X1 _12608_ (
    .A(_3450_),
    .B(vdd),
    .C(_3451_),
    .Y(_3425_[13])
);

FILL SFILL109400x43050 (
);

FILL FILL_4__12271_ (
);

FILL SFILL44040x11050 (
);

FILL FILL_3__16129_ (
);

FILL FILL_2__6851_ (
);

FILL FILL_5__9721_ (
);

FILL FILL_3__11684_ (
);

FILL FILL_5__9301_ (
);

FILL FILL_3__11264_ (
);

DFFSR _16441_ (
    .Q(\datapath_1.regfile_1.regOut[0] [24]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_6769_[24])
);

FILL FILL_0__16156_ (
);

NOR2X1 _16021_ (
    .A(_6476_),
    .B(_6468_),
    .Y(_6477_)
);

FILL FILL_2__10677_ (
);

FILL FILL_2__10257_ (
);

FILL FILL_0__11291_ (
);

FILL FILL_6__15490_ (
);

FILL FILL_3__9639_ (
);

FILL FILL_3_BUFX2_insert550 (
);

FILL FILL_3__9219_ (
);

FILL FILL_3_BUFX2_insert551 (
);

FILL FILL_3_BUFX2_insert552 (
);

FILL FILL_3_BUFX2_insert553 (
);

FILL FILL_5__14483_ (
);

FILL FILL_5__14063_ (
);

FILL FILL_3_BUFX2_insert554 (
);

OAI21X1 _8783_ (
    .A(_970_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .C(_971_),
    .Y(_913_[29])
);

FILL FILL_3_BUFX2_insert555 (
);

FILL FILL_3_BUFX2_insert556 (
);

FILL FILL_6__7224_ (
);

OAI21X1 _8363_ (
    .A(_751_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_752_),
    .Y(_718_[17])
);

FILL FILL_3_BUFX2_insert557 (
);

FILL FILL_3_BUFX2_insert558 (
);

FILL FILL_3_BUFX2_insert559 (
);

FILL FILL_4__13896_ (
);

FILL FILL_4__13476_ (
);

FILL SFILL69160x67050 (
);

FILL FILL_2__14090_ (
);

FILL FILL_3__12889_ (
);

FILL FILL_2__7636_ (
);

FILL FILL_3__12469_ (
);

FILL FILL_2__7216_ (
);

FILL FILL_3__12049_ (
);

FILL FILL_1__13083_ (
);

OAI21X1 _12781_ (
    .A(_3545_),
    .B(IRWrite_bF$buf7),
    .C(_3546_),
    .Y(_3490_[28])
);

FILL FILL_0__12496_ (
);

INVX1 _12361_ (
    .A(ALUOut[6]),
    .Y(_3306_)
);

FILL FILL_0__12076_ (
);

FILL FILL_3__13830_ (
);

FILL FILL_3__13410_ (
);

FILL FILL_4__8503_ (
);

FILL FILL_5__15688_ (
);

FILL FILL_2__12823_ (
);

FILL FILL_2__12403_ (
);

FILL FILL_5__15268_ (
);

OAI21X1 _9988_ (
    .A(_1570_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1571_),
    .Y(_1563_[4])
);

DFFSR _9568_ (
    .Q(\datapath_1.regfile_1.regOut[21] [10]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_1303_[10])
);

NAND2X1 _9148_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1154_)
);

FILL FILL_6__8009_ (
);

FILL FILL_1__11816_ (
);

FILL FILL_2__15295_ (
);

FILL FILL_3__6920_ (
);

FILL FILL_0__8823_ (
);

FILL FILL_0__10809_ (
);

FILL FILL_0__8403_ (
);

FILL FILL_1__14288_ (
);

FILL FILL_5__6846_ (
);

FILL FILL_0_BUFX2_insert680 (
);

FILL FILL_4__15622_ (
);

FILL FILL_0_BUFX2_insert681 (
);

FILL FILL_4__15202_ (
);

FILL FILL_0_BUFX2_insert682 (
);

FILL FILL_0_BUFX2_insert683 (
);

FILL FILL_0_BUFX2_insert684 (
);

NOR2X1 _13986_ (
    .A(_4486_),
    .B(_4483_),
    .Y(_4487_)
);

FILL FILL_3__9392_ (
);

FILL FILL_0_BUFX2_insert685 (
);

OAI22X1 _13566_ (
    .A(_4074_),
    .B(_3905__bF$buf3),
    .C(_3909_),
    .D(_4075_),
    .Y(_4076_)
);

NAND2X1 _13146_ (
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [22]),
    .Y(_3729_)
);

FILL FILL_0_BUFX2_insert686 (
);

FILL FILL_0_BUFX2_insert687 (
);

FILL FILL_3__14615_ (
);

FILL FILL_0_BUFX2_insert688 (
);

FILL FILL_0_BUFX2_insert689 (
);

FILL FILL_1__6838_ (
);

FILL FILL_2__13608_ (
);

FILL SFILL99320x54050 (
);

FILL FILL_0__14642_ (
);

FILL FILL_0__14222_ (
);

FILL FILL_5__11188_ (
);

FILL SFILL28760x74050 (
);

FILL FILL_0__9608_ (
);

FILL FILL_3__7705_ (
);

FILL SFILL59160x65050 (
);

FILL FILL_4__16407_ (
);

FILL FILL_4__11962_ (
);

FILL FILL_4__11542_ (
);

FILL SFILL64120x48050 (
);

FILL FILL_4__11122_ (
);

FILL FILL_1__16014_ (
);

FILL FILL_3__10955_ (
);

FILL FILL_3__10535_ (
);

FILL FILL_3__10115_ (
);

FILL FILL_0__15847_ (
);

INVX1 _15712_ (
    .A(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_6176_)
);

FILL FILL_0__15427_ (
);

FILL FILL_0__15007_ (
);

FILL FILL_0__10982_ (
);

FILL FILL_2__8594_ (
);

FILL FILL_0__10562_ (
);

FILL FILL_0__10142_ (
);

FILL SFILL49640x70050 (
);

FILL FILL_5__13754_ (
);

FILL FILL_5__13334_ (
);

OAI21X1 _7634_ (
    .A(_387_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .C(_388_),
    .Y(_328_[30])
);

FILL SFILL59160x20050 (
);

OAI21X1 _7214_ (
    .A(_168_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .C(_169_),
    .Y(_133_[18])
);

FILL FILL_4__9881_ (
);

FILL FILL_4__12747_ (
);

FILL FILL_4__9041_ (
);

FILL FILL_2__13781_ (
);

FILL FILL_4__12327_ (
);

FILL FILL_2__13361_ (
);

FILL FILL_2__6907_ (
);

FILL FILL_1__12774_ (
);

FILL FILL_1__12354_ (
);

FILL SFILL49560x77050 (
);

FILL FILL_0__9781_ (
);

FILL FILL_2__9799_ (
);

FILL FILL_2__9379_ (
);

FILL FILL_0__11767_ (
);

FILL FILL_0__9361_ (
);

FILL FILL_0__11347_ (
);

OAI22X1 _11632_ (
    .A(_2257_),
    .B(_2344__bF$buf1),
    .C(_2480_),
    .D(_2256_),
    .Y(_2736_)
);

OAI21X1 _11212_ (
    .A(_2326_),
    .B(_2330_),
    .C(_2117_),
    .Y(_2331_)
);

FILL FILL_6__15966_ (
);

FILL FILL_6__15546_ (
);

FILL FILL_4__16160_ (
);

FILL FILL_5__14959_ (
);

FILL FILL_3__15993_ (
);

FILL FILL_5__14539_ (
);

FILL FILL_3__15573_ (
);

FILL FILL_5__14119_ (
);

FILL FILL_3__15153_ (
);

OAI21X1 _8839_ (
    .A(_987_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .C(_988_),
    .Y(_978_[5])
);

FILL SFILL18760x72050 (
);

DFFSR _8419_ (
    .Q(\datapath_1.regfile_1.regOut[12] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_718_[13])
);

FILL FILL_1__7376_ (
);

FILL FILL_2__14986_ (
);

FILL FILL_2__14566_ (
);

FILL FILL_2__14146_ (
);

FILL FILL_0__15180_ (
);

FILL FILL_5__15900_ (
);

FILL SFILL89240x59050 (
);

FILL SFILL54120x46050 (
);

FILL FILL_1__13979_ (
);

FILL FILL_1__13559_ (
);

FILL FILL_1__13139_ (
);

OAI21X1 _12837_ (
    .A(_3562_),
    .B(vdd),
    .C(_3563_),
    .Y(_3555_[4])
);

FILL FILL_3__8243_ (
);

OAI21X1 _12417_ (
    .A(_3342_),
    .B(MemToReg_bF$buf1),
    .C(_3343_),
    .Y(\datapath_1.mux_wd3.dout [24])
);

FILL SFILL18680x79050 (
);

FILL FILL_5__8589_ (
);

FILL FILL_1__14920_ (
);

FILL FILL_1__14500_ (
);

FILL FILL_6__11886_ (
);

FILL FILL_6__11466_ (
);

FILL FILL_4__12080_ (
);

FILL FILL_0__13913_ (
);

FILL FILL_3__16358_ (
);

FILL FILL_5__10879_ (
);

FILL FILL_5__10039_ (
);

FILL FILL_5__9530_ (
);

FILL FILL_3__11493_ (
);

FILL FILL_3__11073_ (
);

FILL FILL_5__9110_ (
);

FILL FILL_0__16385_ (
);

AOI22X1 _16250_ (
    .A(_5562_),
    .B(\datapath_1.regfile_1.regOut[25] [30]),
    .C(\datapath_1.regfile_1.regOut[26] [30]),
    .D(_5484_),
    .Y(_6700_)
);

FILL FILL_2__10486_ (
);

FILL FILL_2__10066_ (
);

FILL FILL_5__11820_ (
);

FILL FILL_1__9522_ (
);

FILL FILL_5__11400_ (
);

FILL FILL_1__9102_ (
);

FILL SFILL89240x14050 (
);

FILL FILL_3__9868_ (
);

FILL FILL_4__10813_ (
);

FILL FILL_3__9028_ (
);

FILL FILL_5__14292_ (
);

OAI21X1 _8592_ (
    .A(_863_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_864_),
    .Y(_848_[8])
);

FILL FILL_1__15705_ (
);

DFFSR _8172_ (
    .Q(\datapath_1.regfile_1.regOut[10] [22]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_588_[22])
);

FILL FILL_6__7033_ (
);

FILL SFILL18680x34050 (
);

FILL FILL_4__13285_ (
);

FILL FILL_1__10420_ (
);

FILL FILL_1__10000_ (
);

FILL FILL_2__7865_ (
);

FILL FILL_3__12698_ (
);

FILL FILL_2__7445_ (
);

FILL FILL_3__12278_ (
);

FILL FILL111960x63050 (
);

OAI21X1 _12590_ (
    .A(_3438_),
    .B(vdd),
    .C(_3439_),
    .Y(_3425_[7])
);

NAND2X1 _12170_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.a [18]),
    .Y(_3167_)
);

FILL FILL_5__12605_ (
);

FILL FILL_6__16084_ (
);

INVX1 _6905_ (
    .A(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_4_)
);

FILL SFILL79240x57050 (
);

FILL FILL_4__8732_ (
);

FILL FILL_4__8312_ (
);

FILL FILL_2__12632_ (
);

FILL FILL_5__15497_ (
);

FILL FILL_5__15077_ (
);

FILL FILL_2__12212_ (
);

NAND2X1 _9797_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1485_)
);

NAND2X1 _9377_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1266_)
);

FILL FILL_1__11625_ (
);

FILL FILL_1__11205_ (
);

FILL FILL_0__8632_ (
);

NAND2X1 _10903_ (
    .A(_2048_),
    .B(_2050_),
    .Y(_2051_)
);

FILL FILL_0__10618_ (
);

FILL FILL_0__8212_ (
);

FILL FILL_1__14097_ (
);

FILL FILL_4__15851_ (
);

FILL FILL_4__15431_ (
);

FILL FILL_4__15011_ (
);

OAI22X1 _13795_ (
    .A(_4299_),
    .B(_3972__bF$buf1),
    .C(_3920_),
    .D(_4298_),
    .Y(_4300_)
);

INVX1 _13375_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_3887_)
);

FILL FILL_3__14844_ (
);

FILL FILL_3__14424_ (
);

FILL FILL_3__14004_ (
);

FILL FILL_4__9937_ (
);

FILL FILL_4__9517_ (
);

FILL FILL_2__13837_ (
);

FILL SFILL79240x12050 (
);

FILL FILL_0__14871_ (
);

FILL FILL_2__13417_ (
);

FILL FILL_0__14451_ (
);

FILL FILL_0__14031_ (
);

FILL FILL111880x25050 (
);

FILL FILL_3__7934_ (
);

FILL FILL_0__9417_ (
);

FILL FILL_4__16216_ (
);

FILL FILL_4__11771_ (
);

FILL FILL_4__11351_ (
);

FILL FILL_3__15629_ (
);

FILL FILL_3__15209_ (
);

FILL FILL_1__16243_ (
);

FILL FILL_3__10764_ (
);

FILL SFILL69240x55050 (
);

FILL FILL_0__15656_ (
);

AOI21X1 _15941_ (
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .B(_5649_),
    .C(_6398_),
    .Y(_6399_)
);

FILL FILL_0__15236_ (
);

OAI22X1 _15521_ (
    .A(_5485__bF$buf3),
    .B(_4484_),
    .C(_5483__bF$buf2),
    .D(_4495_),
    .Y(_5990_)
);

AOI22X1 _15101_ (
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .B(_5579_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_5580_)
);

FILL FILL_0__10791_ (
);

FILL FILL_0__10371_ (
);

FILL FILL_6__14150_ (
);

FILL FILL_3__8719_ (
);

FILL SFILL100120x5050 (
);

FILL FILL_5__13983_ (
);

FILL FILL_5__13563_ (
);

FILL FILL_5__13143_ (
);

OAI21X1 _7863_ (
    .A(_499_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_500_),
    .Y(_458_[21])
);

OAI21X1 _7443_ (
    .A(_280_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .C(_281_),
    .Y(_263_[9])
);

FILL FILL_4_BUFX2_insert910 (
);

DFFSR _7023_ (
    .Q(\datapath_1.regfile_1.regOut[1] [25]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_3_[25])
);

FILL FILL_4_BUFX2_insert911 (
);

FILL FILL_4__12976_ (
);

FILL FILL_4__9270_ (
);

FILL FILL_4_BUFX2_insert912 (
);

FILL FILL_4_BUFX2_insert913 (
);

FILL FILL_2__13590_ (
);

FILL FILL_4__12136_ (
);

FILL FILL_4_BUFX2_insert914 (
);

FILL FILL_2__13170_ (
);

FILL FILL_4_BUFX2_insert915 (
);

FILL FILL_4_BUFX2_insert916 (
);

FILL FILL_4_BUFX2_insert917 (
);

FILL FILL_4_BUFX2_insert918 (
);

FILL FILL_3__11969_ (
);

FILL FILL_4_BUFX2_insert919 (
);

FILL FILL_3__11549_ (
);

FILL FILL_1__12583_ (
);

FILL FILL_3__11129_ (
);

FILL FILL_1__12163_ (
);

OAI22X1 _16306_ (
    .A(_5485__bF$buf2),
    .B(_6754_),
    .C(_5483__bF$buf0),
    .D(_5413_),
    .Y(_6755_)
);

FILL FILL_0__11996_ (
);

FILL FILL_0__9590_ (
);

NOR3X1 _11861_ (
    .A(\datapath_1.ALUResult [10]),
    .B(\datapath_1.ALUResult [6]),
    .C(\datapath_1.ALUResult [16]),
    .Y(_2948_)
);

FILL FILL_0__9170_ (
);

FILL FILL_0__11576_ (
);

FILL SFILL69240x10050 (
);

OAI21X1 _11441_ (
    .A(_2555_),
    .B(_2556_),
    .C(_2323_),
    .Y(_2557_)
);

FILL FILL_0__11156_ (
);

OAI22X1 _11021_ (
    .A(_2136_),
    .B(_2137_),
    .C(_2138_),
    .D(_2139_),
    .Y(_2140_)
);

FILL FILL_3__12910_ (
);

FILL FILL_5__7193_ (
);

FILL FILL_2__11903_ (
);

FILL FILL_5__14768_ (
);

FILL FILL_5__14348_ (
);

FILL FILL_3__15382_ (
);

NAND2X1 _8648_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_902_)
);

NAND2X1 _8228_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_683_)
);

FILL FILL_1__7185_ (
);

FILL FILL_2__14795_ (
);

FILL FILL_2__14375_ (
);

FILL SFILL99400x42050 (
);

FILL SFILL69160x17050 (
);

FILL FILL_1__13788_ (
);

FILL FILL_1__13368_ (
);

FILL FILL_4__14702_ (
);

FILL FILL_3__8892_ (
);

FILL FILL_3__8472_ (
);

NAND2X1 _12646_ (
    .A(vdd),
    .B(memoryOutData[26]),
    .Y(_3477_)
);

NAND3X1 _12226_ (
    .A(_3206_),
    .B(_3207_),
    .C(_3208_),
    .Y(\datapath_1.alu_1.ALUInB [2])
);

FILL FILL_5__8398_ (
);

FILL SFILL99320x49050 (
);

FILL FILL_0__13722_ (
);

FILL FILL_0__13302_ (
);

FILL FILL_3__16167_ (
);

FILL FILL_5__10688_ (
);

FILL FILL_5__10268_ (
);

FILL FILL_0_BUFX2_insert1030 (
);

FILL FILL_0_BUFX2_insert1031 (
);

FILL FILL_0_BUFX2_insert1032 (
);

FILL FILL_0_BUFX2_insert1033 (
);

FILL FILL_0__16194_ (
);

FILL FILL_0_BUFX2_insert1034 (
);

FILL SFILL28760x69050 (
);

FILL FILL_0_BUFX2_insert1035 (
);

FILL FILL_0_BUFX2_insert1036 (
);

FILL FILL_2__10295_ (
);

FILL FILL_0_BUFX2_insert1037 (
);

FILL FILL_0_BUFX2_insert1038 (
);

FILL FILL_0_BUFX2_insert1039 (
);

FILL FILL_1__9751_ (
);

FILL FILL_4__15907_ (
);

FILL FILL_3__9677_ (
);

FILL FILL_2__16101_ (
);

FILL FILL_3_BUFX2_insert930 (
);

FILL FILL_3__9257_ (
);

FILL FILL_3_BUFX2_insert931 (
);

FILL FILL_3_BUFX2_insert932 (
);

FILL FILL_4__10622_ (
);

FILL FILL_3_BUFX2_insert933 (
);

FILL FILL_3_BUFX2_insert934 (
);

FILL FILL_3_BUFX2_insert935 (
);

FILL FILL_1__15934_ (
);

FILL FILL_1__15514_ (
);

FILL FILL_3_BUFX2_insert936 (
);

FILL FILL_3_BUFX2_insert937 (
);

FILL FILL_3_BUFX2_insert938 (
);

FILL FILL_3_BUFX2_insert939 (
);

FILL FILL_4__13094_ (
);

FILL FILL_0__14927_ (
);

FILL FILL_0__14507_ (
);

FILL FILL_2__7674_ (
);

FILL FILL_3__12087_ (
);

FILL FILL_6__13001_ (
);

FILL FILL_5__12834_ (
);

FILL SFILL89400x40050 (
);

FILL FILL_5__12414_ (
);

FILL SFILL59160x15050 (
);

FILL FILL_4__8961_ (
);

FILL FILL_4__8121_ (
);

FILL FILL_4__11827_ (
);

FILL FILL_2__12861_ (
);

FILL FILL_4__11407_ (
);

FILL FILL_2__12441_ (
);

FILL FILL_2__12021_ (
);

DFFSR _9186_ (
    .Q(\datapath_1.regfile_1.regOut[18] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_1108_[12])
);

FILL FILL_1__11854_ (
);

FILL FILL_4__14299_ (
);

FILL FILL_1__11434_ (
);

FILL FILL_1__11014_ (
);

FILL FILL_2__8879_ (
);

FILL FILL_0__8861_ (
);

FILL FILL_2__8459_ (
);

FILL FILL_0__8441_ (
);

FILL FILL_0__10427_ (
);

FILL FILL_0__8021_ (
);

DFFSR _10712_ (
    .Q(\datapath_1.regfile_1.regOut[30] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_1888_[2])
);

FILL FILL_0__10007_ (
);

FILL FILL_6__14626_ (
);

FILL FILL_5__6884_ (
);

FILL FILL_4__15660_ (
);

FILL FILL_6__14206_ (
);

FILL FILL_4__15240_ (
);

DFFSR _13184_ (
    .Q(\datapath_1.mux_iord.din0 [9]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3685_[9])
);

FILL FILL_5__13619_ (
);

FILL SFILL79400x83050 (
);

FILL FILL_2__9400_ (
);

FILL FILL_3__14653_ (
);

FILL SFILL18760x67050 (
);

FILL FILL_3__14233_ (
);

DFFSR _7919_ (
    .Q(\datapath_1.regfile_1.regOut[8] [25]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_458_[25])
);

FILL FILL_1__6876_ (
);

FILL FILL_4__9746_ (
);

FILL FILL_2__13646_ (
);

FILL FILL_2__13226_ (
);

FILL FILL_0__14680_ (
);

FILL FILL_0__14260_ (
);

FILL FILL_1__12639_ (
);

FILL FILL_1__12219_ (
);

FILL FILL_3__7743_ (
);

FILL FILL_0__9646_ (
);

FILL FILL_0__9226_ (
);

FILL FILL_3__7323_ (
);

INVX1 _11917_ (
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_2986_)
);

FILL FILL_5__7249_ (
);

FILL FILL_4__16025_ (
);

FILL FILL_6__10966_ (
);

FILL FILL_4__11580_ (
);

AOI22X1 _14389_ (
    .A(\datapath_1.regfile_1.regOut[28] [19]),
    .B(_3894_),
    .C(_4038__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_4882_)
);

FILL FILL_4__11160_ (
);

FILL FILL_3__15858_ (
);

FILL FILL_3__15438_ (
);

FILL FILL_3__15018_ (
);

FILL FILL_1__16052_ (
);

FILL FILL_3__10993_ (
);

FILL FILL_3__10573_ (
);

FILL FILL_5__8610_ (
);

FILL FILL_3__10153_ (
);

FILL SFILL18760x22050 (
);

FILL FILL_0__15885_ (
);

FILL FILL_6_BUFX2_insert444 (
);

OAI22X1 _15750_ (
    .A(_5530__bF$buf0),
    .B(_4787_),
    .C(_5532__bF$buf1),
    .D(_6212_),
    .Y(_6213_)
);

FILL FILL_0__15465_ (
);

INVX1 _15330_ (
    .A(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_5804_)
);

FILL FILL_0__15045_ (
);

FILL FILL_6_BUFX2_insert449 (
);

FILL FILL_0__10180_ (
);

FILL FILL_5__10900_ (
);

FILL FILL_1__8602_ (
);

FILL FILL_3__8528_ (
);

FILL FILL_3__8108_ (
);

FILL FILL_5__13792_ (
);

FILL FILL_5__13372_ (
);

OAI21X1 _7672_ (
    .A(_456_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_457_),
    .Y(_393_[0])
);

NAND2X1 _7252_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_195_)
);

FILL SFILL79320x45050 (
);

FILL SFILL18680x29050 (
);

FILL SFILL64040x50 (
);

FILL FILL_4__12785_ (
);

FILL FILL_4__12365_ (
);

FILL FILL_2__6945_ (
);

FILL FILL_3__11778_ (
);

FILL FILL111960x58050 (
);

FILL FILL_3__11358_ (
);

FILL FILL_1__12392_ (
);

OAI22X1 _16115_ (
    .A(_6568_),
    .B(_5548__bF$buf1),
    .C(_5489__bF$buf0),
    .D(_5185_),
    .Y(_6569_)
);

FILL FILL_0__11385_ (
);

NOR2X1 _11670_ (
    .A(_2771_),
    .B(_2769_),
    .Y(_2772_)
);

NAND2X1 _11250_ (
    .A(_2367_),
    .B(_2368_),
    .Y(_2369_)
);

FILL FILL_1__9807_ (
);

FILL FILL_4__7812_ (
);

FILL FILL_5__14997_ (
);

FILL FILL_5__14577_ (
);

FILL FILL_2__11712_ (
);

FILL FILL_5__14157_ (
);

FILL FILL_3__15191_ (
);

NAND2X1 _8877_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1014_)
);

NAND2X1 _8457_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_795_)
);

DFFSR _8037_ (
    .Q(\datapath_1.regfile_1.regOut[9] [15]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_523_[15])
);

FILL FILL_1__10705_ (
);

FILL FILL_2__14184_ (
);

FILL FILL_0__7712_ (
);

FILL FILL_1__13597_ (
);

FILL FILL_4__14931_ (
);

FILL FILL_4__14511_ (
);

FILL FILL111960x13050 (
);

NAND2X1 _12875_ (
    .A(vdd),
    .B(\datapath_1.rd1 [17]),
    .Y(_3589_)
);

NAND2X1 _12455_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [5]),
    .Y(_3370_)
);

NAND3X1 _12035_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[12]),
    .C(_3032__bF$buf3),
    .Y(_3072_)
);

FILL FILL_3__13924_ (
);

FILL FILL_3__13504_ (
);

FILL FILL_5_BUFX2_insert460 (
);

FILL FILL_5_BUFX2_insert461 (
);

FILL FILL_2__12917_ (
);

FILL FILL_5_BUFX2_insert462 (
);

FILL FILL_0__13951_ (
);

FILL FILL_5_BUFX2_insert463 (
);

FILL FILL_0__13531_ (
);

FILL FILL_3__16396_ (
);

FILL FILL_0__13111_ (
);

FILL FILL_5_BUFX2_insert464 (
);

FILL FILL_5_BUFX2_insert465 (
);

FILL FILL_5__10497_ (
);

FILL FILL_5_BUFX2_insert466 (
);

FILL FILL_5_BUFX2_insert467 (
);

FILL FILL_1__8199_ (
);

FILL FILL_5_BUFX2_insert468 (
);

FILL FILL_5_BUFX2_insert469 (
);

FILL FILL_2__15389_ (
);

FILL FILL_5__16303_ (
);

FILL FILL_0__8917_ (
);

FILL FILL_1__9980_ (
);

FILL FILL_1__9140_ (
);

FILL FILL_4__15716_ (
);

FILL FILL_2__16330_ (
);

FILL FILL_3__9486_ (
);

FILL FILL_4__10431_ (
);

FILL FILL_4__10011_ (
);

FILL FILL_3__14709_ (
);

FILL FILL_1__15743_ (
);

FILL FILL_1__15323_ (
);

FILL FILL_0__14736_ (
);

INVX1 _14601_ (
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_5089_)
);

FILL FILL_0__14316_ (
);

FILL FILL_2__7483_ (
);

FILL FILL_2__7063_ (
);

FILL FILL_5__12643_ (
);

FILL FILL_5__12223_ (
);

OAI21X1 _6943_ (
    .A(_28_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_29_),
    .Y(_3_[13])
);

FILL FILL_2_BUFX2_insert590 (
);

FILL FILL_2_BUFX2_insert591 (
);

FILL FILL_2_BUFX2_insert592 (
);

FILL FILL_4__8770_ (
);

FILL FILL_2_BUFX2_insert593 (
);

FILL FILL_4__8350_ (
);

FILL FILL_2_BUFX2_insert594 (
);

FILL FILL_4__11636_ (
);

FILL FILL_2_BUFX2_insert595 (
);

FILL FILL_4__11216_ (
);

FILL FILL_2_BUFX2_insert596 (
);

FILL FILL_2__12250_ (
);

FILL FILL_2_BUFX2_insert597 (
);

FILL FILL_2_BUFX2_insert598 (
);

FILL FILL_1__16108_ (
);

FILL FILL_2_BUFX2_insert599 (
);

FILL FILL_3__10629_ (
);

FILL FILL_1__11663_ (
);

FILL FILL_1__11243_ (
);

INVX1 _15806_ (
    .A(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_6268_)
);

FILL SFILL104360x75050 (
);

NAND2X1 _10941_ (
    .A(\control_1.op [0]),
    .B(\control_1.op [1]),
    .Y(_2075_)
);

FILL FILL_2__8268_ (
);

FILL FILL_0__8250_ (
);

FILL FILL_0__10656_ (
);

OAI21X1 _10521_ (
    .A(_1844_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .C(_1845_),
    .Y(_1823_[11])
);

FILL FILL_0__10236_ (
);

DFFSR _10101_ (
    .Q(\datapath_1.regfile_1.regOut[25] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_1563_[31])
);

FILL FILL_5__13848_ (
);

FILL FILL_5__13428_ (
);

FILL FILL_3__14882_ (
);

FILL FILL_3__14462_ (
);

FILL FILL_5__13008_ (
);

FILL FILL_3__14042_ (
);

NAND2X1 _7728_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_431_)
);

NAND2X1 _7308_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_212_)
);

FILL FILL_4__9975_ (
);

FILL FILL_4__9555_ (
);

FILL FILL_4__9135_ (
);

FILL FILL_2__13875_ (
);

FILL FILL_2__13455_ (
);

FILL SFILL99400x37050 (
);

FILL FILL_2__13035_ (
);

FILL FILL_1__12868_ (
);

FILL FILL_1__12448_ (
);

FILL FILL_1__12028_ (
);

FILL FILL_3__7972_ (
);

FILL FILL_0__9875_ (
);

FILL FILL_3__7552_ (
);

FILL FILL112440x81050 (
);

FILL FILL_0__9035_ (
);

OAI21X1 _11726_ (
    .A(_2172_),
    .B(_2811_),
    .C(_2823_),
    .Y(_2824_)
);

OAI21X1 _11306_ (
    .A(_2246_),
    .B(_2240_),
    .C(_2245_),
    .Y(_2425_)
);

FILL FILL_5__7478_ (
);

FILL SFILL104360x30050 (
);

FILL FILL112360x50 (
);

FILL FILL_4__16254_ (
);

FILL FILL_5__7058_ (
);

INVX1 _14198_ (
    .A(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_4695_)
);

FILL FILL_3__15667_ (
);

FILL FILL_3__15247_ (
);

FILL FILL_1__16281_ (
);

FILL FILL_3__10382_ (
);

FILL FILL_0__15694_ (
);

FILL FILL_0__15274_ (
);

FILL FILL_1__8831_ (
);

FILL SFILL104280x37050 (
);

FILL FILL_2__15601_ (
);

FILL FILL_3__8757_ (
);

FILL FILL_3__8337_ (
);

NAND2X1 _7481_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_307_)
);

NAND2X1 _7061_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_88_)
);

FILL FILL_4__12594_ (
);

FILL FILL_4__12174_ (
);

FILL SFILL114520x1050 (
);

FILL FILL_5__9624_ (
);

FILL FILL_3__11587_ (
);

FILL FILL_3__11167_ (
);

FILL SFILL114440x6050 (
);

OAI21X1 _16344_ (
    .A(_6782_),
    .B(gnd),
    .C(_6783_),
    .Y(_6769_[7])
);

FILL FILL_0__16059_ (
);

FILL FILL_0__11194_ (
);

FILL SFILL89400x35050 (
);

FILL FILL_5__11914_ (
);

FILL SFILL28760x19050 (
);

FILL FILL_1__9616_ (
);

FILL FILL_6__15393_ (
);

FILL FILL_4__7621_ (
);

FILL FILL_4__10907_ (
);

FILL FILL_4__7201_ (
);

FILL FILL_2__11941_ (
);

FILL FILL_5__14386_ (
);

FILL FILL_2__11521_ (
);

FILL FILL_2__11101_ (
);

DFFSR _8686_ (
    .Q(\datapath_1.regfile_1.regOut[14] [24]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_848_[24])
);

FILL SFILL113720x8050 (
);

INVX1 _8266_ (
    .A(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_708_)
);

FILL FILL_4__13799_ (
);

FILL FILL_1__10934_ (
);

FILL FILL_4__13379_ (
);

FILL FILL_1__10514_ (
);

FILL FILL_2__7959_ (
);

FILL FILL_0__7941_ (
);

BUFX2 BUFX2_insert280 (
    .A(_3931_),
    .Y(_3931__bF$buf0)
);

FILL FILL_0__7101_ (
);

FILL FILL_2__7119_ (
);

BUFX2 BUFX2_insert281 (
    .A(_5483_),
    .Y(_5483__bF$buf4)
);

BUFX2 BUFX2_insert282 (
    .A(_5483_),
    .Y(_5483__bF$buf3)
);

BUFX2 BUFX2_insert283 (
    .A(_5483_),
    .Y(_5483__bF$buf2)
);

BUFX2 BUFX2_insert284 (
    .A(_5483_),
    .Y(_5483__bF$buf1)
);

BUFX2 BUFX2_insert285 (
    .A(_5483_),
    .Y(_5483__bF$buf0)
);

FILL FILL_4__14740_ (
);

BUFX2 BUFX2_insert286 (
    .A(_5539_),
    .Y(_5539__bF$buf4)
);

FILL FILL_4__14320_ (
);

BUFX2 BUFX2_insert287 (
    .A(_5539_),
    .Y(_5539__bF$buf3)
);

BUFX2 BUFX2_insert288 (
    .A(_5539_),
    .Y(_5539__bF$buf2)
);

FILL FILL_3__8090_ (
);

DFFSR _12684_ (
    .Q(\datapath_1.Data [21]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[21])
);

FILL FILL_0__12399_ (
);

BUFX2 BUFX2_insert289 (
    .A(_5539_),
    .Y(_5539__bF$buf1)
);

NAND3X1 _12264_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [14]),
    .C(_3198__bF$buf2),
    .Y(_3237_)
);

FILL FILL_2__8900_ (
);

FILL FILL_3__13733_ (
);

FILL FILL_3__13313_ (
);

FILL FILL_4__8826_ (
);

FILL SFILL94280x41050 (
);

FILL FILL_2__12726_ (
);

FILL FILL_0__13760_ (
);

FILL FILL_2__12306_ (
);

FILL FILL_0__13340_ (
);

FILL FILL_1__11719_ (
);

FILL FILL_2__15198_ (
);

FILL FILL_5__16112_ (
);

FILL FILL_0__8726_ (
);

FILL SFILL33960x37050 (
);

FILL FILL_4__15945_ (
);

FILL FILL_4__15525_ (
);

FILL FILL_4__15105_ (
);

FILL FILL_3__9295_ (
);

INVX1 _13889_ (
    .A(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_4392_)
);

FILL FILL_4__10660_ (
);

INVX1 _13469_ (
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_3981_)
);

FILL FILL_4__10240_ (
);

DFFSR _13049_ (
    .Q(_2_[2]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3620_[2])
);

FILL FILL_3__14938_ (
);

FILL FILL_1__15972_ (
);

FILL FILL_3__14518_ (
);

FILL FILL_1__15552_ (
);

FILL FILL_1__15132_ (
);

FILL SFILL18760x17050 (
);

FILL FILL_0__14965_ (
);

OAI22X1 _14830_ (
    .A(_5312_),
    .B(_3955__bF$buf1),
    .C(_3971__bF$buf4),
    .D(_5313_),
    .Y(_5314_)
);

FILL FILL_0__14545_ (
);

FILL FILL_0__14125_ (
);

OAI22X1 _14410_ (
    .A(_3947__bF$buf2),
    .B(_4901_),
    .C(_3935__bF$buf1),
    .D(_4900_),
    .Y(_4902_)
);

FILL FILL_2__7292_ (
);

FILL FILL_3__7608_ (
);

FILL FILL_5__12872_ (
);

FILL FILL_5__12452_ (
);

FILL FILL_5__12032_ (
);

FILL SFILL33800x2050 (
);

FILL FILL_4__11865_ (
);

FILL FILL_4__11445_ (
);

FILL SFILL74280x2050 (
);

FILL FILL_4__11025_ (
);

FILL FILL_1__16337_ (
);

FILL FILL_3__10438_ (
);

FILL FILL_1__11892_ (
);

FILL SFILL84200x82050 (
);

FILL FILL_3__10018_ (
);

FILL FILL_1__11472_ (
);

FILL FILL_1__11052_ (
);

NOR2X1 _15615_ (
    .A(_6077_),
    .B(_6080_),
    .Y(_6081_)
);

FILL FILL_0__10885_ (
);

FILL FILL_2__8497_ (
);

FILL FILL_2__8077_ (
);

OAI21X1 _10750_ (
    .A(_1956_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .C(_1957_),
    .Y(_1953_[2])
);

FILL FILL_0__10045_ (
);

DFFSR _10330_ (
    .Q(\datapath_1.regfile_1.regOut[27] [4]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_1693_[4])
);

FILL FILL_5__13657_ (
);

FILL FILL_5__13237_ (
);

FILL FILL_3__14691_ (
);

FILL FILL_3__14271_ (
);

NAND2X1 _7957_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_543_)
);

DFFSR _7537_ (
    .Q(\datapath_1.regfile_1.regOut[5] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_263_[27])
);

INVX1 _7117_ (
    .A(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_125_)
);

FILL FILL_4__9784_ (
);

FILL FILL_4__9364_ (
);

FILL FILL_2__13684_ (
);

FILL FILL_2__13264_ (
);

FILL FILL_1__12257_ (
);

FILL FILL_0__9684_ (
);

OAI21X1 _11955_ (
    .A(_3010_),
    .B(IorD_bF$buf7),
    .C(_3011_),
    .Y(_1_[22])
);

FILL FILL_0__9264_ (
);

FILL FILL_3__7361_ (
);

NAND3X1 _11535_ (
    .A(_2218_),
    .B(_2411_),
    .C(_2645_),
    .Y(_2646_)
);

NOR2X1 _11115_ (
    .A(_2232_),
    .B(_2233_),
    .Y(_2234_)
);

FILL FILL_6__15869_ (
);

FILL FILL_6__15449_ (
);

FILL FILL_5__7287_ (
);

FILL FILL_4__16063_ (
);

FILL SFILL29240x42050 (
);

FILL SFILL110120x12050 (
);

FILL FILL_3__15896_ (
);

FILL FILL_0__12611_ (
);

FILL FILL_3__15476_ (
);

FILL FILL_3__15056_ (
);

FILL FILL_1__16090_ (
);

FILL FILL_1__7699_ (
);

FILL FILL_3__10191_ (
);

FILL FILL_6_BUFX2_insert822 (
);

FILL FILL_2__14889_ (
);

FILL FILL_2__14469_ (
);

FILL FILL_2__14049_ (
);

FILL FILL_0__15083_ (
);

FILL FILL_5__15803_ (
);

FILL FILL_6_BUFX2_insert827 (
);

FILL SFILL114440x20050 (
);

FILL FILL_1__8640_ (
);

FILL FILL_1__8220_ (
);

FILL FILL_2__15830_ (
);

FILL FILL_2__15410_ (
);

FILL FILL_3__8986_ (
);

FILL FILL_3__8566_ (
);

FILL FILL_3__8146_ (
);

FILL FILL_6__6991_ (
);

FILL FILL_1__14823_ (
);

FILL FILL_1__14403_ (
);

NAND2X1 _7290_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_200_)
);

FILL FILL_6__11789_ (
);

FILL FILL_6__11369_ (
);

FILL SFILL104840x77050 (
);

FILL FILL_0__13816_ (
);

FILL FILL_2__6983_ (
);

FILL FILL_5__9853_ (
);

FILL FILL_3__11396_ (
);

FILL FILL_5__9013_ (
);

FILL FILL_0__16288_ (
);

FILL FILL_6__12310_ (
);

NAND2X1 _16153_ (
    .A(_6600_),
    .B(_6605_),
    .Y(_6606_)
);

FILL FILL_2__10389_ (
);

FILL FILL_5__11723_ (
);

FILL FILL_1__9425_ (
);

FILL FILL_5__11303_ (
);

FILL FILL_1__9005_ (
);

FILL FILL_4__7850_ (
);

FILL SFILL104520x50 (
);

FILL FILL_4__7430_ (
);

FILL FILL_2__11750_ (
);

FILL FILL_5__14195_ (
);

FILL FILL_2__11330_ (
);

INVX1 _8495_ (
    .A(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_820_)
);

FILL FILL_1__15608_ (
);

INVX1 _8075_ (
    .A(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_601_)
);

FILL FILL_1__10743_ (
);

FILL FILL_1__10323_ (
);

FILL FILL_0__7750_ (
);

FILL FILL_0__7330_ (
);

FILL FILL_2__7348_ (
);

FILL FILL_6__13935_ (
);

FILL FILL_6__13515_ (
);

INVX1 _12493_ (
    .A(ALUOut[18]),
    .Y(_3395_)
);

AOI22X1 _12073_ (
    .A(\datapath_1.ALUResult [21]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3101_)
);

FILL FILL_5__12508_ (
);

FILL FILL_3__13962_ (
);

FILL FILL_3__13542_ (
);

FILL FILL_3__13122_ (
);

FILL SFILL8600x9050 (
);

FILL FILL_4__8635_ (
);

FILL FILL_4__8215_ (
);

FILL FILL_5_BUFX2_insert840 (
);

FILL FILL_5_BUFX2_insert841 (
);

FILL FILL_2__12955_ (
);

FILL FILL_5_BUFX2_insert842 (
);

FILL FILL_2__12115_ (
);

FILL FILL_5_BUFX2_insert843 (
);

FILL FILL_5_BUFX2_insert844 (
);

FILL FILL_5_BUFX2_insert845 (
);

FILL FILL_5_BUFX2_insert846 (
);

FILL FILL_5_BUFX2_insert847 (
);

FILL FILL_1__11948_ (
);

FILL FILL_5_BUFX2_insert848 (
);

FILL FILL_5_BUFX2_insert849 (
);

FILL FILL_1__11528_ (
);

FILL FILL_1__11108_ (
);

FILL FILL_5__16341_ (
);

FILL FILL_0__8955_ (
);

FILL FILL112440x76050 (
);

NAND2X1 _10806_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1995_)
);

FILL FILL_0__8115_ (
);

FILL FILL_5__6978_ (
);

FILL FILL_4__15754_ (
);

FILL FILL_4__15334_ (
);

NAND3X1 _13698_ (
    .A(_4194_),
    .B(_4197_),
    .C(_4204_),
    .Y(_4205_)
);

NAND2X1 _13278_ (
    .A(_3817_),
    .B(_3803_),
    .Y(_3818_)
);

FILL FILL_2__9914_ (
);

FILL FILL_3__14747_ (
);

FILL FILL_1__15781_ (
);

FILL FILL_3__14327_ (
);

FILL FILL_1__15361_ (
);

FILL FILL112040x62050 (
);

FILL FILL_0__14774_ (
);

FILL FILL_0__14354_ (
);

FILL FILL_3__7837_ (
);

FILL FILL_3__7417_ (
);

FILL SFILL73400x76050 (
);

FILL FILL_5__12261_ (
);

NAND2X1 _6981_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_55_)
);

FILL FILL112440x31050 (
);

FILL FILL_2_BUFX2_insert970 (
);

FILL FILL_2_BUFX2_insert971 (
);

FILL FILL_4__16119_ (
);

FILL FILL_2_BUFX2_insert972 (
);

FILL FILL_2_BUFX2_insert973 (
);

FILL FILL_2_BUFX2_insert974 (
);

FILL FILL_4__11674_ (
);

FILL FILL_2_BUFX2_insert975 (
);

FILL FILL_4__11254_ (
);

FILL FILL_2_BUFX2_insert976 (
);

FILL FILL_2_BUFX2_insert977 (
);

FILL FILL_2_BUFX2_insert978 (
);

FILL FILL_2_BUFX2_insert979 (
);

FILL FILL_1__16146_ (
);

FILL FILL_5__8704_ (
);

FILL FILL_3__10667_ (
);

FILL FILL_3__10247_ (
);

FILL FILL_1__11281_ (
);

FILL FILL_0__15979_ (
);

FILL FILL_0__15559_ (
);

INVX1 _15844_ (
    .A(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_6305_)
);

OAI22X1 _15424_ (
    .A(_5472__bF$buf0),
    .B(_4415_),
    .C(_4414_),
    .D(_5552__bF$buf1),
    .Y(_5895_)
);

FILL FILL_0__15139_ (
);

INVX2 _15004_ (
    .A(_5483__bF$buf0),
    .Y(_5484_)
);

FILL FILL_0__10694_ (
);

FILL FILL_0__10274_ (
);

FILL FILL_6__14053_ (
);

FILL FILL_5__13886_ (
);

FILL FILL_5__13466_ (
);

FILL FILL_5__13046_ (
);

DFFSR _7766_ (
    .Q(\datapath_1.regfile_1.regOut[7] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_393_[0])
);

FILL FILL_3__14080_ (
);

INVX1 _7346_ (
    .A(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_237_)
);

FILL FILL_4__9593_ (
);

FILL FILL_4__12879_ (
);

FILL FILL_4__9173_ (
);

FILL FILL_4__12459_ (
);

FILL FILL_4__12039_ (
);

FILL FILL_2__13493_ (
);

FILL FILL_5__9909_ (
);

FILL FILL_1__12486_ (
);

FILL FILL_1__12066_ (
);

FILL FILL_4__13820_ (
);

NOR2X1 _16209_ (
    .A(_6659_),
    .B(_6657_),
    .Y(_6660_)
);

FILL FILL_4__13400_ (
);

FILL FILL_3__7590_ (
);

FILL FILL_0__11899_ (
);

FILL FILL_0__9493_ (
);

FILL FILL_3__7170_ (
);

AOI22X1 _11764_ (
    .A(_2478_),
    .B(_2364_),
    .C(_2137_),
    .D(_2341__bF$buf3),
    .Y(_2859_)
);

FILL FILL_0__11479_ (
);

INVX8 _11344_ (
    .A(_2337_),
    .Y(_2462_)
);

FILL FILL_0__11059_ (
);

FILL FILL_5__7096_ (
);

FILL FILL_4__16292_ (
);

FILL SFILL94280x36050 (
);

FILL FILL_6__10393_ (
);

FILL FILL_2__11806_ (
);

FILL FILL_0__12840_ (
);

FILL FILL_0__12420_ (
);

FILL FILL_3__15285_ (
);

FILL FILL_0__12000_ (
);

FILL FILL_1__7088_ (
);

FILL FILL_2__14698_ (
);

FILL FILL_2__14278_ (
);

FILL FILL_5__15612_ (
);

FILL FILL_0__7806_ (
);

INVX1 _9912_ (
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_1541_)
);

FILL SFILL13560x2050 (
);

FILL FILL_4__14605_ (
);

FILL FILL_1_BUFX2_insert990 (
);

FILL FILL_1_BUFX2_insert991 (
);

FILL FILL_3__8375_ (
);

FILL FILL_1_BUFX2_insert992 (
);

INVX1 _12969_ (
    .A(_2_[6]),
    .Y(_3631_)
);

FILL FILL_1_BUFX2_insert993 (
);

DFFSR _12549_ (
    .Q(ALUOut[14]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3360_[14])
);

FILL FILL_1_BUFX2_insert994 (
);

OAI21X1 _12129_ (
    .A(_3138_),
    .B(ALUSrcA_bF$buf4),
    .C(_3139_),
    .Y(\datapath_1.alu_1.ALUInA [4])
);

FILL FILL_1_BUFX2_insert995 (
);

FILL FILL_1_BUFX2_insert996 (
);

FILL FILL_1__14632_ (
);

FILL FILL_1_BUFX2_insert997 (
);

FILL FILL_1__14212_ (
);

FILL FILL_1_BUFX2_insert998 (
);

FILL FILL_1_BUFX2_insert999 (
);

FILL FILL_0__13625_ (
);

AOI22X1 _13910_ (
    .A(\datapath_1.regfile_1.regOut[4] [9]),
    .B(_3891__bF$buf1),
    .C(_3998__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_4413_)
);

FILL FILL_5__9662_ (
);

FILL FILL_5__9242_ (
);

FILL SFILL105240x62050 (
);

NAND2X1 _16382_ (
    .A(gnd),
    .B(gnd),
    .Y(_6809_)
);

FILL FILL_0__16097_ (
);

FILL FILL_5__11952_ (
);

FILL FILL_1__9654_ (
);

FILL FILL_5__11532_ (
);

FILL FILL_5__11112_ (
);

FILL FILL_1__9234_ (
);

FILL SFILL8680x53050 (
);

FILL FILL_2__16004_ (
);

FILL FILL_4__10945_ (
);

FILL FILL_4__10525_ (
);

FILL FILL_4__10105_ (
);

FILL FILL_1__15837_ (
);

FILL FILL_1__15417_ (
);

FILL FILL_1__10972_ (
);

FILL FILL_1__10552_ (
);

FILL FILL_1__10132_ (
);

FILL FILL_2__7997_ (
);

BUFX2 BUFX2_insert660 (
    .A(_3037_),
    .Y(_3037__bF$buf1)
);

FILL FILL_2__7577_ (
);

BUFX2 BUFX2_insert661 (
    .A(_3037_),
    .Y(_3037__bF$buf0)
);

BUFX2 BUFX2_insert662 (
    .A(_2481_),
    .Y(_2481__bF$buf3)
);

BUFX2 BUFX2_insert663 (
    .A(_2481_),
    .Y(_2481__bF$buf2)
);

BUFX2 BUFX2_insert664 (
    .A(_2481_),
    .Y(_2481__bF$buf1)
);

BUFX2 BUFX2_insert665 (
    .A(_2481_),
    .Y(_2481__bF$buf0)
);

BUFX2 BUFX2_insert666 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf4 )
);

BUFX2 BUFX2_insert667 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf3 )
);

BUFX2 BUFX2_insert668 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf2 )
);

BUFX2 BUFX2_insert669 (
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf1 )
);

FILL FILL_5__12737_ (
);

FILL FILL_3__13771_ (
);

FILL FILL_5__12317_ (
);

FILL FILL_3__13351_ (
);

FILL SFILL8600x51050 (
);

FILL FILL_4__8864_ (
);

FILL FILL_4__8444_ (
);

FILL FILL_2__12764_ (
);

FILL FILL_2__12344_ (
);

OAI21X1 _9089_ (
    .A(_1113_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .C(_1114_),
    .Y(_1108_[3])
);

FILL FILL_1__11757_ (
);

FILL FILL_1__11337_ (
);

FILL FILL_0__8764_ (
);

FILL FILL_3__6861_ (
);

FILL FILL_5__16150_ (
);

FILL FILL_6__9731_ (
);

FILL FILL_0__8344_ (
);

NAND2X1 _10615_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .Y(_1952_)
);

FILL FILL_4__15983_ (
);

FILL FILL_4__15563_ (
);

FILL FILL_6__14109_ (
);

FILL FILL_4__15143_ (
);

FILL SFILL13640x52050 (
);

OAI21X1 _13087_ (
    .A(_3688_),
    .B(PCEn_bF$buf5),
    .C(_3689_),
    .Y(_3685_[2])
);

FILL FILL_3__14976_ (
);

FILL FILL_2__9723_ (
);

FILL FILL_3__14556_ (
);

FILL FILL_3__14136_ (
);

FILL FILL_1__15590_ (
);

FILL SFILL109480x32050 (
);

FILL FILL_1__15170_ (
);

FILL FILL_4__9649_ (
);

FILL FILL_4__9229_ (
);

FILL FILL_2__13969_ (
);

FILL FILL_2__13549_ (
);

FILL FILL_0__14583_ (
);

FILL FILL_2__13129_ (
);

FILL FILL_0__14163_ (
);

FILL FILL_1__7720_ (
);

FILL FILL_1__7300_ (
);

FILL FILL_2__14910_ (
);

FILL SFILL74200x75050 (
);

FILL FILL_0__9549_ (
);

FILL FILL_3__7226_ (
);

FILL FILL_0__9129_ (
);

FILL FILL_5__12490_ (
);

FILL FILL_5__12070_ (
);

FILL FILL_1__13903_ (
);

FILL FILL_4__16348_ (
);

FILL FILL_6__10449_ (
);

FILL FILL_4__11483_ (
);

FILL FILL_4__11063_ (
);

FILL FILL_1__16375_ (
);

FILL SFILL99480x81050 (
);

FILL FILL_3__10896_ (
);

FILL FILL_5__8513_ (
);

FILL FILL_3__10056_ (
);

FILL FILL_1__11090_ (
);

FILL SFILL59800x38050 (
);

FILL FILL_0__15788_ (
);

INVX1 _15653_ (
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_6118_)
);

FILL FILL_0__15368_ (
);

OAI22X1 _15233_ (
    .A(_5466__bF$buf3),
    .B(_5708_),
    .C(_4178_),
    .D(_5483__bF$buf4),
    .Y(_5709_)
);

FILL FILL_5__10803_ (
);

FILL FILL_1__8505_ (
);

FILL FILL_4__6930_ (
);

FILL FILL_2__10830_ (
);

FILL FILL_5__13695_ (
);

FILL FILL_5__13275_ (
);

FILL FILL_2__10410_ (
);

FILL SFILL74200x30050 (
);

INVX1 _7995_ (
    .A(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_568_)
);

INVX1 _7575_ (
    .A(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_349_)
);

DFFSR _7155_ (
    .Q(\datapath_1.regfile_1.regOut[2] [29]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_68_[29])
);

FILL FILL_4__12268_ (
);

FILL FILL_2__6848_ (
);

FILL FILL_5__9718_ (
);

FILL FILL_1__12295_ (
);

DFFSR _16438_ (
    .Q(\datapath_1.regfile_1.regOut[0] [21]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_6769_[21])
);

OAI22X1 _16018_ (
    .A(_6473_),
    .B(_5503__bF$buf0),
    .C(_5504__bF$buf4),
    .D(_5130_),
    .Y(_6474_)
);

AOI22X1 _11993_ (
    .A(\datapath_1.ALUResult [1]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3041_)
);

FILL SFILL43720x46050 (
);

AOI22X1 _11573_ (
    .A(_2234_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf1),
    .D(_2235_),
    .Y(_2681_)
);

FILL FILL_0__11288_ (
);

NOR2X1 _11153_ (
    .A(\datapath_1.alu_1.ALUInB [18]),
    .B(_2271_),
    .Y(_2272_)
);

FILL FILL_3__12622_ (
);

FILL FILL_3__12202_ (
);

FILL FILL_4__7715_ (
);

FILL FILL_2__11615_ (
);

FILL SFILL33800x82050 (
);

FILL FILL_3__15094_ (
);

FILL FILL112120x50050 (
);

FILL FILL_2__14087_ (
);

FILL FILL_5__15841_ (
);

FILL FILL_5__15421_ (
);

FILL FILL_5__15001_ (
);

FILL FILL_0__7615_ (
);

INVX1 _9721_ (
    .A(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_1434_)
);

OAI21X1 _9301_ (
    .A(_1234_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .C(_1235_),
    .Y(_1173_[31])
);

FILL FILL_4__14834_ (
);

FILL FILL_4__14414_ (
);

OAI21X1 _12778_ (
    .A(_3543_),
    .B(IRWrite_bF$buf7),
    .C(_3544_),
    .Y(_3490_[27])
);

FILL FILL_3__8184_ (
);

INVX1 _12358_ (
    .A(ALUOut[5]),
    .Y(_3304_)
);

FILL FILL_3__13827_ (
);

FILL FILL_1__14861_ (
);

FILL FILL_3__13407_ (
);

FILL FILL_1__14441_ (
);

FILL FILL112040x57050 (
);

FILL FILL_1__14021_ (
);

FILL FILL_0__13854_ (
);

FILL FILL_0__13434_ (
);

FILL FILL_3__16299_ (
);

FILL FILL_0__13014_ (
);

FILL FILL_5__9891_ (
);

FILL FILL_5__9471_ (
);

NAND3X1 _16191_ (
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .B(_5477_),
    .C(_5531__bF$buf4),
    .Y(_6643_)
);

FILL FILL_5__16206_ (
);

FILL FILL_3__6917_ (
);

FILL FILL_1__9883_ (
);

FILL FILL_5__11761_ (
);

FILL FILL_1__9463_ (
);

FILL FILL_5__11341_ (
);

FILL FILL112440x26050 (
);

FILL FILL_1__9043_ (
);

FILL FILL_4__15619_ (
);

FILL FILL_2__16233_ (
);

FILL FILL_3__9389_ (
);

FILL FILL_4__10754_ (
);

FILL FILL_1__15646_ (
);

FILL FILL_1__15226_ (
);

FILL FILL_1__10781_ (
);

FILL FILL_1__10361_ (
);

FILL FILL112040x12050 (
);

FILL FILL_0__14639_ (
);

NOR2X1 _14924_ (
    .A(_5402_),
    .B(_5405_),
    .Y(_5406_)
);

FILL FILL_0__14219_ (
);

INVX1 _14504_ (
    .A(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_4994_)
);

FILL FILL_5__12966_ (
);

FILL FILL_5__12126_ (
);

FILL FILL_3__13580_ (
);

BUFX2 _6846_ (
    .A(_1_[8]),
    .Y(memoryAddress[8])
);

FILL FILL_3__13160_ (
);

FILL FILL_4__8253_ (
);

FILL FILL_4__11959_ (
);

FILL FILL_2__12993_ (
);

FILL FILL_4__11539_ (
);

FILL FILL_2__12573_ (
);

FILL FILL_4__11119_ (
);

FILL FILL_2__12153_ (
);

FILL FILL_6__8599_ (
);

FILL FILL_1__11986_ (
);

FILL FILL_1__11566_ (
);

FILL FILL_1__11146_ (
);

INVX1 _15709_ (
    .A(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_6173_)
);

FILL FILL_4__12900_ (
);

FILL FILL_0__8993_ (
);

FILL FILL_0__10979_ (
);

FILL FILL_0__8573_ (
);

FILL FILL_0__10559_ (
);

DFFSR _10844_ (
    .Q(\datapath_1.regfile_1.regOut[31] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_1953_[6])
);

INVX1 _10424_ (
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_1801_)
);

FILL FILL_0__10139_ (
);

INVX1 _10004_ (
    .A(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_1582_)
);

FILL FILL_4__15792_ (
);

FILL FILL_4__15372_ (
);

FILL FILL_2__9532_ (
);

FILL FILL_0__11920_ (
);

FILL FILL_3__14785_ (
);

FILL FILL_2__9112_ (
);

FILL FILL_3__14365_ (
);

FILL FILL_0__11500_ (
);

FILL FILL_4__9878_ (
);

FILL FILL_4__9038_ (
);

FILL FILL_2__13778_ (
);

FILL FILL_2__13358_ (
);

FILL FILL_0__14392_ (
);

FILL SFILL23720x42050 (
);

FILL FILL_0__9778_ (
);

FILL FILL_3__7875_ (
);

FILL FILL_0__9358_ (
);

FILL FILL_3__7455_ (
);

INVX1 _11629_ (
    .A(_2733_),
    .Y(\datapath_1.ALUResult [17])
);

FILL FILL_3__7035_ (
);

NOR2X1 _11209_ (
    .A(\datapath_1.alu_1.ALUInB [28]),
    .B(_2327_),
    .Y(_2328_)
);

FILL FILL_1__13712_ (
);

FILL FILL_4__16157_ (
);

FILL FILL_4__11292_ (
);

FILL FILL_0__12705_ (
);

FILL FILL_1__16184_ (
);

FILL FILL_5__8742_ (
);

FILL FILL_5__8322_ (
);

FILL FILL_3__10285_ (
);

NOR2X1 _15882_ (
    .A(_6341_),
    .B(_6339_),
    .Y(_6342_)
);

FILL FILL_0__15597_ (
);

FILL FILL_0__15177_ (
);

NOR3X1 _15462_ (
    .A(_5928_),
    .B(_5930_),
    .C(_5931_),
    .Y(_5932_)
);

NOR3X1 _15042_ (
    .A(_5515__bF$buf1),
    .B(_3928_),
    .C(_5521__bF$buf0),
    .Y(_5522_)
);

FILL FILL_1__8734_ (
);

FILL FILL_1__8314_ (
);

FILL SFILL8680x48050 (
);

FILL FILL_2__15924_ (
);

FILL SFILL44120x76050 (
);

FILL FILL_2__15504_ (
);

FILL FILL_5__13084_ (
);

FILL FILL_1__14917_ (
);

DFFSR _7384_ (
    .Q(\datapath_1.regfile_1.regOut[4] [2]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_198_[2])
);

FILL FILL_4__12497_ (
);

FILL FILL_4__12077_ (
);

FILL FILL_3__9601_ (
);

FILL SFILL84280x29050 (
);

FILL FILL_5__9527_ (
);

FILL FILL_5__9107_ (
);

OAI22X1 _16247_ (
    .A(_5400_),
    .B(_5544__bF$buf1),
    .C(_5485__bF$buf0),
    .D(_6696_),
    .Y(_6697_)
);

OAI21X1 _11382_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(_2149_),
    .C(_2498_),
    .Y(_2499_)
);

FILL FILL_0__11097_ (
);

FILL FILL_1__9939_ (
);

FILL FILL_5__11817_ (
);

FILL FILL_1__9519_ (
);

FILL FILL_3__12851_ (
);

FILL SFILL8600x46050 (
);

FILL FILL_3__12431_ (
);

FILL FILL_6__15296_ (
);

FILL FILL_3__12011_ (
);

FILL FILL_4__7944_ (
);

FILL FILL_4__7104_ (
);

FILL FILL_2__11844_ (
);

FILL SFILL13720x40050 (
);

FILL FILL_5__14289_ (
);

FILL FILL_2__11424_ (
);

FILL FILL_2__11004_ (
);

OAI21X1 _8589_ (
    .A(_861_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .C(_862_),
    .Y(_848_[7])
);

FILL SFILL27960x12050 (
);

DFFSR _8169_ (
    .Q(\datapath_1.regfile_1.regOut[10] [19]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_588_[19])
);

FILL FILL_1__10837_ (
);

FILL FILL_1__10417_ (
);

FILL SFILL84200x27050 (
);

FILL FILL_5__15650_ (
);

FILL FILL_0__7844_ (
);

FILL FILL_5__15230_ (
);

FILL FILL_0__7424_ (
);

DFFSR _9950_ (
    .Q(\datapath_1.regfile_1.regOut[24] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_1498_[8])
);

OAI21X1 _9530_ (
    .A(_1346_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1347_),
    .Y(_1303_[22])
);

OAI21X1 _9110_ (
    .A(_1127_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1128_),
    .Y(_1108_[10])
);

FILL FILL_4__14643_ (
);

FILL FILL_4__14223_ (
);

FILL SFILL13640x47050 (
);

OAI21X1 _12587_ (
    .A(_3436_),
    .B(vdd),
    .C(_3437_),
    .Y(_3425_[6])
);

NAND2X1 _12167_ (
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [17]),
    .Y(_3165_)
);

FILL FILL_3__13636_ (
);

FILL SFILL109480x27050 (
);

FILL FILL_3__13216_ (
);

FILL FILL_1__14670_ (
);

FILL FILL_1__14250_ (
);

FILL FILL_0_BUFX2_insert300 (
);

FILL FILL_4__8729_ (
);

FILL FILL_0_BUFX2_insert301 (
);

FILL FILL_0_BUFX2_insert302 (
);

FILL FILL_0_BUFX2_insert303 (
);

FILL FILL_2__12629_ (
);

FILL SFILL19320x68050 (
);

FILL FILL_0__13663_ (
);

FILL FILL_0_BUFX2_insert304 (
);

FILL FILL_2__12209_ (
);

FILL FILL_0__13243_ (
);

FILL FILL_0_BUFX2_insert305 (
);

FILL FILL_0_BUFX2_insert306 (
);

FILL FILL_0_BUFX2_insert307 (
);

FILL FILL_0_BUFX2_insert308 (
);

FILL FILL_5__9280_ (
);

FILL FILL_0_BUFX2_insert309 (
);

FILL FILL_0__8629_ (
);

FILL FILL_5__16015_ (
);

FILL FILL_0__8209_ (
);

FILL FILL_5__11990_ (
);

FILL FILL_5__11570_ (
);

FILL SFILL74280x27050 (
);

FILL FILL_1__9272_ (
);

FILL FILL_5__11150_ (
);

FILL FILL_4__15848_ (
);

FILL FILL_4__15428_ (
);

FILL FILL_4__15008_ (
);

FILL FILL_2__16042_ (
);

FILL FILL_4__10983_ (
);

FILL FILL_4__10563_ (
);

FILL FILL_4__10143_ (
);

FILL FILL112200x83050 (
);

FILL FILL_1__15875_ (
);

FILL FILL_1__15455_ (
);

FILL FILL_1__15035_ (
);

FILL FILL_1__10170_ (
);

FILL SFILL74600x39050 (
);

FILL FILL_0__14868_ (
);

OAI22X1 _14733_ (
    .A(_5217_),
    .B(_3893__bF$buf1),
    .C(_3944__bF$buf3),
    .D(_5218_),
    .Y(_5219_)
);

FILL FILL_0__14448_ (
);

FILL FILL_0__14028_ (
);

AOI22X1 _14313_ (
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .B(_4154_),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_4807_)
);

FILL FILL_2__7195_ (
);

FILL FILL_6__13362_ (
);

FILL SFILL43800x34050 (
);

FILL FILL_5__12775_ (
);

FILL FILL_5__12355_ (
);

FILL FILL_4__8482_ (
);

FILL FILL_4__11768_ (
);

FILL FILL_4__8062_ (
);

FILL FILL_4__11348_ (
);

FILL FILL_2__12382_ (
);

FILL FILL_1__11795_ (
);

FILL FILL_1__11375_ (
);

FILL SFILL99480x31050 (
);

AOI21X1 _15938_ (
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .B(_5606_),
    .C(_6395_),
    .Y(_6396_)
);

NOR2X1 _15518_ (
    .A(_5983_),
    .B(_5986_),
    .Y(_5987_)
);

FILL FILL_0__10788_ (
);

FILL FILL_0__8382_ (
);

FILL FILL_0__10368_ (
);

INVX1 _10653_ (
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_1913_)
);

INVX1 _10233_ (
    .A(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_1694_)
);

FILL FILL_3__11702_ (
);

FILL FILL_4__15181_ (
);

FILL SFILL33800x77050 (
);

FILL FILL_2__9761_ (
);

FILL SFILL64200x68050 (
);

FILL FILL_3__14594_ (
);

FILL FILL_2__9341_ (
);

FILL FILL_3__14174_ (
);

FILL FILL_4_BUFX2_insert880 (
);

FILL FILL_4_BUFX2_insert881 (
);

FILL FILL_4_BUFX2_insert882 (
);

FILL FILL_4__9267_ (
);

FILL FILL_4_BUFX2_insert883 (
);

FILL FILL_2__13587_ (
);

FILL FILL_4_BUFX2_insert884 (
);

FILL FILL_2__13167_ (
);

FILL FILL_4_BUFX2_insert885 (
);

FILL FILL_4_BUFX2_insert886 (
);

FILL FILL_4_BUFX2_insert887 (
);

FILL FILL_5__14921_ (
);

FILL FILL_5__14501_ (
);

FILL FILL_4_BUFX2_insert888 (
);

FILL FILL_4_BUFX2_insert889 (
);

DFFSR _8801_ (
    .Q(\datapath_1.regfile_1.regOut[15] [11]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_913_[11])
);

FILL SFILL68520x76050 (
);

FILL FILL_4__13914_ (
);

FILL FILL_3__7684_ (
);

FILL FILL_0__9167_ (
);

NOR3X1 _11858_ (
    .A(_2942_),
    .B(\datapath_1.ALUResult [25]),
    .C(_2944_),
    .Y(_2945_)
);

AOI21X1 _11438_ (
    .A(_2551_),
    .B(_2427_),
    .C(_2553_),
    .Y(_2554_)
);

NOR2X1 _11018_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2137_)
);

FILL FILL_3__12907_ (
);

FILL FILL_1__13941_ (
);

FILL FILL_4__16386_ (
);

FILL FILL_1__13521_ (
);

FILL FILL_1__13101_ (
);

FILL FILL_6__10067_ (
);

FILL FILL_3__15799_ (
);

FILL FILL_3__15379_ (
);

FILL FILL_0__12514_ (
);

FILL FILL_5__8971_ (
);

FILL SFILL33800x32050 (
);

FILL SFILL64200x23050 (
);

FILL FILL_5__8131_ (
);

AOI21X1 _15691_ (
    .A(_6155_),
    .B(_6133_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [15])
);

OAI22X1 _15271_ (
    .A(_4227_),
    .B(_5503__bF$buf1),
    .C(_5504__bF$buf0),
    .D(_5745_),
    .Y(_5746_)
);

FILL FILL_5__15706_ (
);

FILL FILL_3__16320_ (
);

FILL FILL_1__8963_ (
);

FILL FILL_5__10421_ (
);

FILL FILL_1__8123_ (
);

FILL FILL_5__10001_ (
);

FILL FILL_2__15733_ (
);

FILL FILL_2__15313_ (
);

FILL FILL_3__8889_ (
);

FILL FILL_3__8469_ (
);

FILL FILL_6__6894_ (
);

FILL FILL_1__14726_ (
);

OAI21X1 _7193_ (
    .A(_154_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_155_),
    .Y(_133_[11])
);

FILL FILL_1__14306_ (
);

FILL FILL_0__13719_ (
);

FILL FILL_3__9410_ (
);

FILL FILL_2__6886_ (
);

FILL FILL_5__9756_ (
);

FILL FILL_5__9336_ (
);

FILL FILL_3__11299_ (
);

FILL FILL_6__12213_ (
);

OAI22X1 _16056_ (
    .A(_5530__bF$buf1),
    .B(_6510_),
    .C(_5532__bF$buf2),
    .D(_6509_),
    .Y(_6511_)
);

NOR2X1 _11191_ (
    .A(_2309_),
    .B(_2293_),
    .Y(_2310_)
);

FILL FILL_5__11626_ (
);

FILL FILL_1__9748_ (
);

FILL FILL_3__12660_ (
);

FILL FILL_5__11206_ (
);

FILL FILL_3__12240_ (
);

FILL FILL_4__7753_ (
);

FILL FILL_4__7333_ (
);

FILL FILL_4__10619_ (
);

FILL FILL_2__11653_ (
);

FILL FILL_2__11233_ (
);

FILL FILL_5__14098_ (
);

FILL FILL_6__7679_ (
);

NAND2X1 _8398_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_776_)
);

FILL FILL_1__10646_ (
);

FILL FILL_0__7233_ (
);

FILL FILL_6__13838_ (
);

FILL FILL_4__14872_ (
);

FILL FILL_6__13418_ (
);

FILL FILL_4__14452_ (
);

FILL FILL_4__14032_ (
);

OAI21X1 _12396_ (
    .A(_3328_),
    .B(MemToReg_bF$buf4),
    .C(_3329_),
    .Y(\datapath_1.mux_wd3.dout [17])
);

FILL FILL_3__13865_ (
);

FILL FILL_2__8612_ (
);

FILL FILL_3__13445_ (
);

FILL FILL_3__13025_ (
);

FILL FILL_4__8958_ (
);

FILL FILL_4__8118_ (
);

FILL FILL_2__12858_ (
);

FILL FILL_2__12438_ (
);

FILL FILL_0__13892_ (
);

FILL FILL_2__12018_ (
);

FILL FILL_0__13472_ (
);

FILL SFILL23720x37050 (
);

FILL FILL_5__16244_ (
);

FILL FILL_0__8858_ (
);

FILL FILL_3__6955_ (
);

FILL FILL_0__8438_ (
);

FILL FILL_6__9405_ (
);

OAI21X1 _10709_ (
    .A(_1949_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .C(_1950_),
    .Y(_1888_[31])
);

FILL FILL_0__8018_ (
);

FILL FILL_1__9081_ (
);

FILL FILL_4__15657_ (
);

FILL FILL_4__15237_ (
);

FILL FILL_2__16271_ (
);

FILL FILL_4__10792_ (
);

FILL FILL_4__10372_ (
);

FILL SFILL109640x53050 (
);

FILL FILL_1__15684_ (
);

FILL FILL_1__15264_ (
);

FILL SFILL59800x5050 (
);

FILL FILL_5__7822_ (
);

OAI22X1 _14962_ (
    .A(_5441_),
    .B(_3905__bF$buf0),
    .C(_3977__bF$buf4),
    .D(_5442_),
    .Y(_5443_)
);

FILL FILL_0__14677_ (
);

FILL FILL_0__14257_ (
);

OAI22X1 _14542_ (
    .A(_5030_),
    .B(_3982__bF$buf1),
    .C(_3978_),
    .D(_5031_),
    .Y(_5032_)
);

AOI21X1 _14122_ (
    .A(_4620_),
    .B(_4595_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [13])
);

FILL FILL_1__7814_ (
);

FILL FILL_6__13171_ (
);

FILL SFILL99640x2050 (
);

FILL FILL_5__12584_ (
);

FILL FILL_5__12164_ (
);

BUFX2 _6884_ (
    .A(_2_[14]),
    .Y(memoryWriteData[14])
);

FILL FILL_4__11997_ (
);

FILL FILL_4__11577_ (
);

FILL FILL_4__11157_ (
);

FILL SFILL48920x41050 (
);

FILL FILL_2__12191_ (
);

FILL FILL_1__16049_ (
);

FILL SFILL99240x1050 (
);

FILL FILL_5__8607_ (
);

FILL FILL_1__11184_ (
);

INVX1 _15747_ (
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_6210_)
);

INVX1 _15327_ (
    .A(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_5801_)
);

FILL FILL_0__8191_ (
);

NOR2X1 _10882_ (
    .A(_2023_),
    .B(_2029_),
    .Y(ALUControl[0])
);

DFFSR _10462_ (
    .Q(\datapath_1.regfile_1.regOut[28] [8]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_1758_[8])
);

FILL FILL_0__10177_ (
);

OAI21X1 _10042_ (
    .A(_1606_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1607_),
    .Y(_1563_[22])
);

FILL FILL_3__11931_ (
);

FILL FILL_3__11511_ (
);

FILL FILL_0__16403_ (
);

FILL SFILL13720x35050 (
);

FILL FILL_2__10924_ (
);

FILL FILL_5__13789_ (
);

FILL FILL_2__9990_ (
);

FILL FILL_5__13369_ (
);

FILL FILL_2__10504_ (
);

FILL SFILL88600x23050 (
);

FILL FILL_2__9150_ (
);

DFFSR _7669_ (
    .Q(\datapath_1.regfile_1.regOut[6] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_328_[31])
);

FILL SFILL109560x15050 (
);

NAND2X1 _7249_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_193_)
);

FILL FILL_4__9496_ (
);

FILL SFILL109400x4050 (
);

FILL FILL_2__13396_ (
);

FILL FILL_5__14730_ (
);

FILL FILL_0__6924_ (
);

FILL FILL_5__14310_ (
);

OAI21X1 _8610_ (
    .A(_875_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_876_),
    .Y(_848_[14])
);

FILL FILL_1__12389_ (
);

FILL FILL_4__13723_ (
);

FILL FILL_4__13303_ (
);

FILL FILL_3__7493_ (
);

FILL FILL_0__9396_ (
);

FILL FILL_3__7073_ (
);

OAI21X1 _11667_ (
    .A(_2752_),
    .B(_2344__bF$buf1),
    .C(_2768_),
    .Y(_2769_)
);

NAND2X1 _11247_ (
    .A(_2364_),
    .B(_2365_),
    .Y(_2366_)
);

FILL FILL_3__12716_ (
);

FILL FILL_1__13750_ (
);

FILL FILL_1__13330_ (
);

FILL FILL_4__16195_ (
);

FILL FILL_4__7809_ (
);

FILL FILL_2__11709_ (
);

FILL FILL_0__12743_ (
);

FILL FILL_3__15188_ (
);

FILL FILL_0__12323_ (
);

FILL FILL_5__8780_ (
);

FILL FILL_5__8360_ (
);

FILL SFILL28920x50 (
);

FILL SFILL3560x83050 (
);

FILL FILL_5__15935_ (
);

AOI22X1 _15080_ (
    .A(_5557_),
    .B(\datapath_1.regfile_1.regOut[17] [1]),
    .C(\datapath_1.regfile_1.regOut[18] [1]),
    .D(_5558_),
    .Y(_5559_)
);

FILL FILL_5__15515_ (
);

FILL FILL_0__7709_ (
);

DFFSR _9815_ (
    .Q(\datapath_1.regfile_1.regOut[23] [1]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_1433_[1])
);

FILL FILL_1__8772_ (
);

FILL FILL_5__10650_ (
);

FILL FILL_1__8352_ (
);

FILL FILL_5__10230_ (
);

FILL FILL_4__14928_ (
);

FILL FILL_4__14508_ (
);

FILL FILL_2__15962_ (
);

FILL FILL_2__15542_ (
);

FILL FILL_2__15122_ (
);

FILL FILL_3__8698_ (
);

FILL FILL112200x78050 (
);

FILL FILL_1__14955_ (
);

FILL FILL_1__14535_ (
);

FILL FILL_1__14115_ (
);

FILL FILL_0__13948_ (
);

OAI22X1 _13813_ (
    .A(_4316_),
    .B(_3936__bF$buf0),
    .C(_3935__bF$buf4),
    .D(_4317_),
    .Y(_4318_)
);

FILL FILL_0__13528_ (
);

FILL FILL_0__13108_ (
);

FILL SFILL38840x46050 (
);

FILL FILL_5__9985_ (
);

FILL FILL_5__9145_ (
);

FILL FILL_6__12862_ (
);

AOI22X1 _16285_ (
    .A(_5490_),
    .B(\datapath_1.regfile_1.regOut[7] [31]),
    .C(\datapath_1.regfile_1.regOut[10] [31]),
    .D(_6314_),
    .Y(_6734_)
);

FILL SFILL28920x82050 (
);

FILL FILL_5__11855_ (
);

FILL FILL_1__9977_ (
);

FILL FILL_1__9557_ (
);

FILL FILL_5__11435_ (
);

FILL FILL_1__9137_ (
);

FILL FILL_5__11015_ (
);

FILL FILL_4__7982_ (
);

FILL FILL_2__16327_ (
);

FILL FILL_4__7562_ (
);

FILL FILL_4__10428_ (
);

FILL FILL_2__11882_ (
);

FILL FILL_4__10008_ (
);

FILL FILL_2__11462_ (
);

FILL FILL_2__11042_ (
);

FILL FILL112200x33050 (
);

FILL FILL_1__10875_ (
);

FILL SFILL99480x26050 (
);

FILL FILL_1__10035_ (
);

FILL FILL_0__7882_ (
);

FILL FILL_0__7462_ (
);

FILL SFILL3480x45050 (
);

FILL FILL_0__7042_ (
);

FILL SFILL24120x67050 (
);

FILL FILL_4__14681_ (
);

FILL FILL_4__14261_ (
);

FILL FILL_2__8841_ (
);

FILL FILL_3__13674_ (
);

FILL FILL_3__13254_ (
);

FILL FILL_2__8001_ (
);

FILL FILL_4__8767_ (
);

FILL FILL_4__8347_ (
);

FILL FILL_2__12247_ (
);

FILL FILL_0__13281_ (
);

FILL FILL_5__16053_ (
);

NOR2X1 _10938_ (
    .A(_2054_),
    .B(_2057_),
    .Y(_2072_)
);

FILL FILL_0__8247_ (
);

FILL FILL_6__9214_ (
);

OAI21X1 _10518_ (
    .A(_1842_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .C(_1843_),
    .Y(_1823_[10])
);

FILL FILL_4__15886_ (
);

FILL FILL_1__12601_ (
);

FILL FILL_4__15466_ (
);

FILL FILL_4__15046_ (
);

FILL FILL_2__16080_ (
);

FILL FILL_4__10181_ (
);

FILL FILL_3__14879_ (
);

FILL FILL_2__9626_ (
);

FILL FILL_3__14459_ (
);

FILL FILL_2__9206_ (
);

FILL FILL_3__14039_ (
);

FILL FILL_1__15493_ (
);

FILL FILL_1__15073_ (
);

FILL SFILL33800x27050 (
);

FILL SFILL64200x18050 (
);

FILL FILL_5__7631_ (
);

FILL FILL_5__7211_ (
);

FILL FILL_0__14486_ (
);

OAI22X1 _14771_ (
    .A(_5254_),
    .B(_3884__bF$buf2),
    .C(_3924__bF$buf2),
    .D(_5255_),
    .Y(_5256_)
);

FILL FILL_0__14066_ (
);

OAI22X1 _14351_ (
    .A(_4844_),
    .B(_3941_),
    .C(_3967__bF$buf2),
    .D(_4843_),
    .Y(_4845_)
);

FILL FILL_3__15820_ (
);

FILL FILL_3__15400_ (
);

FILL FILL_1__7623_ (
);

FILL FILL_1__7203_ (
);

FILL FILL_2__14813_ (
);

FILL FILL_3__7969_ (
);

FILL FILL_3__7549_ (
);

FILL FILL_5__12393_ (
);

FILL FILL_1__13806_ (
);

FILL FILL_4__11386_ (
);

FILL FILL_3__8910_ (
);

FILL FILL_1__16278_ (
);

FILL FILL_5__8836_ (
);

FILL FILL_3__10799_ (
);

FILL FILL_3__10379_ (
);

NAND3X1 _15976_ (
    .A(_6426_),
    .B(_6427_),
    .C(_6432_),
    .Y(_6433_)
);

FILL SFILL18680x50 (
);

NAND3X1 _15556_ (
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf0),
    .Y(_6024_)
);

NAND3X1 _15136_ (
    .A(_5607_),
    .B(_5608_),
    .C(_5613_),
    .Y(_5614_)
);

FILL SFILL113560x15050 (
);

OAI21X1 _10691_ (
    .A(_1937_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .C(_1938_),
    .Y(_1888_[25])
);

OAI21X1 _10271_ (
    .A(_1718_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .C(_1719_),
    .Y(_1693_[13])
);

FILL FILL_5__10706_ (
);

FILL FILL_1__8828_ (
);

FILL FILL_3__11740_ (
);

FILL FILL_3__11320_ (
);

FILL FILL_0__16212_ (
);

FILL FILL_5__13598_ (
);

FILL FILL_2__10313_ (
);

DFFSR _7898_ (
    .Q(\datapath_1.regfile_1.regOut[8] [4]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_458_[4])
);

NAND2X1 _7478_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_305_)
);

NAND2X1 _7058_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_86_)
);

FILL SFILL18840x42050 (
);

FILL FILL_1__12198_ (
);

FILL FILL_6__12918_ (
);

FILL FILL_4__13952_ (
);

FILL FILL_4__13532_ (
);

FILL FILL_4__13112_ (
);

INVX1 _11896_ (
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_2972_)
);

AOI21X1 _11476_ (
    .A(_2446_),
    .B(_2590_),
    .C(_2289_),
    .Y(_2591_)
);

NOR2X1 _11056_ (
    .A(_2167_),
    .B(_2174_),
    .Y(_2175_)
);

FILL FILL_3__12525_ (
);

FILL FILL_3__12105_ (
);

FILL FILL_4__7618_ (
);

FILL FILL_2__11938_ (
);

FILL FILL_0__12972_ (
);

FILL FILL_2__11518_ (
);

FILL FILL_0__12132_ (
);

FILL SFILL38920x2050 (
);

FILL FILL_5__15744_ (
);

FILL SFILL38840x7050 (
);

FILL FILL_0__7938_ (
);

FILL FILL_5__15324_ (
);

NAND2X1 _9624_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1390_)
);

DFFSR _9204_ (
    .Q(\datapath_1.regfile_1.regOut[18] [30]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_1108_[30])
);

FILL FILL_1__8581_ (
);

FILL FILL_4__14737_ (
);

FILL FILL_4__14317_ (
);

FILL FILL_2__15771_ (
);

FILL FILL_2__15351_ (
);

FILL SFILL110200x82050 (
);

FILL FILL_3__8087_ (
);

FILL FILL_1__14764_ (
);

FILL FILL_1__14344_ (
);

FILL FILL_5__6902_ (
);

FILL FILL_0__13757_ (
);

FILL FILL_0__13337_ (
);

NAND3X1 _13622_ (
    .A(_4128_),
    .B(_4130_),
    .C(_4127_),
    .Y(_4131_)
);

DFFSR _13202_ (
    .Q(\datapath_1.mux_iord.din0 [27]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[27])
);

FILL FILL_5__9794_ (
);

FILL FILL_5__9374_ (
);

AOI22X1 _16094_ (
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .B(_5785_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_6548_)
);

FILL FILL_5__16109_ (
);

FILL FILL_1__9786_ (
);

FILL FILL_5__11664_ (
);

FILL FILL_5__11244_ (
);

FILL FILL_1__9366_ (
);

FILL SFILL69080x51050 (
);

FILL FILL_2__16136_ (
);

FILL FILL_4__7371_ (
);

FILL FILL_4__10657_ (
);

FILL SFILL48920x36050 (
);

FILL FILL_4__10237_ (
);

FILL FILL_2__11691_ (
);

FILL FILL_2__11271_ (
);

FILL FILL_1__15969_ (
);

FILL FILL_1__15549_ (
);

FILL FILL_1__15129_ (
);

FILL FILL_1__10684_ (
);

FILL FILL_1__10264_ (
);

OAI22X1 _14827_ (
    .A(_3890_),
    .B(_5310_),
    .C(_5309_),
    .D(_3931__bF$buf0),
    .Y(_5311_)
);

OAI22X1 _14407_ (
    .A(_4898_),
    .B(_3936__bF$buf1),
    .C(_3905__bF$buf0),
    .D(_4897_),
    .Y(_4899_)
);

FILL FILL_0__7691_ (
);

FILL FILL_2__7289_ (
);

FILL FILL_4__14490_ (
);

FILL FILL_4__14070_ (
);

FILL FILL_0__15903_ (
);

FILL FILL_5__12869_ (
);

FILL FILL_2__8650_ (
);

FILL FILL_5__12449_ (
);

FILL FILL_2__8230_ (
);

FILL FILL_5__12029_ (
);

FILL FILL_3__13483_ (
);

FILL FILL_4__8996_ (
);

FILL FILL_4__8576_ (
);

FILL FILL_2__12896_ (
);

FILL FILL_2__12476_ (
);

FILL FILL_2__12056_ (
);

FILL SFILL34200x57050 (
);

FILL FILL_0__13090_ (
);

FILL FILL_5__13810_ (
);

FILL FILL_1__11889_ (
);

FILL FILL_1__11469_ (
);

FILL FILL_1__11049_ (
);

FILL SFILL3640x71050 (
);

FILL FILL_0__8896_ (
);

FILL FILL_3__6993_ (
);

FILL FILL_5__16282_ (
);

FILL FILL_0__8476_ (
);

FILL FILL_0__8056_ (
);

OAI21X1 _10747_ (
    .A(_1954_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .C(_1955_),
    .Y(_1953_[1])
);

DFFSR _10327_ (
    .Q(\datapath_1.regfile_1.regOut[27] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_1693_[1])
);

FILL FILL_4__15695_ (
);

FILL FILL_1__12830_ (
);

FILL FILL_1__12410_ (
);

FILL FILL_4__15275_ (
);

FILL FILL_2__9855_ (
);

FILL FILL_0__11823_ (
);

FILL FILL_3__14688_ (
);

FILL FILL_2__9015_ (
);

FILL FILL_3__14268_ (
);

FILL FILL_0__11403_ (
);

FILL FILL_5__7860_ (
);

FILL FILL_5__7440_ (
);

NAND3X1 _14580_ (
    .A(_5060_),
    .B(_5061_),
    .C(_5068_),
    .Y(_5069_)
);

FILL FILL_0__14295_ (
);

OAI22X1 _14160_ (
    .A(_4656_),
    .B(_3930__bF$buf1),
    .C(_3971__bF$buf1),
    .D(_4657_),
    .Y(_4658_)
);

FILL SFILL38920x34050 (
);

FILL FILL_1__7852_ (
);

FILL FILL_1__7432_ (
);

FILL FILL_2__14622_ (
);

FILL FILL_2__14202_ (
);

FILL FILL_3__7358_ (
);

FILL FILL_1__13615_ (
);

FILL FILL_4__11195_ (
);

FILL FILL_1_BUFX2_insert230 (
);

FILL FILL_1_BUFX2_insert231 (
);

FILL FILL_0__12608_ (
);

FILL FILL_1_BUFX2_insert232 (
);

FILL FILL_1_BUFX2_insert233 (
);

FILL FILL_1__16087_ (
);

FILL FILL_1_BUFX2_insert234 (
);

FILL FILL_1_BUFX2_insert235 (
);

FILL FILL_5__8645_ (
);

FILL FILL_1_BUFX2_insert236 (
);

FILL FILL_3__10188_ (
);

FILL FILL_5__8225_ (
);

FILL FILL_1_BUFX2_insert237 (
);

FILL FILL_6_BUFX2_insert792 (
);

FILL FILL_1_BUFX2_insert238 (
);

FILL FILL_6__11942_ (
);

FILL FILL_1_BUFX2_insert239 (
);

NAND3X1 _15785_ (
    .A(_6240_),
    .B(_6241_),
    .C(_6246_),
    .Y(_6247_)
);

INVX1 _15365_ (
    .A(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_5838_)
);

FILL FILL_6_BUFX2_insert797 (
);

FILL FILL_3__16414_ (
);

FILL SFILL28920x77050 (
);

FILL SFILL3560x33050 (
);

FILL FILL_5__10935_ (
);

DFFSR _10080_ (
    .Q(\datapath_1.regfile_1.regOut[25] [10]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_1563_[10])
);

FILL FILL_1__8637_ (
);

FILL FILL_5__10515_ (
);

FILL FILL_1__8217_ (
);

FILL FILL_2__15827_ (
);

FILL SFILL104440x50050 (
);

FILL FILL_2__15407_ (
);

FILL FILL_0__16021_ (
);

FILL FILL_2__10962_ (
);

FILL FILL_2__10542_ (
);

FILL FILL_2__10122_ (
);

NAND2X1 _7287_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .Y(_262_)
);

FILL FILL112200x28050 (
);

FILL FILL_3__9924_ (
);

FILL FILL_3__9504_ (
);

FILL FILL_0__6962_ (
);

FILL FILL_6__12727_ (
);

FILL FILL_4__13761_ (
);

FILL FILL_4__13341_ (
);

INVX2 _11285_ (
    .A(_2403_),
    .Y(_2404_)
);

FILL FILL_2__7501_ (
);

FILL FILL_3__12754_ (
);

FILL FILL_6__15199_ (
);

FILL FILL_3__12334_ (
);

FILL SFILL28920x32050 (
);

FILL FILL_4__7847_ (
);

FILL FILL_4__7427_ (
);

FILL FILL_2__11747_ (
);

FILL SFILL89160x43050 (
);

FILL FILL_0__12781_ (
);

FILL FILL_2__11327_ (
);

FILL FILL_0__12361_ (
);

FILL FILL_6__16140_ (
);

FILL FILL_5__15973_ (
);

FILL FILL_5__15553_ (
);

FILL FILL_5__15133_ (
);

FILL FILL_0__7747_ (
);

FILL FILL_0__7327_ (
);

NAND2X1 _9853_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1502_)
);

DFFSR _9433_ (
    .Q(\datapath_1.regfile_1.regOut[20] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_1238_[3])
);

INVX1 _9013_ (
    .A(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_1084_)
);

FILL FILL_1__8390_ (
);

FILL SFILL28840x39050 (
);

FILL FILL_4__14966_ (
);

FILL FILL_4__14546_ (
);

FILL FILL_4__14126_ (
);

FILL FILL_2__15580_ (
);

FILL FILL_2__15160_ (
);

FILL FILL_2__8706_ (
);

FILL FILL_3__13959_ (
);

FILL FILL_1__14993_ (
);

FILL FILL_3__13539_ (
);

FILL FILL_1__14573_ (
);

FILL FILL_3__13119_ (
);

FILL FILL_1__14153_ (
);

FILL FILL_0__13986_ (
);

AOI21X1 _13851_ (
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .B(_3894_),
    .C(_4354_),
    .Y(_4355_)
);

FILL FILL_0__13566_ (
);

FILL FILL_0__13146_ (
);

INVX1 _13431_ (
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_3943_)
);

INVX1 _13011_ (
    .A(_2_[20]),
    .Y(_3659_)
);

FILL FILL_3__14900_ (
);

FILL FILL_6__12060_ (
);

FILL FILL_5__16338_ (
);

FILL FILL_5__11893_ (
);

FILL FILL_1__9595_ (
);

FILL FILL_5__11473_ (
);

FILL FILL_5__11053_ (
);

FILL FILL_2__16365_ (
);

FILL FILL_4__7180_ (
);

FILL FILL_4__10886_ (
);

FILL SFILL94360x61050 (
);

FILL FILL_4__10046_ (
);

FILL FILL_2__11080_ (
);

FILL FILL_1__15778_ (
);

FILL FILL_1__15358_ (
);

FILL FILL_1__10493_ (
);

OAI22X1 _14636_ (
    .A(_3972__bF$buf0),
    .B(_5123_),
    .C(_3944__bF$buf0),
    .D(_5122_),
    .Y(_5124_)
);

NOR2X1 _14216_ (
    .A(_4702_),
    .B(_4712_),
    .Y(_4713_)
);

FILL FILL_0__7080_ (
);

FILL FILL_2__7098_ (
);

FILL SFILL79160x41050 (
);

FILL FILL_3__10820_ (
);

FILL FILL_6__13265_ (
);

FILL FILL_3__10400_ (
);

FILL FILL_0__15712_ (
);

FILL SFILL103640x46050 (
);

FILL FILL_5__12258_ (
);

FILL FILL_3__13292_ (
);

NAND2X1 _6978_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_53_)
);

FILL FILL_4__8385_ (
);

FILL SFILL18680x2050 (
);

FILL SFILL18840x37050 (
);

FILL FILL_2__12285_ (
);

FILL FILL_1__11698_ (
);

FILL FILL_1__11278_ (
);

FILL FILL_4__12612_ (
);

FILL FILL_5__16091_ (
);

NAND2X1 _10976_ (
    .A(vdd),
    .B(\control_1.next [1]),
    .Y(_2102_)
);

NAND2X1 _10556_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1869_)
);

NAND2X1 _10136_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1650_)
);

FILL FILL_3__11605_ (
);

FILL FILL_4__15084_ (
);

FILL FILL_2__9664_ (
);

FILL FILL_3__14497_ (
);

FILL FILL_2__9244_ (
);

FILL FILL_0__11632_ (
);

FILL FILL_0__11212_ (
);

FILL FILL_3__14077_ (
);

FILL FILL_5__14824_ (
);

FILL FILL_5__14404_ (
);

NAND2X1 _8704_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_919_)
);

FILL FILL_1__7241_ (
);

FILL FILL_4__13817_ (
);

FILL FILL_2__14851_ (
);

FILL FILL_2__14431_ (
);

FILL FILL_3__7587_ (
);

FILL FILL_2__14011_ (
);

FILL FILL_3__7167_ (
);

FILL FILL_1__13844_ (
);

FILL FILL_1__13424_ (
);

FILL FILL_4__16289_ (
);

FILL FILL_1__13004_ (
);

FILL FILL_0__12837_ (
);

NAND2X1 _12702_ (
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[2]),
    .Y(_3494_)
);

FILL FILL_0__12417_ (
);

FILL FILL_5__8874_ (
);

FILL FILL_5__8454_ (
);

NAND3X1 _15594_ (
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf3),
    .Y(_6061_)
);

AOI22X1 _15174_ (
    .A(_5649_),
    .B(\datapath_1.regfile_1.regOut[23] [3]),
    .C(\datapath_1.regfile_1.regOut[22] [3]),
    .D(_5650_),
    .Y(_5651_)
);

FILL FILL_5__15609_ (
);

INVX1 _9909_ (
    .A(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_1539_)
);

FILL FILL_3__16223_ (
);

FILL FILL_1__8866_ (
);

FILL FILL_5__10744_ (
);

FILL FILL_5__10324_ (
);

FILL FILL_1__8446_ (
);

FILL SFILL69080x46050 (
);

FILL FILL_2__15636_ (
);

FILL FILL_2__15216_ (
);

FILL FILL_4__6871_ (
);

FILL FILL_0__16250_ (
);

FILL FILL_2__10771_ (
);

FILL FILL_1__14629_ (
);

FILL FILL_1__14209_ (
);

INVX1 _7096_ (
    .A(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_111_)
);

FILL FILL_3__9733_ (
);

NAND3X1 _13907_ (
    .A(_4401_),
    .B(_4402_),
    .C(_4409_),
    .Y(_4410_)
);

FILL SFILL74760x71050 (
);

FILL FILL_5__9659_ (
);

FILL FILL_5__9239_ (
);

FILL FILL_4__13990_ (
);

FILL FILL_6__12116_ (
);

NAND2X1 _16379_ (
    .A(gnd),
    .B(gnd),
    .Y(_6807_)
);

FILL FILL_4__13570_ (
);

FILL FILL_4__13150_ (
);

FILL FILL_5__11949_ (
);

NOR2X1 _11094_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(_2212_),
    .Y(_2213_)
);

FILL FILL_2__7730_ (
);

FILL FILL_3__12983_ (
);

FILL FILL_5__11529_ (
);

FILL FILL_2__7310_ (
);

FILL FILL_5__11109_ (
);

FILL FILL_3__12143_ (
);

FILL FILL_4__7236_ (
);

FILL FILL_2__11976_ (
);

FILL FILL_2__11556_ (
);

FILL FILL_0__12590_ (
);

FILL FILL_2__11136_ (
);

FILL FILL_0__12170_ (
);

FILL FILL_1__10969_ (
);

FILL FILL_1__10549_ (
);

FILL FILL_1__10129_ (
);

FILL FILL_5_CLKBUF1_insert1080 (
);

FILL SFILL3640x66050 (
);

FILL FILL_5_CLKBUF1_insert1081 (
);

FILL FILL_5__15782_ (
);

FILL FILL_0__7976_ (
);

FILL FILL_5__15362_ (
);

FILL FILL_5_CLKBUF1_insert1082 (
);

FILL FILL_5_CLKBUF1_insert1083 (
);

FILL FILL_0__7556_ (
);

INVX1 _9662_ (
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_1415_)
);

INVX1 _9242_ (
    .A(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_1196_)
);

FILL SFILL43880x73050 (
);

FILL FILL_1__11910_ (
);

FILL FILL_4__14775_ (
);

FILL FILL_4__14355_ (
);

NAND3X1 _12299_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3263_)
);

FILL FILL_0__10903_ (
);

FILL FILL_3__13768_ (
);

FILL FILL_2__8515_ (
);

FILL SFILL3560x4050 (
);

FILL FILL_3__13348_ (
);

FILL FILL_1__14382_ (
);

FILL FILL_5__6940_ (
);

FILL FILL_0__13795_ (
);

INVX1 _13660_ (
    .A(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_4168_)
);

FILL FILL_0__13375_ (
);

NAND2X1 _13240_ (
    .A(\datapath_1.a3 [4]),
    .B(_3777_),
    .Y(_3783_)
);

FILL SFILL38920x29050 (
);

FILL FILL_1__6932_ (
);

FILL FILL_4__9802_ (
);

FILL FILL_2__13702_ (
);

FILL FILL_3__6858_ (
);

FILL FILL_5__16147_ (
);

FILL SFILL3640x21050 (
);

FILL FILL_5__11282_ (
);

FILL FILL_2__16174_ (
);

FILL FILL_4__10695_ (
);

FILL FILL_4__10275_ (
);

FILL FILL_1__15587_ (
);

FILL FILL_1__15167_ (
);

FILL FILL_5__7725_ (
);

FILL FILL_5__7305_ (
);

FILL SFILL59000x42050 (
);

OAI22X1 _14865_ (
    .A(_5346_),
    .B(_3910_),
    .C(_3977__bF$buf3),
    .D(_5347_),
    .Y(_5348_)
);

NOR2X1 _14445_ (
    .A(_4933_),
    .B(_4936_),
    .Y(_4937_)
);

INVX1 _14025_ (
    .A(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_4525_)
);

FILL FILL_3__15914_ (
);

FILL SFILL3560x28050 (
);

FILL FILL_1__7717_ (
);

FILL SFILL104440x45050 (
);

FILL FILL_2__14907_ (
);

FILL FILL_0__15941_ (
);

FILL FILL_0__15521_ (
);

FILL FILL_0__15101_ (
);

FILL FILL_5__12487_ (
);

FILL FILL_5__12067_ (
);

FILL FILL_4__8194_ (
);

FILL SFILL33880x71050 (
);

FILL FILL_2__12094_ (
);

FILL FILL_1__11087_ (
);

FILL FILL_4__12841_ (
);

FILL FILL_4__12421_ (
);

FILL FILL_4__12001_ (
);

NAND2X1 _10785_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1981_)
);

FILL FILL_0__8094_ (
);

FILL SFILL49080x42050 (
);

NAND2X1 _10365_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1762_)
);

FILL FILL_3__11834_ (
);

FILL FILL_3__11414_ (
);

FILL SFILL28920x27050 (
);

FILL FILL_4__6927_ (
);

FILL FILL_0__16306_ (
);

FILL FILL_2__9893_ (
);

FILL FILL_2__10827_ (
);

FILL FILL_2__9473_ (
);

FILL FILL_2__10407_ (
);

FILL FILL_0__11861_ (
);

FILL FILL_0__11441_ (
);

FILL FILL_0__11021_ (
);

FILL FILL_4__9399_ (
);

FILL FILL_2__13299_ (
);

FILL FILL_5__14633_ (
);

FILL FILL_5__14213_ (
);

DFFSR _8933_ (
    .Q(\datapath_1.regfile_1.regOut[16] [15]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_978_[15])
);

INVX1 _8513_ (
    .A(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_832_)
);

FILL FILL_1__7890_ (
);

FILL FILL_1__7470_ (
);

FILL FILL_1__7050_ (
);

FILL FILL_4__13626_ (
);

FILL FILL_2__14660_ (
);

FILL FILL_2__14240_ (
);

FILL FILL_0__9299_ (
);

FILL FILL_3__12619_ (
);

FILL FILL_3_BUFX2_insert50 (
);

FILL FILL_1__13653_ (
);

FILL FILL_3_BUFX2_insert51 (
);

FILL FILL_1__13233_ (
);

FILL FILL_4__16098_ (
);

FILL FILL_3_BUFX2_insert52 (
);

FILL FILL_3_BUFX2_insert53 (
);

FILL FILL_3_BUFX2_insert54 (
);

FILL FILL_3_BUFX2_insert55 (
);

FILL FILL_1_BUFX2_insert610 (
);

FILL FILL_3_BUFX2_insert56 (
);

FILL FILL_3_BUFX2_insert57 (
);

FILL FILL_1_BUFX2_insert611 (
);

FILL FILL_0__12646_ (
);

FILL FILL_1_BUFX2_insert612 (
);

DFFSR _12931_ (
    .Q(\datapath_1.a [12]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3555_[12])
);

FILL FILL_3_BUFX2_insert58 (
);

INVX1 _12511_ (
    .A(ALUOut[24]),
    .Y(_3407_)
);

FILL FILL_3_BUFX2_insert59 (
);

FILL FILL_1_BUFX2_insert613 (
);

FILL FILL_0__12226_ (
);

FILL FILL_1_BUFX2_insert614 (
);

FILL FILL_1_BUFX2_insert615 (
);

FILL FILL_1_BUFX2_insert616 (
);

FILL FILL_1_BUFX2_insert617 (
);

FILL FILL_5__8263_ (
);

FILL FILL_1_BUFX2_insert618 (
);

FILL FILL_1_BUFX2_insert619 (
);

FILL FILL_5__15838_ (
);

FILL FILL_5__15418_ (
);

FILL SFILL39480x54050 (
);

FILL SFILL54280x60050 (
);

FILL FILL_3__16032_ (
);

INVX1 _9718_ (
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_1496_)
);

FILL FILL_5__10973_ (
);

FILL FILL_5__10553_ (
);

FILL FILL_1__8255_ (
);

FILL FILL_5__10133_ (
);

FILL FILL_2__15865_ (
);

FILL FILL_2__15445_ (
);

FILL FILL_2__15025_ (
);

FILL SFILL39000x83050 (
);

FILL SFILL94360x56050 (
);

FILL FILL_2__10580_ (
);

FILL FILL_2__10160_ (
);

FILL FILL_1__14858_ (
);

FILL FILL_1__14438_ (
);

FILL FILL_1__14018_ (
);

FILL FILL_3__9542_ (
);

FILL FILL_3__9122_ (
);

NOR2X1 _13716_ (
    .A(_4222_),
    .B(_3971__bF$buf3),
    .Y(_4223_)
);

FILL FILL_5__9888_ (
);

FILL FILL_5__9468_ (
);

OAI22X1 _16188_ (
    .A(_5485__bF$buf4),
    .B(_6639_),
    .C(_5483__bF$buf3),
    .D(_5281_),
    .Y(_6640_)
);

FILL FILL_5__11758_ (
);

FILL FILL_5__11338_ (
);

FILL FILL_3__12372_ (
);

FILL FILL_4__7885_ (
);

FILL FILL_4__7465_ (
);

FILL FILL_4__7045_ (
);

FILL FILL_2__11785_ (
);

FILL FILL_2__11365_ (
);

FILL SFILL94360x11050 (
);

FILL FILL_1__10778_ (
);

FILL FILL_1__10358_ (
);

FILL FILL_5__15591_ (
);

FILL FILL_5__15171_ (
);

INVX1 _9891_ (
    .A(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_1527_)
);

FILL FILL_0__7365_ (
);

INVX1 _9471_ (
    .A(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_1308_)
);

DFFSR _9051_ (
    .Q(\datapath_1.regfile_1.regOut[17] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_1043_[5])
);

FILL FILL_4__14584_ (
);

FILL FILL_4__14164_ (
);

FILL SFILL8760x73050 (
);

FILL FILL_2__8744_ (
);

FILL FILL_3__13997_ (
);

FILL FILL_2__8324_ (
);

FILL FILL_3__13577_ (
);

FILL FILL_3__13157_ (
);

FILL FILL_1__14191_ (
);

FILL SFILL114600x73050 (
);

FILL FILL_5__13904_ (
);

FILL SFILL53960x63050 (
);

FILL SFILL29000x81050 (
);

FILL FILL_4__9611_ (
);

FILL FILL_2__13931_ (
);

FILL FILL_5__16376_ (
);

FILL FILL_2__13511_ (
);

FILL FILL_5__11091_ (
);

FILL FILL_4__15789_ (
);

FILL FILL_4__15369_ (
);

FILL FILL_1__12504_ (
);

FILL FILL_0__9931_ (
);

FILL FILL_0__9511_ (
);

FILL FILL_0__11917_ (
);

FILL FILL_2__9529_ (
);

FILL FILL_2__9109_ (
);

FILL FILL_1__15396_ (
);

FILL FILL_5__7954_ (
);

FILL FILL_5__7114_ (
);

FILL FILL_4__16310_ (
);

FILL FILL_0__14389_ (
);

INVX1 _14674_ (
    .A(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_5161_)
);

INVX1 _14254_ (
    .A(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_4750_)
);

FILL FILL_3__15723_ (
);

FILL FILL_3__15303_ (
);

FILL FILL_1__7946_ (
);

FILL FILL_1__7106_ (
);

FILL FILL_2__14716_ (
);

FILL FILL_0__15750_ (
);

FILL FILL_0__15330_ (
);

FILL SFILL114920x49050 (
);

FILL FILL_5__12296_ (
);

FILL FILL_1__13709_ (
);

FILL FILL_4__11289_ (
);

FILL FILL_5__8739_ (
);

FILL SFILL114520x35050 (
);

FILL FILL_5__8319_ (
);

OAI22X1 _15879_ (
    .A(_5485__bF$buf1),
    .B(_6338_),
    .C(_5526__bF$buf1),
    .D(_4920_),
    .Y(_6339_)
);

FILL FILL_4__12650_ (
);

INVX1 _15459_ (
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_5929_)
);

NAND3X1 _15039_ (
    .A(_5475_),
    .B(\datapath_1.PCJump [23]),
    .C(_5477_),
    .Y(_5519_)
);

FILL FILL_4__12230_ (
);

DFFSR _10594_ (
    .Q(\datapath_1.regfile_1.regOut[29] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_1823_[12])
);

INVX1 _10174_ (
    .A(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_1675_)
);

FILL FILL_3__11643_ (
);

FILL SFILL43960x61050 (
);

FILL FILL_3__11223_ (
);

FILL FILL_6__14088_ (
);

NAND2X1 _16400_ (
    .A(gnd),
    .B(gnd),
    .Y(_6821_)
);

FILL FILL_0__16115_ (
);

FILL FILL_2__10636_ (
);

FILL FILL_2__9282_ (
);

FILL FILL_0__11670_ (
);

FILL FILL_0__11250_ (
);

FILL SFILL78680x60050 (
);

FILL FILL_5__14862_ (
);

FILL FILL_5__14442_ (
);

FILL FILL_5__14022_ (
);

INVX1 _8742_ (
    .A(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_944_)
);

FILL SFILL104520x78050 (
);

INVX1 _8322_ (
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_725_)
);

FILL SFILL43880x68050 (
);

FILL FILL_4__13855_ (
);

FILL FILL_4__13435_ (
);

FILL FILL_4__13015_ (
);

NOR2X1 _11799_ (
    .A(_2891_),
    .B(_2883_),
    .Y(_2892_)
);

OAI21X1 _11379_ (
    .A(_2494_),
    .B(_2488_),
    .C(_2495_),
    .Y(_2496_)
);

FILL FILL_3__12848_ (
);

FILL FILL_3__12428_ (
);

FILL FILL_1__13882_ (
);

FILL FILL_1__13462_ (
);

FILL FILL_3__12008_ (
);

FILL FILL_1__13042_ (
);

FILL SFILL59080x39050 (
);

FILL FILL_0__12875_ (
);

INVX1 _12740_ (
    .A(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3519_)
);

FILL FILL_0__12455_ (
);

FILL FILL_0__12035_ (
);

NAND3X1 _12320_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf0),
    .Y(_3279_)
);

FILL FILL_5__8492_ (
);

FILL FILL_5__8072_ (
);

FILL FILL_5__15647_ (
);

FILL FILL_5__15227_ (
);

FILL FILL_3__16261_ (
);

DFFSR _9947_ (
    .Q(\datapath_1.regfile_1.regOut[24] [5]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_1498_[5])
);

OAI21X1 _9527_ (
    .A(_1344_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .C(_1345_),
    .Y(_1303_[21])
);

FILL SFILL3640x16050 (
);

OAI21X1 _9107_ (
    .A(_1125_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1126_),
    .Y(_1108_[9])
);

FILL FILL_5__10782_ (
);

FILL FILL_1__8484_ (
);

FILL FILL_5__10362_ (
);

FILL FILL_1__8064_ (
);

FILL FILL_2__15674_ (
);

FILL SFILL104520x33050 (
);

FILL FILL_2__15254_ (
);

FILL SFILL43880x23050 (
);

FILL FILL_1__14667_ (
);

FILL FILL_1__14247_ (
);

FILL FILL_0_BUFX2_insert270 (
);

FILL FILL_0_BUFX2_insert271 (
);

FILL SFILL59000x37050 (
);

FILL FILL_0_BUFX2_insert272 (
);

FILL FILL_0_BUFX2_insert273 (
);

FILL FILL_3__9771_ (
);

FILL FILL_0_BUFX2_insert274 (
);

FILL FILL_3__9351_ (
);

OAI22X1 _13945_ (
    .A(_4446_),
    .B(_3909_),
    .C(_3881_),
    .D(_4445_),
    .Y(_4447_)
);

FILL FILL_0_BUFX2_insert275 (
);

OAI22X1 _13525_ (
    .A(_3947__bF$buf3),
    .B(_4035_),
    .C(_3944__bF$buf4),
    .D(_4034_),
    .Y(_4036_)
);

OAI21X1 _13105_ (
    .A(_3700_),
    .B(PCEn_bF$buf6),
    .C(_3701_),
    .Y(_3685_[8])
);

FILL FILL_0_BUFX2_insert276 (
);

FILL FILL_0_BUFX2_insert277 (
);

FILL FILL_0_BUFX2_insert278 (
);

FILL FILL_5__9277_ (
);

FILL FILL_0_BUFX2_insert279 (
);

FILL FILL_0__14601_ (
);

FILL FILL_5__11987_ (
);

FILL FILL_5__11567_ (
);

FILL FILL_1__9269_ (
);

FILL FILL_5__11147_ (
);

FILL FILL_3__12181_ (
);

FILL FILL_4__7694_ (
);

FILL FILL_2__16039_ (
);

FILL FILL_2__11594_ (
);

FILL FILL_2__11174_ (
);

FILL FILL_1__10167_ (
);

FILL FILL_4__11921_ (
);

FILL FILL_4__11501_ (
);

FILL FILL_0__7594_ (
);

FILL FILL_6__8981_ (
);

FILL SFILL49080x37050 (
);

FILL FILL_0__7174_ (
);

OAI21X1 _9280_ (
    .A(_1220_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .C(_1221_),
    .Y(_1173_[24])
);

FILL FILL_3__10914_ (
);

FILL FILL_4__14393_ (
);

FILL FILL_0__15806_ (
);

FILL FILL_2__8973_ (
);

FILL FILL_0__10941_ (
);

FILL FILL_3__13386_ (
);

FILL FILL_0__10521_ (
);

FILL FILL_2__8133_ (
);

FILL FILL_4__8899_ (
);

FILL FILL_4__8479_ (
);

FILL FILL_4__8059_ (
);

FILL FILL_2__12379_ (
);

FILL SFILL33880x21050 (
);

FILL FILL_5__13713_ (
);

FILL SFILL115000x5050 (
);

FILL FILL_1__6970_ (
);

FILL FILL_4__9420_ (
);

FILL FILL_4__9000_ (
);

FILL FILL_4__12706_ (
);

FILL FILL_2__13740_ (
);

FILL SFILL18600x44050 (
);

FILL FILL_2__13320_ (
);

FILL FILL_5__16185_ (
);

FILL FILL_3__6896_ (
);

FILL FILL_0__8379_ (
);

FILL FILL_1__12733_ (
);

FILL FILL_4__15598_ (
);

FILL FILL_4__15178_ (
);

FILL FILL_1__12313_ (
);

FILL SFILL94440x44050 (
);

FILL FILL_0__9740_ (
);

FILL FILL_2__9758_ (
);

FILL FILL_2__9338_ (
);

FILL FILL_0__11726_ (
);

FILL FILL_0__11306_ (
);

FILL FILL_6__15925_ (
);

FILL FILL_5__7763_ (
);

FILL FILL_5__7343_ (
);

FILL FILL_0__14198_ (
);

NAND3X1 _14483_ (
    .A(_4972_),
    .B(_4973_),
    .C(_4971_),
    .Y(_4974_)
);

NAND2X1 _14063_ (
    .A(_4562_),
    .B(_4555_),
    .Y(_4563_)
);

FILL FILL_5__14918_ (
);

FILL SFILL23880x64050 (
);

FILL FILL_3__15952_ (
);

FILL FILL_3__15532_ (
);

FILL SFILL98760x52050 (
);

FILL FILL_3__15112_ (
);

FILL FILL_1__7755_ (
);

FILL FILL_1__7335_ (
);

FILL FILL_2__14945_ (
);

FILL FILL_2__14525_ (
);

FILL FILL_2__14105_ (
);

FILL SFILL103720x29050 (
);

FILL FILL_1__13938_ (
);

FILL FILL_1__13518_ (
);

FILL FILL_4__11098_ (
);

FILL FILL_3__8622_ (
);

FILL FILL_3__8202_ (
);

FILL FILL_5__8968_ (
);

FILL FILL_5__8128_ (
);

FILL FILL_6__11845_ (
);

NOR2X1 _15688_ (
    .A(_6151_),
    .B(_6152_),
    .Y(_6153_)
);

FILL FILL_6__11425_ (
);

INVX1 _15268_ (
    .A(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_5743_)
);

FILL FILL_3__16317_ (
);

FILL FILL_3__11872_ (
);

FILL FILL_5__10418_ (
);

FILL FILL_3__11452_ (
);

FILL FILL_3__11032_ (
);

FILL FILL_4__6965_ (
);

FILL FILL_0__16344_ (
);

FILL FILL_2__10445_ (
);

FILL FILL_2__9091_ (
);

FILL FILL_2__10025_ (
);

FILL SFILL39000x33050 (
);

FILL FILL_1__9901_ (
);

FILL FILL112360x1050 (
);

FILL FILL_3__9407_ (
);

FILL FILL_5__14671_ (
);

FILL FILL_5__14251_ (
);

FILL FILL_0__6865_ (
);

FILL FILL112280x6050 (
);

INVX1 _8971_ (
    .A(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_1056_)
);

DFFSR _8551_ (
    .Q(\datapath_1.regfile_1.regOut[13] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_783_[17])
);

OAI21X1 _8131_ (
    .A(_637_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_638_),
    .Y(_588_[25])
);

FILL FILL_4__13664_ (
);

FILL SFILL8760x68050 (
);

FILL FILL_4__13244_ (
);

NAND2X1 _11188_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(_2306_),
    .Y(_2307_)
);

FILL FILL_2__7824_ (
);

FILL FILL_3__12657_ (
);

FILL FILL_3__12237_ (
);

FILL FILL_1__13691_ (
);

FILL FILL_1__13271_ (
);

FILL SFILL114600x68050 (
);

FILL FILL_0__12264_ (
);

FILL SFILL53960x58050 (
);

FILL FILL_6__16043_ (
);

FILL FILL_5__15876_ (
);

FILL FILL_5__15456_ (
);

FILL FILL_5__15036_ (
);

OAI21X1 _9756_ (
    .A(_1456_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1457_),
    .Y(_1433_[12])
);

FILL FILL_3__16070_ (
);

OAI21X1 _9336_ (
    .A(_1301_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1302_),
    .Y(_1238_[0])
);

FILL FILL_5__10171_ (
);

FILL FILL_4__14869_ (
);

FILL FILL_4__14449_ (
);

FILL FILL_4__14029_ (
);

FILL FILL_2__15483_ (
);

FILL FILL_2__15063_ (
);

FILL SFILL8760x23050 (
);

FILL FILL_2__8609_ (
);

FILL SFILL13800x60050 (
);

FILL FILL_1__14896_ (
);

FILL FILL_1__14476_ (
);

FILL FILL_1__14056_ (
);

FILL FILL_4__15810_ (
);

FILL FILL_0__13889_ (
);

INVX1 _13754_ (
    .A(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_4260_)
);

FILL FILL_0__13469_ (
);

FILL FILL_3__9160_ (
);

NOR2X1 _13334_ (
    .A(_3798_),
    .B(_3800_),
    .Y(\datapath_1.regfile_1.regEn [20])
);

FILL FILL_3__14803_ (
);

FILL FILL_5__9086_ (
);

FILL SFILL114600x23050 (
);

FILL SFILL53960x13050 (
);

FILL FILL_0__14830_ (
);

FILL FILL_0__14410_ (
);

FILL FILL_5__11796_ (
);

FILL FILL_1__9498_ (
);

FILL FILL_5__11376_ (
);

FILL FILL_1__9078_ (
);

FILL FILL_2__16268_ (
);

FILL FILL_4__10789_ (
);

FILL FILL_4__7083_ (
);

FILL FILL_4__10369_ (
);

FILL FILL_5__7819_ (
);

FILL FILL_1__10396_ (
);

OAI22X1 _14959_ (
    .A(_3947__bF$buf3),
    .B(_5439_),
    .C(_3909_),
    .D(_5438_),
    .Y(_5440_)
);

AOI22X1 _14539_ (
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .B(_4005__bF$buf2),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_5029_)
);

FILL FILL_4__11730_ (
);

FILL SFILL3720x49050 (
);

FILL FILL_4__11310_ (
);

NOR2X1 _14119_ (
    .A(_4614_),
    .B(_4617_),
    .Y(_4618_)
);

FILL FILL_1__16202_ (
);

FILL FILL_3__10303_ (
);

OAI22X1 _15900_ (
    .A(_5472__bF$buf1),
    .B(_4983_),
    .C(_4982_),
    .D(_5552__bF$buf0),
    .Y(_6359_)
);

FILL FILL_0__15615_ (
);

FILL FILL_2__8782_ (
);

FILL FILL_2__8362_ (
);

FILL FILL_0__10750_ (
);

FILL FILL112360x60050 (
);

FILL FILL_2__12188_ (
);

FILL FILL_5__13942_ (
);

FILL FILL_5__13522_ (
);

FILL FILL_5__13102_ (
);

INVX1 _7822_ (
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_473_)
);

DFFSR _7402_ (
    .Q(\datapath_1.regfile_1.regOut[4] [20]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_198_[20])
);

FILL FILL_4_BUFX2_insert500 (
);

FILL FILL_4_BUFX2_insert501 (
);

FILL FILL_4_BUFX2_insert502 (
);

FILL FILL_4_BUFX2_insert503 (
);

FILL FILL_4__12515_ (
);

FILL FILL_4_BUFX2_insert504 (
);

FILL FILL_4_BUFX2_insert505 (
);

FILL FILL_4_BUFX2_insert506 (
);

NOR2X1 _10879_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2027_)
);

FILL FILL_0__8188_ (
);

FILL FILL_4_BUFX2_insert507 (
);

DFFSR _10459_ (
    .Q(\datapath_1.regfile_1.regOut[28] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_1758_[5])
);

OAI21X1 _10039_ (
    .A(_1604_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1605_),
    .Y(_1563_[21])
);

FILL FILL_4_BUFX2_insert508 (
);

FILL FILL_3__11928_ (
);

FILL FILL_4_BUFX2_insert509 (
);

FILL FILL_1__12962_ (
);

FILL FILL_3__11508_ (
);

FILL FILL_1__12122_ (
);

FILL SFILL43960x11050 (
);

FILL FILL112280x67050 (
);

FILL FILL_2__9987_ (
);

FILL FILL_0__11955_ (
);

FILL FILL_2__9147_ (
);

OAI21X1 _11820_ (
    .A(_2903_),
    .B(_2902_),
    .C(_2910_),
    .Y(\datapath_1.ALUResult [3])
);

FILL FILL_0__11535_ (
);

FILL FILL_0__11115_ (
);

AOI21X1 _11400_ (
    .A(_2163_),
    .B(_2515_),
    .C(_2516_),
    .Y(_2517_)
);

FILL FILL_5__7992_ (
);

FILL FILL_5__7572_ (
);

INVX1 _14292_ (
    .A(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_4787_)
);

FILL FILL_5__14727_ (
);

FILL FILL_5__14307_ (
);

FILL FILL_3__15761_ (
);

FILL FILL_3__15341_ (
);

FILL SFILL44520x3050 (
);

OAI21X1 _8607_ (
    .A(_873_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_874_),
    .Y(_848_[13])
);

FILL FILL_1__7984_ (
);

FILL SFILL64760x59050 (
);

FILL FILL_1__7564_ (
);

FILL SFILL104520x28050 (
);

FILL FILL_2__14754_ (
);

FILL SFILL43880x18050 (
);

FILL FILL_2__14334_ (
);

FILL FILL_1__13747_ (
);

FILL FILL_1__13327_ (
);

FILL FILL_3__8851_ (
);

OAI21X1 _12605_ (
    .A(_3448_),
    .B(vdd),
    .C(_3449_),
    .Y(_3425_[12])
);

FILL FILL_3__8011_ (
);

FILL FILL112280x22050 (
);

FILL SFILL84280x5050 (
);

FILL FILL_5__8777_ (
);

FILL FILL_5__8357_ (
);

AOI21X1 _15497_ (
    .A(_5966_),
    .B(_5943_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [10])
);

AOI21X1 _15077_ (
    .A(_5508_),
    .B(_5556_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [0])
);

FILL FILL_3__16126_ (
);

FILL FILL_5__10647_ (
);

FILL FILL_1__8769_ (
);

FILL FILL_3__11681_ (
);

FILL FILL_1__8349_ (
);

FILL FILL_3__11261_ (
);

FILL FILL_2__15959_ (
);

FILL FILL_2__15539_ (
);

FILL FILL_2__15119_ (
);

FILL FILL_0__16153_ (
);

FILL FILL_2__10674_ (
);

FILL FILL_2__10254_ (
);

FILL FILL_3__9636_ (
);

FILL FILL_3_BUFX2_insert520 (
);

FILL FILL_3__9216_ (
);

FILL FILL_3_BUFX2_insert521 (
);

FILL FILL_3_BUFX2_insert522 (
);

FILL FILL_5__14480_ (
);

FILL FILL_3_BUFX2_insert523 (
);

FILL FILL_5__14060_ (
);

FILL FILL_3_BUFX2_insert524 (
);

OAI21X1 _8780_ (
    .A(_968_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_969_),
    .Y(_913_[28])
);

FILL FILL_3_BUFX2_insert525 (
);

OAI21X1 _8360_ (
    .A(_749_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .C(_750_),
    .Y(_718_[16])
);

FILL FILL_3_BUFX2_insert526 (
);

FILL FILL_3_BUFX2_insert527 (
);

FILL FILL_3_BUFX2_insert528 (
);

FILL FILL_3_BUFX2_insert529 (
);

FILL FILL_4__13893_ (
);

FILL FILL_6__12019_ (
);

FILL FILL_4__13473_ (
);

FILL FILL_3__12886_ (
);

FILL FILL_2__7633_ (
);

FILL FILL_3__12466_ (
);

FILL FILL_2__7213_ (
);

FILL FILL_3__12046_ (
);

FILL FILL_1__13080_ (
);

FILL FILL_4__7979_ (
);

FILL FILL_4__7559_ (
);

FILL FILL_2__11879_ (
);

FILL FILL_2__11459_ (
);

FILL FILL_0__12493_ (
);

FILL FILL_2__11039_ (
);

FILL SFILL33880x16050 (
);

FILL FILL_0__12073_ (
);

FILL SFILL53880x50 (
);

FILL FILL_4__8500_ (
);

FILL SFILL18600x39050 (
);

FILL FILL_5__15685_ (
);

FILL FILL_2__12400_ (
);

FILL FILL_0__7879_ (
);

FILL FILL_5__15265_ (
);

OAI21X1 _9985_ (
    .A(_1568_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .C(_1569_),
    .Y(_1563_[3])
);

FILL FILL_0__7459_ (
);

DFFSR _9565_ (
    .Q(\datapath_1.regfile_1.regOut[21] [7]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1303_[7])
);

FILL FILL_0__7039_ (
);

NAND2X1 _9145_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1152_)
);

FILL FILL_1__11813_ (
);

FILL FILL_4__14678_ (
);

FILL FILL_4__14258_ (
);

FILL FILL_2__15292_ (
);

FILL FILL_2__8838_ (
);

FILL FILL_0__10806_ (
);

FILL FILL_0__8400_ (
);

FILL FILL_1__14285_ (
);

FILL FILL_0_BUFX2_insert650 (
);

FILL FILL_5__6843_ (
);

FILL FILL_0_BUFX2_insert651 (
);

FILL FILL_0_BUFX2_insert652 (
);

FILL FILL_0_BUFX2_insert653 (
);

FILL FILL_0_BUFX2_insert654 (
);

INVX1 _13983_ (
    .A(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_4484_)
);

FILL FILL_0__13698_ (
);

FILL FILL_0__13278_ (
);

FILL FILL_0_BUFX2_insert655 (
);

OAI22X1 _13563_ (
    .A(_4071_),
    .B(_3893__bF$buf0),
    .C(_3972__bF$buf3),
    .D(_4072_),
    .Y(_4073_)
);

FILL FILL_0_BUFX2_insert656 (
);

NAND2X1 _13143_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_pcsrc.dout [21]),
    .Y(_3727_)
);

FILL FILL_0_BUFX2_insert657 (
);

FILL FILL_3__14612_ (
);

FILL FILL_0_BUFX2_insert658 (
);

FILL FILL_0_BUFX2_insert659 (
);

FILL FILL_2__13605_ (
);

FILL FILL_5__11185_ (
);

FILL FILL_2__16077_ (
);

FILL FILL_4__10178_ (
);

FILL FILL_3__7702_ (
);

FILL FILL_0__9605_ (
);

FILL FILL_5__7628_ (
);

FILL FILL_5__7208_ (
);

FILL FILL_4__16404_ (
);

FILL FILL_6__10925_ (
);

OAI22X1 _14768_ (
    .A(_3902__bF$buf3),
    .B(_5252_),
    .C(_5251_),
    .D(_3955__bF$buf2),
    .Y(_5253_)
);

FILL SFILL23800x57050 (
);

FILL SFILL79400x1050 (
);

OAI22X1 _14348_ (
    .A(_4840_),
    .B(_3944__bF$buf0),
    .C(_3959_),
    .D(_4841_),
    .Y(_4842_)
);

FILL FILL_3__15817_ (
);

FILL SFILL84040x68050 (
);

FILL FILL_1__16011_ (
);

FILL FILL_3__10952_ (
);

FILL FILL_3__10532_ (
);

FILL FILL_3__10112_ (
);

FILL FILL_0__15844_ (
);

FILL FILL_0__15424_ (
);

FILL FILL_0__15004_ (
);

FILL FILL_2__8591_ (
);

FILL SFILL39000x28050 (
);

FILL FILL_4__8097_ (
);

FILL FILL_3__8907_ (
);

FILL FILL_5__13751_ (
);

FILL FILL_5__13331_ (
);

OAI21X1 _7631_ (
    .A(_385_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_386_),
    .Y(_328_[29])
);

OAI21X1 _7211_ (
    .A(_166_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .C(_167_),
    .Y(_133_[17])
);

FILL FILL_4__12744_ (
);

FILL FILL_4__12324_ (
);

OAI21X1 _10688_ (
    .A(_1935_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .C(_1936_),
    .Y(_1888_[24])
);

FILL FILL_6__9384_ (
);

OAI21X1 _10268_ (
    .A(_1716_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1717_),
    .Y(_1693_[12])
);

FILL SFILL23800x12050 (
);

FILL FILL_2__6904_ (
);

FILL FILL_3__11737_ (
);

FILL FILL_1__12771_ (
);

FILL FILL_3__11317_ (
);

FILL FILL_1__12351_ (
);

FILL FILL_0__16209_ (
);

FILL FILL_2__9796_ (
);

FILL FILL_2__9376_ (
);

FILL FILL_0__11764_ (
);

FILL FILL_0__11344_ (
);

FILL SFILL78840x81050 (
);

FILL FILL_5__7381_ (
);

FILL SFILL13480x43050 (
);

FILL FILL_5__14956_ (
);

FILL FILL_3__15990_ (
);

FILL FILL_5__14536_ (
);

FILL FILL_3__15570_ (
);

FILL FILL_5__14116_ (
);

OAI21X1 _8836_ (
    .A(_985_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_986_),
    .Y(_978_[4])
);

FILL FILL_3__15150_ (
);

DFFSR _8416_ (
    .Q(\datapath_1.regfile_1.regOut[12] [10]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_718_[10])
);

FILL FILL_1__7373_ (
);

FILL FILL_4__13949_ (
);

FILL FILL_2__14983_ (
);

FILL FILL_4__13529_ (
);

FILL FILL_2__14563_ (
);

FILL FILL_4__13109_ (
);

FILL FILL_2__14143_ (
);

FILL SFILL103640x1050 (
);

FILL FILL_3__7299_ (
);

FILL SFILL13800x55050 (
);

FILL FILL_1__13976_ (
);

FILL FILL_1__13556_ (
);

FILL FILL_1__13136_ (
);

FILL SFILL74040x66050 (
);

FILL FILL_0__12969_ (
);

FILL FILL_3__8660_ (
);

OAI21X1 _12834_ (
    .A(_3560_),
    .B(vdd),
    .C(_3561_),
    .Y(_3555_[3])
);

FILL FILL_3__8240_ (
);

OAI21X1 _12414_ (
    .A(_3340_),
    .B(MemToReg_bF$buf2),
    .C(_3341_),
    .Y(\datapath_1.mux_wd3.dout [23])
);

FILL FILL_0__12129_ (
);

FILL FILL_5__8586_ (
);

FILL FILL_0__13910_ (
);

FILL FILL_3__16355_ (
);

FILL FILL_1__8998_ (
);

FILL FILL_5__10876_ (
);

FILL FILL_1__8578_ (
);

FILL FILL_3__11490_ (
);

FILL FILL_5__10036_ (
);

FILL FILL_3__11070_ (
);

FILL FILL_2__15768_ (
);

FILL FILL_2__15348_ (
);

FILL FILL_0__16382_ (
);

FILL FILL_2__10063_ (
);

FILL SFILL13800x10050 (
);

FILL FILL_3__9865_ (
);

AOI22X1 _13619_ (
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .B(_3942__bF$buf1),
    .C(_4051__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_4128_)
);

FILL FILL_4__10810_ (
);

FILL FILL_3__9025_ (
);

FILL FILL_6__7870_ (
);

FILL FILL_1__15702_ (
);

FILL FILL_4__13282_ (
);

FILL FILL_2__7862_ (
);

FILL FILL_3__12695_ (
);

FILL FILL_2__7442_ (
);

FILL FILL_3__12275_ (
);

FILL FILL_4__7368_ (
);

FILL FILL112360x55050 (
);

FILL FILL_2__11688_ (
);

FILL FILL_2__11268_ (
);

FILL FILL_5__12602_ (
);

INVX1 _6902_ (
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_66_)
);

FILL SFILL64040x64050 (
);

FILL FILL_5__15494_ (
);

FILL FILL_0__7688_ (
);

FILL FILL_5__15074_ (
);

FILL FILL_6__8655_ (
);

NAND2X1 _9794_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1483_)
);

NAND2X1 _9374_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1264_)
);

FILL FILL_4__14487_ (
);

FILL FILL_1__11622_ (
);

FILL FILL_4__14067_ (
);

FILL FILL_1__11202_ (
);

FILL FILL_2__8647_ (
);

FILL FILL_2__8227_ (
);

NAND2X1 _10900_ (
    .A(\control_1.reg_state.dout [0]),
    .B(_2048_),
    .Y(_2049_)
);

FILL FILL_0__10615_ (
);

FILL FILL_1__14094_ (
);

OAI21X1 _13792_ (
    .A(_4295_),
    .B(_3967__bF$buf0),
    .C(_4296_),
    .Y(_4297_)
);

NAND3X1 _13372_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3880_),
    .C(_3883_),
    .Y(_3884_)
);

FILL FILL_0__13087_ (
);

FILL FILL_5__13807_ (
);

FILL FILL_3__14841_ (
);

FILL FILL112360x10050 (
);

FILL FILL_3__14421_ (
);

FILL FILL_3__14001_ (
);

FILL FILL_4__9934_ (
);

FILL FILL_4__9514_ (
);

FILL FILL_2__13834_ (
);

FILL FILL_2__13414_ (
);

FILL FILL_5__16279_ (
);

FILL FILL_1__12827_ (
);

FILL FILL_1__12407_ (
);

CLKBUF1 CLKBUF1_insert200 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert201 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert202 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert203 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf21)
);

FILL FILL_3__7931_ (
);

FILL FILL_0__9414_ (
);

CLKBUF1 CLKBUF1_insert204 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert205 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert206 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf18)
);

FILL FILL_1__15299_ (
);

CLKBUF1 CLKBUF1_insert207 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert208 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf16)
);

FILL FILL_5__7857_ (
);

FILL FILL_5__7437_ (
);

CLKBUF1 CLKBUF1_insert209 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf15)
);

FILL FILL_4__16213_ (
);

NOR2X1 _14997_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5477_)
);

INVX1 _14577_ (
    .A(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_5066_)
);

OAI22X1 _14157_ (
    .A(_3884__bF$buf0),
    .B(_4653_),
    .C(_4654_),
    .D(_3925_),
    .Y(_4655_)
);

FILL FILL_3__15626_ (
);

FILL FILL_3__15206_ (
);

FILL FILL_1__16240_ (
);

FILL FILL_1__7849_ (
);

FILL FILL_3__10761_ (
);

FILL FILL_1__7429_ (
);

FILL FILL_2__14619_ (
);

FILL FILL_0__15653_ (
);

FILL FILL_0__15233_ (
);

FILL FILL_5__12199_ (
);

FILL SFILL54040x62050 (
);

FILL FILL_3__8716_ (
);

FILL FILL_5__13980_ (
);

FILL FILL_5__13560_ (
);

FILL FILL_5__13140_ (
);

OAI21X1 _7860_ (
    .A(_497_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_498_),
    .Y(_458_[20])
);

OAI21X1 _7440_ (
    .A(_278_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_279_),
    .Y(_263_[8])
);

DFFSR _7020_ (
    .Q(\datapath_1.regfile_1.regOut[1] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_3_[22])
);

FILL FILL_4__12973_ (
);

FILL FILL_4__12133_ (
);

OAI21X1 _10497_ (
    .A(_1828_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .C(_1829_),
    .Y(_1823_[3])
);

DFFSR _10077_ (
    .Q(\datapath_1.regfile_1.regOut[25] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_1563_[7])
);

FILL FILL_3__11966_ (
);

FILL FILL_3__11546_ (
);

FILL FILL_1__12580_ (
);

FILL FILL_3__11126_ (
);

FILL FILL_1__12160_ (
);

FILL FILL_0__16018_ (
);

NAND3X1 _16303_ (
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf0),
    .Y(_6752_)
);

FILL FILL_2__10959_ (
);

FILL FILL_2__10539_ (
);

FILL FILL_0__11993_ (
);

FILL FILL_0__11573_ (
);

FILL FILL_2__10119_ (
);

FILL FILL_0__11153_ (
);

FILL FILL_6__15772_ (
);

FILL FILL_6__15352_ (
);

FILL FILL_5__7190_ (
);

FILL FILL_2__11900_ (
);

FILL FILL_5__14765_ (
);

FILL FILL_0__6959_ (
);

FILL FILL_5__14345_ (
);

NAND2X1 _8645_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_900_)
);

NAND2X1 _8225_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_681_)
);

FILL FILL_1__7182_ (
);

FILL FILL_4__13758_ (
);

FILL FILL_4__13338_ (
);

FILL FILL_2__14792_ (
);

FILL FILL_2__14372_ (
);

FILL FILL_1__13785_ (
);

FILL FILL_1__13365_ (
);

FILL FILL_0__12778_ (
);

NAND2X1 _12643_ (
    .A(vdd),
    .B(memoryOutData[25]),
    .Y(_3475_)
);

FILL FILL_0__12358_ (
);

NAND3X1 _12223_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(vdd),
    .C(_3196__bF$buf0),
    .Y(_3206_)
);

FILL FILL_5__8395_ (
);

FILL SFILL79160x73050 (
);

FILL SFILL44040x60050 (
);

FILL FILL_6__11272_ (
);

FILL FILL_3__16164_ (
);

FILL FILL_5__10685_ (
);

FILL FILL_5__10265_ (
);

FILL FILL_1__8387_ (
);

FILL FILL_2__15997_ (
);

FILL FILL_0_BUFX2_insert1000 (
);

FILL FILL_0_BUFX2_insert1001 (
);

FILL FILL_2__15577_ (
);

FILL FILL_0_BUFX2_insert1002 (
);

FILL FILL_2__15157_ (
);

FILL FILL_0_BUFX2_insert1003 (
);

FILL FILL_0__16191_ (
);

FILL FILL_0_BUFX2_insert1004 (
);

FILL FILL_0_BUFX2_insert1005 (
);

FILL FILL_0_BUFX2_insert1006 (
);

FILL FILL_2__10292_ (
);

FILL FILL_0_BUFX2_insert1007 (
);

FILL FILL_0_BUFX2_insert1008 (
);

FILL FILL_0_BUFX2_insert1009 (
);

FILL FILL_4__15904_ (
);

FILL FILL_3__9674_ (
);

FILL FILL_3_BUFX2_insert900 (
);

AOI22X1 _13848_ (
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .B(_4005__bF$buf3),
    .C(_4001__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_4352_)
);

FILL FILL_3__9254_ (
);

FILL FILL_3_BUFX2_insert901 (
);

NOR2X1 _13428_ (
    .A(_3913_),
    .B(_3939_),
    .Y(_3940_)
);

FILL FILL_3_BUFX2_insert902 (
);

FILL SFILL109480x7050 (
);

FILL FILL_3_BUFX2_insert903 (
);

INVX1 _13008_ (
    .A(_2_[19]),
    .Y(_3657_)
);

FILL FILL_3_BUFX2_insert904 (
);

FILL FILL_3_BUFX2_insert905 (
);

FILL FILL_1__15931_ (
);

FILL FILL_3_BUFX2_insert906 (
);

FILL FILL_1__15511_ (
);

FILL FILL_3_BUFX2_insert907 (
);

FILL FILL_3_BUFX2_insert908 (
);

FILL FILL_3_BUFX2_insert909 (
);

FILL FILL_4__13091_ (
);

FILL FILL_0__14924_ (
);

FILL FILL_0__14504_ (
);

FILL SFILL109720x68050 (
);

FILL FILL_2__7671_ (
);

FILL FILL_2__7251_ (
);

FILL FILL_3__12084_ (
);

FILL FILL_4__7597_ (
);

FILL FILL_4__7177_ (
);

FILL FILL_2__11497_ (
);

FILL FILL_2__11077_ (
);

FILL FILL_5__12831_ (
);

FILL FILL_5__12411_ (
);

FILL FILL_4__11824_ (
);

FILL FILL_4__11404_ (
);

FILL FILL_0__7497_ (
);

FILL FILL_0__7077_ (
);

FILL FILL_6__8464_ (
);

DFFSR _9183_ (
    .Q(\datapath_1.regfile_1.regOut[18] [9]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_1108_[9])
);

FILL FILL_3__10817_ (
);

FILL FILL_1__11851_ (
);

FILL FILL_4__14296_ (
);

FILL FILL_1__11431_ (
);

FILL SFILL38760x80050 (
);

FILL FILL_1__11011_ (
);

FILL SFILL69160x71050 (
);

FILL FILL_0__15709_ (
);

FILL FILL_2__8876_ (
);

FILL FILL_2__8456_ (
);

FILL FILL_3__13289_ (
);

FILL FILL_0__10424_ (
);

FILL FILL_0__10004_ (
);

FILL FILL_5__6881_ (
);

DFFSR _13181_ (
    .Q(\datapath_1.mux_iord.din0 [6]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3685_[6])
);

FILL FILL_5__13616_ (
);

FILL FILL_3__14650_ (
);

FILL FILL_3__14230_ (
);

DFFSR _7916_ (
    .Q(\datapath_1.regfile_1.regOut[8] [22]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_458_[22])
);

FILL FILL_1__6873_ (
);

FILL FILL_4__9743_ (
);

FILL FILL_4__12609_ (
);

FILL FILL_2__13643_ (
);

FILL FILL_2__13223_ (
);

FILL FILL_5__16088_ (
);

FILL FILL_1__12636_ (
);

FILL FILL_1__12216_ (
);

FILL FILL_3__7740_ (
);

FILL FILL_0__9643_ (
);

FILL FILL_3__7320_ (
);

INVX1 _11914_ (
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_2984_)
);

FILL FILL_0__11629_ (
);

FILL FILL_0__9223_ (
);

FILL FILL_0__11209_ (
);

FILL FILL_6__15828_ (
);

FILL FILL_6__15408_ (
);

FILL FILL_5__7246_ (
);

FILL FILL_4__16022_ (
);

FILL FILL_6__10543_ (
);

OAI22X1 _14386_ (
    .A(_4877_),
    .B(_3936__bF$buf1),
    .C(_3902__bF$buf3),
    .D(_4878_),
    .Y(_4879_)
);

FILL FILL_3__15855_ (
);

FILL FILL_3__15435_ (
);

FILL FILL_3__15015_ (
);

FILL FILL_3__10990_ (
);

FILL FILL_1__7238_ (
);

FILL FILL_3__10570_ (
);

FILL FILL_3__10150_ (
);

FILL SFILL28840x3050 (
);

FILL FILL_2__14848_ (
);

FILL FILL_6_BUFX2_insert413 (
);

FILL FILL_0__15882_ (
);

FILL FILL_2__14428_ (
);

FILL FILL_2__14008_ (
);

FILL FILL_0__15462_ (
);

FILL FILL_0__15042_ (
);

FILL SFILL28760x8050 (
);

FILL FILL_6_BUFX2_insert418 (
);

FILL SFILL99640x79050 (
);

FILL FILL_3__8525_ (
);

FILL FILL_3__8105_ (
);

FILL FILL_6__6950_ (
);

FILL SFILL8680x4050 (
);

FILL FILL_6__11748_ (
);

FILL FILL_4__12782_ (
);

FILL FILL_6__11328_ (
);

FILL FILL_4__12362_ (
);

FILL SFILL64120x52050 (
);

FILL FILL_2__6942_ (
);

FILL FILL_5__9812_ (
);

FILL FILL_3__11775_ (
);

FILL FILL_3__11355_ (
);

FILL FILL_4__6868_ (
);

FILL FILL_0__16247_ (
);

NAND3X1 _16112_ (
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6566_)
);

FILL FILL_2__10768_ (
);

FILL FILL_0__11382_ (
);

FILL FILL_1__9804_ (
);

FILL FILL_5__14994_ (
);

FILL FILL_5__14574_ (
);

FILL FILL_5__14154_ (
);

FILL FILL_6__7735_ (
);

NAND2X1 _8874_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1012_)
);

NAND2X1 _8454_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_793_)
);

DFFSR _8034_ (
    .Q(\datapath_1.regfile_1.regOut[9] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_523_[12])
);

FILL FILL_4__13987_ (
);

FILL FILL_1__10702_ (
);

FILL FILL_4__13567_ (
);

FILL FILL_4__13147_ (
);

FILL FILL_2__14181_ (
);

FILL FILL_2__7727_ (
);

FILL FILL_2__7307_ (
);

FILL FILL_1__13594_ (
);

FILL SFILL54920x78050 (
);

FILL FILL_1__13174_ (
);

FILL FILL_0__12587_ (
);

NAND2X1 _12872_ (
    .A(vdd),
    .B(\datapath_1.rd1 [16]),
    .Y(_3587_)
);

NAND2X1 _12452_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [4]),
    .Y(_3368_)
);

FILL FILL_0__12167_ (
);

NAND3X1 _12032_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [11]),
    .C(_3034__bF$buf3),
    .Y(_3070_)
);

FILL FILL_3__13921_ (
);

FILL FILL_3__13501_ (
);

FILL SFILL89640x77050 (
);

FILL FILL_5_BUFX2_insert430 (
);

FILL FILL_5_BUFX2_insert431 (
);

FILL FILL_5__15779_ (
);

FILL FILL_2__12914_ (
);

FILL FILL_5__15359_ (
);

FILL FILL_5_BUFX2_insert432 (
);

FILL FILL_5_BUFX2_insert433 (
);

FILL FILL_3__16393_ (
);

INVX1 _9659_ (
    .A(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_1413_)
);

FILL FILL_5_BUFX2_insert434 (
);

INVX1 _9239_ (
    .A(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_1194_)
);

FILL FILL_5_BUFX2_insert435 (
);

FILL SFILL64040x14050 (
);

FILL FILL_5_BUFX2_insert436 (
);

FILL FILL_5__10494_ (
);

FILL FILL_1__8196_ (
);

FILL FILL_5_BUFX2_insert437 (
);

FILL FILL_5_BUFX2_insert438 (
);

FILL FILL_1__11907_ (
);

FILL FILL_5_BUFX2_insert439 (
);

FILL FILL_2__15386_ (
);

FILL FILL_5__16300_ (
);

FILL FILL_0__8914_ (
);

FILL SFILL89240x63050 (
);

FILL FILL_1__14799_ (
);

FILL FILL_1__14379_ (
);

FILL FILL_5__6937_ (
);

FILL SFILL68360x22050 (
);

FILL FILL_4__15713_ (
);

FILL FILL_3__9483_ (
);

INVX1 _13657_ (
    .A(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_4165_)
);

OAI21X1 _13237_ (
    .A(_3775_),
    .B(_3779_),
    .C(\datapath_1.a3 [4]),
    .Y(_3780_)
);

FILL FILL_3__14706_ (
);

FILL SFILL18680x83050 (
);

FILL FILL_1__15740_ (
);

FILL FILL_1__15320_ (
);

FILL FILL_1__6929_ (
);

FILL FILL_0__14733_ (
);

FILL FILL_0__14313_ (
);

FILL SFILL58760x79050 (
);

FILL FILL_5__11699_ (
);

FILL FILL_2__7480_ (
);

FILL FILL_5__11279_ (
);

FILL FILL_2__7060_ (
);

FILL FILL_5__12640_ (
);

FILL FILL_5__12220_ (
);

OAI21X1 _6940_ (
    .A(_26_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .C(_27_),
    .Y(_3_[12])
);

FILL FILL_2_BUFX2_insert560 (
);

FILL FILL_1__10299_ (
);

FILL FILL_2_BUFX2_insert561 (
);

FILL FILL_2_BUFX2_insert562 (
);

FILL FILL_2_BUFX2_insert563 (
);

FILL FILL_2_BUFX2_insert564 (
);

FILL FILL_4__11633_ (
);

FILL FILL_2_BUFX2_insert565 (
);

FILL FILL_4__11213_ (
);

FILL FILL_2_BUFX2_insert566 (
);

FILL FILL_2_BUFX2_insert567 (
);

FILL FILL_2_BUFX2_insert568 (
);

FILL FILL_6__8273_ (
);

FILL FILL_2_BUFX2_insert569 (
);

FILL FILL_1__16105_ (
);

FILL FILL_3__10626_ (
);

FILL FILL_1__11660_ (
);

FILL FILL_1__11240_ (
);

FILL FILL_0__15938_ (
);

FILL FILL_0__15518_ (
);

NOR2X1 _15803_ (
    .A(_6263_),
    .B(_6264_),
    .Y(_6265_)
);

FILL FILL_2__8265_ (
);

FILL FILL_0__10653_ (
);

FILL FILL_3__13098_ (
);

FILL FILL_0__10233_ (
);

FILL SFILL54040x12050 (
);

FILL FILL_6__14012_ (
);

FILL FILL_5__13845_ (
);

FILL FILL_5__13425_ (
);

FILL FILL_5__13005_ (
);

NAND2X1 _7725_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_429_)
);

NAND2X1 _7305_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_210_)
);

FILL SFILL79240x61050 (
);

FILL FILL_4__9552_ (
);

FILL FILL_4__9132_ (
);

FILL FILL_4__12838_ (
);

FILL FILL_2__13872_ (
);

FILL FILL_4__12418_ (
);

FILL FILL_2__13452_ (
);

FILL FILL_2__13032_ (
);

FILL FILL_6__9478_ (
);

FILL FILL_1__12865_ (
);

FILL FILL_1__12445_ (
);

FILL FILL_1__12025_ (
);

FILL FILL_0__9872_ (
);

FILL FILL_0__11858_ (
);

FILL FILL_0__9032_ (
);

OAI21X1 _11723_ (
    .A(_2800_),
    .B(_2344__bF$buf1),
    .C(_2820_),
    .Y(_2821_)
);

FILL FILL_0__11438_ (
);

FILL FILL_0__11018_ (
);

NOR2X1 _11303_ (
    .A(_2421_),
    .B(_2415_),
    .Y(_2422_)
);

FILL FILL_5__7475_ (
);

FILL SFILL44040x55050 (
);

FILL FILL_5__7055_ (
);

FILL FILL_4__16251_ (
);

NOR2X1 _14195_ (
    .A(_4691_),
    .B(_4679_),
    .Y(_4692_)
);

FILL FILL_3__15664_ (
);

FILL FILL_3__15244_ (
);

FILL FILL_1__7887_ (
);

FILL FILL_1__7467_ (
);

FILL FILL_1__7047_ (
);

FILL FILL_2__14657_ (
);

FILL FILL_0__15691_ (
);

FILL FILL_2__14237_ (
);

FILL FILL_0__15271_ (
);

FILL FILL_1_BUFX2_insert580 (
);

FILL FILL_1_BUFX2_insert581 (
);

FILL FILL_3__8754_ (
);

FILL FILL_1_BUFX2_insert582 (
);

FILL FILL_3__8334_ (
);

DFFSR _12928_ (
    .Q(\datapath_1.a [9]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_3555_[9])
);

FILL FILL_1_BUFX2_insert583 (
);

INVX1 _12508_ (
    .A(ALUOut[23]),
    .Y(_3405_)
);

FILL FILL_1_BUFX2_insert584 (
);

FILL FILL_1_BUFX2_insert585 (
);

FILL FILL_1_BUFX2_insert586 (
);

FILL FILL_1_BUFX2_insert587 (
);

FILL FILL_1_BUFX2_insert588 (
);

FILL FILL_1_BUFX2_insert589 (
);

FILL FILL_4__12591_ (
);

FILL FILL_4__12171_ (
);

FILL SFILL44040x10050 (
);

FILL FILL_3__16449_ (
);

FILL FILL_3__16029_ (
);

FILL FILL_5__9621_ (
);

FILL FILL_3__11584_ (
);

FILL FILL_3__11164_ (
);

OAI21X1 _16341_ (
    .A(_6780_),
    .B(gnd),
    .C(_6781_),
    .Y(_6769_[6])
);

FILL FILL_0__16056_ (
);

FILL FILL_2__10997_ (
);

FILL FILL_2__10577_ (
);

FILL FILL_2__10157_ (
);

FILL FILL_0__11191_ (
);

FILL FILL_5__11911_ (
);

FILL FILL_1__9613_ (
);

FILL FILL_3__9539_ (
);

FILL FILL_4__10904_ (
);

FILL FILL_3__9119_ (
);

FILL FILL_0__6997_ (
);

FILL FILL_5__14383_ (
);

DFFSR _8683_ (
    .Q(\datapath_1.regfile_1.regOut[14] [21]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_848_[21])
);

INVX1 _8263_ (
    .A(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_706_)
);

FILL FILL_1__10931_ (
);

FILL FILL_4__13796_ (
);

FILL FILL_1__10511_ (
);

FILL FILL_4__13376_ (
);

FILL SFILL69160x66050 (
);

FILL SFILL34040x53050 (
);

FILL FILL_2__7956_ (
);

FILL FILL_3__12789_ (
);

BUFX2 BUFX2_insert250 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf4)
);

FILL FILL_2__7116_ (
);

FILL FILL_3__12369_ (
);

BUFX2 BUFX2_insert251 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf3)
);

BUFX2 BUFX2_insert252 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf2)
);

BUFX2 BUFX2_insert253 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf1)
);

BUFX2 BUFX2_insert254 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf0)
);

FILL SFILL74120x49050 (
);

BUFX2 BUFX2_insert255 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf4 )
);

BUFX2 BUFX2_insert256 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf3 )
);

BUFX2 BUFX2_insert257 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf2 )
);

BUFX2 BUFX2_insert258 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf1 )
);

DFFSR _12681_ (
    .Q(\datapath_1.Data [18]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[18])
);

BUFX2 BUFX2_insert259 (
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf0 )
);

FILL FILL_0__12396_ (
);

AOI22X1 _12261_ (
    .A(_2_[11]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [11]),
    .Y(_3235_)
);

FILL FILL_3__13730_ (
);

FILL FILL_3__13310_ (
);

FILL FILL_4__8823_ (
);

FILL FILL_4__8403_ (
);

FILL FILL_2__12723_ (
);

FILL FILL_5__15588_ (
);

FILL FILL_5__15168_ (
);

FILL FILL_2__12303_ (
);

INVX1 _9888_ (
    .A(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_1525_)
);

INVX1 _9468_ (
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_1306_)
);

DFFSR _9048_ (
    .Q(\datapath_1.regfile_1.regOut[17] [2]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_1043_[2])
);

FILL FILL_1__11716_ (
);

FILL FILL_2__15195_ (
);

FILL FILL_0__8723_ (
);

FILL FILL_0__10709_ (
);

FILL FILL_1__14188_ (
);

FILL FILL_4__15942_ (
);

FILL FILL_4__15522_ (
);

FILL FILL_4__15102_ (
);

NOR2X1 _13886_ (
    .A(_4377_),
    .B(_4389_),
    .Y(_4390_)
);

FILL FILL_3__9292_ (
);

NAND3X1 _13466_ (
    .A(_3898_),
    .B(_3880_),
    .C(_3879_),
    .Y(_3978_)
);

OAI21X1 _13046_ (
    .A(_3681_),
    .B(vdd),
    .C(_3682_),
    .Y(_3620_[31])
);

FILL FILL_3__14935_ (
);

FILL FILL_3__14515_ (
);

FILL FILL_4__9608_ (
);

FILL FILL_2__13928_ (
);

FILL FILL_0__14962_ (
);

FILL FILL_2__13508_ (
);

FILL SFILL99320x53050 (
);

FILL FILL_0__14542_ (
);

FILL FILL_0__14122_ (
);

FILL FILL_5__11088_ (
);

FILL FILL_0__9928_ (
);

FILL FILL_0__9508_ (
);

FILL FILL_3__7605_ (
);

FILL SFILL59160x64050 (
);

FILL FILL_4__16307_ (
);

FILL SFILL68840x69050 (
);

FILL FILL_6__10408_ (
);

FILL FILL_4__11862_ (
);

FILL FILL_4__11442_ (
);

FILL SFILL64120x47050 (
);

FILL FILL_4__11022_ (
);

FILL FILL_1__16334_ (
);

FILL FILL_6__8082_ (
);

FILL FILL_3__10435_ (
);

FILL FILL_3__10015_ (
);

FILL FILL_0__15747_ (
);

FILL FILL_0__15327_ (
);

INVX1 _15612_ (
    .A(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_6078_)
);

FILL FILL_0__10882_ (
);

FILL FILL_2__8494_ (
);

FILL FILL_2__8074_ (
);

FILL FILL_0__10042_ (
);

FILL FILL_6__14661_ (
);

FILL FILL_5__13654_ (
);

FILL FILL_5__13234_ (
);

NAND2X1 _7954_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_541_)
);

DFFSR _7534_ (
    .Q(\datapath_1.regfile_1.regOut[5] [24]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_263_[24])
);

INVX1 _7114_ (
    .A(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_123_)
);

FILL FILL_4__9781_ (
);

FILL FILL_4__9361_ (
);

FILL FILL_4__12647_ (
);

FILL FILL_2__13681_ (
);

FILL FILL_4__12227_ (
);

FILL FILL_2__13261_ (
);

FILL FILL_1__12254_ (
);

FILL FILL_0__9681_ (
);

FILL FILL_2__9279_ (
);

OAI21X1 _11952_ (
    .A(_3008_),
    .B(IorD_bF$buf5),
    .C(_3009_),
    .Y(_1_[21])
);

FILL FILL_0__9261_ (
);

FILL FILL_0__11667_ (
);

FILL FILL_0__11247_ (
);

OAI21X1 _11532_ (
    .A(_2547_),
    .B(_2548_),
    .C(_2567_),
    .Y(_2643_)
);

FILL SFILL89320x51050 (
);

NOR2X1 _11112_ (
    .A(_2230_),
    .B(_2229_),
    .Y(_2231_)
);

FILL FILL_4__16060_ (
);

FILL FILL_5__14859_ (
);

FILL FILL_3__15893_ (
);

FILL FILL_5__14439_ (
);

FILL FILL_5__14019_ (
);

FILL FILL_3__15473_ (
);

INVX1 _8739_ (
    .A(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_942_)
);

FILL FILL_3__15053_ (
);

FILL SFILL18760x71050 (
);

INVX1 _8319_ (
    .A(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_723_)
);

FILL FILL_1__7696_ (
);

FILL FILL_2__14886_ (
);

FILL FILL_2__14466_ (
);

FILL FILL_2__14046_ (
);

FILL FILL_0__15080_ (
);

FILL FILL_5__15800_ (
);

FILL SFILL89240x58050 (
);

FILL SFILL54120x45050 (
);

FILL FILL_1__13879_ (
);

FILL FILL_1__13459_ (
);

FILL FILL_1__13039_ (
);

FILL FILL_3__8983_ (
);

FILL FILL_3__8143_ (
);

INVX1 _12737_ (
    .A(\datapath_1.PCJump [16]),
    .Y(_3517_)
);

AOI22X1 _12317_ (
    .A(_2_[25]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3277_)
);

FILL FILL_1__14820_ (
);

FILL FILL_5__8489_ (
);

FILL FILL_1__14400_ (
);

FILL FILL_5__8069_ (
);

FILL FILL_0__13813_ (
);

FILL FILL_3__16258_ (
);

FILL FILL_5__10779_ (
);

FILL FILL_2__6980_ (
);

FILL FILL_5__10359_ (
);

FILL FILL_5__9850_ (
);

FILL FILL_3__11393_ (
);

FILL FILL_5__9010_ (
);

FILL FILL_0__16285_ (
);

INVX1 _16150_ (
    .A(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_6603_)
);

FILL FILL_2__10386_ (
);

FILL FILL_5__11720_ (
);

FILL FILL_1__9422_ (
);

FILL FILL_5__11300_ (
);

FILL FILL_1__9002_ (
);

FILL SFILL89240x13050 (
);

FILL FILL_3__9768_ (
);

FILL FILL_3__9348_ (
);

FILL FILL_5__14192_ (
);

FILL FILL_6__7353_ (
);

INVX1 _8492_ (
    .A(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_818_)
);

FILL FILL_1__15605_ (
);

INVX1 _8072_ (
    .A(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_599_)
);

FILL SFILL18680x33050 (
);

FILL FILL_1__10320_ (
);

FILL FILL_2__7765_ (
);

FILL FILL_3__12598_ (
);

FILL FILL_2__7345_ (
);

FILL FILL_3__12178_ (
);

FILL FILL111960x62050 (
);

INVX1 _12490_ (
    .A(ALUOut[17]),
    .Y(_3393_)
);

NAND3X1 _12070_ (
    .A(_3096_),
    .B(_3097_),
    .C(_3098_),
    .Y(\datapath_1.mux_pcsrc.dout [20])
);

FILL FILL_5__12505_ (
);

FILL SFILL79240x56050 (
);

FILL FILL_4__8632_ (
);

FILL FILL_4__11918_ (
);

FILL FILL_5_BUFX2_insert810 (
);

FILL FILL_4__8212_ (
);

FILL FILL_5_BUFX2_insert811 (
);

FILL FILL_2__12952_ (
);

FILL FILL_5__15397_ (
);

FILL FILL_2__12532_ (
);

FILL FILL_5_BUFX2_insert812 (
);

FILL FILL_2__12112_ (
);

FILL FILL_5_BUFX2_insert813 (
);

FILL FILL_5_BUFX2_insert814 (
);

DFFSR _9697_ (
    .Q(\datapath_1.regfile_1.regOut[22] [11]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_1368_[11])
);

OAI21X1 _9277_ (
    .A(_1218_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1219_),
    .Y(_1173_[23])
);

FILL FILL_6__8138_ (
);

FILL FILL_5_BUFX2_insert815 (
);

FILL FILL_5_BUFX2_insert816 (
);

FILL FILL111880x69050 (
);

FILL FILL_5_BUFX2_insert817 (
);

FILL FILL_1__11945_ (
);

FILL FILL_5_BUFX2_insert818 (
);

FILL FILL_1__11525_ (
);

FILL FILL_5_BUFX2_insert819 (
);

FILL FILL_1__11105_ (
);

FILL FILL_0__8952_ (
);

FILL FILL_0__10938_ (
);

FILL FILL_0__8532_ (
);

FILL FILL_0__8112_ (
);

NAND2X1 _10803_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1993_)
);

FILL FILL_0__10518_ (
);

FILL FILL_5__6975_ (
);

FILL FILL_4__15751_ (
);

FILL FILL_4__15331_ (
);

INVX1 _13695_ (
    .A(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_4202_)
);

OR2X2 _13275_ (
    .A(_3796_),
    .B(_3815_),
    .Y(_3816_)
);

FILL FILL_2__9911_ (
);

FILL FILL_3__14744_ (
);

FILL FILL_3__14324_ (
);

FILL FILL_1__6967_ (
);

FILL FILL_4__9417_ (
);

FILL FILL_2__13737_ (
);

FILL SFILL79240x11050 (
);

FILL FILL_2__13317_ (
);

FILL FILL_0__14771_ (
);

FILL FILL_0__14351_ (
);

FILL FILL_0__9737_ (
);

FILL FILL_3__7834_ (
);

FILL FILL_3__7414_ (
);

FILL SFILL69640x68050 (
);

FILL FILL_2_BUFX2_insert940 (
);

FILL FILL_4__16116_ (
);

FILL FILL_2_BUFX2_insert941 (
);

FILL SFILL109400x37050 (
);

FILL FILL_2_BUFX2_insert942 (
);

FILL FILL_2_BUFX2_insert943 (
);

FILL FILL_2_BUFX2_insert944 (
);

FILL FILL_4__11671_ (
);

FILL FILL_2_BUFX2_insert945 (
);

FILL FILL_4__11251_ (
);

FILL FILL_2_BUFX2_insert946 (
);

FILL FILL_3__15949_ (
);

FILL FILL_2_BUFX2_insert947 (
);

FILL FILL_3__15529_ (
);

FILL FILL_2_BUFX2_insert948 (
);

FILL FILL_3__15109_ (
);

FILL FILL_2_BUFX2_insert949 (
);

FILL FILL_1__16143_ (
);

FILL FILL_3__10664_ (
);

FILL FILL_5__8701_ (
);

FILL FILL_3__10244_ (
);

FILL FILL_0__15976_ (
);

FILL SFILL69240x54050 (
);

FILL FILL_0__15556_ (
);

OAI22X1 _15841_ (
    .A(_4856_),
    .B(_5548__bF$buf1),
    .C(_5526__bF$buf1),
    .D(_4875_),
    .Y(_6302_)
);

NOR3X1 _15421_ (
    .A(_5887_),
    .B(_5889_),
    .C(_5891_),
    .Y(_5892_)
);

FILL FILL_0__15136_ (
);

INVX4 _15001_ (
    .A(_5480__bF$buf3),
    .Y(_5481_)
);

FILL FILL_0__10691_ (
);

FILL FILL_0__10271_ (
);

FILL FILL_3__8619_ (
);

FILL FILL_5__13883_ (
);

FILL FILL_5__13463_ (
);

FILL FILL_5__13043_ (
);

INVX1 _7763_ (
    .A(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_454_)
);

INVX1 _7343_ (
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_235_)
);

FILL FILL_4__9590_ (
);

FILL FILL_4__12876_ (
);

FILL FILL_4__9170_ (
);

FILL FILL_4__12456_ (
);

FILL FILL_2__13490_ (
);

FILL FILL_4__12036_ (
);

FILL FILL_3__11869_ (
);

FILL FILL_5__9906_ (
);

FILL FILL_3__11449_ (
);

FILL FILL_1__12483_ (
);

FILL FILL_3__11029_ (
);

FILL FILL_1__12063_ (
);

OAI22X1 _16206_ (
    .A(_5489__bF$buf2),
    .B(_5354_),
    .C(_5527__bF$buf1),
    .D(_5319_),
    .Y(_6657_)
);

FILL FILL_0__11896_ (
);

FILL FILL_0__9490_ (
);

FILL FILL_2__9088_ (
);

AOI21X1 _11761_ (
    .A(_2854_),
    .B(_2855_),
    .C(_2364_),
    .Y(_2856_)
);

FILL FILL_0__11476_ (
);

OAI21X1 _11341_ (
    .A(_2110_),
    .B(_2457_),
    .C(_2459_),
    .Y(_2460_)
);

FILL FILL_0__11056_ (
);

FILL FILL_6__15255_ (
);

FILL FILL_5__7093_ (
);

FILL FILL_2__11803_ (
);

FILL FILL_5__14668_ (
);

FILL FILL_5__14248_ (
);

INVX1 _8968_ (
    .A(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_1054_)
);

FILL FILL_3__15282_ (
);

FILL FILL_6__7829_ (
);

DFFSR _8548_ (
    .Q(\datapath_1.regfile_1.regOut[13] [14]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_783_[14])
);

OAI21X1 _8128_ (
    .A(_635_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .C(_636_),
    .Y(_588_[24])
);

FILL FILL_1__7085_ (
);

FILL FILL_2__14695_ (
);

FILL FILL_2__14275_ (
);

FILL SFILL99400x41050 (
);

FILL SFILL69160x16050 (
);

FILL FILL_0__7803_ (
);

FILL FILL_1__13688_ (
);

FILL FILL_1__13268_ (
);

FILL FILL_4__14602_ (
);

FILL FILL_1_BUFX2_insert960 (
);

FILL FILL_1_BUFX2_insert961 (
);

FILL FILL_1_BUFX2_insert962 (
);

INVX1 _12966_ (
    .A(_2_[5]),
    .Y(_3629_)
);

FILL FILL_3__8372_ (
);

FILL FILL_1_BUFX2_insert963 (
);

DFFSR _12546_ (
    .Q(ALUOut[11]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3360_[11])
);

FILL SFILL59240x52050 (
);

OAI21X1 _12126_ (
    .A(_3136_),
    .B(ALUSrcA_bF$buf7),
    .C(_3137_),
    .Y(\datapath_1.alu_1.ALUInA [3])
);

FILL FILL_1_BUFX2_insert964 (
);

FILL FILL_1_BUFX2_insert965 (
);

FILL FILL_1_BUFX2_insert966 (
);

FILL FILL_1_BUFX2_insert967 (
);

FILL FILL_1_BUFX2_insert968 (
);

FILL FILL_1_BUFX2_insert969 (
);

FILL FILL_6__11175_ (
);

FILL SFILL99320x48050 (
);

FILL FILL_0__13622_ (
);

FILL FILL_3__16067_ (
);

FILL FILL_5__10168_ (
);

FILL FILL_0__16094_ (
);

FILL SFILL28760x68050 (
);

FILL SFILL59160x59050 (
);

FILL FILL_2__10195_ (
);

FILL FILL_1__9651_ (
);

FILL FILL_1__9231_ (
);

FILL FILL_4__15807_ (
);

FILL FILL_3__9997_ (
);

FILL FILL_2__16001_ (
);

FILL FILL_4__10942_ (
);

FILL FILL_3__9157_ (
);

FILL FILL_4__10522_ (
);

FILL FILL_4__10102_ (
);

FILL FILL_1__15834_ (
);

FILL FILL_1__15414_ (
);

FILL FILL_6__7162_ (
);

FILL SFILL89800x53050 (
);

FILL FILL_0__14827_ (
);

FILL FILL_0__14407_ (
);

FILL FILL_2__7994_ (
);

BUFX2 BUFX2_insert630 (
    .A(_3977_),
    .Y(_3977__bF$buf1)
);

FILL FILL_2__7574_ (
);

BUFX2 BUFX2_insert631 (
    .A(_3977_),
    .Y(_3977__bF$buf0)
);

BUFX2 BUFX2_insert632 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf4 )
);

BUFX2 BUFX2_insert633 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf3 )
);

BUFX2 BUFX2_insert634 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf2 )
);

FILL FILL_6__13741_ (
);

BUFX2 BUFX2_insert635 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf1 )
);

FILL FILL_6__13321_ (
);

BUFX2 BUFX2_insert636 (
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf0 )
);

BUFX2 BUFX2_insert637 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf4 )
);

BUFX2 BUFX2_insert638 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf3 )
);

FILL SFILL49640x64050 (
);

BUFX2 BUFX2_insert639 (
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf2 )
);

FILL FILL_5__12734_ (
);

FILL FILL_5__12314_ (
);

FILL SFILL28760x23050 (
);

FILL SFILL59160x14050 (
);

FILL FILL_4__8861_ (
);

FILL FILL_4__8441_ (
);

FILL FILL_4__8021_ (
);

FILL FILL_4__11727_ (
);

FILL FILL_2__12761_ (
);

FILL FILL_4__11307_ (
);

FILL FILL_2__12341_ (
);

OAI21X1 _9086_ (
    .A(_1111_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .C(_1112_),
    .Y(_1108_[2])
);

FILL FILL_1__11754_ (
);

FILL FILL_4__14199_ (
);

FILL FILL_1__11334_ (
);

FILL FILL_2__8779_ (
);

FILL FILL_0__8761_ (
);

FILL FILL_2__8359_ (
);

FILL FILL_0__10747_ (
);

FILL FILL_0__8341_ (
);

FILL SFILL89320x46050 (
);

DFFSR _10612_ (
    .Q(\datapath_1.regfile_1.regOut[29] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_1823_[30])
);

FILL FILL_4__15980_ (
);

FILL FILL_4__15560_ (
);

FILL FILL_4__15140_ (
);

OAI21X1 _13084_ (
    .A(_3686_),
    .B(PCEn_bF$buf3),
    .C(_3687_),
    .Y(_3685_[1])
);

FILL FILL_5__13939_ (
);

FILL FILL_2__9720_ (
);

FILL FILL_3__14973_ (
);

FILL FILL_5__13519_ (
);

FILL FILL_3__14553_ (
);

FILL FILL_2__9300_ (
);

INVX1 _7819_ (
    .A(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_471_)
);

FILL FILL_3__14133_ (
);

FILL FILL_4_BUFX2_insert470 (
);

FILL FILL_4_BUFX2_insert471 (
);

FILL FILL_4__9646_ (
);

FILL FILL_4__9226_ (
);

FILL FILL_4_BUFX2_insert472 (
);

FILL FILL_4_BUFX2_insert473 (
);

FILL FILL_2__13966_ (
);

FILL FILL_4_BUFX2_insert474 (
);

FILL FILL_2__13546_ (
);

FILL FILL_0__14580_ (
);

FILL FILL_2__13126_ (
);

FILL FILL_4_BUFX2_insert475 (
);

FILL FILL_0__14160_ (
);

FILL FILL_4_BUFX2_insert476 (
);

FILL FILL_4_BUFX2_insert477 (
);

FILL FILL_4_BUFX2_insert478 (
);

FILL FILL_4_BUFX2_insert479 (
);

FILL FILL_1__12959_ (
);

FILL FILL_1__12119_ (
);

FILL FILL_0__9546_ (
);

FILL FILL_3__7223_ (
);

FILL FILL_0__9126_ (
);

AOI21X1 _11817_ (
    .A(_2124_),
    .B(_2907_),
    .C(_2458_),
    .Y(_2908_)
);

FILL SFILL33960x41050 (
);

FILL FILL_5__7989_ (
);

FILL FILL_5__7569_ (
);

FILL FILL_1__13900_ (
);

FILL FILL_4__16345_ (
);

AOI22X1 _14289_ (
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .B(_4102_),
    .C(_3995__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_4784_)
);

FILL FILL_6__10026_ (
);

FILL FILL_4__11480_ (
);

FILL FILL_4__11060_ (
);

FILL FILL_3__15758_ (
);

FILL FILL_3__15338_ (
);

FILL FILL_1__16372_ (
);

FILL FILL_3__10893_ (
);

FILL FILL_5__8510_ (
);

FILL FILL_3__10053_ (
);

FILL SFILL18760x21050 (
);

FILL FILL_0__15785_ (
);

FILL FILL_0__15365_ (
);

NOR3X1 _15650_ (
    .A(_6107_),
    .B(_6096_),
    .C(_6115_),
    .Y(_6116_)
);

NOR2X1 _15230_ (
    .A(_5705_),
    .B(_5695_),
    .Y(_5706_)
);

FILL FILL_5__10800_ (
);

FILL FILL_1__8502_ (
);

FILL FILL_3__8848_ (
);

FILL FILL_3__8008_ (
);

FILL FILL_5__13692_ (
);

FILL FILL_5__13272_ (
);

FILL FILL_6__6853_ (
);

INVX1 _7992_ (
    .A(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_566_)
);

INVX1 _7572_ (
    .A(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_347_)
);

DFFSR _7152_ (
    .Q(\datapath_1.regfile_1.regOut[2] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_68_[26])
);

FILL SFILL79320x44050 (
);

FILL SFILL18680x28050 (
);

FILL SFILL99240x50 (
);

FILL FILL_4__12265_ (
);

FILL FILL_2__6845_ (
);

FILL FILL_3__11678_ (
);

FILL FILL111960x57050 (
);

FILL FILL_3__11258_ (
);

FILL FILL_1__12292_ (
);

DFFSR _16435_ (
    .Q(\datapath_1.regfile_1.regOut[0] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_6769_[18])
);

INVX1 _16015_ (
    .A(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_6471_)
);

NAND3X1 _11990_ (
    .A(_3033_),
    .B(_3035_),
    .C(_3038_),
    .Y(\datapath_1.mux_pcsrc.dout [0])
);

INVX1 _11570_ (
    .A(_2677_),
    .Y(_2678_)
);

FILL FILL_0__11285_ (
);

OAI21X1 _11150_ (
    .A(_2266_),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .C(_2268_),
    .Y(_2269_)
);

FILL FILL_4__7712_ (
);

FILL FILL_3_BUFX2_insert490 (
);

FILL FILL_3_BUFX2_insert491 (
);

FILL FILL_3_BUFX2_insert492 (
);

FILL FILL_5__14897_ (
);

FILL FILL_5__14477_ (
);

FILL FILL_3_BUFX2_insert493 (
);

FILL FILL_2__11612_ (
);

FILL FILL_5__14057_ (
);

FILL FILL_3_BUFX2_insert494 (
);

FILL FILL_3__15091_ (
);

OAI21X1 _8777_ (
    .A(_966_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .C(_967_),
    .Y(_913_[27])
);

FILL FILL_3_BUFX2_insert495 (
);

FILL FILL_3_BUFX2_insert496 (
);

OAI21X1 _8357_ (
    .A(_747_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_748_),
    .Y(_718_[15])
);

FILL FILL_6__7218_ (
);

FILL FILL_3_BUFX2_insert497 (
);

FILL FILL_3_BUFX2_insert498 (
);

FILL FILL_3_BUFX2_insert499 (
);

FILL SFILL39560x24050 (
);

FILL FILL_2__14084_ (
);

FILL FILL_0__7612_ (
);

FILL SFILL94440x6050 (
);

FILL FILL_1__13497_ (
);

FILL FILL_4__14831_ (
);

FILL FILL_4__14411_ (
);

FILL FILL111960x12050 (
);

OAI21X1 _12775_ (
    .A(_3541_),
    .B(IRWrite_bF$buf4),
    .C(_3542_),
    .Y(_3490_[26])
);

INVX1 _12355_ (
    .A(ALUOut[4]),
    .Y(_3302_)
);

FILL FILL_3__13824_ (
);

FILL FILL_3__13404_ (
);

FILL FILL_4__8917_ (
);

FILL FILL_0__13851_ (
);

FILL FILL_0__13431_ (
);

FILL FILL_3__16296_ (
);

FILL FILL_0__13011_ (
);

FILL FILL_5__10397_ (
);

FILL FILL_1__8099_ (
);

FILL SFILL104600x9050 (
);

FILL FILL_2__15289_ (
);

FILL SFILL69320x42050 (
);

FILL FILL_3__6914_ (
);

FILL FILL_5__16203_ (
);

FILL FILL_1__9880_ (
);

FILL FILL_1__9040_ (
);

FILL FILL_4__15616_ (
);

FILL FILL_2__16230_ (
);

FILL FILL_3__9386_ (
);

FILL FILL_4__10751_ (
);

FILL FILL_3__14609_ (
);

FILL FILL_1__15643_ (
);

FILL FILL_1__15223_ (
);

FILL SFILL69240x49050 (
);

FILL FILL_0__14636_ (
);

INVX1 _14921_ (
    .A(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_5403_)
);

FILL FILL_0__14216_ (
);

INVX1 _14501_ (
    .A(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_4991_)
);

FILL FILL_6__13130_ (
);

FILL FILL_5__12963_ (
);

FILL FILL_5__12123_ (
);

BUFX2 _6843_ (
    .A(_1_[5]),
    .Y(memoryAddress[5])
);

FILL FILL_4__8250_ (
);

FILL FILL_4__11956_ (
);

FILL FILL_2__12990_ (
);

FILL FILL_4__11536_ (
);

FILL FILL_2__12570_ (
);

FILL FILL_4__11116_ (
);

FILL FILL_2__12150_ (
);

FILL FILL_1__16008_ (
);

FILL FILL_3__10949_ (
);

FILL FILL_1__11983_ (
);

FILL FILL_3__10529_ (
);

FILL FILL_1__11563_ (
);

FILL FILL_3__10109_ (
);

FILL FILL_1__11143_ (
);

FILL SFILL59720x54050 (
);

NOR2X1 _15706_ (
    .A(_6161_),
    .B(_6169_),
    .Y(_6170_)
);

FILL FILL_0__8990_ (
);

FILL FILL_2__8588_ (
);

FILL FILL_0__10976_ (
);

FILL FILL_0__8570_ (
);

DFFSR _10841_ (
    .Q(\datapath_1.regfile_1.regOut[31] [3]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_1953_[3])
);

FILL FILL_0__10556_ (
);

INVX1 _10421_ (
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .Y(_1799_)
);

FILL FILL_0__10136_ (
);

INVX1 _10001_ (
    .A(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_1580_)
);

FILL FILL_5__13748_ (
);

FILL FILL_5__13328_ (
);

FILL FILL_3__14782_ (
);

FILL FILL_3__14362_ (
);

FILL FILL_6__6909_ (
);

OAI21X1 _7628_ (
    .A(_383_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .C(_384_),
    .Y(_328_[28])
);

OAI21X1 _7208_ (
    .A(_164_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .C(_165_),
    .Y(_133_[16])
);

FILL FILL_4__9875_ (
);

FILL FILL_4__9035_ (
);

FILL FILL_2__13775_ (
);

FILL FILL_2__13355_ (
);

FILL FILL_1__12768_ (
);

FILL FILL_1__12348_ (
);

FILL FILL_3__7872_ (
);

FILL FILL_0__9775_ (
);

FILL FILL_0__9355_ (
);

FILL FILL_3__7452_ (
);

FILL FILL112440x80050 (
);

FILL FILL_3__7032_ (
);

NAND3X1 _11626_ (
    .A(_2268_),
    .B(_2462__bF$buf0),
    .C(_2688_),
    .Y(_2731_)
);

OAI21X1 _11206_ (
    .A(_2319_),
    .B(_2320_),
    .C(_2324_),
    .Y(_2325_)
);

FILL FILL_5__7798_ (
);

FILL FILL_5__7378_ (
);

FILL FILL_4__16154_ (
);

FILL SFILL64440x5050 (
);

AOI22X1 _14098_ (
    .A(_4051__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [13]),
    .C(\datapath_1.regfile_1.regOut[25] [13]),
    .D(_4040_),
    .Y(_4597_)
);

FILL FILL_3__15987_ (
);

FILL FILL_0__12702_ (
);

FILL FILL_3__15567_ (
);

FILL FILL_3__15147_ (
);

FILL FILL_1__16181_ (
);

FILL FILL_3__10282_ (
);

FILL FILL_0__15594_ (
);

FILL FILL_0__15174_ (
);

FILL FILL_1__8731_ (
);

FILL FILL_1__8311_ (
);

FILL FILL_2__15921_ (
);

FILL FILL_2__15501_ (
);

FILL FILL_3__8657_ (
);

FILL FILL_3__8237_ (
);

FILL FILL_5__13081_ (
);

FILL FILL_1__14914_ (
);

FILL SFILL12760x64050 (
);

OAI21X1 _7381_ (
    .A(_259_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .C(_260_),
    .Y(_198_[31])
);

FILL FILL_4__12494_ (
);

FILL FILL_4__12074_ (
);

FILL FILL_0__13907_ (
);

FILL FILL_5__9524_ (
);

FILL FILL_3__11487_ (
);

FILL FILL_5__9104_ (
);

FILL FILL_3__11067_ (
);

FILL FILL_0__16379_ (
);

AOI21X1 _16244_ (
    .A(_6671_),
    .B(_6694_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [29])
);

FILL FILL_0__11094_ (
);

FILL SFILL89400x34050 (
);

FILL FILL_1__9936_ (
);

FILL FILL_5__11814_ (
);

FILL SFILL28760x18050 (
);

FILL FILL_1__9516_ (
);

FILL FILL_4__7941_ (
);

FILL SFILL113800x2050 (
);

FILL FILL_4__7101_ (
);

FILL FILL_4__10807_ (
);

FILL FILL_2__11841_ (
);

FILL FILL_5__14286_ (
);

FILL FILL_2__11421_ (
);

FILL FILL_2__11001_ (
);

OAI21X1 _8586_ (
    .A(_859_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_860_),
    .Y(_848_[6])
);

DFFSR _8166_ (
    .Q(\datapath_1.regfile_1.regOut[10] [16]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_588_[16])
);

FILL SFILL49240x45050 (
);

FILL FILL_1__10834_ (
);

FILL FILL_4__13699_ (
);

FILL SFILL89000x20050 (
);

FILL FILL_4__13279_ (
);

FILL FILL_1__10414_ (
);

FILL FILL_0__7841_ (
);

FILL FILL_2__7859_ (
);

FILL FILL_2__7439_ (
);

FILL FILL_0__7421_ (
);

FILL FILL_4__14640_ (
);

FILL FILL_4__14220_ (
);

OAI21X1 _12584_ (
    .A(_3434_),
    .B(vdd),
    .C(_3435_),
    .Y(_3425_[5])
);

FILL FILL_0__12299_ (
);

NAND2X1 _12164_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.a [16]),
    .Y(_3163_)
);

FILL FILL_3__13633_ (
);

FILL FILL_3__13213_ (
);

FILL FILL_6__16078_ (
);

FILL FILL_4__8726_ (
);

FILL SFILL94280x40050 (
);

FILL FILL_2__12626_ (
);

FILL FILL_0__13660_ (
);

FILL FILL_2__12206_ (
);

FILL FILL_0__13240_ (
);

FILL FILL_1__11619_ (
);

FILL FILL_2__15098_ (
);

FILL FILL_5__16012_ (
);

FILL FILL_0__8626_ (
);

FILL FILL_0__8206_ (
);

FILL SFILL33960x36050 (
);

FILL FILL_4__15845_ (
);

FILL FILL_4__15425_ (
);

FILL FILL_4__15005_ (
);

FILL FILL_4__10980_ (
);

AOI21X1 _13789_ (
    .A(_4267_),
    .B(_4294_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [6])
);

FILL FILL_4__10560_ (
);

NAND3X1 _13369_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3880_),
    .C(_3879_),
    .Y(_3881_)
);

FILL FILL_4__10140_ (
);

FILL FILL_3__14838_ (
);

FILL FILL_3__14418_ (
);

FILL FILL_1__15872_ (
);

FILL FILL_1__15452_ (
);

FILL FILL_1__15032_ (
);

FILL SFILL18760x16050 (
);

FILL SFILL84280x83050 (
);

FILL SFILL33560x22050 (
);

FILL FILL_0__14865_ (
);

NAND2X1 _14730_ (
    .A(_5215_),
    .B(_5208_),
    .Y(_5216_)
);

FILL FILL_0__14445_ (
);

FILL FILL_0__14025_ (
);

NAND3X1 _14310_ (
    .A(_4801_),
    .B(_4804_),
    .C(_4800_),
    .Y(_4805_)
);

FILL FILL_2__7192_ (
);

CLKBUF1 CLKBUF1_insert170 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert171 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert172 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert173 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf51)
);

FILL FILL_3__7928_ (
);

FILL FILL_3__7508_ (
);

CLKBUF1 CLKBUF1_insert174 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert175 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf49)
);

FILL FILL_5__12772_ (
);

CLKBUF1 CLKBUF1_insert176 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf48)
);

FILL FILL_5__12352_ (
);

CLKBUF1 CLKBUF1_insert177 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert178 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf46)
);

FILL SFILL33800x1050 (
);

CLKBUF1 CLKBUF1_insert179 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf45)
);

FILL FILL_4__11765_ (
);

FILL FILL_4__11345_ (
);

FILL SFILL74280x1050 (
);

FILL FILL_1__16237_ (
);

FILL FILL_3__10758_ (
);

FILL FILL_1__11792_ (
);

FILL SFILL84200x81050 (
);

FILL FILL_1__11372_ (
);

AOI22X1 _15935_ (
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .B(_5577_),
    .C(_5479_),
    .D(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_6393_)
);

INVX1 _15515_ (
    .A(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_5984_)
);

FILL FILL_2__8397_ (
);

FILL FILL_0__10785_ (
);

INVX1 _10650_ (
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_1911_)
);

FILL FILL_0__10365_ (
);

INVX1 _10230_ (
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_1756_)
);

FILL FILL_6__14984_ (
);

FILL FILL_6__14564_ (
);

FILL FILL_5__13977_ (
);

FILL FILL_5__13557_ (
);

FILL FILL_3__14591_ (
);

FILL FILL_5__13137_ (
);

FILL FILL_3__14171_ (
);

OAI21X1 _7857_ (
    .A(_495_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_496_),
    .Y(_458_[19])
);

OAI21X1 _7437_ (
    .A(_276_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_277_),
    .Y(_263_[7])
);

DFFSR _7017_ (
    .Q(\datapath_1.regfile_1.regOut[1] [19]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_3_[19])
);

FILL FILL_4_BUFX2_insert850 (
);

FILL FILL_4_BUFX2_insert851 (
);

FILL FILL_4__9684_ (
);

FILL FILL_4_BUFX2_insert852 (
);

FILL FILL_4__9264_ (
);

FILL FILL_4_BUFX2_insert853 (
);

FILL FILL_4_BUFX2_insert854 (
);

FILL FILL_2__13584_ (
);

FILL SFILL114440x64050 (
);

FILL FILL_2__13164_ (
);

FILL FILL_4_BUFX2_insert855 (
);

FILL FILL_4_BUFX2_insert856 (
);

FILL FILL_4_BUFX2_insert857 (
);

FILL FILL_4_BUFX2_insert858 (
);

FILL FILL_4_BUFX2_insert859 (
);

FILL FILL_1__12997_ (
);

FILL FILL_1__12577_ (
);

FILL FILL_1__12157_ (
);

FILL FILL_4__13911_ (
);

FILL FILL_3__7681_ (
);

FILL SFILL74280x81050 (
);

FILL FILL_0__9164_ (
);

NAND3X1 _11855_ (
    .A(_2799_),
    .B(_2941_),
    .C(_2733_),
    .Y(_2942_)
);

NOR2X1 _11435_ (
    .A(_2550_),
    .B(_2413_),
    .Y(_2551_)
);

AOI22X1 _11015_ (
    .A(_2133_),
    .B(_2132_),
    .C(_2122_),
    .D(_2123_),
    .Y(_2134_)
);

FILL FILL_3__12904_ (
);

FILL FILL_4__16383_ (
);

FILL FILL_5__7187_ (
);

FILL FILL_3__15796_ (
);

FILL FILL_3__15376_ (
);

FILL FILL_0__12511_ (
);

FILL FILL_1__7599_ (
);

FILL FILL_1__7179_ (
);

FILL FILL_2__14789_ (
);

FILL FILL_2__14369_ (
);

FILL FILL_5__15703_ (
);

FILL FILL_1__8960_ (
);

FILL FILL_1__8120_ (
);

FILL FILL_2__15730_ (
);

FILL FILL_3__8886_ (
);

FILL FILL_2__15310_ (
);

FILL FILL_3__8466_ (
);

FILL FILL_1__14723_ (
);

FILL FILL_1__14303_ (
);

OAI21X1 _7190_ (
    .A(_152_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_153_),
    .Y(_133_[10])
);

FILL FILL_0__13716_ (
);

FILL FILL_2__6883_ (
);

FILL FILL_5__9753_ (
);

FILL FILL_3__11296_ (
);

FILL FILL_0__16188_ (
);

NOR3X1 _16053_ (
    .A(_6503_),
    .B(_6505_),
    .C(_6507_),
    .Y(_6508_)
);

FILL FILL_2__10289_ (
);

FILL FILL_1__9745_ (
);

FILL FILL_5__11623_ (
);

FILL FILL_5__11203_ (
);

FILL FILL_3_BUFX2_insert870 (
);

FILL FILL_4__7750_ (
);

FILL FILL_4__7330_ (
);

FILL FILL_3_BUFX2_insert871 (
);

FILL FILL_4__10616_ (
);

FILL FILL_3_BUFX2_insert872 (
);

FILL FILL_3_BUFX2_insert873 (
);

FILL FILL_2__11650_ (
);

FILL FILL_3_BUFX2_insert874 (
);

FILL FILL_2__11230_ (
);

FILL FILL_5__14095_ (
);

FILL FILL_1__15928_ (
);

FILL FILL_3_BUFX2_insert875 (
);

NAND2X1 _8395_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_774_)
);

FILL FILL_1__15508_ (
);

FILL FILL_3_BUFX2_insert876 (
);

FILL FILL_3_BUFX2_insert877 (
);

FILL FILL_3_BUFX2_insert878 (
);

FILL FILL_3_BUFX2_insert879 (
);

FILL FILL_1__10643_ (
);

FILL FILL_4__13088_ (
);

FILL SFILL104360x69050 (
);

FILL FILL_0__7230_ (
);

FILL FILL_2__7248_ (
);

FILL SFILL43880x8050 (
);

OAI21X1 _12393_ (
    .A(_3326_),
    .B(MemToReg_bF$buf5),
    .C(_3327_),
    .Y(\datapath_1.mux_wd3.dout [16])
);

FILL FILL_5__12828_ (
);

FILL FILL_5__12408_ (
);

FILL FILL_3__13862_ (
);

FILL FILL_3__13442_ (
);

FILL FILL_3__13022_ (
);

FILL FILL_4__8955_ (
);

FILL SFILL8600x8050 (
);

FILL FILL_4__8115_ (
);

FILL FILL_2__12855_ (
);

FILL FILL_2__12435_ (
);

FILL FILL_2__12015_ (
);

FILL FILL_1__11848_ (
);

FILL FILL_1__11428_ (
);

FILL FILL_1__11008_ (
);

FILL FILL_3__6952_ (
);

FILL FILL_5__16241_ (
);

FILL FILL_0__8855_ (
);

FILL FILL112440x75050 (
);

FILL FILL_0__8015_ (
);

OAI21X1 _10706_ (
    .A(_1947_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .C(_1948_),
    .Y(_1888_[30])
);

FILL FILL_5__6878_ (
);

FILL SFILL104360x24050 (
);

FILL FILL_4__15654_ (
);

FILL FILL_4__15234_ (
);

OAI22X1 _13598_ (
    .A(_4106_),
    .B(_3936__bF$buf2),
    .C(_3966__bF$buf3),
    .D(_4105_),
    .Y(_4107_)
);

DFFSR _13178_ (
    .Q(\datapath_1.mux_iord.din0 [3]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3685_[3])
);

FILL FILL_3__14647_ (
);

FILL FILL_1__15681_ (
);

FILL FILL_3__14227_ (
);

FILL FILL_1__15261_ (
);

FILL FILL112040x61050 (
);

FILL FILL_0__14674_ (
);

FILL FILL_0__14254_ (
);

FILL FILL_1__7811_ (
);

FILL FILL_3__7737_ (
);

FILL FILL_3__7317_ (
);

FILL FILL_5__12581_ (
);

FILL FILL_5__12161_ (
);

BUFX2 _6881_ (
    .A(_2_[11]),
    .Y(memoryWriteData[11])
);

FILL FILL112440x30050 (
);

FILL FILL_4__16019_ (
);

FILL FILL_4__11994_ (
);

FILL FILL_4__11574_ (
);

FILL FILL_4__11154_ (
);

FILL FILL_1__16046_ (
);

FILL FILL_5__8604_ (
);

FILL FILL_3__10567_ (
);

FILL FILL_3__10147_ (
);

FILL FILL_6_BUFX2_insert382 (
);

FILL FILL_1__11181_ (
);

FILL FILL_6__11901_ (
);

FILL FILL_0__15879_ (
);

AOI22X1 _15744_ (
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .B(_5579_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_6207_)
);

FILL FILL_0__15459_ (
);

NAND3X1 _15324_ (
    .A(_5786_),
    .B(_5792_),
    .C(_5797_),
    .Y(_5798_)
);

FILL FILL_0__15039_ (
);

FILL FILL_6_BUFX2_insert388 (
);

FILL FILL_0__10174_ (
);

FILL FILL_0__16400_ (
);

FILL FILL_2__10921_ (
);

FILL FILL_5__13786_ (
);

FILL FILL_5__13366_ (
);

FILL FILL_2__10501_ (
);

DFFSR _7666_ (
    .Q(\datapath_1.regfile_1.regOut[6] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_328_[28])
);

FILL SFILL33640x55050 (
);

NAND2X1 _7246_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_191_)
);

FILL FILL_4__9493_ (
);

FILL FILL_4__12779_ (
);

FILL FILL_4__12359_ (
);

FILL FILL_2__13393_ (
);

FILL FILL_0__6921_ (
);

FILL FILL_2__6939_ (
);

FILL FILL_5__9809_ (
);

FILL FILL_1__12386_ (
);

FILL FILL_4__13720_ (
);

FILL FILL_4__13300_ (
);

OAI22X1 _16109_ (
    .A(_6561_),
    .B(_5545__bF$buf2),
    .C(_5485__bF$buf1),
    .D(_6562_),
    .Y(_6563_)
);

FILL FILL_0__9393_ (
);

FILL FILL_0__11799_ (
);

FILL FILL_3__7490_ (
);

FILL FILL_0__11379_ (
);

FILL FILL_3__7070_ (
);

NOR2X1 _11664_ (
    .A(_2752_),
    .B(_2765_),
    .Y(_2766_)
);

NAND2X1 _11244_ (
    .A(_2362_),
    .B(_2360_),
    .Y(_2363_)
);

FILL FILL_3__12713_ (
);

FILL FILL_6__15158_ (
);

FILL FILL_4__16192_ (
);

FILL FILL_4__7806_ (
);

FILL SFILL94280x35050 (
);

FILL FILL_2__11706_ (
);

FILL FILL_0__12740_ (
);

FILL FILL_3__15185_ (
);

FILL FILL_0__12320_ (
);

FILL SFILL79000x58050 (
);

FILL SFILL13880x7050 (
);

FILL FILL_2__14598_ (
);

FILL FILL_2__14178_ (
);

FILL FILL_5__15932_ (
);

FILL FILL_5__15512_ (
);

FILL FILL_0__7706_ (
);

NAND2X1 _9812_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1495_)
);

FILL FILL_4__14925_ (
);

FILL FILL_4__14505_ (
);

FILL FILL_3__8695_ (
);

NAND2X1 _12869_ (
    .A(vdd),
    .B(\datapath_1.rd1 [15]),
    .Y(_3585_)
);

FILL FILL_3__8275_ (
);

NAND2X1 _12449_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [3]),
    .Y(_3366_)
);

AOI22X1 _12029_ (
    .A(\datapath_1.ALUResult [10]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3068_)
);

FILL FILL_3__13918_ (
);

FILL FILL_1__14952_ (
);

FILL FILL_1__14532_ (
);

FILL FILL_1__14112_ (
);

FILL SFILL79400x27050 (
);

FILL SFILL84280x78050 (
);

FILL FILL_6__11078_ (
);

FILL FILL_0__13945_ (
);

OAI22X1 _13810_ (
    .A(_4313_),
    .B(_3944__bF$buf3),
    .C(_3959_),
    .D(_4314_),
    .Y(_4315_)
);

FILL FILL_0__13525_ (
);

FILL FILL_0__13105_ (
);

FILL FILL_5__9982_ (
);

FILL FILL_5__9142_ (
);

NOR2X1 _16282_ (
    .A(_6717_),
    .B(_6731_),
    .Y(_6732_)
);

FILL SFILL79000x13050 (
);

FILL FILL_1__9974_ (
);

FILL FILL_5__11852_ (
);

FILL FILL_1__9554_ (
);

FILL FILL_5__11432_ (
);

FILL FILL_1__9134_ (
);

FILL FILL_5__11012_ (
);

FILL SFILL8680x52050 (
);

FILL FILL_2__16324_ (
);

FILL FILL_4__10425_ (
);

FILL FILL_4__10005_ (
);

FILL FILL_1__15737_ (
);

FILL FILL_1__15317_ (
);

FILL SFILL84200x76050 (
);

FILL FILL_1__10872_ (
);

FILL FILL_1__10452_ (
);

FILL FILL_1__10032_ (
);

FILL SFILL84280x33050 (
);

FILL FILL_2__7477_ (
);

FILL FILL_2__7057_ (
);

FILL FILL_6__13224_ (
);

FILL SFILL109480x76050 (
);

FILL FILL_5__12637_ (
);

FILL FILL_3__13671_ (
);

FILL FILL_5__12217_ (
);

FILL FILL_3__13251_ (
);

OAI21X1 _6937_ (
    .A(_24_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_25_),
    .Y(_3_[11])
);

FILL FILL_4__8764_ (
);

FILL FILL_4__8344_ (
);

FILL FILL_2__12244_ (
);

FILL FILL_1__11657_ (
);

FILL FILL_1__11237_ (
);

FILL SFILL84200x31050 (
);

FILL FILL_5__16050_ (
);

NOR2X1 _10935_ (
    .A(_2065_),
    .B(_2068_),
    .Y(_2069_)
);

FILL FILL_0__8244_ (
);

OAI21X1 _10515_ (
    .A(_1840_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1841_),
    .Y(_1823_[9])
);

FILL FILL_4__15883_ (
);

FILL FILL_4__15463_ (
);

FILL FILL_4__15043_ (
);

FILL SFILL13640x51050 (
);

FILL FILL_3__14876_ (
);

FILL FILL_2__9623_ (
);

FILL FILL_3__14456_ (
);

FILL FILL_3__14036_ (
);

FILL FILL_1__15490_ (
);

FILL FILL_1__15070_ (
);

FILL FILL_4__9549_ (
);

FILL FILL_4__9129_ (
);

FILL FILL_2__13869_ (
);

FILL FILL_2__13449_ (
);

FILL FILL_0__14483_ (
);

FILL FILL_2__13029_ (
);

FILL FILL_0__14063_ (
);

FILL FILL_1__7620_ (
);

FILL FILL_1__7200_ (
);

FILL FILL_2__14810_ (
);

FILL FILL_0__9869_ (
);

FILL FILL_3__7966_ (
);

FILL SFILL13560x58050 (
);

FILL FILL_3__7546_ (
);

FILL FILL_0__9029_ (
);

FILL FILL_5__12390_ (
);

FILL FILL_1__13803_ (
);

FILL FILL_4__16248_ (
);

FILL FILL_4__11383_ (
);

FILL FILL_1__16275_ (
);

FILL SFILL99480x80050 (
);

FILL FILL_5__8833_ (
);

FILL FILL_3__10796_ (
);

FILL FILL_3__10376_ (
);

INVX1 _15973_ (
    .A(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_6430_)
);

FILL FILL_0__15688_ (
);

INVX1 _15553_ (
    .A(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_6021_)
);

FILL FILL_0__15268_ (
);

INVX1 _15133_ (
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_5611_)
);

FILL FILL_5__10703_ (
);

FILL FILL_1__8825_ (
);

FILL FILL_1__8405_ (
);

FILL FILL_5__13595_ (
);

FILL FILL_2__10310_ (
);

DFFSR _7895_ (
    .Q(\datapath_1.regfile_1.regOut[8] [1]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_458_[1])
);

NAND2X1 _7475_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_303_)
);

NAND2X1 _7055_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_84_)
);

FILL FILL_4__12588_ (
);

FILL FILL_4__12168_ (
);

FILL FILL_5__9618_ (
);

FILL FILL_1__12195_ (
);

OAI21X1 _16338_ (
    .A(_6778_),
    .B(gnd),
    .C(_6779_),
    .Y(_6769_[5])
);

INVX1 _11893_ (
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_2970_)
);

FILL FILL_0__11188_ (
);

NAND3X1 _11473_ (
    .A(_2286_),
    .B(_2439_),
    .C(_2587_),
    .Y(_2588_)
);

FILL FILL_5__11908_ (
);

XOR2X1 _11053_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2172_)
);

FILL FILL_3__12522_ (
);

FILL FILL_3__12102_ (
);

FILL SFILL104440x12050 (
);

FILL FILL_4__7615_ (
);

FILL FILL_2__11935_ (
);

FILL FILL_2__11515_ (
);

FILL SFILL33800x81050 (
);

FILL FILL_1__10928_ (
);

FILL FILL_1__10508_ (
);

FILL FILL_5__15741_ (
);

FILL FILL_0__7935_ (
);

FILL FILL_5__15321_ (
);

NAND2X1 _9621_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1388_)
);

DFFSR _9201_ (
    .Q(\datapath_1.regfile_1.regOut[18] [27]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_1108_[27])
);

FILL SFILL104360x19050 (
);

FILL FILL_4__14734_ (
);

FILL FILL_4__14314_ (
);

DFFSR _12678_ (
    .Q(\datapath_1.Data [15]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3425_[15])
);

FILL FILL_3__8084_ (
);

NAND3X1 _12258_ (
    .A(_3230_),
    .B(_3231_),
    .C(_3232_),
    .Y(\datapath_1.alu_1.ALUInB [10])
);

FILL FILL_3__13727_ (
);

FILL FILL_3__13307_ (
);

FILL FILL_1__14761_ (
);

FILL FILL_1__14341_ (
);

FILL FILL112040x56050 (
);

FILL FILL_0__13754_ (
);

FILL FILL_0__13334_ (
);

FILL FILL_3__16199_ (
);

FILL FILL_5__9791_ (
);

FILL FILL_5__9371_ (
);

INVX1 _16091_ (
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_6545_)
);

FILL FILL_5__16106_ (
);

FILL FILL_1__9783_ (
);

FILL FILL_5__11661_ (
);

FILL FILL_5__11241_ (
);

FILL FILL_1__9363_ (
);

FILL FILL112440x25050 (
);

FILL FILL_4__15939_ (
);

FILL FILL_4__15519_ (
);

FILL FILL_2__16133_ (
);

FILL FILL_3__9289_ (
);

FILL FILL_4__10654_ (
);

FILL FILL_4__10234_ (
);

FILL FILL_1__15966_ (
);

FILL FILL_1__15546_ (
);

FILL FILL_1__15126_ (
);

FILL SFILL49320x28050 (
);

FILL FILL_1__10681_ (
);

FILL FILL_1__10261_ (
);

FILL FILL_0__14959_ (
);

FILL FILL112040x11050 (
);

AOI22X1 _14824_ (
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .B(_3942__bF$buf1),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_5308_)
);

FILL FILL_0__14539_ (
);

AOI22X1 _14404_ (
    .A(_3995__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [20]),
    .C(\datapath_1.regfile_1.regOut[6] [20]),
    .D(_4001__bF$buf3),
    .Y(_4896_)
);

FILL FILL_0__14119_ (
);

FILL FILL_2__7286_ (
);

FILL FILL_0__15900_ (
);

FILL FILL_5__12866_ (
);

FILL FILL_5__12446_ (
);

FILL FILL_5__12026_ (
);

FILL FILL_3__13480_ (
);

FILL FILL_4__8993_ (
);

FILL FILL_4__8573_ (
);

FILL FILL_4__11859_ (
);

FILL FILL_2__12893_ (
);

FILL FILL_4__11439_ (
);

FILL FILL_2__12473_ (
);

FILL FILL_4__11019_ (
);

FILL FILL_2__12053_ (
);

FILL FILL_1__11886_ (
);

FILL SFILL98600x74050 (
);

FILL FILL_1__11466_ (
);

FILL FILL_1__11046_ (
);

NOR3X1 _15609_ (
    .A(_6065_),
    .B(_6054_),
    .C(_6075_),
    .Y(_6076_)
);

FILL FILL_3__6990_ (
);

FILL FILL_0__8893_ (
);

FILL FILL_6__9860_ (
);

FILL FILL_0__8473_ (
);

FILL FILL_0__10879_ (
);

OAI21X1 _10744_ (
    .A(_2016_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_2017_),
    .Y(_1953_[0])
);

FILL FILL_0__10039_ (
);

NAND2X1 _10324_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1755_)
);

FILL FILL_4__15692_ (
);

FILL FILL_4__15272_ (
);

FILL SFILL23320x72050 (
);

FILL FILL_2__9852_ (
);

FILL FILL_0__11820_ (
);

FILL FILL_3__14685_ (
);

FILL FILL_3__14265_ (
);

FILL FILL_2__9012_ (
);

FILL FILL_0__11400_ (
);

FILL FILL_4__9778_ (
);

FILL FILL_4__9358_ (
);

FILL FILL_2__13678_ (
);

FILL FILL_2__13258_ (
);

FILL FILL_0__14292_ (
);

FILL SFILL23720x41050 (
);

FILL FILL_0__9678_ (
);

FILL FILL_3__7355_ (
);

OAI21X1 _11949_ (
    .A(_3006_),
    .B(IorD_bF$buf7),
    .C(_3007_),
    .Y(_1_[20])
);

FILL FILL_0__9258_ (
);

AOI22X1 _11529_ (
    .A(_2223_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf0),
    .D(_2224_),
    .Y(_2640_)
);

INVX1 _11109_ (
    .A(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2228_)
);

FILL FILL_1__13612_ (
);

FILL FILL_4__16057_ (
);

FILL FILL_4__11192_ (
);

FILL FILL_0__12605_ (
);

FILL FILL_1__16084_ (
);

FILL FILL_5__8642_ (
);

FILL FILL_6_BUFX2_insert761 (
);

FILL FILL_3__10185_ (
);

FILL FILL_5__8222_ (
);

INVX1 _15782_ (
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_6244_)
);

FILL FILL_0__15497_ (
);

NAND3X1 _15362_ (
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5835_)
);

FILL FILL_0__15077_ (
);

FILL FILL_6_BUFX2_insert766 (
);

FILL FILL_3__16411_ (
);

FILL FILL_5__10932_ (
);

FILL FILL_5__10512_ (
);

FILL FILL_1__8634_ (
);

FILL FILL_1__8214_ (
);

FILL SFILL8680x47050 (
);

FILL FILL_2__15824_ (
);

FILL FILL_2__15404_ (
);

FILL SFILL109560x64050 (
);

FILL FILL_1__14817_ (
);

DFFSR _7284_ (
    .Q(\datapath_1.regfile_1.regOut[3] [30]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_133_[30])
);

FILL FILL_4__12397_ (
);

FILL FILL_3__9921_ (
);

FILL FILL_3__9501_ (
);

FILL SFILL84280x28050 (
);

FILL FILL_2__6977_ (
);

FILL FILL_5__9847_ (
);

FILL FILL_5__9427_ (
);

FILL FILL_5__9007_ (
);

NOR2X1 _16147_ (
    .A(_6596_),
    .B(_6599_),
    .Y(_6600_)
);

INVX1 _11282_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .Y(_2401_)
);

FILL FILL_5__11717_ (
);

FILL FILL_3__12751_ (
);

FILL FILL_1__9419_ (
);

FILL SFILL8600x45050 (
);

FILL FILL_3__12331_ (
);

FILL FILL_4__7844_ (
);

FILL FILL_4__7424_ (
);

FILL FILL_2__11744_ (
);

FILL FILL_5__14189_ (
);

FILL FILL_2__11324_ (
);

INVX1 _8489_ (
    .A(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_816_)
);

INVX1 _8069_ (
    .A(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_597_)
);

FILL FILL_1__10317_ (
);

FILL SFILL84200x26050 (
);

FILL FILL_5__15970_ (
);

FILL FILL_5__15550_ (
);

FILL FILL_0__7744_ (
);

FILL FILL_5__15130_ (
);

FILL FILL_0__7324_ (
);

NAND2X1 _9850_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1500_)
);

DFFSR _9430_ (
    .Q(\datapath_1.regfile_1.regOut[20] [0]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1238_[0])
);

INVX1 _9010_ (
    .A(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_1082_)
);

FILL FILL_4__14963_ (
);

FILL FILL_4__14543_ (
);

FILL FILL_4__14123_ (
);

FILL SFILL13640x46050 (
);

INVX1 _12487_ (
    .A(ALUOut[16]),
    .Y(_3391_)
);

NAND3X1 _12067_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[20]),
    .C(_3032__bF$buf2),
    .Y(_3096_)
);

FILL FILL_2__8703_ (
);

FILL FILL_3__13956_ (
);

FILL FILL_1__14990_ (
);

FILL FILL_3__13536_ (
);

FILL FILL_1__14570_ (
);

FILL FILL_3__13116_ (
);

FILL FILL_1__14150_ (
);

FILL FILL_4__8629_ (
);

FILL FILL_5_BUFX2_insert780 (
);

FILL FILL_4__8209_ (
);

FILL FILL_5_BUFX2_insert781 (
);

FILL FILL_0__13983_ (
);

FILL FILL_2__12529_ (
);

FILL FILL_5_BUFX2_insert782 (
);

FILL FILL_2__12109_ (
);

FILL FILL_5_BUFX2_insert783 (
);

FILL FILL_0__13563_ (
);

FILL FILL_0__13143_ (
);

FILL FILL_5_BUFX2_insert784 (
);

FILL FILL_5_BUFX2_insert785 (
);

FILL FILL_5_BUFX2_insert786 (
);

FILL FILL_5_BUFX2_insert787 (
);

FILL FILL_5_BUFX2_insert788 (
);

FILL FILL_5_BUFX2_insert789 (
);

FILL SFILL74200x69050 (
);

FILL FILL_5__16335_ (
);

FILL FILL_6__9916_ (
);

FILL FILL_0__8529_ (
);

FILL FILL_0__8109_ (
);

FILL FILL_5__11890_ (
);

FILL FILL_1__9592_ (
);

FILL FILL_5__11470_ (
);

FILL SFILL74280x26050 (
);

FILL FILL_1__9172_ (
);

FILL FILL_5__11050_ (
);

FILL FILL_4__15748_ (
);

FILL FILL_4__15328_ (
);

FILL FILL_2__16362_ (
);

FILL FILL_3__9098_ (
);

FILL FILL_4__10883_ (
);

FILL FILL_4__10043_ (
);

FILL FILL_2__9908_ (
);

FILL FILL_1__15775_ (
);

FILL SFILL99480x75050 (
);

FILL FILL_1__15355_ (
);

FILL FILL_1__10490_ (
);

FILL FILL_0__14768_ (
);

OAI22X1 _14633_ (
    .A(_3967__bF$buf3),
    .B(_5119_),
    .C(_3966__bF$buf3),
    .D(_5120_),
    .Y(_5121_)
);

FILL FILL_0__14348_ (
);

AOI22X1 _14213_ (
    .A(_4038__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[23] [15]),
    .C(\datapath_1.regfile_1.regOut[27] [15]),
    .D(_4129_),
    .Y(_4710_)
);

FILL SFILL38840x50050 (
);

FILL FILL_2__7095_ (
);

FILL SFILL74200x24050 (
);

FILL FILL_5__12255_ (
);

NAND2X1 _6975_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_51_)
);

FILL FILL_4__8382_ (
);

FILL FILL_4__11668_ (
);

FILL FILL_4__11248_ (
);

FILL FILL_2__12282_ (
);

FILL FILL_1__11695_ (
);

FILL FILL_1__11275_ (
);

FILL SFILL99480x30050 (
);

OAI22X1 _15838_ (
    .A(_5485__bF$buf1),
    .B(_6298_),
    .C(_5483__bF$buf2),
    .D(_4869_),
    .Y(_6299_)
);

NOR3X1 _15418_ (
    .A(_5888_),
    .B(_5509_),
    .C(_5688_),
    .Y(_5889_)
);

FILL FILL_0__10688_ (
);

NAND2X1 _10973_ (
    .A(\control_1.next [0]),
    .B(vdd),
    .Y(_2100_)
);

NAND2X1 _10553_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1867_)
);

FILL FILL_0__10268_ (
);

NAND2X1 _10133_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1648_)
);

FILL FILL_6__14467_ (
);

FILL FILL_3__11602_ (
);

FILL FILL_6__14047_ (
);

FILL FILL_4__15081_ (
);

FILL SFILL33800x76050 (
);

FILL FILL_2__9661_ (
);

FILL SFILL64200x67050 (
);

FILL FILL_3__14494_ (
);

FILL FILL_2__9241_ (
);

FILL FILL_3__14074_ (
);

FILL FILL112120x44050 (
);

FILL FILL_4__9167_ (
);

FILL FILL_2__13487_ (
);

FILL FILL_5__14821_ (
);

FILL FILL_5__14401_ (
);

NAND2X1 _8701_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_917_)
);

FILL FILL_4__13814_ (
);

FILL SFILL89800x5050 (
);

FILL FILL_0__9487_ (
);

FILL FILL_3__7584_ (
);

NOR2X1 _11758_ (
    .A(_2156_),
    .B(_2852_),
    .Y(_2853_)
);

FILL FILL_3__7164_ (
);

OAI21X1 _11338_ (
    .A(_2456_),
    .B(_2115_),
    .C(_2350_),
    .Y(_2457_)
);

FILL FILL_1__13841_ (
);

FILL FILL_1__13421_ (
);

FILL FILL_4__16286_ (
);

FILL FILL_1__13001_ (
);

FILL FILL_3__15699_ (
);

FILL FILL_0__12834_ (
);

FILL FILL_0__12414_ (
);

FILL FILL_3__15279_ (
);

FILL FILL_5__8871_ (
);

FILL FILL_5__8451_ (
);

INVX1 _15591_ (
    .A(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_6058_)
);

NOR2X1 _15171_ (
    .A(_5646_),
    .B(_5647_),
    .Y(_5648_)
);

FILL FILL_5__15606_ (
);

FILL FILL_3__16220_ (
);

INVX1 _9906_ (
    .A(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_1537_)
);

FILL FILL_1__8863_ (
);

FILL FILL_1__8443_ (
);

FILL FILL_5__10321_ (
);

FILL FILL_2__15633_ (
);

FILL FILL_2__15213_ (
);

FILL FILL_3__8789_ (
);

FILL FILL_3__8369_ (
);

FILL FILL_1__14626_ (
);

INVX1 _7093_ (
    .A(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_109_)
);

FILL FILL_1__14206_ (
);

FILL FILL_3__9730_ (
);

FILL FILL_0__13619_ (
);

INVX1 _13904_ (
    .A(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_4407_)
);

FILL FILL_5__9656_ (
);

FILL FILL_3__11199_ (
);

FILL FILL_5__9236_ (
);

NAND2X1 _16376_ (
    .A(gnd),
    .B(gnd),
    .Y(_6805_)
);

FILL FILL_5__11946_ (
);

INVX1 _11091_ (
    .A(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2210_)
);

FILL FILL_1__9648_ (
);

FILL FILL_3__12980_ (
);

FILL FILL_5__11526_ (
);

FILL FILL_1__9228_ (
);

FILL FILL_5__11106_ (
);

FILL FILL_3__12140_ (
);

FILL FILL_4__10939_ (
);

FILL FILL_4__7233_ (
);

FILL FILL_2__11973_ (
);

FILL FILL_4__10519_ (
);

FILL FILL_2__11553_ (
);

FILL FILL_6__7999_ (
);

FILL FILL_2__11133_ (
);

DFFSR _8298_ (
    .Q(\datapath_1.regfile_1.regOut[11] [20]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_653_[20])
);

FILL FILL_1__10966_ (
);

FILL FILL_1__10546_ (
);

FILL FILL_1__10126_ (
);

FILL FILL_0__7973_ (
);

FILL FILL_0__7553_ (
);

FILL FILL_4__14772_ (
);

FILL FILL_4__14352_ (
);

FILL SFILL54200x20050 (
);

NAND3X1 _12296_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3198__bF$buf1),
    .Y(_3261_)
);

FILL FILL_0__10900_ (
);

FILL FILL_2__8512_ (
);

FILL FILL_3__13765_ (
);

FILL FILL_3__13345_ (
);

FILL FILL_4__8858_ (
);

FILL FILL_4__8438_ (
);

FILL FILL_4__8018_ (
);

FILL FILL_2__12758_ (
);

FILL FILL_0__13792_ (
);

FILL FILL_2__12338_ (
);

FILL FILL_0__13372_ (
);

FILL SFILL23720x36050 (
);

FILL FILL_0__8758_ (
);

FILL FILL_3__6855_ (
);

FILL FILL_5__16144_ (
);

FILL FILL_0__8338_ (
);

DFFSR _10609_ (
    .Q(\datapath_1.regfile_1.regOut[29] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1823_[27])
);

FILL FILL_4__15977_ (
);

FILL FILL_4__15557_ (
);

FILL FILL_4__15137_ (
);

FILL FILL_2__16171_ (
);

FILL FILL_4__10692_ (
);

FILL FILL_4__10272_ (
);

FILL FILL_1__15584_ (
);

FILL FILL_1__15164_ (
);

FILL FILL_5__7722_ (
);

FILL FILL_5__7302_ (
);

FILL FILL_0__14997_ (
);

FILL FILL_0__14577_ (
);

OAI22X1 _14862_ (
    .A(_5344_),
    .B(_3982__bF$buf3),
    .C(_3983__bF$buf4),
    .D(_5343_),
    .Y(_5345_)
);

FILL FILL_0__14157_ (
);

INVX1 _14442_ (
    .A(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_4934_)
);

FILL SFILL48520x71050 (
);

FILL SFILL99960x7050 (
);

NAND3X1 _14022_ (
    .A(_4521_),
    .B(_4522_),
    .C(_4520_),
    .Y(_4523_)
);

FILL FILL_3__15911_ (
);

FILL FILL_1__7714_ (
);

FILL FILL_2__14904_ (
);

FILL SFILL109560x59050 (
);

FILL FILL_5__12484_ (
);

FILL FILL_5__12064_ (
);

FILL SFILL99560x6050 (
);

FILL FILL_4__8191_ (
);

FILL FILL_4__11897_ (
);

FILL FILL_4__11477_ (
);

FILL FILL_4__11057_ (
);

FILL FILL_2__12091_ (
);

FILL FILL_1__16369_ (
);

FILL FILL_5__8507_ (
);

FILL FILL_1__11084_ (
);

FILL FILL_6__11804_ (
);

OAI22X1 _15647_ (
    .A(_5549__bF$buf4),
    .B(_4625_),
    .C(_5466__bF$buf3),
    .D(_4622_),
    .Y(_6113_)
);

OAI22X1 _15227_ (
    .A(_4167_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf0),
    .D(_4165_),
    .Y(_5703_)
);

FILL FILL_0__10497_ (
);

FILL FILL_0__8091_ (
);

NAND2X1 _10782_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1979_)
);

NAND2X1 _10362_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1760_)
);

FILL FILL_3__11831_ (
);

FILL FILL_3__11411_ (
);

FILL FILL_4__6924_ (
);

FILL FILL_0__16303_ (
);

FILL SFILL13720x34050 (
);

FILL FILL_2__9890_ (
);

FILL FILL_2__10824_ (
);

FILL FILL_5__13689_ (
);

FILL FILL_5__13269_ (
);

FILL FILL_2__10404_ (
);

FILL FILL_2__9470_ (
);

INVX1 _7989_ (
    .A(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_564_)
);

INVX1 _7569_ (
    .A(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_345_)
);

DFFSR _7149_ (
    .Q(\datapath_1.regfile_1.regOut[2] [23]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_68_[23])
);

FILL FILL_4__9396_ (
);

FILL SFILL109400x3050 (
);

FILL FILL_2__13296_ (
);

FILL SFILL38920x83050 (
);

FILL FILL_5__14630_ (
);

FILL FILL_5__14210_ (
);

DFFSR _8930_ (
    .Q(\datapath_1.regfile_1.regOut[16] [12]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_978_[12])
);

INVX1 _8510_ (
    .A(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_830_)
);

FILL FILL_1__12289_ (
);

FILL FILL_4__13623_ (
);

NOR2X1 _11987_ (
    .A(ALUOp_0_bF$buf1),
    .B(PCSource_1_bF$buf3),
    .Y(_3036_)
);

FILL FILL_0__9296_ (
);

OAI21X1 _11567_ (
    .A(_2661_),
    .B(_2662_),
    .C(_2675_),
    .Y(\datapath_1.ALUResult [21])
);

INVX1 _11147_ (
    .A(\datapath_1.alu_1.ALUInA [17]),
    .Y(_2266_)
);

FILL FILL_3__12616_ (
);

FILL FILL_3_BUFX2_insert20 (
);

FILL FILL_1__13650_ (
);

FILL FILL_3_BUFX2_insert21 (
);

FILL FILL_1__13230_ (
);

FILL FILL_4__16095_ (
);

FILL FILL_3_BUFX2_insert22 (
);

FILL FILL_3_BUFX2_insert23 (
);

FILL FILL_3_BUFX2_insert24 (
);

FILL FILL_4__7709_ (
);

FILL FILL_6__10196_ (
);

FILL FILL_3_BUFX2_insert25 (
);

FILL FILL_3_BUFX2_insert26 (
);

FILL FILL_3_BUFX2_insert27 (
);

FILL FILL_2__11609_ (
);

FILL FILL_0__12643_ (
);

FILL FILL_3_BUFX2_insert28 (
);

FILL FILL_3_BUFX2_insert29 (
);

FILL FILL_3__15088_ (
);

FILL FILL_0__12223_ (
);

FILL FILL_6__16002_ (
);

FILL FILL_5__8260_ (
);

FILL FILL_5__15835_ (
);

FILL FILL_5__15415_ (
);

FILL FILL_0__7609_ (
);

DFFSR _9715_ (
    .Q(\datapath_1.regfile_1.regOut[22] [29]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_1368_[29])
);

FILL FILL_5__10970_ (
);

FILL FILL_5__10550_ (
);

FILL FILL_1__8252_ (
);

FILL FILL_5__10130_ (
);

FILL FILL_4__14828_ (
);

FILL FILL_4__14408_ (
);

FILL FILL_2__15862_ (
);

FILL FILL_2__15442_ (
);

FILL FILL_2__15022_ (
);

FILL FILL_3__8598_ (
);

FILL FILL_1__14855_ (
);

FILL FILL_1__14435_ (
);

FILL FILL_1__14015_ (
);

FILL SFILL38040x62050 (
);

FILL FILL_0__13848_ (
);

FILL FILL_0__13428_ (
);

NAND2X1 _13713_ (
    .A(_4212_),
    .B(_4219_),
    .Y(_4220_)
);

FILL FILL_0__13008_ (
);

FILL FILL_5__9885_ (
);

FILL FILL_5__9465_ (
);

FILL FILL_5__9045_ (
);

NAND3X1 _16185_ (
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf0),
    .Y(_6637_)
);

FILL SFILL28920x81050 (
);

FILL SFILL74200x19050 (
);

FILL FILL_5__11755_ (
);

FILL FILL_1__9877_ (
);

FILL FILL_5__11335_ (
);

FILL FILL_1__9037_ (
);

FILL FILL_2__16227_ (
);

FILL FILL_4__7882_ (
);

FILL FILL_4__7462_ (
);

FILL FILL_4__7042_ (
);

FILL FILL_4__10748_ (
);

FILL FILL_2__11782_ (
);

FILL FILL_2__11362_ (
);

FILL FILL112200x32050 (
);

FILL FILL_1__10775_ (
);

FILL SFILL99480x25050 (
);

INVX1 _14918_ (
    .A(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_5400_)
);

FILL FILL_0__7362_ (
);

FILL FILL_4__14581_ (
);

FILL FILL_4__14161_ (
);

FILL FILL_2__8741_ (
);

FILL FILL_3__13994_ (
);

FILL FILL_2__8321_ (
);

FILL FILL_3__13574_ (
);

FILL FILL_3__13154_ (
);

FILL FILL_4__8247_ (
);

FILL FILL_2__12987_ (
);

FILL FILL_2__12567_ (
);

FILL FILL_2__12147_ (
);

FILL FILL_5__13901_ (
);

FILL SFILL89960x30050 (
);

FILL FILL_0__8987_ (
);

FILL FILL_5__16373_ (
);

FILL FILL_0__8567_ (
);

FILL FILL_6__9534_ (
);

DFFSR _10838_ (
    .Q(\datapath_1.regfile_1.regOut[31] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_1953_[0])
);

FILL FILL_0__8147_ (
);

INVX1 _10418_ (
    .A(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_1797_)
);

FILL FILL_4__15786_ (
);

FILL FILL_4__15366_ (
);

FILL FILL_1__12501_ (
);

FILL FILL_2__9526_ (
);

FILL FILL_0__11914_ (
);

FILL FILL_3__14779_ (
);

FILL FILL_3__14359_ (
);

FILL FILL_2__9106_ (
);

FILL FILL_1__15393_ (
);

FILL SFILL33800x26050 (
);

FILL FILL_5__7951_ (
);

FILL SFILL64200x17050 (
);

FILL FILL_5__7111_ (
);

FILL FILL_0__14386_ (
);

NOR2X1 _14671_ (
    .A(_5157_),
    .B(_3983__bF$buf1),
    .Y(_5158_)
);

AOI22X1 _14251_ (
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .B(_4038__bF$buf3),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_4747_)
);

FILL FILL_3__15720_ (
);

FILL FILL_3__15300_ (
);

FILL FILL_1__7943_ (
);

FILL FILL_1__7103_ (
);

FILL FILL_2__14713_ (
);

FILL FILL_3__7869_ (
);

FILL FILL_3__7449_ (
);

FILL FILL_5__12293_ (
);

FILL FILL_1__13706_ (
);

FILL FILL_4__11286_ (
);

FILL FILL_1__16178_ (
);

FILL FILL_3__10699_ (
);

FILL FILL_5__8736_ (
);

FILL FILL_3__10279_ (
);

FILL FILL_5__8316_ (
);

NOR2X1 _15876_ (
    .A(_6333_),
    .B(_6335_),
    .Y(_6336_)
);

AOI21X1 _15456_ (
    .A(_5926_),
    .B(_5905_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [9])
);

NOR2X1 _15036_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(\datapath_1.PCJump [26]),
    .Y(_5516_)
);

DFFSR _10591_ (
    .Q(\datapath_1.regfile_1.regOut[29] [9]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_1823_[9])
);

INVX1 _10171_ (
    .A(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_1673_)
);

FILL FILL_1__8728_ (
);

FILL FILL_3__11640_ (
);

FILL FILL_3__11220_ (
);

FILL FILL_2__15918_ (
);

FILL FILL_0__16112_ (
);

FILL FILL_2__10633_ (
);

FILL FILL_5__13498_ (
);

INVX1 _7798_ (
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_521_)
);

OAI21X1 _7378_ (
    .A(_257_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .C(_258_),
    .Y(_198_[30])
);

FILL SFILL18840x41050 (
);

FILL FILL_3_BUFX2_insert110 (
);

FILL FILL_1__12098_ (
);

FILL FILL_4__13852_ (
);

FILL FILL_4__13432_ (
);

FILL FILL_4__13012_ (
);

AND2X2 _11796_ (
    .A(_2888_),
    .B(_2148_),
    .Y(_2889_)
);

OAI22X1 _11376_ (
    .A(_2351_),
    .B(_2352_),
    .C(_2354_),
    .D(_2355_),
    .Y(_2493_)
);

FILL FILL_3__12845_ (
);

FILL FILL_3__12425_ (
);

FILL FILL_3__12005_ (
);

FILL FILL_4__7938_ (
);

FILL FILL_2__11838_ (
);

FILL FILL_0__12872_ (
);

FILL FILL_2__11418_ (
);

FILL FILL_0__12452_ (
);

FILL FILL_0__12032_ (
);

FILL FILL_5__15644_ (
);

FILL SFILL38840x6050 (
);

FILL FILL_5__15224_ (
);

FILL FILL_0__7838_ (
);

FILL FILL_0__7418_ (
);

DFFSR _9944_ (
    .Q(\datapath_1.regfile_1.regOut[24] [2]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1498_[2])
);

OAI21X1 _9524_ (
    .A(_1342_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1343_),
    .Y(_1303_[20])
);

OAI21X1 _9104_ (
    .A(_1123_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .C(_1124_),
    .Y(_1108_[8])
);

FILL FILL_1__8481_ (
);

FILL FILL_1__8061_ (
);

FILL FILL_4__14637_ (
);

FILL FILL_2__15671_ (
);

FILL FILL_4__14217_ (
);

FILL FILL_2__15251_ (
);

FILL FILL_1__14664_ (
);

FILL FILL_1__14244_ (
);

FILL FILL_0_BUFX2_insert240 (
);

FILL FILL_0_BUFX2_insert241 (
);

FILL FILL_0_BUFX2_insert242 (
);

FILL FILL_0_BUFX2_insert243 (
);

FILL FILL_0__13657_ (
);

FILL FILL_0_BUFX2_insert244 (
);

NAND3X1 _13942_ (
    .A(_4433_),
    .B(_4436_),
    .C(_4443_),
    .Y(_4444_)
);

FILL FILL_0__13237_ (
);

FILL FILL_0_BUFX2_insert245 (
);

OAI22X1 _13522_ (
    .A(_4031_),
    .B(_3982__bF$buf2),
    .C(_3978_),
    .D(_4032_),
    .Y(_4033_)
);

OAI21X1 _13102_ (
    .A(_3698_),
    .B(PCEn_bF$buf4),
    .C(_3699_),
    .Y(_3685_[7])
);

FILL FILL_0_BUFX2_insert246 (
);

FILL FILL_0_BUFX2_insert247 (
);

FILL FILL_0_BUFX2_insert248 (
);

FILL FILL_5__9274_ (
);

FILL FILL_0_BUFX2_insert249 (
);

FILL FILL_6__12991_ (
);

FILL FILL_5__16009_ (
);

FILL FILL_5__11984_ (
);

FILL FILL_5__11564_ (
);

FILL FILL_1__9266_ (
);

FILL FILL_5__11144_ (
);

FILL SFILL69080x50050 (
);

FILL FILL_4__7691_ (
);

FILL FILL_2__16036_ (
);

FILL FILL_4__10977_ (
);

FILL FILL_4__10557_ (
);

FILL FILL_4__10137_ (
);

FILL FILL_2__11591_ (
);

FILL FILL_2__11171_ (
);

FILL FILL_1__15869_ (
);

FILL FILL_1__15449_ (
);

FILL FILL_1__15029_ (
);

FILL FILL_1__10164_ (
);

INVX1 _14727_ (
    .A(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_5213_)
);

INVX1 _14307_ (
    .A(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_4802_)
);

FILL FILL_0__7591_ (
);

BUFX2 BUFX2_insert980 (
    .A(_3967_),
    .Y(_3967__bF$buf2)
);

FILL FILL_0__7171_ (
);

BUFX2 BUFX2_insert981 (
    .A(_3967_),
    .Y(_3967__bF$buf1)
);

FILL FILL_2__7189_ (
);

BUFX2 BUFX2_insert982 (
    .A(_3967_),
    .Y(_3967__bF$buf0)
);

BUFX2 BUFX2_insert983 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf7 )
);

FILL FILL_3__10911_ (
);

FILL FILL_6__13776_ (
);

BUFX2 BUFX2_insert984 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf6 )
);

BUFX2 BUFX2_insert985 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf5 )
);

BUFX2 BUFX2_insert986 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf4 )
);

FILL FILL_4__14390_ (
);

BUFX2 BUFX2_insert987 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf3 )
);

BUFX2 BUFX2_insert988 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf2 )
);

FILL FILL_0__15803_ (
);

BUFX2 BUFX2_insert989 (
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf1 )
);

FILL SFILL13720x29050 (
);

FILL FILL_5__12769_ (
);

FILL FILL_2__8970_ (
);

FILL FILL_5__12349_ (
);

FILL FILL_3__13383_ (
);

FILL FILL_2__8130_ (
);

FILL FILL_4__8896_ (
);

FILL FILL_4__8476_ (
);

FILL FILL_4__8056_ (
);

FILL FILL_2__12376_ (
);

FILL FILL_5__13710_ (
);

FILL FILL_1__11789_ (
);

FILL FILL_1__11369_ (
);

FILL FILL_4__12703_ (
);

FILL SFILL3640x70050 (
);

FILL FILL_3__6893_ (
);

FILL FILL_5__16182_ (
);

FILL FILL_0__8376_ (
);

FILL FILL_6__9343_ (
);

INVX1 _10647_ (
    .A(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_1909_)
);

DFFSR _10227_ (
    .Q(\datapath_1.regfile_1.regOut[26] [29]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1628_[29])
);

FILL FILL_1__12730_ (
);

FILL FILL_4__15595_ (
);

FILL FILL_4__15175_ (
);

FILL FILL_1__12310_ (
);

FILL FILL_2__9755_ (
);

FILL FILL_3__14588_ (
);

FILL FILL_2__9335_ (
);

FILL FILL_0__11723_ (
);

FILL FILL_3__14168_ (
);

FILL FILL_0__11303_ (
);

FILL FILL_5__7760_ (
);

FILL FILL_5__7340_ (
);

FILL SFILL3560x77050 (
);

NOR2X1 _14480_ (
    .A(_4967_),
    .B(_4970_),
    .Y(_4971_)
);

FILL FILL_0__14195_ (
);

INVX1 _14060_ (
    .A(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_4560_)
);

FILL FILL_5__14915_ (
);

FILL SFILL38920x33050 (
);

FILL FILL_1__7752_ (
);

FILL FILL_1__7332_ (
);

FILL FILL_4__13908_ (
);

FILL FILL_2__14942_ (
);

FILL FILL_2__14522_ (
);

FILL FILL_3__7678_ (
);

FILL FILL_2__14102_ (
);

FILL SFILL44120x9050 (
);

FILL FILL_1__13935_ (
);

FILL FILL_1__13515_ (
);

FILL FILL_4__11095_ (
);

FILL FILL_0__12508_ (
);

FILL FILL_5__8965_ (
);

FILL FILL_5__8125_ (
);

INVX1 _15685_ (
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_6150_)
);

NAND3X1 _15265_ (
    .A(_5735_),
    .B(_5736_),
    .C(_5739_),
    .Y(_5740_)
);

FILL FILL_3__16314_ (
);

FILL SFILL28920x76050 (
);

FILL SFILL3560x32050 (
);

FILL FILL_5__10835_ (
);

FILL FILL_1__8957_ (
);

FILL FILL_5__10415_ (
);

FILL FILL_1__8117_ (
);

FILL FILL_2__15727_ (
);

FILL FILL_2__15307_ (
);

FILL FILL_4__6962_ (
);

FILL FILL_0__16341_ (
);

FILL FILL_2__10442_ (
);

FILL FILL_2__10022_ (
);

FILL FILL_6__6888_ (
);

OAI21X1 _7187_ (
    .A(_150_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_151_),
    .Y(_133_[9])
);

FILL FILL112200x27050 (
);

FILL FILL_3__9404_ (
);

FILL FILL_0__6862_ (
);

FILL FILL_4__13661_ (
);

FILL FILL_4__13241_ (
);

FILL SFILL113720x40050 (
);

OAI21X1 _11185_ (
    .A(_2261_),
    .B(_2284_),
    .C(_2303_),
    .Y(_2304_)
);

FILL FILL_2__7821_ (
);

FILL FILL_3__12654_ (
);

FILL FILL_3__12234_ (
);

FILL SFILL28920x31050 (
);

FILL FILL_4__7747_ (
);

FILL FILL_4__7327_ (
);

FILL FILL_2__11647_ (
);

FILL FILL_2__11227_ (
);

FILL FILL_0__12261_ (
);

FILL FILL_5__15873_ (
);

FILL FILL_5__15453_ (
);

FILL FILL_5__15033_ (
);

FILL FILL_0__7227_ (
);

FILL FILL_6__8614_ (
);

OAI21X1 _9753_ (
    .A(_1454_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1455_),
    .Y(_1433_[11])
);

DFFSR _9333_ (
    .Q(\datapath_1.regfile_1.regOut[19] [31]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_1173_[31])
);

FILL FILL_4__14866_ (
);

FILL FILL_4__14446_ (
);

FILL FILL_4__14026_ (
);

FILL FILL_2__15480_ (
);

FILL FILL_2__15060_ (
);

FILL FILL_3__13859_ (
);

FILL FILL_2__8606_ (
);

FILL FILL_3__13439_ (
);

FILL FILL_1__14893_ (
);

FILL FILL_1__14473_ (
);

FILL FILL_3__13019_ (
);

FILL FILL_1__14053_ (
);

FILL FILL_0__13886_ (
);

AOI22X1 _13751_ (
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .B(_4038__bF$buf1),
    .C(_4079__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_4257_)
);

FILL FILL_0__13466_ (
);

AND2X2 _13331_ (
    .A(_3813_),
    .B(_3856_),
    .Y(\datapath_1.regfile_1.regEn [18])
);

FILL FILL_0__13046_ (
);

FILL FILL_3__14800_ (
);

FILL FILL_5__9083_ (
);

FILL FILL_5__16238_ (
);

FILL FILL_3__6949_ (
);

FILL FILL_5__11793_ (
);

FILL FILL_1__9495_ (
);

FILL FILL_5__11373_ (
);

FILL SFILL14120x59050 (
);

FILL FILL_2__16265_ (
);

FILL FILL_4__7080_ (
);

FILL FILL_4__10786_ (
);

FILL FILL_4__10366_ (
);

FILL SFILL94360x60050 (
);

FILL FILL_4_BUFX2_insert70 (
);

FILL FILL_4_BUFX2_insert71 (
);

FILL FILL_4_BUFX2_insert72 (
);

FILL FILL_1__15678_ (
);

FILL FILL_4_BUFX2_insert73 (
);

FILL FILL_1__15258_ (
);

FILL FILL_4_BUFX2_insert74 (
);

FILL FILL_4_BUFX2_insert75 (
);

FILL FILL_5__7816_ (
);

FILL FILL_4_BUFX2_insert76 (
);

FILL FILL_4_BUFX2_insert77 (
);

FILL FILL_1__10393_ (
);

FILL FILL_4_BUFX2_insert78 (
);

FILL FILL_4_BUFX2_insert79 (
);

AOI22X1 _14956_ (
    .A(_4129_),
    .B(\datapath_1.regfile_1.regOut[27] [31]),
    .C(\datapath_1.regfile_1.regOut[31] [31]),
    .D(_3995__bF$buf0),
    .Y(_5437_)
);

NOR2X1 _14536_ (
    .A(_5025_),
    .B(_5022_),
    .Y(_5026_)
);

INVX1 _14116_ (
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_4615_)
);

FILL FILL_1__7808_ (
);

FILL FILL_3__10300_ (
);

FILL FILL_0__15612_ (
);

FILL FILL_5__12998_ (
);

FILL FILL_5__12578_ (
);

FILL FILL_5__12158_ (
);

BUFX2 _6878_ (
    .A(_2_[8]),
    .Y(memoryWriteData[8])
);

FILL SFILL18680x1050 (
);

FILL SFILL18840x36050 (
);

FILL FILL_2__12185_ (
);

FILL FILL_1__11598_ (
);

FILL FILL_1__11178_ (
);

FILL FILL_4__12512_ (
);

NAND2X1 _10876_ (
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2024_)
);

FILL FILL_0__8185_ (
);

DFFSR _10456_ (
    .Q(\datapath_1.regfile_1.regOut[28] [2]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_1758_[2])
);

OAI21X1 _10036_ (
    .A(_1602_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1603_),
    .Y(_1563_[20])
);

FILL FILL_3__11925_ (
);

FILL FILL_3__11505_ (
);

FILL FILL_2__9984_ (
);

FILL FILL_2__10918_ (
);

FILL SFILL80040x50050 (
);

FILL FILL_0__11952_ (
);

FILL FILL_2__9144_ (
);

FILL FILL_3__14397_ (
);

FILL FILL_0__11532_ (
);

FILL FILL_0__11112_ (
);

FILL FILL_6__15731_ (
);

FILL FILL_6__15311_ (
);

FILL FILL_5__14724_ (
);

FILL FILL_5__14304_ (
);

FILL FILL_0__6918_ (
);

OAI21X1 _8604_ (
    .A(_871_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_872_),
    .Y(_848_[12])
);

FILL FILL_1__7981_ (
);

FILL FILL_1__7561_ (
);

FILL FILL_4__13717_ (
);

FILL FILL_2__14751_ (
);

FILL FILL_2__14331_ (
);

FILL FILL_3__7487_ (
);

FILL FILL_3__7067_ (
);

FILL FILL_1__13744_ (
);

FILL FILL_1__13324_ (
);

FILL FILL_4__16189_ (
);

FILL FILL_0__12737_ (
);

OAI21X1 _12602_ (
    .A(_3446_),
    .B(vdd),
    .C(_3447_),
    .Y(_3425_[11])
);

FILL FILL_0__12317_ (
);

FILL SFILL69480x59050 (
);

FILL FILL_5__8774_ (
);

FILL FILL_5__8354_ (
);

FILL FILL_6__11651_ (
);

FILL FILL_6__11231_ (
);

NOR2X1 _15494_ (
    .A(_5960_),
    .B(_5963_),
    .Y(_5964_)
);

FILL FILL_5__15929_ (
);

NOR2X1 _15074_ (
    .A(_5553_),
    .B(_5550_),
    .Y(_5554_)
);

FILL FILL_5__15509_ (
);

FILL FILL_3__16123_ (
);

NAND2X1 _9809_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1493_)
);

FILL FILL_1__8766_ (
);

FILL FILL_5__10644_ (
);

FILL FILL_1__8346_ (
);

FILL FILL_2__15956_ (
);

FILL FILL_2__15536_ (
);

FILL FILL_2__15116_ (
);

FILL FILL_0__16150_ (
);

FILL FILL_2__10671_ (
);

FILL FILL_2__10251_ (
);

FILL FILL_1__14949_ (
);

FILL FILL_1__14529_ (
);

FILL FILL_1__14109_ (
);

FILL FILL_3__9633_ (
);

AOI22X1 _13807_ (
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .B(_4038__bF$buf2),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_4312_)
);

FILL FILL_3__9213_ (
);

FILL FILL_5__9979_ (
);

FILL FILL_5__9139_ (
);

FILL FILL_4__13890_ (
);

FILL FILL_4__13470_ (
);

OAI22X1 _16279_ (
    .A(_5463__bF$buf2),
    .B(_6728_),
    .C(_6727_),
    .D(_5504__bF$buf2),
    .Y(_6729_)
);

FILL FILL_5__11849_ (
);

FILL FILL_2__7630_ (
);

FILL FILL_3__12883_ (
);

FILL FILL_5__11429_ (
);

FILL FILL_3__12463_ (
);

FILL FILL_2__7210_ (
);

FILL FILL_5__11009_ (
);

FILL FILL_3__12043_ (
);

FILL FILL_4__7976_ (
);

FILL FILL_4__7556_ (
);

FILL FILL_2__11876_ (
);

FILL FILL_2__11456_ (
);

FILL FILL_0__12490_ (
);

FILL FILL_2__11036_ (
);

FILL FILL_0__12070_ (
);

FILL FILL_1__10449_ (
);

FILL FILL_1__10029_ (
);

FILL SFILL3640x65050 (
);

FILL FILL_5__15682_ (
);

FILL FILL_0__7876_ (
);

FILL FILL_5__15262_ (
);

FILL FILL_0__7456_ (
);

OAI21X1 _9982_ (
    .A(_1566_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1567_),
    .Y(_1563_[2])
);

DFFSR _9562_ (
    .Q(\datapath_1.regfile_1.regOut[21] [4]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1303_[4])
);

FILL FILL_0__7036_ (
);

NAND2X1 _9142_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1150_)
);

FILL SFILL104520x82050 (
);

FILL SFILL43880x72050 (
);

FILL FILL_1__11810_ (
);

FILL FILL_4__14675_ (
);

FILL FILL_4__14255_ (
);

INVX1 _12199_ (
    .A(\datapath_1.PCJump [28]),
    .Y(_3186_)
);

FILL FILL_2__8835_ (
);

FILL FILL_3__13668_ (
);

FILL FILL_0__10803_ (
);

FILL SFILL3560x3050 (
);

FILL FILL_3__13248_ (
);

FILL FILL_1__14282_ (
);

FILL FILL_0_BUFX2_insert620 (
);

FILL FILL_5__6840_ (
);

FILL FILL_0_BUFX2_insert621 (
);

FILL SFILL38120x45050 (
);

FILL SFILL3480x8050 (
);

FILL FILL_0_BUFX2_insert622 (
);

FILL FILL_0_BUFX2_insert623 (
);

FILL FILL_0_BUFX2_insert624 (
);

INVX1 _13980_ (
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_4481_)
);

FILL FILL_0__13695_ (
);

FILL FILL_0__13275_ (
);

FILL FILL_0_BUFX2_insert625 (
);

NOR2X1 _13560_ (
    .A(_4069_),
    .B(_4054_),
    .Y(_4070_)
);

FILL FILL_0_BUFX2_insert626 (
);

NAND2X1 _13140_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [20]),
    .Y(_3725_)
);

FILL FILL_0_BUFX2_insert627 (
);

FILL SFILL38920x28050 (
);

FILL FILL_0_BUFX2_insert628 (
);

FILL FILL_0_BUFX2_insert629 (
);

FILL SFILL83560x54050 (
);

FILL FILL_2__13602_ (
);

FILL FILL_5__16047_ (
);

FILL SFILL3640x20050 (
);

FILL FILL_5__11182_ (
);

FILL FILL_2__16074_ (
);

FILL FILL_4__10175_ (
);

FILL FILL_0__9602_ (
);

FILL FILL_1__15487_ (
);

FILL FILL_1__15067_ (
);

FILL FILL_5__7625_ (
);

FILL FILL_5__7205_ (
);

FILL FILL_4__16401_ (
);

FILL SFILL28600x50050 (
);

FILL SFILL59000x41050 (
);

NOR2X1 _14765_ (
    .A(_5239_),
    .B(_5249_),
    .Y(_5250_)
);

FILL FILL_6__10502_ (
);

NAND3X1 _14345_ (
    .A(_4837_),
    .B(_4838_),
    .C(_4834_),
    .Y(_4839_)
);

FILL FILL_3__15814_ (
);

FILL FILL_1__7617_ (
);

FILL SFILL104440x44050 (
);

FILL FILL_2__14807_ (
);

FILL FILL_0__15841_ (
);

FILL FILL_0__15421_ (
);

FILL FILL_0__15001_ (
);

FILL FILL_5__12387_ (
);

FILL FILL_4__8094_ (
);

FILL SFILL33880x70050 (
);

FILL FILL_3__8904_ (
);

FILL FILL_6__11707_ (
);

FILL FILL_4__12741_ (
);

FILL FILL_4__12321_ (
);

OAI21X1 _10685_ (
    .A(_1933_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1934_),
    .Y(_1888_[23])
);

FILL SFILL49080x41050 (
);

OAI21X1 _10265_ (
    .A(_1714_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .C(_1715_),
    .Y(_1693_[11])
);

FILL FILL_2__6901_ (
);

FILL FILL_3__11734_ (
);

FILL FILL_3__11314_ (
);

FILL SFILL28920x26050 (
);

FILL FILL_0__16206_ (
);

FILL FILL_2__9793_ (
);

FILL FILL_0__11761_ (
);

FILL FILL_2__10307_ (
);

FILL FILL_2__9373_ (
);

FILL FILL_0__11341_ (
);

FILL FILL_4__9299_ (
);

FILL FILL_5__14953_ (
);

FILL FILL_5__14533_ (
);

FILL FILL_5__14113_ (
);

OAI21X1 _8833_ (
    .A(_983_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .C(_984_),
    .Y(_978_[3])
);

DFFSR _8413_ (
    .Q(\datapath_1.regfile_1.regOut[12] [7]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_718_[7])
);

FILL FILL_1__7370_ (
);

FILL FILL_4__13946_ (
);

FILL FILL_2__14980_ (
);

FILL FILL_4__13526_ (
);

FILL FILL_2__14560_ (
);

FILL FILL_4__13106_ (
);

FILL FILL_2__14140_ (
);

FILL FILL_3__7296_ (
);

FILL FILL_3__12519_ (
);

FILL FILL_1__13973_ (
);

FILL FILL_1__13553_ (
);

FILL FILL_1__13133_ (
);

FILL FILL_0__12966_ (
);

OAI21X1 _12831_ (
    .A(_3558_),
    .B(vdd),
    .C(_3559_),
    .Y(_3555_[2])
);

FILL FILL_0__12126_ (
);

OAI21X1 _12411_ (
    .A(_3338_),
    .B(MemToReg_bF$buf3),
    .C(_3339_),
    .Y(\datapath_1.mux_wd3.dout [22])
);

FILL FILL_5__8583_ (
);

FILL FILL_5__15738_ (
);

FILL FILL_5__15318_ (
);

FILL SFILL39480x53050 (
);

FILL FILL_3__16352_ (
);

NAND2X1 _9618_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1386_)
);

FILL FILL_1__8995_ (
);

FILL FILL_5__10873_ (
);

FILL FILL_1__8575_ (
);

FILL FILL_5__10453_ (
);

FILL FILL_5__10033_ (
);

FILL FILL_2__15765_ (
);

FILL FILL_2__15345_ (
);

FILL SFILL39000x82050 (
);

FILL SFILL94360x55050 (
);

FILL FILL_2__10060_ (
);

FILL FILL_1__14758_ (
);

FILL FILL_1__14338_ (
);

FILL FILL_3__9862_ (
);

INVX1 _13616_ (
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_4125_)
);

FILL FILL_3__9022_ (
);

FILL FILL_5__9788_ (
);

FILL FILL_5__9368_ (
);

AOI22X1 _16088_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [26]),
    .C(\datapath_1.regfile_1.regOut[22] [26]),
    .D(_5650_),
    .Y(_6542_)
);

FILL FILL_5__11658_ (
);

FILL FILL_5__11238_ (
);

FILL FILL_3__12272_ (
);

FILL FILL_4__7365_ (
);

FILL FILL_2__11685_ (
);

FILL FILL_2__11265_ (
);

FILL SFILL94360x10050 (
);

FILL FILL_1__10678_ (
);

FILL FILL_1__10258_ (
);

FILL FILL_5__15491_ (
);

FILL FILL_5__15071_ (
);

FILL FILL_0__7685_ (
);

NAND2X1 _9791_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1481_)
);

FILL FILL_6__8232_ (
);

NAND2X1 _9371_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1262_)
);

FILL FILL112440x50 (
);

FILL FILL_4__14484_ (
);

FILL FILL_4__14064_ (
);

FILL FILL_2__8644_ (
);

FILL FILL_3__13897_ (
);

FILL FILL_2__8224_ (
);

FILL FILL_3__13477_ (
);

FILL FILL_1__14091_ (
);

FILL FILL_0__13084_ (
);

FILL SFILL114600x72050 (
);

FILL FILL_5__13804_ (
);

FILL SFILL53960x62050 (
);

FILL SFILL84360x53050 (
);

FILL FILL_4__9931_ (
);

FILL FILL_4__9511_ (
);

FILL FILL_2__13831_ (
);

FILL FILL_3__6987_ (
);

FILL FILL_2__13411_ (
);

FILL FILL_5__16276_ (
);

FILL FILL_6__9017_ (
);

FILL FILL_4__15689_ (
);

FILL FILL_1__12824_ (
);

FILL FILL_1__12404_ (
);

FILL FILL_4__15269_ (
);

FILL FILL_2__9849_ (
);

FILL SFILL114520x79050 (
);

FILL FILL_2__9429_ (
);

FILL FILL_0__11817_ (
);

FILL FILL_0__9411_ (
);

FILL FILL_2__9009_ (
);

FILL FILL_1__15296_ (
);

FILL FILL_5__7854_ (
);

FILL FILL_5__7434_ (
);

FILL FILL_4__16210_ (
);

NOR2X1 _14994_ (
    .A(_5473_),
    .B(_5467_),
    .Y(_5474_)
);

INVX1 _14574_ (
    .A(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_5063_)
);

FILL FILL_0__14289_ (
);

NAND3X1 _14154_ (
    .A(_4643_),
    .B(_4644_),
    .C(_4651_),
    .Y(_4652_)
);

FILL FILL_3__15623_ (
);

FILL FILL_3__15203_ (
);

FILL FILL_1__7846_ (
);

FILL SFILL114120x65050 (
);

FILL FILL_1__7426_ (
);

FILL FILL_2__14616_ (
);

FILL FILL_0__15650_ (
);

FILL FILL_0__15230_ (
);

FILL FILL_5__12196_ (
);

FILL FILL_1__13609_ (
);

FILL FILL_4__11189_ (
);

FILL FILL_3__8713_ (
);

FILL FILL_5__8639_ (
);

FILL FILL_5__8219_ (
);

FILL SFILL53880x24050 (
);

FILL FILL_4__12970_ (
);

AOI22X1 _15779_ (
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_6241_)
);

OAI22X1 _15359_ (
    .A(_5466__bF$buf3),
    .B(_5831_),
    .C(_4313_),
    .D(_5483__bF$buf4),
    .Y(_5832_)
);

FILL FILL_4__12130_ (
);

FILL FILL_3__16408_ (
);

OAI21X1 _10494_ (
    .A(_1826_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1827_),
    .Y(_1823_[2])
);

FILL FILL_5__10929_ (
);

DFFSR _10074_ (
    .Q(\datapath_1.regfile_1.regOut[25] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_1563_[4])
);

FILL FILL_5__10509_ (
);

FILL FILL_3__11963_ (
);

FILL FILL_3__11543_ (
);

FILL SFILL43960x60050 (
);

FILL FILL_3__11123_ (
);

FILL FILL_0__16015_ (
);

INVX1 _16300_ (
    .A(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_6749_)
);

FILL FILL_2__10956_ (
);

FILL FILL_2__10536_ (
);

FILL FILL_0__11990_ (
);

FILL FILL_2__10116_ (
);

FILL FILL_0__11570_ (
);

FILL FILL_0__11150_ (
);

FILL FILL_3__9918_ (
);

FILL FILL_5__14762_ (
);

FILL FILL_0__6956_ (
);

FILL FILL_5__14342_ (
);

NAND2X1 _8642_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_898_)
);

NAND2X1 _8222_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_679_)
);

FILL FILL_4__13755_ (
);

FILL FILL_4__13335_ (
);

NOR2X1 _11699_ (
    .A(_2792_),
    .B(_2798_),
    .Y(_2799_)
);

NOR2X1 _11279_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2398_)
);

FILL FILL_3__12748_ (
);

FILL FILL_1__13782_ (
);

FILL FILL_3__12328_ (
);

FILL FILL_1__13362_ (
);

FILL FILL112280x71050 (
);

FILL FILL_0__12775_ (
);

NAND2X1 _12640_ (
    .A(vdd),
    .B(memoryOutData[24]),
    .Y(_3473_)
);

FILL FILL_0__12355_ (
);

NAND3X1 _12220_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [1]),
    .C(_3198__bF$buf4),
    .Y(_3204_)
);

FILL FILL_5__8392_ (
);

FILL SFILL83560x49050 (
);

FILL FILL_5__15967_ (
);

FILL FILL_5__15547_ (
);

FILL FILL_5__15127_ (
);

NAND2X1 _9847_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .Y(_1562_)
);

FILL FILL_3__16161_ (
);

INVX1 _9427_ (
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_1299_)
);

FILL SFILL3640x15050 (
);

FILL FILL_5__10682_ (
);

INVX1 _9007_ (
    .A(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_1080_)
);

FILL FILL_1__8384_ (
);

FILL FILL_5__10262_ (
);

FILL FILL_2__15994_ (
);

FILL FILL_2__15574_ (
);

FILL SFILL104520x32050 (
);

FILL FILL_2__15154_ (
);

FILL SFILL43880x22050 (
);

FILL FILL_1__14987_ (
);

FILL FILL_1__14567_ (
);

FILL FILL_1__14147_ (
);

FILL FILL_4__15901_ (
);

FILL SFILL59000x36050 (
);

FILL FILL_3__9671_ (
);

INVX1 _13845_ (
    .A(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_4349_)
);

FILL FILL_3__9251_ (
);

OAI22X1 _13425_ (
    .A(_3933_),
    .B(_3936__bF$buf3),
    .C(_3935__bF$buf3),
    .D(_3934_),
    .Y(_3937_)
);

INVX1 _13005_ (
    .A(_2_[18]),
    .Y(_3655_)
);

FILL FILL_5__9597_ (
);

FILL FILL_6__12474_ (
);

FILL SFILL104440x39050 (
);

FILL FILL_0__14921_ (
);

FILL FILL_0__14501_ (
);

FILL FILL_5__11887_ (
);

FILL FILL_5__11467_ (
);

FILL FILL_1__9169_ (
);

FILL FILL_5__11047_ (
);

FILL FILL_3__12081_ (
);

FILL FILL_2__16359_ (
);

FILL FILL_4__7594_ (
);

FILL SFILL33880x65050 (
);

FILL FILL_4__7174_ (
);

FILL FILL_2__11494_ (
);

FILL FILL_2__11074_ (
);

FILL FILL_1__10487_ (
);

FILL SFILL49000x79050 (
);

FILL FILL_1__10067_ (
);

FILL FILL_4__11821_ (
);

FILL FILL_4__11401_ (
);

FILL FILL_0__7494_ (
);

FILL SFILL49080x36050 (
);

FILL FILL_0__7074_ (
);

DFFSR _9180_ (
    .Q(\datapath_1.regfile_1.regOut[18] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_1108_[6])
);

FILL FILL_3__10814_ (
);

FILL FILL_6__13679_ (
);

FILL FILL_4__14293_ (
);

FILL FILL_0__15706_ (
);

FILL FILL_2__8873_ (
);

FILL FILL_2__8453_ (
);

FILL FILL_0__10421_ (
);

FILL FILL_3__13286_ (
);

FILL FILL_0__10001_ (
);

FILL FILL_6__14620_ (
);

FILL FILL_4__8379_ (
);

FILL FILL_2__12699_ (
);

FILL FILL_2__12279_ (
);

FILL FILL_5__13613_ (
);

DFFSR _7913_ (
    .Q(\datapath_1.regfile_1.regOut[8] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_458_[19])
);

FILL FILL_1__6870_ (
);

FILL FILL_4__9740_ (
);

FILL FILL_4__12606_ (
);

FILL FILL_2__13640_ (
);

FILL FILL_2__13220_ (
);

FILL FILL_5__16085_ (
);

FILL FILL_0__8699_ (
);

FILL SFILL49000x34050 (
);

FILL FILL_1__12633_ (
);

FILL FILL_4__15498_ (
);

FILL FILL_1__12213_ (
);

FILL FILL_4__15078_ (
);

FILL SFILL94440x43050 (
);

FILL FILL_0__9640_ (
);

FILL FILL_2__9658_ (
);

FILL FILL_0__9220_ (
);

INVX1 _11911_ (
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_2982_)
);

FILL FILL_2__9238_ (
);

FILL FILL_0__11626_ (
);

FILL FILL_0__11206_ (
);

FILL FILL_5__7243_ (
);

OAI22X1 _14383_ (
    .A(_4874_),
    .B(_3935__bF$buf1),
    .C(_3971__bF$buf0),
    .D(_4875_),
    .Y(_4876_)
);

FILL FILL_0__14098_ (
);

FILL FILL_5__14818_ (
);

FILL FILL_3__15852_ (
);

FILL FILL_3__15432_ (
);

FILL FILL_3__15012_ (
);

FILL FILL_1__7235_ (
);

FILL FILL_2__14845_ (
);

FILL FILL_2__14425_ (
);

FILL FILL_2__14005_ (
);

FILL FILL_1__13838_ (
);

FILL FILL_1__13418_ (
);

FILL FILL_3__8522_ (
);

FILL FILL_3__8102_ (
);

FILL FILL_5__8868_ (
);

FILL FILL_5__8448_ (
);

NAND3X1 _15588_ (
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf1),
    .Y(_6055_)
);

INVX1 _15168_ (
    .A(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_5645_)
);

FILL SFILL23800x61050 (
);

FILL FILL_3__16217_ (
);

FILL SFILL84040x72050 (
);

FILL FILL_5__10318_ (
);

FILL FILL_3__11772_ (
);

FILL FILL_3__11352_ (
);

FILL FILL_4__6865_ (
);

FILL FILL_0__16244_ (
);

FILL FILL_2__10765_ (
);

FILL FILL_1__9801_ (
);

FILL SFILL4440x59050 (
);

FILL FILL_3__9727_ (
);

FILL FILL_5__14991_ (
);

FILL FILL_5__14571_ (
);

FILL FILL_5__14151_ (
);

FILL FILL112280x5050 (
);

NAND2X1 _8871_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1010_)
);

FILL FILL_6__7312_ (
);

NAND2X1 _8451_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_791_)
);

DFFSR _8031_ (
    .Q(\datapath_1.regfile_1.regOut[9] [9]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_523_[9])
);

FILL FILL_4__13984_ (
);

FILL FILL_4__13564_ (
);

FILL SFILL8760x67050 (
);

FILL FILL_4__13144_ (
);

NOR2X1 _11088_ (
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(_2206_),
    .Y(_2207_)
);

FILL FILL_3__12977_ (
);

FILL FILL_2__7724_ (
);

FILL FILL_2__7304_ (
);

FILL FILL_1__13591_ (
);

FILL FILL_3__12137_ (
);

FILL FILL_1__13171_ (
);

FILL FILL_0__12584_ (
);

FILL FILL_0__12164_ (
);

FILL SFILL84360x48050 (
);

FILL FILL_5_BUFX2_insert400 (
);

FILL FILL_5_BUFX2_insert401 (
);

FILL FILL_2__12911_ (
);

FILL FILL_5__15776_ (
);

FILL FILL_5_BUFX2_insert402 (
);

FILL FILL_5__15356_ (
);

FILL FILL_3__16390_ (
);

FILL FILL_5_BUFX2_insert403 (
);

FILL FILL_5_BUFX2_insert404 (
);

INVX1 _9656_ (
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_1411_)
);

FILL FILL_5_BUFX2_insert405 (
);

INVX1 _9236_ (
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_1192_)
);

FILL FILL_5_BUFX2_insert406 (
);

FILL FILL_5__10491_ (
);

FILL FILL_1__8193_ (
);

FILL FILL_5_BUFX2_insert407 (
);

FILL FILL_5_BUFX2_insert408 (
);

FILL FILL_1__11904_ (
);

FILL FILL_4__14769_ (
);

FILL FILL_5_BUFX2_insert409 (
);

FILL FILL_4__14349_ (
);

FILL FILL_2__15383_ (
);

FILL FILL_0__8911_ (
);

FILL SFILL8760x22050 (
);

FILL FILL_2__8509_ (
);

FILL SFILL84760x17050 (
);

FILL FILL_1__14796_ (
);

FILL FILL_1__14376_ (
);

FILL FILL_5__6934_ (
);

FILL FILL_4__15710_ (
);

FILL FILL_0__13789_ (
);

FILL FILL_3__9480_ (
);

OAI22X1 _13654_ (
    .A(_4161_),
    .B(_3972__bF$buf1),
    .C(_3924__bF$buf0),
    .D(_4160_),
    .Y(_4162_)
);

FILL FILL_0__13369_ (
);

NOR2X1 _13234_ (
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_3777_)
);

FILL FILL_3__14703_ (
);

FILL SFILL114600x22050 (
);

FILL FILL_1__6926_ (
);

FILL SFILL53960x12050 (
);

FILL FILL_0__14730_ (
);

FILL FILL_0__14310_ (
);

FILL FILL_5__11696_ (
);

FILL FILL_1__9398_ (
);

FILL FILL_5__11276_ (
);

FILL FILL_2__16168_ (
);

FILL FILL_4__10689_ (
);

FILL FILL_4__10269_ (
);

FILL FILL_5__7719_ (
);

FILL SFILL53880x19050 (
);

FILL FILL_2_BUFX2_insert530 (
);

FILL FILL_1__10296_ (
);

FILL FILL_2_BUFX2_insert531 (
);

FILL FILL_2_BUFX2_insert532 (
);

NOR2X1 _14859_ (
    .A(_5341_),
    .B(_5329_),
    .Y(_5342_)
);

FILL FILL_2_BUFX2_insert533 (
);

FILL FILL_2_BUFX2_insert534 (
);

INVX1 _14439_ (
    .A(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_4931_)
);

FILL FILL_4__11630_ (
);

FILL FILL_2_BUFX2_insert535 (
);

NOR2X1 _14019_ (
    .A(_4516_),
    .B(_4519_),
    .Y(_4520_)
);

FILL FILL_4__11210_ (
);

FILL FILL_3__15908_ (
);

FILL FILL_2_BUFX2_insert536 (
);

FILL FILL_2_BUFX2_insert537 (
);

FILL FILL_2_BUFX2_insert538 (
);

FILL FILL_2_BUFX2_insert539 (
);

FILL FILL_1__16102_ (
);

FILL SFILL43960x55050 (
);

FILL FILL_3__10623_ (
);

FILL FILL_0__15935_ (
);

FILL FILL_0__15515_ (
);

NAND2X1 _15800_ (
    .A(_6255_),
    .B(_6261_),
    .Y(_6262_)
);

FILL FILL_0__10650_ (
);

FILL FILL_2__8262_ (
);

FILL FILL_0__10230_ (
);

FILL FILL_3__13095_ (
);

FILL FILL_4__8188_ (
);

FILL FILL_2__12088_ (
);

FILL FILL_5__13842_ (
);

FILL FILL_5__13422_ (
);

FILL FILL_5__13002_ (
);

NAND2X1 _7722_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_427_)
);

NAND2X1 _7302_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_208_)
);

FILL FILL_4__12835_ (
);

FILL FILL_4__12415_ (
);

FILL FILL_0__8088_ (
);

NAND2X1 _10779_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1977_)
);

NAND2X1 _10359_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .Y(_1822_)
);

FILL FILL_3__11828_ (
);

FILL FILL_1__12862_ (
);

FILL FILL_3__11408_ (
);

FILL FILL_1__12442_ (
);

FILL FILL_1__12022_ (
);

FILL SFILL43960x10050 (
);

FILL FILL112280x66050 (
);

FILL FILL_2__9887_ (
);

FILL FILL_0__11855_ (
);

FILL FILL_2__9467_ (
);

NAND2X1 _11720_ (
    .A(_2172_),
    .B(_2817_),
    .Y(_2818_)
);

FILL FILL_0__11435_ (
);

FILL FILL_0__11015_ (
);

NAND2X1 _11300_ (
    .A(_2250_),
    .B(_2418_),
    .Y(_2419_)
);

FILL FILL_5__7892_ (
);

FILL FILL_6__15214_ (
);

FILL FILL_5__7472_ (
);

FILL FILL_5__7052_ (
);

OAI22X1 _14192_ (
    .A(_4687_),
    .B(_3936__bF$buf2),
    .C(_3935__bF$buf3),
    .D(_4688_),
    .Y(_4689_)
);

FILL FILL_5__14627_ (
);

FILL FILL_3__15661_ (
);

FILL FILL_5__14207_ (
);

FILL FILL_3__15241_ (
);

DFFSR _8927_ (
    .Q(\datapath_1.regfile_1.regOut[16] [9]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_978_[9])
);

INVX1 _8507_ (
    .A(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_828_)
);

FILL FILL_1__7884_ (
);

FILL FILL_1__7464_ (
);

FILL FILL_1__7044_ (
);

FILL FILL_2__14654_ (
);

FILL SFILL43880x17050 (
);

FILL FILL_2__14234_ (
);

FILL FILL_1__13647_ (
);

FILL FILL_1__13227_ (
);

FILL SFILL43800x4050 (
);

FILL FILL_1_BUFX2_insert550 (
);

FILL FILL_3__8751_ (
);

FILL FILL_1_BUFX2_insert551 (
);

FILL FILL_3__8331_ (
);

DFFSR _12925_ (
    .Q(\datapath_1.a [6]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_3555_[6])
);

FILL FILL_1_BUFX2_insert552 (
);

FILL FILL_1_BUFX2_insert553 (
);

INVX1 _12505_ (
    .A(ALUOut[22]),
    .Y(_3403_)
);

FILL FILL_1_BUFX2_insert554 (
);

FILL FILL112280x21050 (
);

FILL FILL_1_BUFX2_insert555 (
);

FILL SFILL84280x4050 (
);

FILL FILL_1_BUFX2_insert556 (
);

FILL FILL_1_BUFX2_insert557 (
);

FILL FILL_5__8257_ (
);

FILL FILL_1_BUFX2_insert558 (
);

FILL FILL_1_BUFX2_insert559 (
);

AOI21X1 _15397_ (
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .B(_5570__bF$buf3),
    .C(_5868_),
    .Y(_5869_)
);

FILL FILL_6__11134_ (
);

FILL FILL_3__16026_ (
);

FILL FILL_5__10967_ (
);

FILL FILL_5__10547_ (
);

FILL FILL_5__10127_ (
);

FILL FILL_1__8249_ (
);

FILL FILL_3__11581_ (
);

FILL FILL_3__11161_ (
);

FILL FILL_2__15859_ (
);

FILL FILL_2__15439_ (
);

FILL FILL_2__15019_ (
);

FILL FILL_0__16053_ (
);

FILL FILL_2__10994_ (
);

FILL FILL_2__10574_ (
);

FILL FILL_2__10154_ (
);

FILL FILL_1__9610_ (
);

FILL FILL_3__9536_ (
);

FILL FILL_4__10901_ (
);

FILL FILL_3__9116_ (
);

FILL FILL_5__14380_ (
);

FILL FILL_0__6994_ (
);

DFFSR _8680_ (
    .Q(\datapath_1.regfile_1.regOut[14] [18]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_848_[18])
);

INVX1 _8260_ (
    .A(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_704_)
);

FILL FILL_4__13793_ (
);

FILL FILL_4__13373_ (
);

FILL SFILL18200x69050 (
);

FILL FILL_2__7953_ (
);

FILL FILL_3__12786_ (
);

FILL FILL_3__12366_ (
);

FILL FILL_2__7113_ (
);

FILL FILL_4__7879_ (
);

FILL FILL_6__13700_ (
);

BUFX2 BUFX2_insert225 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf4 )
);

FILL FILL_4__7459_ (
);

FILL FILL_4__7039_ (
);

BUFX2 BUFX2_insert226 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf3 )
);

BUFX2 BUFX2_insert227 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf2 )
);

FILL FILL_2__11779_ (
);

BUFX2 BUFX2_insert228 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf1 )
);

FILL FILL_2__11359_ (
);

BUFX2 BUFX2_insert229 (
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf0 )
);

FILL FILL_0__12393_ (
);

FILL SFILL33880x15050 (
);

FILL FILL_4__8400_ (
);

FILL FILL_2__12720_ (
);

FILL FILL_5__15585_ (
);

FILL SFILL33400x44050 (
);

FILL SFILL49000x29050 (
);

FILL FILL_2__12300_ (
);

FILL FILL_5__15165_ (
);

FILL FILL_0__7359_ (
);

INVX1 _9885_ (
    .A(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_1523_)
);

INVX1 _9465_ (
    .A(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_1304_)
);

OAI21X1 _9045_ (
    .A(_1104_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1105_),
    .Y(_1043_[31])
);

FILL FILL_4__14998_ (
);

FILL FILL_4__14578_ (
);

FILL FILL_1__11713_ (
);

FILL FILL_4__14158_ (
);

FILL FILL_2__15192_ (
);

FILL SFILL94440x38050 (
);

FILL FILL_0__8720_ (
);

FILL FILL_2__8738_ (
);

FILL FILL_0__10706_ (
);

FILL FILL_2__8318_ (
);

FILL FILL_1__14185_ (
);

FILL FILL_0__13598_ (
);

AOI21X1 _13883_ (
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .B(_4225_),
    .C(_4386_),
    .Y(_4387_)
);

FILL SFILL84520x74050 (
);

INVX1 _13463_ (
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_3975_)
);

FILL SFILL23880x58050 (
);

OAI21X1 _13043_ (
    .A(_3679_),
    .B(vdd),
    .C(_3680_),
    .Y(_3620_[30])
);

FILL FILL_3__14932_ (
);

FILL FILL_3__14512_ (
);

FILL FILL_4__9605_ (
);

FILL FILL_2__13925_ (
);

FILL FILL_2__13505_ (
);

FILL FILL_5__11085_ (
);

FILL SFILL84120x60050 (
);

FILL FILL_1__12918_ (
);

FILL FILL_2__16397_ (
);

FILL FILL_4__10498_ (
);

FILL FILL_0__9925_ (
);

FILL FILL_0__9505_ (
);

FILL FILL_3__7602_ (
);

FILL FILL_5__7948_ (
);

FILL FILL_5__7108_ (
);

FILL FILL_4__16304_ (
);

NOR2X1 _14668_ (
    .A(_5144_),
    .B(_5154_),
    .Y(_5155_)
);

INVX1 _14248_ (
    .A(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_4744_)
);

FILL FILL_3__15717_ (
);

FILL SFILL8040x72050 (
);

FILL FILL_1__16331_ (
);

FILL SFILL79320x5050 (
);

FILL SFILL23880x13050 (
);

FILL FILL_3__10432_ (
);

FILL FILL_3__10012_ (
);

FILL FILL_0__15744_ (
);

FILL FILL_0__15324_ (
);

FILL SFILL53960x6050 (
);

FILL FILL_2__8491_ (
);

FILL FILL_2__8071_ (
);

FILL FILL_5__13651_ (
);

FILL FILL_5__13231_ (
);

NAND2X1 _7951_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_539_)
);

DFFSR _7531_ (
    .Q(\datapath_1.regfile_1.regOut[5] [21]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_263_[21])
);

INVX1 _7111_ (
    .A(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_121_)
);

FILL FILL_4__12644_ (
);

FILL FILL_4__12224_ (
);

DFFSR _10588_ (
    .Q(\datapath_1.regfile_1.regOut[29] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_1823_[6])
);

INVX1 _10168_ (
    .A(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_1671_)
);

FILL SFILL23800x11050 (
);

FILL FILL_3__11637_ (
);

FILL FILL_3__11217_ (
);

FILL FILL_1__12251_ (
);

FILL FILL_0__16109_ (
);

FILL FILL_2__9276_ (
);

FILL FILL_0__11664_ (
);

FILL FILL_0__11244_ (
);

FILL FILL_5__14856_ (
);

FILL FILL_3__15890_ (
);

FILL FILL_5__14436_ (
);

FILL FILL_5__14016_ (
);

FILL FILL_3__15470_ (
);

INVX1 _8736_ (
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_940_)
);

FILL FILL_3__15050_ (
);

INVX1 _8316_ (
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_721_)
);

FILL FILL_1__7693_ (
);

FILL FILL_4__13849_ (
);

FILL FILL_4__13429_ (
);

FILL FILL_2__14883_ (
);

FILL FILL_2__14463_ (
);

FILL FILL_4__13009_ (
);

FILL FILL_2__14043_ (
);

FILL FILL_3__7199_ (
);

FILL SFILL8760x17050 (
);

FILL SFILL13800x54050 (
);

FILL FILL_1__13876_ (
);

FILL FILL_1__13456_ (
);

FILL FILL_1__13036_ (
);

FILL FILL_3__8980_ (
);

FILL FILL_0__12869_ (
);

INVX1 _12734_ (
    .A(\datapath_1.PCJump [15]),
    .Y(_3515_)
);

FILL FILL_0__12449_ (
);

FILL FILL_3__8140_ (
);

FILL FILL_0__12029_ (
);

NAND3X1 _12314_ (
    .A(_3272_),
    .B(_3273_),
    .C(_3274_),
    .Y(\datapath_1.alu_1.ALUInB [24])
);

FILL FILL_5__8486_ (
);

FILL SFILL114600x17050 (
);

FILL FILL_5__8066_ (
);

FILL FILL_0__13810_ (
);

FILL FILL_3__16255_ (
);

FILL FILL_5__10776_ (
);

FILL FILL_1__8898_ (
);

FILL FILL_1__8478_ (
);

FILL FILL_3__11390_ (
);

FILL FILL_1__8058_ (
);

FILL FILL_2__15668_ (
);

FILL FILL_2__15248_ (
);

FILL FILL_0__16282_ (
);

FILL FILL_2__10383_ (
);

FILL FILL_3__9765_ (
);

FILL FILL_3__9345_ (
);

INVX1 _13939_ (
    .A(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_4441_)
);

NAND2X1 _13519_ (
    .A(_4029_),
    .B(_4022_),
    .Y(_4030_)
);

FILL FILL_1__15602_ (
);

FILL FILL_6__12568_ (
);

FILL FILL_2__7762_ (
);

FILL FILL_3__12595_ (
);

FILL FILL_2__7342_ (
);

FILL FILL_3__12175_ (
);

FILL FILL_4__7688_ (
);

FILL FILL112360x54050 (
);

FILL FILL_2__11588_ (
);

FILL FILL_2__11168_ (
);

FILL FILL_5__12502_ (
);

FILL SFILL89480x7050 (
);

FILL FILL_4__11915_ (
);

FILL FILL_5__15394_ (
);

FILL FILL_0__7588_ (
);

DFFSR _9694_ (
    .Q(\datapath_1.regfile_1.regOut[22] [8]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_1368_[8])
);

FILL FILL_0__7168_ (
);

OAI21X1 _9274_ (
    .A(_1216_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .C(_1217_),
    .Y(_1173_[22])
);

FILL FILL_3__10908_ (
);

FILL FILL_1__11942_ (
);

FILL SFILL88840x4050 (
);

FILL FILL_4__14387_ (
);

FILL FILL_1__11522_ (
);

FILL FILL_1__11102_ (
);

FILL FILL_2__8967_ (
);

FILL FILL_0__10935_ (
);

FILL FILL_2__8127_ (
);

NAND2X1 _10800_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1991_)
);

FILL FILL_0__10515_ (
);

FILL FILL_5__6972_ (
);

INVX1 _13692_ (
    .A(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_4199_)
);

NOR2X1 _13272_ (
    .A(_3799_),
    .B(_3812_),
    .Y(_3813_)
);

FILL FILL_5__13707_ (
);

FILL FILL_3__14741_ (
);

FILL FILL_3__14321_ (
);

FILL FILL_1__6964_ (
);

FILL FILL_4__9414_ (
);

FILL FILL_2__13734_ (
);

FILL FILL_2__13314_ (
);

FILL FILL_5__16179_ (
);

FILL FILL_1__12727_ (
);

FILL FILL_1__12307_ (
);

FILL FILL_3__7831_ (
);

FILL FILL_0__9734_ (
);

FILL FILL112280x16050 (
);

FILL FILL_1__15199_ (
);

FILL FILL_5__7757_ (
);

FILL FILL_2_BUFX2_insert910 (
);

FILL FILL_5__7337_ (
);

FILL FILL_4__16113_ (
);

FILL FILL_2_BUFX2_insert911 (
);

FILL FILL_2_BUFX2_insert912 (
);

OAI22X1 _14897_ (
    .A(_3916_),
    .B(_5377_),
    .C(_5378_),
    .D(_3972__bF$buf3),
    .Y(_5379_)
);

FILL FILL_2_BUFX2_insert913 (
);

INVX1 _14477_ (
    .A(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_4968_)
);

FILL FILL_2_BUFX2_insert914 (
);

INVX1 _14057_ (
    .A(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_4557_)
);

FILL FILL_2_BUFX2_insert915 (
);

FILL FILL_2_BUFX2_insert916 (
);

FILL FILL_3__15946_ (
);

FILL FILL_3__15526_ (
);

FILL FILL_2_BUFX2_insert917 (
);

FILL FILL_2_BUFX2_insert918 (
);

FILL FILL_3__15106_ (
);

FILL FILL_2_BUFX2_insert919 (
);

FILL FILL_1__16140_ (
);

FILL FILL_1__7749_ (
);

FILL FILL_3__10661_ (
);

FILL FILL_1__7329_ (
);

FILL FILL_3__10241_ (
);

FILL FILL_2__14939_ (
);

FILL FILL_0__15973_ (
);

FILL FILL_2__14519_ (
);

FILL FILL_0__15553_ (
);

FILL FILL_0__15133_ (
);

FILL FILL_5__12099_ (
);

FILL SFILL54040x61050 (
);

FILL FILL_3__8616_ (
);

FILL FILL_5__13880_ (
);

FILL FILL_5__13460_ (
);

FILL SFILL115080x49050 (
);

FILL FILL_5__13040_ (
);

INVX1 _7760_ (
    .A(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_452_)
);

INVX1 _7340_ (
    .A(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_233_)
);

FILL FILL_4__12873_ (
);

FILL FILL_4__12453_ (
);

FILL FILL_4__12033_ (
);

INVX1 _10397_ (
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_1783_)
);

FILL FILL_5__9903_ (
);

FILL FILL_3__11866_ (
);

FILL FILL_3__11446_ (
);

FILL FILL_1__12480_ (
);

FILL FILL_3__11026_ (
);

FILL FILL_1__12060_ (
);

FILL FILL_4__6959_ (
);

FILL FILL_0__16338_ (
);

AOI21X1 _16203_ (
    .A(_6631_),
    .B(_6654_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [28])
);

FILL FILL_0__11893_ (
);

FILL FILL_2__10439_ (
);

FILL FILL_2__10019_ (
);

FILL FILL_2__9085_ (
);

FILL FILL_0__11473_ (
);

FILL FILL_0__11053_ (
);

FILL FILL_5__7090_ (
);

FILL FILL_2__11800_ (
);

FILL FILL_5__14665_ (
);

FILL FILL_0__6859_ (
);

FILL FILL_5__14245_ (
);

INVX1 _8965_ (
    .A(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_1052_)
);

DFFSR _8545_ (
    .Q(\datapath_1.regfile_1.regOut[13] [11]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_783_[11])
);

OAI21X1 _8125_ (
    .A(_633_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .C(_634_),
    .Y(_588_[23])
);

FILL FILL_1__7082_ (
);

FILL FILL_4__13658_ (
);

FILL FILL_4__13238_ (
);

FILL FILL_2__14692_ (
);

FILL FILL_2__14272_ (
);

FILL FILL_2__7818_ (
);

FILL FILL_0__7800_ (
);

FILL FILL_1__13685_ (
);

FILL FILL_1__13265_ (
);

FILL FILL_1_BUFX2_insert930 (
);

FILL FILL_1_BUFX2_insert931 (
);

INVX1 _12963_ (
    .A(_2_[4]),
    .Y(_3627_)
);

FILL FILL_1_BUFX2_insert932 (
);

DFFSR _12543_ (
    .Q(ALUOut[8]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3360_[8])
);

FILL FILL_0__12258_ (
);

FILL FILL_1_BUFX2_insert933 (
);

OAI21X1 _12123_ (
    .A(_3134_),
    .B(ALUSrcA_bF$buf3),
    .C(_3135_),
    .Y(\datapath_1.alu_1.ALUInA [2])
);

FILL FILL_1_BUFX2_insert934 (
);

FILL FILL_1_BUFX2_insert935 (
);

FILL FILL_1_BUFX2_insert936 (
);

FILL SFILL48760x81050 (
);

FILL FILL_1_BUFX2_insert937 (
);

FILL SFILL79160x72050 (
);

FILL FILL_1_BUFX2_insert938 (
);

FILL FILL_1_BUFX2_insert939 (
);

FILL FILL_3__16064_ (
);

FILL FILL_5__10165_ (
);

FILL FILL_2__15897_ (
);

FILL FILL_2__15477_ (
);

FILL FILL_2__15057_ (
);

FILL FILL_0__16091_ (
);

FILL FILL_2__10192_ (
);

FILL FILL_4__15804_ (
);

FILL FILL_3__9994_ (
);

OAI22X1 _13748_ (
    .A(_4253_),
    .B(_3902__bF$buf1),
    .C(_3966__bF$buf3),
    .D(_4252_),
    .Y(_4254_)
);

FILL FILL_3__9154_ (
);

NAND2X1 _13328_ (
    .A(_3777_),
    .B(_3752_),
    .Y(_3855_)
);

FILL SFILL109480x6050 (
);

FILL FILL_1__15831_ (
);

FILL FILL_1__15411_ (
);

FILL FILL_6__12377_ (
);

FILL FILL_0__14824_ (
);

FILL FILL_0__14404_ (
);

FILL FILL_2__7991_ (
);

BUFX2 BUFX2_insert600 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf7)
);

FILL FILL_2__7571_ (
);

BUFX2 BUFX2_insert601 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf6)
);

BUFX2 BUFX2_insert602 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf5)
);

BUFX2 BUFX2_insert603 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf4)
);

BUFX2 BUFX2_insert604 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf3)
);

BUFX2 BUFX2_insert605 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf2)
);

FILL FILL_4__7497_ (
);

FILL FILL_4__7077_ (
);

BUFX2 BUFX2_insert606 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf1)
);

BUFX2 BUFX2_insert607 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf0)
);

BUFX2 BUFX2_insert608 (
    .A(_5515_),
    .Y(_5515__bF$buf3)
);

FILL FILL_2__11397_ (
);

BUFX2 BUFX2_insert609 (
    .A(_5515_),
    .Y(_5515__bF$buf2)
);

FILL FILL_5__12731_ (
);

FILL FILL_5__12311_ (
);

FILL FILL_4__11724_ (
);

FILL FILL_4__11304_ (
);

FILL FILL_6__8784_ (
);

OAI21X1 _9083_ (
    .A(_1109_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .C(_1110_),
    .Y(_1108_[1])
);

FILL FILL_1__11751_ (
);

FILL FILL_4__14196_ (
);

FILL FILL_1__11331_ (
);

FILL FILL_0__15609_ (
);

FILL FILL_2__8776_ (
);

FILL FILL_2__8356_ (
);

FILL FILL_0__10744_ (
);

FILL FILL_0__10324_ (
);

FILL FILL_6__14943_ (
);

FILL FILL_6__14523_ (
);

FILL SFILL74120x53050 (
);

OAI21X1 _13081_ (
    .A(_3748_),
    .B(PCEn_bF$buf4),
    .C(_3749_),
    .Y(_3685_[0])
);

FILL FILL_5__13936_ (
);

FILL FILL_3__14970_ (
);

FILL FILL_5__13516_ (
);

FILL SFILL74920x36050 (
);

FILL FILL_3__14550_ (
);

INVX1 _7816_ (
    .A(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_469_)
);

FILL FILL_3__14130_ (
);

FILL FILL_4_BUFX2_insert440 (
);

FILL FILL_4__9643_ (
);

FILL FILL_4_BUFX2_insert441 (
);

FILL FILL_4_BUFX2_insert442 (
);

FILL FILL_4__9223_ (
);

FILL FILL_4__12509_ (
);

FILL FILL_4_BUFX2_insert443 (
);

FILL FILL_2__13963_ (
);

FILL FILL_4_BUFX2_insert444 (
);

FILL FILL_2__13543_ (
);

FILL FILL_4_BUFX2_insert445 (
);

FILL FILL_2__13123_ (
);

FILL FILL_6__9989_ (
);

FILL FILL_4_BUFX2_insert446 (
);

FILL FILL_4_BUFX2_insert447 (
);

FILL SFILL13800x49050 (
);

FILL FILL_4_BUFX2_insert448 (
);

FILL FILL_4_BUFX2_insert449 (
);

FILL FILL_1__12956_ (
);

FILL FILL_1__12116_ (
);

FILL FILL_0__11949_ (
);

FILL FILL_0__9543_ (
);

FILL FILL_0__9123_ (
);

OAI22X1 _11814_ (
    .A(_2122_),
    .B(_2346_),
    .C(_2347__bF$buf2),
    .D(_2355_),
    .Y(_2905_)
);

FILL FILL_3__7220_ (
);

FILL FILL_0__11529_ (
);

FILL FILL_0__11109_ (
);

FILL FILL_5__7986_ (
);

FILL FILL_5__7566_ (
);

FILL FILL_4__16342_ (
);

AOI21X1 _14286_ (
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .B(_4225_),
    .C(_4780_),
    .Y(_4781_)
);

FILL FILL_3__15755_ (
);

FILL FILL_3__15335_ (
);

FILL FILL_1__7978_ (
);

FILL FILL_3__10890_ (
);

FILL FILL_1__7558_ (
);

FILL FILL_3__10050_ (
);

FILL SFILL28840x2050 (
);

FILL FILL_2__14748_ (
);

FILL FILL_0__15782_ (
);

FILL FILL_2__14328_ (
);

FILL FILL_0__15362_ (
);

FILL SFILL28760x7050 (
);

FILL FILL_3__8845_ (
);

FILL FILL_3__8005_ (
);

FILL SFILL8680x3050 (
);

FILL FILL_4__12262_ (
);

FILL SFILL64120x51050 (
);

FILL FILL_2__6842_ (
);

FILL FILL_3__11675_ (
);

FILL FILL_3__11255_ (
);

DFFSR _16432_ (
    .Q(\datapath_1.regfile_1.regOut[0] [15]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_6769_[15])
);

FILL FILL_0__16147_ (
);

FILL FILL112360x49050 (
);

NAND3X1 _16012_ (
    .A(_6466_),
    .B(_6467_),
    .C(_6465_),
    .Y(_6468_)
);

FILL FILL_2__10668_ (
);

FILL FILL_2__10248_ (
);

FILL FILL_0__11282_ (
);

FILL FILL_3_BUFX2_insert460 (
);

FILL FILL_3_BUFX2_insert461 (
);

FILL SFILL64040x58050 (
);

FILL FILL_3_BUFX2_insert462 (
);

FILL FILL_5__14894_ (
);

FILL FILL_5__14474_ (
);

FILL FILL_3_BUFX2_insert463 (
);

FILL FILL_5__14054_ (
);

FILL FILL_3_BUFX2_insert464 (
);

OAI21X1 _8774_ (
    .A(_964_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_965_),
    .Y(_913_[26])
);

FILL FILL_3_BUFX2_insert465 (
);

FILL FILL_3_BUFX2_insert466 (
);

OAI21X1 _8354_ (
    .A(_745_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_746_),
    .Y(_718_[14])
);

FILL FILL_3_BUFX2_insert467 (
);

FILL FILL_3_BUFX2_insert468 (
);

FILL FILL_4__13887_ (
);

FILL FILL_3_BUFX2_insert469 (
);

FILL FILL_4__13467_ (
);

FILL FILL_2__14081_ (
);

FILL FILL_2__7627_ (
);

FILL FILL_2__7207_ (
);

FILL FILL_1__13494_ (
);

OAI21X1 _12772_ (
    .A(_3539_),
    .B(IRWrite_bF$buf3),
    .C(_3540_),
    .Y(_3490_[25])
);

FILL FILL_0__12487_ (
);

INVX1 _12352_ (
    .A(ALUOut[3]),
    .Y(_3300_)
);

FILL FILL_0__12067_ (
);

FILL FILL_3__13821_ (
);

FILL FILL_3__13401_ (
);

FILL FILL_4__8914_ (
);

FILL FILL_5__15679_ (
);

FILL FILL_5__15259_ (
);

FILL FILL_3__16293_ (
);

OAI21X1 _9979_ (
    .A(_1564_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1565_),
    .Y(_1563_[1])
);

DFFSR _9559_ (
    .Q(\datapath_1.regfile_1.regOut[21] [1]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_1303_[1])
);

NAND2X1 _9139_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1148_)
);

FILL SFILL64040x13050 (
);

FILL FILL_5__10394_ (
);

FILL FILL_1__8096_ (
);

FILL FILL_1__11807_ (
);

FILL FILL_2__15286_ (
);

FILL FILL_3__6911_ (
);

FILL FILL_5__16200_ (
);

FILL SFILL89240x62050 (
);

FILL FILL_1__14699_ (
);

FILL FILL_1__14279_ (
);

FILL FILL_5__6837_ (
);

FILL FILL_0_BUFX2_insert590 (
);

FILL FILL_4__15613_ (
);

FILL FILL_0_BUFX2_insert591 (
);

FILL FILL_0_BUFX2_insert592 (
);

FILL FILL_0_BUFX2_insert593 (
);

FILL FILL_0_BUFX2_insert594 (
);

FILL FILL_3__9383_ (
);

INVX1 _13977_ (
    .A(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_4478_)
);

FILL FILL_0_BUFX2_insert595 (
);

OAI22X1 _13557_ (
    .A(_4065_),
    .B(_3955__bF$buf2),
    .C(_3924__bF$buf1),
    .D(_4066_),
    .Y(_4067_)
);

FILL FILL_0_BUFX2_insert596 (
);

NAND2X1 _13137_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [19]),
    .Y(_3723_)
);

FILL FILL_0_BUFX2_insert597 (
);

FILL FILL_3__14606_ (
);

FILL FILL_0_BUFX2_insert598 (
);

FILL FILL_1__15640_ (
);

FILL FILL_0_BUFX2_insert599 (
);

FILL FILL_1__15220_ (
);

FILL FILL_0__14633_ (
);

FILL FILL_0__14213_ (
);

FILL FILL_5__11599_ (
);

FILL SFILL54040x56050 (
);

FILL FILL_2__7380_ (
);

FILL FILL_5__11179_ (
);

FILL FILL_5__12960_ (
);

FILL FILL_5__12120_ (
);

BUFX2 _6840_ (
    .A(_1_[2]),
    .Y(memoryAddress[2])
);

FILL FILL_4__11953_ (
);

FILL FILL_4__11533_ (
);

FILL FILL_4__11113_ (
);

FILL FILL_1__16005_ (
);

FILL FILL_3__10946_ (
);

FILL FILL_1__11980_ (
);

FILL FILL_3__10526_ (
);

FILL FILL_1__11560_ (
);

FILL FILL_3__10106_ (
);

FILL FILL_1__11140_ (
);

FILL FILL_0__15838_ (
);

AOI22X1 _15703_ (
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .B(_5494_),
    .C(_5479_),
    .D(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_6167_)
);

FILL FILL_0__15418_ (
);

FILL FILL_0__10973_ (
);

FILL FILL_2__8585_ (
);

FILL FILL_0__10553_ (
);

FILL FILL_0__10133_ (
);

FILL SFILL54040x11050 (
);

FILL FILL_5__13745_ (
);

FILL FILL_5__13325_ (
);

OAI21X1 _7625_ (
    .A(_381_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .C(_382_),
    .Y(_328_[27])
);

OAI21X1 _7205_ (
    .A(_162_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .C(_163_),
    .Y(_133_[15])
);

FILL FILL_4__9872_ (
);

FILL FILL_4__12738_ (
);

FILL FILL_4__9032_ (
);

FILL FILL_2__13772_ (
);

FILL FILL_4__12318_ (
);

FILL FILL_2__13352_ (
);

FILL FILL111880x73050 (
);

FILL FILL_1__12765_ (
);

FILL FILL_1__12345_ (
);

FILL FILL_0__9772_ (
);

FILL FILL_0__9352_ (
);

FILL FILL_0__11758_ (
);

FILL FILL_0__11338_ (
);

OAI21X1 _11623_ (
    .A(_2507_),
    .B(_2518_),
    .C(_2257_),
    .Y(_2728_)
);

NOR2X1 _11203_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2322_)
);

FILL FILL_5__7375_ (
);

FILL FILL_6__15117_ (
);

FILL FILL_4__16151_ (
);

FILL FILL_6__10672_ (
);

NAND3X1 _14095_ (
    .A(_4592_),
    .B(_4593_),
    .C(_4591_),
    .Y(_4594_)
);

FILL FILL_3__15984_ (
);

FILL FILL_3__15564_ (
);

FILL FILL_3__15144_ (
);

FILL FILL_1__7367_ (
);

FILL FILL_2__14977_ (
);

FILL FILL_2__14557_ (
);

FILL FILL_2__14137_ (
);

FILL FILL_0__15591_ (
);

FILL FILL_0__15171_ (
);

FILL FILL_3__8654_ (
);

FILL FILL_3__8234_ (
);

OAI21X1 _12828_ (
    .A(_3556_),
    .B(vdd),
    .C(_3557_),
    .Y(_3555_[1])
);

OAI21X1 _12408_ (
    .A(_3336_),
    .B(MemToReg_bF$buf7),
    .C(_3337_),
    .Y(\datapath_1.mux_wd3.dout [21])
);

FILL SFILL8520x24050 (
);

FILL FILL_1__14911_ (
);

FILL FILL_4__12491_ (
);

FILL FILL_6__11037_ (
);

FILL FILL_4__12071_ (
);

FILL FILL_0__13904_ (
);

FILL FILL_3__16349_ (
);

FILL FILL_5__9941_ (
);

FILL FILL_5__9521_ (
);

FILL FILL_3__11484_ (
);

FILL FILL_5__9101_ (
);

FILL FILL_3__11064_ (
);

FILL FILL_4__6997_ (
);

FILL FILL_0__16376_ (
);

NOR2X1 _16241_ (
    .A(_6689_),
    .B(_6691_),
    .Y(_6692_)
);

FILL FILL_2__10897_ (
);

FILL FILL_2__10057_ (
);

FILL FILL_0__11091_ (
);

FILL FILL_1__9933_ (
);

FILL FILL_5__11811_ (
);

FILL FILL_1__9513_ (
);

FILL FILL_3__9859_ (
);

FILL FILL_3__9019_ (
);

FILL FILL_4__10804_ (
);

FILL FILL_0__6897_ (
);

FILL FILL_5__14283_ (
);

FILL FILL_6__7864_ (
);

OAI21X1 _8583_ (
    .A(_857_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .C(_858_),
    .Y(_848_[5])
);

DFFSR _8163_ (
    .Q(\datapath_1.regfile_1.regOut[10] [13]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_588_[13])
);

FILL FILL_1__10831_ (
);

FILL FILL_4__13696_ (
);

FILL FILL_4__13276_ (
);

FILL FILL_1__10411_ (
);

FILL SFILL69160x65050 (
);

FILL SFILL34040x52050 (
);

FILL FILL_2__7856_ (
);

FILL FILL_2__7436_ (
);

FILL FILL_3__12269_ (
);

FILL SFILL74120x48050 (
);

OAI21X1 _12581_ (
    .A(_3432_),
    .B(vdd),
    .C(_3433_),
    .Y(_3425_[4])
);

FILL FILL_0__12296_ (
);

NAND2X1 _12161_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [15]),
    .Y(_3161_)
);

FILL FILL_3__13630_ (
);

FILL FILL_3__13210_ (
);

FILL FILL_4__8723_ (
);

FILL FILL_2__12623_ (
);

FILL FILL_5__15488_ (
);

FILL FILL_2__12203_ (
);

FILL FILL_5__15068_ (
);

NAND2X1 _9788_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1479_)
);

NAND2X1 _9368_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1260_)
);

FILL FILL_1__11616_ (
);

FILL FILL_2__15095_ (
);

FILL FILL_0__8623_ (
);

FILL FILL_0__8203_ (
);

FILL FILL_1__14088_ (
);

FILL FILL_4__15842_ (
);

FILL FILL_4__15422_ (
);

FILL FILL_4__15002_ (
);

NOR2X1 _13786_ (
    .A(_4291_),
    .B(_4288_),
    .Y(_4292_)
);

INVX1 _13366_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_3878_)
);

FILL FILL_3__14835_ (
);

FILL FILL_3__14415_ (
);

FILL FILL_4__9928_ (
);

FILL FILL_4__9508_ (
);

FILL FILL_2__13828_ (
);

FILL FILL_0__14862_ (
);

FILL FILL_2__13408_ (
);

FILL FILL_0__14442_ (
);

FILL FILL_0__14022_ (
);

CLKBUF1 CLKBUF1_insert140 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf84)
);

CLKBUF1 CLKBUF1_insert141 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf83)
);

CLKBUF1 CLKBUF1_insert142 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf82)
);

CLKBUF1 CLKBUF1_insert143 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf81)
);

FILL SFILL28760x72050 (
);

CLKBUF1 CLKBUF1_insert144 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf80)
);

FILL FILL_0__9408_ (
);

FILL FILL_3__7505_ (
);

FILL SFILL59160x63050 (
);

CLKBUF1 CLKBUF1_insert145 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf79)
);

CLKBUF1 CLKBUF1_insert146 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf78)
);

CLKBUF1 CLKBUF1_insert147 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf77)
);

CLKBUF1 CLKBUF1_insert148 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf76)
);

CLKBUF1 CLKBUF1_insert149 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf75)
);

FILL FILL_4__16207_ (
);

FILL FILL_4__11762_ (
);

FILL FILL_4__11342_ (
);

FILL SFILL64120x46050 (
);

FILL FILL_1__16234_ (
);

FILL FILL_3__10755_ (
);

FILL FILL_0__15647_ (
);

OAI22X1 _15932_ (
    .A(_6389_),
    .B(_5544__bF$buf3),
    .C(_5523_),
    .D(_4991_),
    .Y(_6390_)
);

FILL FILL_0__15227_ (
);

NOR3X1 _15512_ (
    .A(_5515__bF$buf3),
    .B(_4481_),
    .C(_5521__bF$buf3),
    .Y(_5981_)
);

FILL SFILL28680x79050 (
);

FILL FILL_2__8394_ (
);

FILL FILL_0__10782_ (
);

FILL FILL_0__10362_ (
);

FILL FILL_5__13974_ (
);

FILL FILL_5__13554_ (
);

FILL FILL_5__13134_ (
);

OAI21X1 _7854_ (
    .A(_493_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .C(_494_),
    .Y(_458_[18])
);

OAI21X1 _7434_ (
    .A(_274_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .C(_275_),
    .Y(_263_[6])
);

DFFSR _7014_ (
    .Q(\datapath_1.regfile_1.regOut[1] [16]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_3_[16])
);

FILL FILL_4_BUFX2_insert820 (
);

FILL FILL_4__9681_ (
);

FILL FILL_4_BUFX2_insert821 (
);

FILL FILL_4__9261_ (
);

FILL FILL_4_BUFX2_insert822 (
);

FILL FILL_4__12967_ (
);

FILL FILL_4_BUFX2_insert823 (
);

FILL FILL_4__12127_ (
);

FILL FILL_4_BUFX2_insert824 (
);

FILL FILL_2__13581_ (
);

FILL FILL_4_BUFX2_insert825 (
);

FILL FILL_2__13161_ (
);

FILL SFILL85000x42050 (
);

FILL FILL_4_BUFX2_insert826 (
);

FILL FILL_4_BUFX2_insert827 (
);

FILL SFILL68840x23050 (
);

FILL FILL_4_BUFX2_insert828 (
);

FILL FILL_4_BUFX2_insert829 (
);

FILL FILL_1__12994_ (
);

FILL FILL_1__12574_ (
);

FILL FILL_1__12154_ (
);

FILL FILL_2__9599_ (
);

FILL FILL_0__11987_ (
);

NOR3X1 _11852_ (
    .A(\datapath_1.ALUResult [4]),
    .B(\datapath_1.ALUResult [3]),
    .C(_2938_),
    .Y(_2939_)
);

FILL FILL_0__11567_ (
);

FILL FILL_0__9161_ (
);

FILL FILL_0__11147_ (
);

INVX2 _11432_ (
    .A(_2407_),
    .Y(_2548_)
);

FILL SFILL89320x50050 (
);

AOI22X1 _11012_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(_2128_),
    .C(_2130_),
    .D(_2129_),
    .Y(_2131_)
);

FILL FILL_3__12901_ (
);

FILL FILL_6__15766_ (
);

FILL FILL_5__7184_ (
);

FILL FILL_4__16380_ (
);

FILL FILL_5__14759_ (
);

FILL FILL_3__15793_ (
);

FILL FILL_5__14339_ (
);

FILL FILL_3__15373_ (
);

NAND2X1 _8639_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_896_)
);

NAND2X1 _8219_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_677_)
);

FILL FILL_1__7596_ (
);

FILL FILL_1__7176_ (
);

FILL FILL_2__14786_ (
);

FILL FILL_2__14366_ (
);

FILL FILL_5__15700_ (
);

FILL SFILL89240x57050 (
);

FILL SFILL54120x44050 (
);

FILL FILL_1__13779_ (
);

FILL FILL_1__13359_ (
);

FILL FILL_3__8883_ (
);

FILL FILL_3__8463_ (
);

NAND2X1 _12637_ (
    .A(vdd),
    .B(memoryOutData[23]),
    .Y(_3471_)
);

AOI22X1 _12217_ (
    .A(_2_[0]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf2),
    .D(gnd),
    .Y(_3202_)
);

FILL SFILL18680x77050 (
);

FILL FILL_5__8389_ (
);

FILL FILL_1__14720_ (
);

FILL FILL_1__14300_ (
);

FILL FILL_6__11686_ (
);

FILL FILL_0__13713_ (
);

FILL FILL_3__16158_ (
);

FILL SFILL89640x26050 (
);

FILL FILL_5__10679_ (
);

FILL FILL_2__6880_ (
);

FILL FILL_5__9750_ (
);

FILL FILL_5__10259_ (
);

FILL FILL_3__11293_ (
);

FILL FILL_0__16185_ (
);

NOR3X1 _16050_ (
    .A(_6504_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6505_)
);

FILL FILL_2__10286_ (
);

FILL FILL_1__9742_ (
);

FILL FILL_5__11620_ (
);

FILL FILL_5__11200_ (
);

FILL SFILL89240x12050 (
);

FILL FILL_3__9668_ (
);

FILL FILL_3_BUFX2_insert840 (
);

FILL FILL_3__9248_ (
);

FILL FILL_3_BUFX2_insert841 (
);

FILL FILL_3_BUFX2_insert842 (
);

FILL FILL_3_BUFX2_insert843 (
);

FILL FILL_3_BUFX2_insert844 (
);

FILL FILL_5__14092_ (
);

FILL FILL_1__15925_ (
);

FILL FILL_3_BUFX2_insert845 (
);

FILL FILL_1__15505_ (
);

NAND2X1 _8392_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_772_)
);

FILL FILL_3_BUFX2_insert846 (
);

FILL FILL_3_BUFX2_insert847 (
);

FILL FILL_3_BUFX2_insert848 (
);

FILL FILL_3_BUFX2_insert849 (
);

FILL SFILL18680x32050 (
);

FILL FILL_1__10640_ (
);

FILL FILL_4__13085_ (
);

FILL FILL_0__14918_ (
);

FILL FILL_2__7245_ (
);

FILL FILL_3__12498_ (
);

FILL FILL_3__12078_ (
);

FILL FILL111960x61050 (
);

OAI21X1 _12390_ (
    .A(_3324_),
    .B(MemToReg_bF$buf5),
    .C(_3325_),
    .Y(\datapath_1.mux_wd3.dout [15])
);

FILL FILL_5__12825_ (
);

FILL FILL_5__12405_ (
);

FILL FILL_4__8952_ (
);

FILL FILL_4__8532_ (
);

FILL FILL_4__8112_ (
);

FILL FILL_4__11818_ (
);

FILL FILL_2__12852_ (
);

FILL FILL_2__12432_ (
);

FILL FILL_5__15297_ (
);

FILL FILL_2__12012_ (
);

FILL FILL_6__8878_ (
);

NAND2X1 _9597_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1372_)
);

DFFSR _9177_ (
    .Q(\datapath_1.regfile_1.regOut[18] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_1108_[3])
);

FILL FILL_1__11845_ (
);

FILL FILL_1__11425_ (
);

FILL FILL_1__11005_ (
);

FILL FILL_0__8852_ (
);

OAI21X1 _10703_ (
    .A(_1945_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1946_),
    .Y(_1888_[29])
);

FILL FILL_0__8012_ (
);

FILL FILL_0__10418_ (
);

FILL FILL_0_BUFX2_insert970 (
);

FILL FILL_5__6875_ (
);

FILL SFILL44040x49050 (
);

FILL FILL_0_BUFX2_insert971 (
);

FILL FILL_4__15651_ (
);

FILL FILL_0_BUFX2_insert972 (
);

FILL FILL_4__15231_ (
);

FILL FILL_0_BUFX2_insert973 (
);

FILL FILL_0_BUFX2_insert974 (
);

NAND3X1 _13595_ (
    .A(_4101_),
    .B(_4103_),
    .C(_4100_),
    .Y(_4104_)
);

FILL FILL_0_BUFX2_insert975 (
);

DFFSR _13175_ (
    .Q(\datapath_1.mux_iord.din0 [0]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3685_[0])
);

FILL FILL_0_BUFX2_insert976 (
);

FILL FILL_0_BUFX2_insert977 (
);

FILL FILL_2__9811_ (
);

FILL FILL_3__14644_ (
);

FILL FILL_0_BUFX2_insert978 (
);

FILL FILL_3__14224_ (
);

FILL FILL_0_BUFX2_insert979 (
);

FILL FILL_1__6867_ (
);

FILL FILL_4__9737_ (
);

FILL FILL_2__13637_ (
);

FILL FILL_2__13217_ (
);

FILL FILL_0__14671_ (
);

FILL FILL_0__14251_ (
);

FILL FILL_3__7734_ (
);

FILL FILL_0__9637_ (
);

FILL FILL_0__9217_ (
);

INVX1 _11908_ (
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_2980_)
);

FILL FILL_3__7314_ (
);

FILL SFILL8520x19050 (
);

FILL FILL_4__16016_ (
);

FILL FILL_4__11991_ (
);

FILL FILL_4__11571_ (
);

FILL FILL_4__11151_ (
);

FILL FILL_3__15849_ (
);

FILL FILL_3__15429_ (
);

FILL FILL_3__15009_ (
);

FILL FILL_1__16043_ (
);

FILL FILL_5__8601_ (
);

FILL FILL_3__10564_ (
);

FILL FILL_3__10144_ (
);

FILL FILL_6_BUFX2_insert352 (
);

FILL FILL_0__15876_ (
);

FILL SFILL69240x53050 (
);

OAI22X1 _15741_ (
    .A(_4795_),
    .B(_5539__bF$buf2),
    .C(_5469__bF$buf2),
    .D(_4765_),
    .Y(_6204_)
);

FILL FILL_0__15456_ (
);

OAI22X1 _15321_ (
    .A(_5530__bF$buf3),
    .B(_5794_),
    .C(_5532__bF$buf0),
    .D(_5793_),
    .Y(_5795_)
);

FILL FILL_0__15036_ (
);

FILL SFILL109000x22050 (
);

FILL FILL_6_BUFX2_insert357 (
);

FILL FILL_0__10171_ (
);

FILL FILL_6__14370_ (
);

FILL SFILL114680x56050 (
);

FILL FILL_3__8519_ (
);

FILL FILL_5__13783_ (
);

FILL FILL_5__13363_ (
);

DFFSR _7663_ (
    .Q(\datapath_1.regfile_1.regOut[6] [25]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_328_[25])
);

NAND2X1 _7243_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_189_)
);

FILL FILL_4__9490_ (
);

FILL FILL_4__12776_ (
);

FILL FILL_4__12356_ (
);

FILL FILL_2__13390_ (
);

FILL FILL_2__6936_ (
);

FILL FILL_5__9806_ (
);

FILL FILL_3__11769_ (
);

FILL FILL_3__11349_ (
);

FILL FILL_1__12383_ (
);

OAI22X1 _16106_ (
    .A(_5480__bF$buf2),
    .B(_5192_),
    .C(_5189_),
    .D(_5569_),
    .Y(_6560_)
);

FILL FILL_0__9390_ (
);

FILL FILL_0__11796_ (
);

FILL FILL_0__11376_ (
);

NAND3X1 _11661_ (
    .A(_2747_),
    .B(_2751_),
    .C(_2763_),
    .Y(\datapath_1.ALUResult [15])
);

NAND3X1 _11241_ (
    .A(_2359_),
    .B(_2353_),
    .C(_2356_),
    .Y(_2360_)
);

FILL FILL_3__12710_ (
);

FILL FILL_4__7803_ (
);

FILL FILL_5__14988_ (
);

FILL FILL_5__14568_ (
);

FILL FILL_2__11703_ (
);

FILL FILL_5__14148_ (
);

NAND2X1 _8868_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1008_)
);

FILL FILL_3__15182_ (
);

NAND2X1 _8448_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_789_)
);

DFFSR _8028_ (
    .Q(\datapath_1.regfile_1.regOut[9] [6]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_523_[6])
);

FILL FILL_2__14595_ (
);

FILL FILL_2__14175_ (
);

FILL SFILL99400x40050 (
);

FILL SFILL69160x15050 (
);

FILL FILL_0__7703_ (
);

FILL FILL_1__13588_ (
);

FILL FILL_1__13168_ (
);

FILL FILL_4__14922_ (
);

FILL FILL_4__14502_ (
);

NAND2X1 _12866_ (
    .A(vdd),
    .B(\datapath_1.rd1 [14]),
    .Y(_3583_)
);

FILL FILL_3__8272_ (
);

NAND2X1 _12446_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [2]),
    .Y(_3364_)
);

NAND3X1 _12026_ (
    .A(_3063_),
    .B(_3064_),
    .C(_3065_),
    .Y(\datapath_1.mux_pcsrc.dout [9])
);

FILL FILL_3__13915_ (
);

FILL FILL_5__8198_ (
);

FILL FILL_5_BUFX2_insert370 (
);

FILL FILL_2__12908_ (
);

FILL FILL_5_BUFX2_insert371 (
);

FILL SFILL99320x47050 (
);

FILL FILL_5_BUFX2_insert372 (
);

FILL FILL_0__13942_ (
);

FILL FILL_5_BUFX2_insert373 (
);

FILL FILL_3__16387_ (
);

FILL FILL_0__13522_ (
);

FILL FILL_0__13102_ (
);

FILL FILL_5_BUFX2_insert374 (
);

FILL FILL_5_BUFX2_insert375 (
);

FILL FILL_5__10488_ (
);

FILL FILL_5_BUFX2_insert376 (
);

FILL FILL_5__10068_ (
);

FILL FILL_5_BUFX2_insert377 (
);

FILL FILL_5_BUFX2_insert378 (
);

FILL FILL_5_BUFX2_insert379 (
);

FILL SFILL89400x83050 (
);

FILL SFILL28760x67050 (
);

FILL FILL_0__8908_ (
);

FILL SFILL59160x58050 (
);

FILL FILL_1__9551_ (
);

FILL FILL_1__9131_ (
);

FILL FILL_4__15707_ (
);

FILL FILL_2__16321_ (
);

FILL FILL_3__9897_ (
);

FILL FILL_3__9477_ (
);

FILL FILL_4__10422_ (
);

FILL FILL_4__10002_ (
);

FILL FILL_6__7482_ (
);

FILL FILL_1__15734_ (
);

FILL FILL_1__15314_ (
);

FILL SFILL89800x52050 (
);

FILL FILL_0__14727_ (
);

FILL FILL_0__14307_ (
);

FILL FILL_2__7474_ (
);

FILL FILL_2__7054_ (
);

FILL FILL_5__12634_ (
);

FILL FILL_5__12214_ (
);

FILL SFILL28760x22050 (
);

OAI21X1 _6934_ (
    .A(_22_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_23_),
    .Y(_3_[10])
);

FILL SFILL59160x13050 (
);

FILL FILL_4__8761_ (
);

FILL FILL_4__8341_ (
);

FILL FILL_4__11627_ (
);

FILL FILL_2__12661_ (
);

FILL FILL_4__11207_ (
);

FILL FILL_2__12241_ (
);

FILL FILL_6__8267_ (
);

FILL FILL_1__11654_ (
);

FILL FILL_1__11234_ (
);

FILL FILL_4__14099_ (
);

FILL FILL_0__8661_ (
);

INVX1 _10932_ (
    .A(\control_1.op [1]),
    .Y(_2066_)
);

FILL FILL_0__10647_ (
);

FILL FILL_0__8241_ (
);

FILL FILL_2__8259_ (
);

FILL SFILL89320x45050 (
);

OAI21X1 _10512_ (
    .A(_1838_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .C(_1839_),
    .Y(_1823_[8])
);

FILL FILL_6__14846_ (
);

FILL FILL_6__14426_ (
);

FILL FILL_4__15880_ (
);

FILL FILL_4__15460_ (
);

FILL FILL_4__15040_ (
);

FILL FILL_5__13839_ (
);

FILL FILL_3__14873_ (
);

FILL FILL_5__13419_ (
);

FILL FILL_2__9620_ (
);

FILL FILL_3__14453_ (
);

FILL SFILL18760x65050 (
);

NAND2X1 _7719_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_425_)
);

FILL FILL_3__14033_ (
);

FILL FILL_4__9546_ (
);

FILL FILL_4__9126_ (
);

FILL FILL_2__13866_ (
);

FILL FILL_2__13446_ (
);

FILL FILL_0__14480_ (
);

FILL FILL_2__13026_ (
);

FILL FILL_0__14060_ (
);

FILL FILL_1__12859_ (
);

FILL FILL_1__12439_ (
);

FILL FILL_1__12019_ (
);

FILL FILL_0__9866_ (
);

FILL FILL_3__7963_ (
);

FILL FILL_3__7543_ (
);

FILL FILL_3__7123_ (
);

FILL FILL_0__9026_ (
);

NOR2X1 _11717_ (
    .A(_2815_),
    .B(_2805_),
    .Y(_2816_)
);

FILL FILL_5__7889_ (
);

FILL FILL_1__13800_ (
);

FILL FILL_5__7469_ (
);

FILL FILL_5__7049_ (
);

FILL FILL_4__16245_ (
);

OAI22X1 _14189_ (
    .A(_4684_),
    .B(_3944__bF$buf0),
    .C(_3959_),
    .D(_4685_),
    .Y(_4686_)
);

FILL FILL_4__11380_ (
);

FILL FILL_3__15658_ (
);

FILL FILL_3__15238_ (
);

FILL FILL_1__16272_ (
);

FILL FILL_3__10793_ (
);

FILL FILL_5__8830_ (
);

FILL FILL_3__10373_ (
);

FILL SFILL18760x20050 (
);

AOI22X1 _15970_ (
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .B(_5567_),
    .C(_5565__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_6427_)
);

FILL FILL_0__15685_ (
);

NOR3X1 _15550_ (
    .A(_5515__bF$buf0),
    .B(_4543_),
    .C(_5521__bF$buf2),
    .Y(_6018_)
);

FILL FILL_0__15265_ (
);

AOI22X1 _15130_ (
    .A(_5481_),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .C(\datapath_1.regfile_1.regOut[6] [2]),
    .D(_5565__bF$buf0),
    .Y(_5608_)
);

FILL FILL_5__10700_ (
);

FILL FILL_1__8822_ (
);

FILL FILL_1__8402_ (
);

FILL FILL_3__8748_ (
);

FILL FILL_3__8328_ (
);

FILL FILL_5__13592_ (
);

FILL FILL_5__13172_ (
);

NAND2X1 _7892_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_520_)
);

NAND2X1 _7472_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_301_)
);

NAND2X1 _7052_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_82_)
);

FILL SFILL79320x43050 (
);

FILL SFILL18680x27050 (
);

FILL FILL_4__12585_ (
);

FILL FILL_4__12165_ (
);

FILL FILL_3__11998_ (
);

FILL FILL_5__9615_ (
);

FILL FILL_3__11578_ (
);

FILL FILL111960x56050 (
);

FILL FILL_3__11158_ (
);

FILL FILL_1__12192_ (
);

OAI21X1 _16335_ (
    .A(_6776_),
    .B(gnd),
    .C(_6777_),
    .Y(_6769_[4])
);

INVX1 _11890_ (
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_2968_)
);

AOI21X1 _11470_ (
    .A(_2582_),
    .B(_2584_),
    .C(_2583_),
    .Y(_2585_)
);

FILL FILL_0__11185_ (
);

FILL FILL_5__11905_ (
);

XOR2X1 _11050_ (
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2169_)
);

FILL FILL_1__9607_ (
);

FILL FILL_4__7612_ (
);

FILL FILL_2__11932_ (
);

FILL FILL_5__14797_ (
);

FILL FILL_5__14377_ (
);

FILL FILL_2__11512_ (
);

FILL FILL_6__7958_ (
);

DFFSR _8677_ (
    .Q(\datapath_1.regfile_1.regOut[14] [15]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_848_[15])
);

INVX1 _8257_ (
    .A(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_702_)
);

FILL FILL_1__10925_ (
);

FILL FILL_1__10505_ (
);

FILL FILL_0__7932_ (
);

FILL FILL_1__13397_ (
);

FILL SFILL79640x19050 (
);

FILL SFILL110040x67050 (
);

FILL FILL_4__14731_ (
);

FILL FILL_4__14311_ (
);

FILL FILL111960x11050 (
);

DFFSR _12675_ (
    .Q(\datapath_1.Data [12]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3425_[12])
);

FILL FILL_3__8081_ (
);

NAND3X1 _12255_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3230_)
);

FILL FILL_3__13724_ (
);

FILL FILL_3__13304_ (
);

FILL SFILL114360x75050 (
);

FILL FILL_2__12717_ (
);

FILL FILL_0__13751_ (
);

FILL FILL_0__13331_ (
);

FILL FILL_3__16196_ (
);

FILL FILL_5__10297_ (
);

FILL FILL_2__15189_ (
);

FILL FILL_0__8717_ (
);

FILL FILL_5__16103_ (
);

FILL FILL_1__9780_ (
);

FILL FILL_1__9360_ (
);

FILL FILL_4__15936_ (
);

FILL FILL_4__15516_ (
);

FILL FILL_2__16130_ (
);

FILL FILL_3__9286_ (
);

FILL FILL_4__10651_ (
);

FILL FILL_4__10231_ (
);

FILL FILL_3__14929_ (
);

FILL FILL_3__14509_ (
);

FILL FILL_1__15963_ (
);

FILL FILL_1__15543_ (
);

FILL FILL_6__7291_ (
);

FILL FILL_1__15123_ (
);

FILL SFILL69240x48050 (
);

FILL FILL_0__14956_ (
);

AOI22X1 _14821_ (
    .A(_3882__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [28]),
    .C(\datapath_1.regfile_1.regOut[13] [28]),
    .D(_4051__bF$buf3),
    .Y(_5305_)
);

FILL FILL_0__14536_ (
);

NOR2X1 _14401_ (
    .A(_4883_),
    .B(_4893_),
    .Y(_4894_)
);

FILL FILL_0__14116_ (
);

FILL FILL_5__12863_ (
);

FILL FILL_5__12443_ (
);

FILL FILL_5__12023_ (
);

FILL FILL_4__8990_ (
);

FILL FILL_4__8570_ (
);

FILL FILL_4__11856_ (
);

FILL FILL_2__12890_ (
);

FILL FILL_4__11436_ (
);

FILL FILL_2__12470_ (
);

FILL FILL_4__11016_ (
);

FILL FILL_2__12050_ (
);

FILL FILL_1__16328_ (
);

FILL FILL_3__10429_ (
);

FILL FILL_1__11883_ (
);

FILL FILL_3__10009_ (
);

FILL FILL_1__11463_ (
);

FILL FILL_1__11043_ (
);

OAI22X1 _15606_ (
    .A(_5549__bF$buf1),
    .B(_6072_),
    .C(_5466__bF$buf1),
    .D(_6071_),
    .Y(_6073_)
);

FILL FILL_0__8890_ (
);

FILL FILL_2__8488_ (
);

FILL FILL_0__10876_ (
);

FILL FILL_0__8470_ (
);

FILL SFILL104360x73050 (
);

FILL FILL_2__8068_ (
);

DFFSR _10741_ (
    .Q(\datapath_1.regfile_1.regOut[30] [31]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_1888_[31])
);

NAND2X1 _10321_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1753_)
);

FILL FILL_0__10036_ (
);

FILL FILL_5__13648_ (
);

FILL FILL_5__13228_ (
);

FILL FILL_3__14682_ (
);

NAND2X1 _7948_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_537_)
);

FILL FILL_3__14262_ (
);

DFFSR _7528_ (
    .Q(\datapath_1.regfile_1.regOut[5] [18]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_263_[18])
);

INVX1 _7108_ (
    .A(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_119_)
);

FILL FILL_4__9775_ (
);

FILL FILL_4__9355_ (
);

FILL FILL_2__13675_ (
);

FILL FILL_2__13255_ (
);

FILL SFILL99400x35050 (
);

FILL FILL_1__12248_ (
);

FILL FILL_0__9675_ (
);

FILL FILL_0__9255_ (
);

OAI21X1 _11946_ (
    .A(_3004_),
    .B(IorD_bF$buf6),
    .C(_3005_),
    .Y(_1_[19])
);

FILL FILL_3__7352_ (
);

AOI21X1 _11526_ (
    .A(_2634_),
    .B(_2636_),
    .C(_2220_),
    .Y(_2637_)
);

NOR2X1 _11106_ (
    .A(_2224_),
    .B(_2223_),
    .Y(_2225_)
);

FILL FILL_5__7698_ (
);

FILL FILL_4__16054_ (
);

FILL FILL_6__10155_ (
);

FILL FILL_3__15887_ (
);

FILL FILL_0__12602_ (
);

FILL FILL_3__15467_ (
);

FILL FILL_3__15047_ (
);

FILL FILL_1__16081_ (
);

FILL FILL_6_BUFX2_insert730 (
);

FILL FILL_3__10182_ (
);

FILL FILL_0__15494_ (
);

FILL SFILL89400x78050 (
);

FILL FILL_0__15074_ (
);

FILL FILL_6_BUFX2_insert735 (
);

FILL SFILL64040x3050 (
);

FILL FILL_1__8631_ (
);

FILL FILL_1__8211_ (
);

FILL FILL_2__15821_ (
);

FILL FILL_2__15401_ (
);

FILL FILL_3__8977_ (
);

FILL FILL_3__8137_ (
);

FILL SFILL49720x51050 (
);

FILL FILL_1__14814_ (
);

DFFSR _7281_ (
    .Q(\datapath_1.regfile_1.regOut[3] [27]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_133_[27])
);

FILL FILL_4__12394_ (
);

FILL FILL_0__13807_ (
);

FILL FILL_2__6974_ (
);

FILL FILL_5__9424_ (
);

FILL FILL_3__11387_ (
);

FILL FILL_5__9004_ (
);

FILL FILL_0__16279_ (
);

INVX1 _16144_ (
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_6597_)
);

FILL FILL_5__11714_ (
);

FILL FILL_1__9416_ (
);

FILL FILL_6__15193_ (
);

FILL FILL_4__7841_ (
);

FILL FILL_4__7421_ (
);

FILL FILL_4__10707_ (
);

FILL FILL_2__11741_ (
);

FILL FILL_5__14186_ (
);

FILL FILL_2__11321_ (
);

INVX1 _8486_ (
    .A(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_814_)
);

INVX1 _8066_ (
    .A(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_595_)
);

FILL FILL_4__13599_ (
);

FILL FILL_1__10314_ (
);

FILL FILL_2__7759_ (
);

FILL FILL_0__7741_ (
);

FILL FILL_0__7321_ (
);

FILL FILL_2__7339_ (
);

FILL SFILL94680x53050 (
);

FILL FILL_4__14960_ (
);

FILL FILL_4__14540_ (
);

FILL FILL_4__14120_ (
);

INVX1 _12484_ (
    .A(ALUOut[15]),
    .Y(_3389_)
);

FILL FILL_0__12199_ (
);

NAND3X1 _12064_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [19]),
    .C(_3034__bF$buf4),
    .Y(_3094_)
);

FILL FILL_3__13953_ (
);

FILL FILL_2__8700_ (
);

FILL SFILL94200x82050 (
);

FILL FILL_3__13533_ (
);

FILL FILL_3__13113_ (
);

FILL FILL_4__8626_ (
);

FILL FILL_4__8206_ (
);

FILL FILL_5_BUFX2_insert750 (
);

FILL FILL_5_BUFX2_insert751 (
);

FILL FILL_5_BUFX2_insert752 (
);

FILL FILL_2__12526_ (
);

FILL FILL_0__13980_ (
);

FILL FILL_2__12106_ (
);

FILL FILL_5_BUFX2_insert753 (
);

FILL FILL_0__13560_ (
);

FILL FILL_0__13140_ (
);

FILL FILL_5_BUFX2_insert754 (
);

FILL FILL_5_BUFX2_insert755 (
);

FILL FILL_5_BUFX2_insert756 (
);

FILL FILL_5_BUFX2_insert757 (
);

FILL FILL_1__11939_ (
);

FILL FILL_5_BUFX2_insert758 (
);

FILL FILL_5_BUFX2_insert759 (
);

FILL FILL_1__11519_ (
);

FILL FILL_5__16332_ (
);

FILL FILL_0__8526_ (
);

FILL FILL_0__8106_ (
);

FILL SFILL33960x35050 (
);

FILL FILL_5__6969_ (
);

FILL FILL_4__15745_ (
);

FILL FILL_4__15325_ (
);

FILL FILL_4__10880_ (
);

NOR2X1 _13689_ (
    .A(_4195_),
    .B(_3935__bF$buf2),
    .Y(_4196_)
);

FILL FILL_3__9095_ (
);

NOR2X1 _13269_ (
    .A(_3781_),
    .B(_3810_),
    .Y(\datapath_1.regfile_1.regEn [2])
);

FILL FILL_4__10040_ (
);

FILL FILL_2__9905_ (
);

FILL FILL_3__14738_ (
);

FILL FILL_3__14318_ (
);

FILL FILL_1__15772_ (
);

FILL FILL_1__15352_ (
);

FILL SFILL18760x15050 (
);

FILL SFILL84280x82050 (
);

FILL FILL_0__14765_ (
);

NAND3X1 _14630_ (
    .A(_5114_),
    .B(_5117_),
    .C(_5113_),
    .Y(_5118_)
);

FILL FILL_0__14345_ (
);

INVX1 _14210_ (
    .A(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_4707_)
);

FILL FILL_2__7092_ (
);

FILL FILL_3__7828_ (
);

FILL FILL_5__12252_ (
);

NAND2X1 _6972_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_49_)
);

FILL FILL_2_BUFX2_insert880 (
);

FILL SFILL79320x38050 (
);

FILL FILL_2_BUFX2_insert881 (
);

FILL FILL_2_BUFX2_insert882 (
);

FILL SFILL59000x9050 (
);

FILL FILL_2_BUFX2_insert883 (
);

FILL FILL_2_BUFX2_insert884 (
);

FILL FILL_4__11665_ (
);

FILL SFILL33720x5050 (
);

FILL FILL_2_BUFX2_insert885 (
);

FILL FILL_4__11245_ (
);

FILL FILL_2_BUFX2_insert886 (
);

FILL FILL_2_BUFX2_insert887 (
);

FILL FILL_2_BUFX2_insert888 (
);

FILL FILL_2_BUFX2_insert889 (
);

FILL FILL_1__16137_ (
);

FILL FILL_3__10658_ (
);

FILL FILL_3__10238_ (
);

FILL FILL_1__11692_ (
);

FILL SFILL84200x80050 (
);

FILL FILL_1__11272_ (
);

NAND3X1 _15835_ (
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf1),
    .Y(_6296_)
);

NAND2X1 _15415_ (
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .B(_5693_),
    .Y(_5886_)
);

FILL FILL_0__10685_ (
);

OAI21X1 _10970_ (
    .A(_2044_),
    .B(_2097_),
    .C(_2063_),
    .Y(_2045_)
);

NAND2X1 _10550_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1865_)
);

FILL FILL_0__10265_ (
);

NAND2X1 _10130_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1646_)
);

FILL SFILL109480x80050 (
);

FILL FILL_5__13877_ (
);

FILL FILL_5__13457_ (
);

FILL FILL_3__14491_ (
);

FILL FILL_5__13037_ (
);

INVX1 _7757_ (
    .A(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_450_)
);

FILL FILL_3__14071_ (
);

INVX1 _7337_ (
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_231_)
);

FILL FILL_4__9164_ (
);

FILL FILL_2__13484_ (
);

FILL SFILL114440x63050 (
);

FILL FILL_1__12897_ (
);

FILL FILL_1__12477_ (
);

FILL FILL_1__12057_ (
);

FILL FILL_4__13811_ (
);

FILL FILL_0__9484_ (
);

FILL FILL_3__7581_ (
);

NOR2X1 _11755_ (
    .A(_2488_),
    .B(_2494_),
    .Y(_2850_)
);

FILL FILL_3__7161_ (
);

OAI21X1 _11335_ (
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .C(_2321_),
    .Y(_2454_)
);

FILL FILL_6__15669_ (
);

FILL FILL_5__7087_ (
);

FILL FILL_4__16283_ (
);

FILL SFILL93400x78050 (
);

FILL FILL_3__15696_ (
);

FILL FILL_0__12831_ (
);

FILL FILL_0__12411_ (
);

FILL FILL_3__15276_ (
);

FILL FILL_1__7499_ (
);

FILL FILL_1__7079_ (
);

FILL FILL_2__14689_ (
);

FILL FILL_2__14269_ (
);

FILL FILL_5__15603_ (
);

INVX1 _9903_ (
    .A(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_1535_)
);

FILL FILL_1__8860_ (
);

FILL FILL_1__8440_ (
);

FILL FILL_1__8020_ (
);

FILL FILL_2__15630_ (
);

FILL FILL_2__15210_ (
);

FILL FILL_3__8786_ (
);

FILL FILL_3__8366_ (
);

FILL FILL_1__14623_ (
);

FILL FILL_1__14203_ (
);

INVX1 _7090_ (
    .A(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_107_)
);

FILL FILL_6__11589_ (
);

FILL FILL_0__13616_ (
);

INVX1 _13901_ (
    .A(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_4404_)
);

FILL FILL_5__9653_ (
);

FILL FILL_3__11196_ (
);

FILL FILL_5__9233_ (
);

FILL FILL_6__12530_ (
);

FILL FILL_0__16088_ (
);

NAND2X1 _16373_ (
    .A(gnd),
    .B(gnd),
    .Y(_6803_)
);

FILL FILL_2__10189_ (
);

FILL FILL_5__11943_ (
);

FILL FILL_1__9645_ (
);

FILL FILL_5__11523_ (
);

FILL FILL_1__9225_ (
);

FILL FILL_5__11103_ (
);

FILL FILL_2__16415_ (
);

FILL FILL_4__10936_ (
);

FILL FILL_4__7230_ (
);

FILL FILL_2__11970_ (
);

FILL FILL_4__10516_ (
);

FILL FILL_2__11550_ (
);

FILL FILL_2__11130_ (
);

FILL FILL_1__15828_ (
);

FILL FILL_1__15408_ (
);

DFFSR _8295_ (
    .Q(\datapath_1.regfile_1.regOut[11] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_653_[17])
);

FILL FILL_1__10963_ (
);

FILL FILL_1__10543_ (
);

FILL FILL_1__10123_ (
);

FILL FILL_0__7970_ (
);

FILL FILL_2__7988_ (
);

FILL SFILL104360x68050 (
);

BUFX2 BUFX2_insert570 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf37)
);

FILL FILL_2__7568_ (
);

FILL FILL_0__7550_ (
);

BUFX2 BUFX2_insert571 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf36)
);

BUFX2 BUFX2_insert572 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf35)
);

BUFX2 BUFX2_insert573 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf34)
);

FILL FILL_6__13735_ (
);

BUFX2 BUFX2_insert574 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf33)
);

BUFX2 BUFX2_insert575 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf32)
);

BUFX2 BUFX2_insert576 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf31)
);

BUFX2 BUFX2_insert577 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf30)
);

BUFX2 BUFX2_insert578 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf29)
);

BUFX2 BUFX2_insert579 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf28)
);

AOI22X1 _12293_ (
    .A(_2_[19]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3259_)
);

FILL FILL_5__12728_ (
);

FILL FILL_3__13762_ (
);

FILL FILL_5__12308_ (
);

FILL FILL_3__13342_ (
);

FILL FILL_4__8855_ (
);

FILL SFILL8600x7050 (
);

FILL FILL_4__8015_ (
);

FILL FILL_2__12755_ (
);

FILL FILL_2__12335_ (
);

FILL FILL_1__11748_ (
);

FILL FILL_1__11328_ (
);

FILL FILL_3__6852_ (
);

FILL FILL_5__16141_ (
);

FILL FILL_0__8755_ (
);

FILL FILL112440x74050 (
);

FILL FILL_0__8335_ (
);

DFFSR _10606_ (
    .Q(\datapath_1.regfile_1.regOut[29] [24]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1823_[24])
);

FILL FILL_0_BUFX2_insert90 (
);

FILL FILL_0_BUFX2_insert91 (
);

FILL FILL_4__15974_ (
);

FILL FILL_0_BUFX2_insert92 (
);

FILL SFILL104360x23050 (
);

FILL FILL_0_BUFX2_insert93 (
);

FILL FILL_4__15554_ (
);

FILL FILL_0_BUFX2_insert94 (
);

FILL FILL_4__15134_ (
);

FILL FILL_0_BUFX2_insert95 (
);

FILL FILL_0_BUFX2_insert96 (
);

FILL FILL_0_BUFX2_insert97 (
);

OAI22X1 _13498_ (
    .A(_4007_),
    .B(_3930__bF$buf2),
    .C(_3967__bF$buf1),
    .D(_4008_),
    .Y(_4009_)
);

FILL FILL_0_BUFX2_insert98 (
);

DFFSR _13078_ (
    .Q(_2_[31]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_3620_[31])
);

FILL FILL_0_BUFX2_insert99 (
);

FILL FILL_3__14967_ (
);

FILL FILL_3__14547_ (
);

FILL FILL_3__14127_ (
);

FILL FILL_1__15581_ (
);

FILL FILL_1__15161_ (
);

FILL FILL_0__14994_ (
);

FILL FILL_0__14574_ (
);

FILL FILL_0__14154_ (
);

FILL FILL_1__7711_ (
);

FILL FILL_2__14901_ (
);

FILL FILL_3__7637_ (
);

FILL FILL_3__7217_ (
);

FILL FILL_5__12481_ (
);

FILL SFILL73400x74050 (
);

FILL FILL_5__12061_ (
);

FILL FILL_4__16339_ (
);

FILL FILL_4__11894_ (
);

FILL FILL_4__11474_ (
);

FILL FILL_4__11054_ (
);

FILL FILL_1__16366_ (
);

FILL FILL_3__10887_ (
);

FILL FILL_5__8504_ (
);

FILL FILL_3__10047_ (
);

FILL FILL_1__11081_ (
);

FILL FILL_0__15779_ (
);

FILL FILL_0__15359_ (
);

OAI22X1 _15644_ (
    .A(_5463__bF$buf1),
    .B(_4660_),
    .C(_6109_),
    .D(_5495__bF$buf3),
    .Y(_6110_)
);

INVX8 _15224_ (
    .A(_5524__bF$buf0),
    .Y(_5700_)
);

FILL FILL_0__10494_ (
);

FILL FILL_1__8916_ (
);

FILL SFILL94280x79050 (
);

FILL FILL_6__14273_ (
);

FILL FILL_4__6921_ (
);

FILL FILL_0__16300_ (
);

FILL FILL_5__13686_ (
);

FILL FILL_2__10821_ (
);

FILL FILL_5__13266_ (
);

FILL FILL_2__10401_ (
);

FILL FILL_6__6847_ (
);

INVX1 _7986_ (
    .A(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_562_)
);

INVX1 _7566_ (
    .A(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_343_)
);

DFFSR _7146_ (
    .Q(\datapath_1.regfile_1.regOut[2] [20]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_68_[20])
);

FILL FILL_4__9393_ (
);

FILL FILL_4__12259_ (
);

FILL FILL_2__13293_ (
);

FILL FILL_2__6839_ (
);

FILL FILL_1__12286_ (
);

FILL SFILL37960x62050 (
);

FILL FILL_4__13620_ (
);

DFFSR _16429_ (
    .Q(\datapath_1.regfile_1.regOut[0] [12]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_6769_[12])
);

NOR2X1 _16009_ (
    .A(_6463_),
    .B(_6464_),
    .Y(_6465_)
);

FILL FILL_0__9293_ (
);

NAND3X1 _11984_ (
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[0]),
    .C(_3032__bF$buf0),
    .Y(_3033_)
);

FILL FILL_0__11699_ (
);

OAI21X1 _11564_ (
    .A(_2231_),
    .B(_2668_),
    .C(_2462__bF$buf0),
    .Y(_2673_)
);

FILL FILL_0__11279_ (
);

NOR2X1 _11144_ (
    .A(_2239_),
    .B(_2241_),
    .Y(_2263_)
);

FILL FILL_3__12613_ (
);

FILL FILL_4__16092_ (
);

FILL FILL_4__7706_ (
);

FILL FILL_2__11606_ (
);

FILL FILL_0__12640_ (
);

FILL FILL_0__12220_ (
);

FILL FILL_3__15085_ (
);

FILL FILL_2__14498_ (
);

FILL FILL_2__14078_ (
);

FILL FILL_5__15832_ (
);

FILL FILL_5__15412_ (
);

FILL FILL_0__7606_ (
);

DFFSR _9712_ (
    .Q(\datapath_1.regfile_1.regOut[22] [26]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_1368_[26])
);

FILL FILL_4__14825_ (
);

FILL FILL_4__14405_ (
);

FILL FILL_3__8595_ (
);

OAI21X1 _12769_ (
    .A(_3537_),
    .B(IRWrite_bF$buf3),
    .C(_3538_),
    .Y(_3490_[24])
);

INVX1 _12349_ (
    .A(ALUOut[2]),
    .Y(_3298_)
);

FILL FILL_3__13818_ (
);

FILL FILL_1__14852_ (
);

FILL FILL_1__14432_ (
);

FILL FILL_1__14012_ (
);

FILL FILL_0__13845_ (
);

FILL FILL_0__13425_ (
);

INVX1 _13710_ (
    .A(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_4217_)
);

FILL FILL_0__13005_ (
);

FILL FILL_5__9882_ (
);

FILL FILL_5__9462_ (
);

FILL FILL_5__9042_ (
);

INVX1 _16182_ (
    .A(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_6634_)
);

FILL FILL_3__6908_ (
);

FILL FILL_5__11752_ (
);

FILL FILL_1__9874_ (
);

FILL FILL_5__11332_ (
);

FILL FILL_1__9034_ (
);

FILL SFILL8680x51050 (
);

FILL FILL_2__16224_ (
);

FILL FILL_4__10745_ (
);

FILL FILL_4__10325_ (
);

FILL FILL_1__15637_ (
);

FILL FILL_1__15217_ (
);

FILL SFILL84200x75050 (
);

FILL FILL_1__10772_ (
);

OAI22X1 _14915_ (
    .A(_3947__bF$buf0),
    .B(_5395_),
    .C(_3977__bF$buf0),
    .D(_5396_),
    .Y(_5397_)
);

FILL FILL_2__7377_ (
);

FILL SFILL109480x75050 (
);

FILL FILL_5__12957_ (
);

FILL FILL_3__13991_ (
);

FILL FILL_5__12117_ (
);

FILL FILL_3__13571_ (
);

BUFX2 _6837_ (
    .A(_0_),
    .Y(MemWrite)
);

FILL FILL_3__13151_ (
);

FILL FILL_4__8244_ (
);

FILL FILL_2__12984_ (
);

FILL FILL_2__12144_ (
);

FILL FILL_1__11977_ (
);

FILL FILL_1__11557_ (
);

FILL FILL_1__11137_ (
);

FILL SFILL109880x44050 (
);

FILL SFILL84200x30050 (
);

FILL FILL_5__16370_ (
);

FILL FILL_0__8984_ (
);

FILL SFILL74280x75050 (
);

FILL SFILL23560x14050 (
);

INVX1 _10835_ (
    .A(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_2014_)
);

FILL FILL_0__8144_ (
);

INVX1 _10415_ (
    .A(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_1795_)
);

FILL FILL_4__15783_ (
);

FILL FILL_6__14329_ (
);

FILL FILL_4__15363_ (
);

FILL SFILL13640x50050 (
);

FILL FILL_0__11911_ (
);

FILL FILL_2__9523_ (
);

FILL FILL_3__14776_ (
);

FILL FILL_2__9103_ (
);

FILL FILL_3__14356_ (
);

FILL FILL_1__15390_ (
);

FILL FILL_4__9869_ (
);

FILL FILL_4__9029_ (
);

FILL FILL_2__13769_ (
);

FILL FILL_2__13349_ (
);

FILL FILL_0__14383_ (
);

FILL SFILL114440x13050 (
);

FILL FILL_1__7940_ (
);

FILL FILL_1__7100_ (
);

FILL FILL_2__14710_ (
);

FILL SFILL74200x73050 (
);

FILL FILL_3__7866_ (
);

FILL FILL_0__9769_ (
);

FILL FILL_0__9349_ (
);

FILL FILL_3__7446_ (
);

FILL FILL_5__12290_ (
);

FILL SFILL74280x30050 (
);

FILL FILL_1__13703_ (
);

FILL FILL_4__16148_ (
);

FILL FILL_4__11283_ (
);

FILL SFILL19240x78050 (
);

FILL FILL_1__16175_ (
);

FILL FILL_3__10696_ (
);

FILL FILL_5__8733_ (
);

FILL FILL_3__10276_ (
);

FILL FILL_5__8313_ (
);

OAI21X1 _15873_ (
    .A(_4897_),
    .B(_5535__bF$buf3),
    .C(_6332_),
    .Y(_6333_)
);

FILL FILL_0__15588_ (
);

FILL FILL_6__11610_ (
);

FILL FILL_0__15168_ (
);

NOR2X1 _15453_ (
    .A(_5920_),
    .B(_5923_),
    .Y(_5924_)
);

NOR2X1 _15033_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5513_)
);

FILL SFILL53960x50 (
);

FILL FILL_1__8725_ (
);

FILL FILL_2__15915_ (
);

FILL FILL_5__13495_ (
);

FILL FILL_2__10630_ (
);

DFFSR _7795_ (
    .Q(\datapath_1.regfile_1.regOut[7] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_393_[29])
);

FILL FILL_1__14908_ (
);

OAI21X1 _7375_ (
    .A(_255_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_256_),
    .Y(_198_[29])
);

FILL FILL_4__12488_ (
);

FILL FILL_4__12068_ (
);

FILL FILL_5__9938_ (
);

FILL FILL_5__9518_ (
);

FILL FILL_1__12095_ (
);

OAI21X1 _16238_ (
    .A(_5338_),
    .B(_5535__bF$buf0),
    .C(_6688_),
    .Y(_6689_)
);

AOI21X1 _11793_ (
    .A(_2371_),
    .B(_2620_),
    .C(_2885_),
    .Y(_2886_)
);

INVX1 _11373_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .Y(_2490_)
);

FILL FILL_0__11088_ (
);

FILL FILL_5__11808_ (
);

FILL FILL_3__12842_ (
);

FILL FILL_3__12422_ (
);

FILL FILL_3__12002_ (
);

FILL SFILL104440x11050 (
);

FILL FILL_4__7935_ (
);

FILL FILL_2__11835_ (
);

FILL FILL_2__11415_ (
);

FILL SFILL33800x80050 (
);

FILL FILL_1__10828_ (
);

FILL FILL_1__10408_ (
);

FILL FILL_5__15641_ (
);

FILL FILL112440x69050 (
);

FILL FILL_5__15221_ (
);

FILL FILL_0__7835_ (
);

FILL FILL_0__7415_ (
);

OAI21X1 _9941_ (
    .A(_1559_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .C(_1560_),
    .Y(_1498_[31])
);

OAI21X1 _9521_ (
    .A(_1340_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1341_),
    .Y(_1303_[19])
);

OAI21X1 _9101_ (
    .A(_1121_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1122_),
    .Y(_1108_[7])
);

FILL SFILL104360x18050 (
);

FILL FILL_4__14634_ (
);

FILL FILL_4__14214_ (
);

OAI21X1 _12998_ (
    .A(_3649_),
    .B(vdd),
    .C(_3650_),
    .Y(_3620_[15])
);

OAI21X1 _12578_ (
    .A(_3430_),
    .B(vdd),
    .C(_3431_),
    .Y(_3425_[3])
);

NAND2X1 _12158_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.a [14]),
    .Y(_3159_)
);

FILL FILL_3__13627_ (
);

FILL FILL_3__13207_ (
);

FILL FILL_1__14661_ (
);

FILL FILL_1__14241_ (
);

FILL SFILL108680x26050 (
);

FILL FILL_0__13654_ (
);

FILL FILL_0__13234_ (
);

FILL FILL_3__16099_ (
);

FILL FILL_5__9271_ (
);

FILL FILL_5__16006_ (
);

FILL FILL_5__11981_ (
);

FILL FILL_1__9683_ (
);

FILL FILL_5__11561_ (
);

FILL FILL_1__9263_ (
);

FILL FILL_5__11141_ (
);

FILL FILL112440x24050 (
);

FILL FILL_4__15839_ (
);

FILL FILL_4__15419_ (
);

FILL FILL_2__16033_ (
);

FILL FILL_4__10974_ (
);

FILL FILL_4__10554_ (
);

FILL FILL_4__10134_ (
);

FILL SFILL13640x50 (
);

FILL FILL_1__15866_ (
);

FILL FILL_1__15446_ (
);

FILL FILL_1__15026_ (
);

FILL SFILL33720x42050 (
);

FILL SFILL49320x27050 (
);

FILL FILL_1__10581_ (
);

FILL FILL_1__10161_ (
);

FILL FILL_0__14859_ (
);

FILL FILL112040x10050 (
);

INVX1 _14724_ (
    .A(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_5210_)
);

FILL FILL_0__14439_ (
);

FILL FILL_0__14019_ (
);

OAI22X1 _14304_ (
    .A(_3983__bF$buf3),
    .B(_4797_),
    .C(_3977__bF$buf4),
    .D(_4798_),
    .Y(_4799_)
);

BUFX2 BUFX2_insert950 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf7 )
);

BUFX2 BUFX2_insert951 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf6 )
);

FILL FILL_2__7186_ (
);

BUFX2 BUFX2_insert952 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf5 )
);

BUFX2 BUFX2_insert953 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf4 )
);

BUFX2 BUFX2_insert954 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf3 )
);

BUFX2 BUFX2_insert955 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf2 )
);

BUFX2 BUFX2_insert956 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf1 )
);

BUFX2 BUFX2_insert957 (
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf0 )
);

FILL FILL_0__15800_ (
);

BUFX2 BUFX2_insert958 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf7 )
);

BUFX2 BUFX2_insert959 (
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf6 )
);

FILL FILL_5__12766_ (
);

FILL FILL_5__12346_ (
);

FILL FILL_3__13380_ (
);

FILL FILL_4__8893_ (
);

FILL FILL_4__8473_ (
);

FILL FILL_4__11759_ (
);

FILL FILL_4__11339_ (
);

FILL FILL_2__12373_ (
);

FILL FILL_1__11786_ (
);

FILL FILL_1__11366_ (
);

AOI21X1 _15929_ (
    .A(_6387_),
    .B(_6369_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [21])
);

FILL FILL_4__12700_ (
);

AOI22X1 _15509_ (
    .A(\datapath_1.regfile_1.regOut[31] [11]),
    .B(_5571_),
    .C(_5570__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_5978_)
);

FILL FILL_3__6890_ (
);

FILL FILL_0__8373_ (
);

FILL FILL_0__10779_ (
);

FILL FILL_0__10359_ (
);

INVX1 _10644_ (
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_1907_)
);

DFFSR _10224_ (
    .Q(\datapath_1.regfile_1.regOut[26] [26]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_1628_[26])
);

FILL FILL_4__15592_ (
);

FILL FILL_4__15172_ (
);

FILL SFILL94280x29050 (
);

FILL FILL_2__9752_ (
);

FILL FILL_3__14585_ (
);

FILL FILL_0__11720_ (
);

FILL FILL_3__14165_ (
);

FILL FILL_0__11300_ (
);

FILL FILL_4_BUFX2_insert790 (
);

FILL FILL_4__9678_ (
);

FILL FILL_4_BUFX2_insert791 (
);

FILL FILL_4_BUFX2_insert792 (
);

FILL FILL_4__9258_ (
);

FILL FILL_2__13998_ (
);

FILL FILL_4_BUFX2_insert793 (
);

FILL FILL_4_BUFX2_insert794 (
);

FILL FILL_2__13578_ (
);

FILL FILL_4_BUFX2_insert795 (
);

FILL FILL_2__13158_ (
);

FILL FILL_0__14192_ (
);

FILL FILL_4_BUFX2_insert796 (
);

FILL FILL_5__14912_ (
);

FILL FILL_4_BUFX2_insert797 (
);

FILL FILL_4_BUFX2_insert798 (
);

FILL FILL_4_BUFX2_insert799 (
);

FILL FILL_4__13905_ (
);

FILL FILL_0__9998_ (
);

FILL FILL_3__7675_ (
);

FILL FILL_0__9158_ (
);

NAND3X1 _11849_ (
    .A(_2934_),
    .B(_2933_),
    .C(_2936_),
    .Y(\datapath_1.ALUResult [0])
);

OAI21X1 _11429_ (
    .A(_2544_),
    .B(_2361_),
    .C(_2370_),
    .Y(_2545_)
);

INVX1 _11009_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2128_)
);

FILL FILL_1__13932_ (
);

FILL FILL_4__16377_ (
);

FILL FILL_1__13512_ (
);

FILL FILL_4__11092_ (
);

FILL FILL_0__12505_ (
);

FILL FILL_5__8962_ (
);

FILL FILL_5__8122_ (
);

INVX1 _15682_ (
    .A(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_6147_)
);

FILL FILL_0__15397_ (
);

OAI22X1 _15262_ (
    .A(_5478__bF$buf2),
    .B(_4217_),
    .C(_5552__bF$buf3),
    .D(_4210_),
    .Y(_5737_)
);

FILL SFILL63400x22050 (
);

FILL FILL_3__16311_ (
);

FILL FILL_5__10832_ (
);

FILL FILL_1__8954_ (
);

FILL FILL_5__10412_ (
);

FILL FILL_1__8114_ (
);

FILL SFILL8680x46050 (
);

FILL SFILL13720x83050 (
);

FILL FILL_2__15724_ (
);

FILL FILL_2__15304_ (
);

FILL FILL_1__14717_ (
);

OAI21X1 _7184_ (
    .A(_148_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .C(_149_),
    .Y(_133_[8])
);

FILL SFILL53800x79050 (
);

FILL FILL_4__12297_ (
);

FILL FILL_3__9401_ (
);

FILL SFILL84280x27050 (
);

FILL FILL_2__6877_ (
);

FILL FILL_5__9747_ (
);

FILL FILL_6__12624_ (
);

NAND2X1 _16047_ (
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .B(_5693_),
    .Y(_6502_)
);

NOR2X1 _11182_ (
    .A(\datapath_1.alu_1.ALUInA [24]),
    .B(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2301_)
);

FILL FILL_1__9739_ (
);

FILL FILL_5__11617_ (
);

FILL FILL_3__12651_ (
);

FILL SFILL8600x44050 (
);

FILL FILL_3__12231_ (
);

FILL FILL_6__15096_ (
);

FILL FILL_4__7744_ (
);

FILL FILL_4__7324_ (
);

FILL FILL_2__11644_ (
);

FILL FILL_2__11224_ (
);

FILL FILL_5__14089_ (
);

NAND2X1 _8389_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_770_)
);

FILL FILL_1__10637_ (
);

FILL SFILL84200x25050 (
);

FILL FILL_5__15870_ (
);

FILL FILL_5__15450_ (
);

FILL FILL_5__15030_ (
);

FILL FILL_0__7224_ (
);

OAI21X1 _9750_ (
    .A(_1452_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .C(_1453_),
    .Y(_1433_[10])
);

FILL SFILL114040x39050 (
);

DFFSR _9330_ (
    .Q(\datapath_1.regfile_1.regOut[19] [28]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_1173_[28])
);

FILL FILL_4__14863_ (
);

FILL FILL_4__14443_ (
);

FILL FILL_4__14023_ (
);

FILL SFILL13640x45050 (
);

OAI21X1 _12387_ (
    .A(_3322_),
    .B(MemToReg_bF$buf3),
    .C(_3323_),
    .Y(\datapath_1.mux_wd3.dout [14])
);

FILL FILL_3__13856_ (
);

FILL FILL_2__8603_ (
);

FILL FILL_3__13436_ (
);

FILL FILL_1__14890_ (
);

FILL FILL_1__14470_ (
);

FILL FILL_3__13016_ (
);

FILL FILL_1__14050_ (
);

FILL FILL_4__8529_ (
);

FILL FILL_4__8109_ (
);

FILL FILL_2__12849_ (
);

FILL FILL_0__13883_ (
);

FILL FILL_2__12429_ (
);

FILL SFILL19320x66050 (
);

FILL FILL_0__13463_ (
);

FILL FILL_2__12009_ (
);

FILL FILL_0__13043_ (
);

FILL FILL_5__9080_ (
);

FILL SFILL74200x68050 (
);

FILL FILL_5__16235_ (
);

FILL FILL_3__6946_ (
);

FILL FILL_0__8849_ (
);

FILL FILL_0__8009_ (
);

FILL FILL_5__11790_ (
);

FILL FILL_5__11370_ (
);

FILL FILL_1__9492_ (
);

FILL FILL_4__15648_ (
);

FILL FILL_4__15228_ (
);

FILL FILL_2__16262_ (
);

FILL FILL_4__10783_ (
);

FILL FILL_4__10363_ (
);

FILL FILL_4_BUFX2_insert40 (
);

FILL FILL_2__9808_ (
);

FILL FILL_4_BUFX2_insert41 (
);

FILL FILL112200x81050 (
);

FILL FILL_1__15675_ (
);

FILL FILL_4_BUFX2_insert42 (
);

FILL FILL_1__15255_ (
);

FILL FILL_4_BUFX2_insert43 (
);

FILL FILL_4_BUFX2_insert44 (
);

FILL FILL_4_BUFX2_insert45 (
);

FILL FILL_5__7813_ (
);

FILL FILL_4_BUFX2_insert46 (
);

FILL FILL_4_BUFX2_insert47 (
);

FILL FILL_1__10390_ (
);

FILL FILL_4_BUFX2_insert48 (
);

FILL FILL_4_BUFX2_insert49 (
);

INVX1 _14953_ (
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_5434_)
);

FILL FILL_0__14668_ (
);

FILL FILL_0__14248_ (
);

INVX1 _14533_ (
    .A(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_5023_)
);

INVX1 _14113_ (
    .A(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_4612_)
);

FILL FILL_1__7805_ (
);

FILL FILL_6__13582_ (
);

FILL FILL_5__12995_ (
);

FILL FILL_5__12575_ (
);

FILL SFILL74200x23050 (
);

FILL FILL_5__12155_ (
);

BUFX2 _6875_ (
    .A(_2_[5]),
    .Y(memoryWriteData[5])
);

FILL SFILL95160x21050 (
);

FILL FILL_4__11988_ (
);

FILL FILL_4__11568_ (
);

FILL FILL_4__11148_ (
);

FILL FILL_2__12182_ (
);

FILL FILL_1__11595_ (
);

FILL FILL_1__11175_ (
);

NAND2X1 _15738_ (
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .B(_5570__bF$buf2),
    .Y(_6201_)
);

NOR3X1 _15318_ (
    .A(_5787_),
    .B(_5791_),
    .C(_5789_),
    .Y(_5792_)
);

FILL FILL_0__8182_ (
);

NAND2X1 _10873_ (
    .A(\aluControl_1.inst [2]),
    .B(_2020_),
    .Y(_2021_)
);

FILL FILL_0__10168_ (
);

OAI21X1 _10453_ (
    .A(_1819_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1820_),
    .Y(_1758_[31])
);

OAI21X1 _10033_ (
    .A(_1600_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1601_),
    .Y(_1563_[19])
);

FILL FILL_3__11922_ (
);

FILL FILL_3__11502_ (
);

FILL FILL_2__10915_ (
);

FILL FILL_2__9981_ (
);

FILL SFILL33800x75050 (
);

FILL SFILL64200x66050 (
);

FILL FILL_2__9141_ (
);

FILL FILL_3__14394_ (
);

FILL SFILL43320x25050 (
);

FILL FILL_4__9487_ (
);

FILL FILL_2__13387_ (
);

FILL FILL_5__14721_ (
);

FILL FILL_0__6915_ (
);

FILL FILL_5__14301_ (
);

OAI21X1 _8601_ (
    .A(_869_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_870_),
    .Y(_848_[11])
);

FILL FILL_4__13714_ (
);

FILL FILL_3__7484_ (
);

FILL FILL_0__9387_ (
);

FILL FILL_3__7064_ (
);

OAI21X1 _11658_ (
    .A(_2402_),
    .B(_2403_),
    .C(_2760_),
    .Y(_2761_)
);

NOR2X1 _11238_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2357_)
);

FILL FILL_3__12707_ (
);

FILL FILL_1__13741_ (
);

FILL FILL_1__13321_ (
);

FILL FILL_4__16186_ (
);

FILL FILL_0__12734_ (
);

FILL FILL_3__15599_ (
);

FILL FILL_3__15179_ (
);

FILL FILL_0__12314_ (
);

FILL SFILL89400x3050 (
);

FILL FILL_5__8771_ (
);

FILL SFILL33800x30050 (
);

FILL FILL_5__8351_ (
);

FILL SFILL64200x21050 (
);

INVX1 _15491_ (
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_5961_)
);

FILL FILL_5__15926_ (
);

NAND3X1 _15071_ (
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf0),
    .Y(_5551_)
);

FILL FILL_5__15506_ (
);

NAND2X1 _9806_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1491_)
);

FILL FILL_3__16120_ (
);

FILL FILL_1__8763_ (
);

FILL FILL_5__10641_ (
);

FILL FILL112440x19050 (
);

FILL FILL_1__8343_ (
);

FILL FILL_4__14919_ (
);

FILL FILL_2__15953_ (
);

FILL FILL_2__15533_ (
);

FILL FILL_2__15113_ (
);

FILL FILL_3__8269_ (
);

FILL FILL_1__14946_ (
);

FILL FILL_1__14526_ (
);

FILL FILL_1__14106_ (
);

FILL FILL_0__13939_ (
);

FILL FILL_3__9630_ (
);

NOR3X1 _13804_ (
    .A(_4303_),
    .B(_4305_),
    .C(_4308_),
    .Y(_4309_)
);

FILL FILL_0__13519_ (
);

FILL FILL_3__9210_ (
);

FILL FILL_5__9976_ (
);

FILL FILL_5__9556_ (
);

FILL FILL_5__9136_ (
);

FILL FILL_3__11099_ (
);

FILL FILL_6__12433_ (
);

OAI22X1 _16276_ (
    .A(_6724_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf3),
    .D(_6725_),
    .Y(_6726_)
);

FILL FILL_5__11846_ (
);

FILL FILL_1__9548_ (
);

FILL FILL_3__12880_ (
);

FILL FILL_5__11426_ (
);

FILL FILL_3__12460_ (
);

FILL FILL_1__9128_ (
);

FILL FILL_5__11006_ (
);

FILL FILL_3__12040_ (
);

FILL FILL_4__7973_ (
);

FILL FILL_2__16318_ (
);

FILL FILL_4__7553_ (
);

FILL FILL_2__11873_ (
);

FILL FILL_4__10419_ (
);

FILL FILL_2__11453_ (
);

FILL FILL_2__11033_ (
);

NAND2X1 _8198_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_663_)
);

FILL FILL_6__7059_ (
);

FILL FILL_1__10446_ (
);

FILL FILL_1__10026_ (
);

FILL FILL_0__7873_ (
);

FILL FILL_0__7453_ (
);

FILL FILL_0__7033_ (
);

FILL FILL_6__13638_ (
);

FILL FILL_4__14672_ (
);

FILL FILL_4__14252_ (
);

INVX1 _12196_ (
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3184_)
);

FILL FILL_2__8832_ (
);

FILL FILL_3__13665_ (
);

FILL FILL_0__10800_ (
);

FILL FILL_3__13245_ (
);

FILL FILL_4__8758_ (
);

FILL FILL_4__8338_ (
);

FILL FILL_2__12658_ (
);

FILL FILL_2__12238_ (
);

FILL FILL_0__13692_ (
);

FILL FILL_0__13272_ (
);

FILL SFILL23720x35050 (
);

FILL FILL_5__16044_ (
);

FILL FILL_0__8658_ (
);

NOR2X1 _10929_ (
    .A(_2049_),
    .B(_2057_),
    .Y(_2063_)
);

FILL FILL_0__8238_ (
);

OAI21X1 _10509_ (
    .A(_1836_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .C(_1837_),
    .Y(_1823_[7])
);

FILL FILL_4__15877_ (
);

FILL FILL_4__15457_ (
);

FILL FILL_4__15037_ (
);

FILL FILL_2__16071_ (
);

FILL FILL_4__10172_ (
);

FILL SFILL58440x34050 (
);

FILL FILL_2__9617_ (
);

FILL FILL_1__15484_ (
);

FILL FILL_1__15064_ (
);

FILL FILL_5__7622_ (
);

FILL FILL_5__7202_ (
);

FILL FILL_0__14897_ (
);

FILL FILL_0__14477_ (
);

AOI22X1 _14762_ (
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .B(_3942__bF$buf3),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_5247_)
);

FILL FILL_0__14057_ (
);

NOR2X1 _14342_ (
    .A(_4835_),
    .B(_3954__bF$buf2),
    .Y(_4836_)
);

FILL FILL_3__15811_ (
);

FILL FILL_1__7614_ (
);

FILL FILL_2__14804_ (
);

FILL FILL_5__12384_ (
);

FILL FILL_4__8091_ (
);

FILL FILL_4__11797_ (
);

FILL FILL_4__11377_ (
);

FILL FILL_3__8901_ (
);

FILL FILL_1__16269_ (
);

FILL FILL_5__8827_ (
);

NOR3X1 _15967_ (
    .A(_6413_),
    .B(_6402_),
    .C(_6424_),
    .Y(_6425_)
);

AOI22X1 _15547_ (
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .B(_5567_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_6015_)
);

AOI21X1 _15127_ (
    .A(_5582_),
    .B(_5605_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [1])
);

OAI21X1 _10682_ (
    .A(_1931_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1932_),
    .Y(_1888_[22])
);

FILL FILL_0__10397_ (
);

OAI21X1 _10262_ (
    .A(_1712_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .C(_1713_),
    .Y(_1693_[10])
);

FILL SFILL8600x39050 (
);

FILL FILL_3__11731_ (
);

FILL FILL_3__11311_ (
);

FILL FILL_0__16203_ (
);

FILL SFILL13720x33050 (
);

FILL FILL_2__9790_ (
);

FILL FILL_5__13589_ (
);

FILL FILL_2__10304_ (
);

FILL FILL_5__13169_ (
);

FILL FILL_2__9370_ (
);

NAND2X1 _7889_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_518_)
);

NAND2X1 _7469_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_299_)
);

FILL SFILL109560x13050 (
);

NAND2X1 _7049_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_80_)
);

FILL FILL_4__9296_ (
);

FILL SFILL109400x2050 (
);

FILL SFILL38920x82050 (
);

FILL FILL_5__14950_ (
);

FILL FILL_5__14530_ (
);

FILL FILL_5__14110_ (
);

OAI21X1 _8830_ (
    .A(_981_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .C(_982_),
    .Y(_978_[2])
);

DFFSR _8410_ (
    .Q(\datapath_1.regfile_1.regOut[12] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_718_[4])
);

FILL FILL_1__12189_ (
);

FILL FILL_4__13943_ (
);

FILL FILL_4__13523_ (
);

FILL FILL_4__13103_ (
);

INVX1 _11887_ (
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3030_)
);

FILL FILL_3__7293_ (
);

INVX1 _11467_ (
    .A(_2292_),
    .Y(_2582_)
);

FILL SFILL88520x28050 (
);

NOR2X1 _11047_ (
    .A(_2164_),
    .B(_2165_),
    .Y(_2166_)
);

FILL FILL_3__12516_ (
);

FILL FILL_1__13970_ (
);

FILL FILL_1__13550_ (
);

FILL FILL_1__13130_ (
);

FILL FILL_4__7609_ (
);

FILL FILL_2__11929_ (
);

FILL FILL_0__12963_ (
);

FILL FILL_2__11509_ (
);

FILL FILL_0__12123_ (
);

FILL FILL_5__8580_ (
);

FILL SFILL3560x81050 (
);

FILL FILL_5__15735_ (
);

FILL FILL_5__15315_ (
);

FILL FILL_0__7929_ (
);

FILL FILL_0__7509_ (
);

NAND2X1 _9615_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1384_)
);

FILL FILL_1__8992_ (
);

FILL FILL_5__10870_ (
);

FILL FILL_1__8572_ (
);

FILL FILL_5__10450_ (
);

FILL FILL_5__10030_ (
);

FILL FILL_4__14728_ (
);

FILL FILL_4__14308_ (
);

FILL FILL_2__15762_ (
);

FILL FILL_2__15342_ (
);

FILL FILL_3__8498_ (
);

FILL FILL_3__8078_ (
);

FILL FILL112200x76050 (
);

FILL SFILL99480x69050 (
);

FILL FILL_1__14755_ (
);

FILL FILL_1__14335_ (
);

FILL FILL_0__13748_ (
);

INVX1 _13613_ (
    .A(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_4122_)
);

FILL FILL_0__13328_ (
);

FILL SFILL38840x44050 (
);

FILL FILL_5__9785_ (
);

FILL FILL_5__9365_ (
);

NAND3X1 _16085_ (
    .A(_6535_),
    .B(_6539_),
    .C(_6531_),
    .Y(_6540_)
);

FILL SFILL43800x27050 (
);

FILL SFILL28920x80050 (
);

FILL SFILL74200x18050 (
);

FILL FILL_1__9777_ (
);

FILL FILL_5__11655_ (
);

FILL FILL_1__9357_ (
);

FILL FILL_5__11235_ (
);

FILL FILL_2__16127_ (
);

FILL FILL_4__7362_ (
);

FILL FILL_4__10648_ (
);

FILL FILL_2__11682_ (
);

FILL FILL_2__11262_ (
);

FILL FILL112200x31050 (
);

FILL FILL_1__10675_ (
);

FILL SFILL99480x24050 (
);

FILL FILL_1__10255_ (
);

OAI22X1 _14818_ (
    .A(_5300_),
    .B(_3930__bF$buf0),
    .C(_3924__bF$buf3),
    .D(_5301_),
    .Y(_5302_)
);

FILL FILL_0__7682_ (
);

FILL FILL_4__14481_ (
);

FILL FILL_6__13027_ (
);

FILL FILL_4__14061_ (
);

FILL FILL_3__13894_ (
);

FILL FILL_2__8641_ (
);

FILL FILL_3__13474_ (
);

FILL FILL_2__8221_ (
);

FILL SFILL68840x6050 (
);

FILL FILL112120x38050 (
);

FILL FILL_4__8987_ (
);

FILL FILL_4__8567_ (
);

FILL FILL_4__8147_ (
);

FILL FILL_2__12887_ (
);

FILL FILL_2__12467_ (
);

FILL FILL_2__12047_ (
);

FILL FILL_0__13081_ (
);

FILL FILL_5__13801_ (
);

FILL SFILL24520x34050 (
);

FILL SFILL89480x67050 (
);

FILL FILL_0__8887_ (
);

FILL FILL_5__16273_ (
);

FILL FILL_3__6984_ (
);

FILL FILL_0__8467_ (
);

DFFSR _10738_ (
    .Q(\datapath_1.regfile_1.regOut[30] [28]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_1888_[28])
);

NAND2X1 _10318_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1751_)
);

FILL FILL_4__15686_ (
);

FILL FILL_1__12401_ (
);

FILL FILL_4__15266_ (
);

FILL FILL_2__9846_ (
);

FILL FILL_2__9426_ (
);

FILL FILL_0__11814_ (
);

FILL FILL_3__14679_ (
);

FILL FILL_3__14259_ (
);

FILL FILL_2__9006_ (
);

FILL FILL_1__15293_ (
);

FILL SFILL33800x25050 (
);

FILL FILL_5__7851_ (
);

FILL FILL_5__7431_ (
);

NOR2X1 _14991_ (
    .A(\datapath_1.PCJump [26]),
    .B(_5470_),
    .Y(_5471_)
);

AOI22X1 _14571_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [23]),
    .C(\datapath_1.regfile_1.regOut[6] [23]),
    .D(_4001__bF$buf0),
    .Y(_5060_)
);

FILL FILL_0__14286_ (
);

INVX1 _14151_ (
    .A(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_4649_)
);

FILL FILL_3__15620_ (
);

FILL FILL_3__15200_ (
);

FILL FILL_1__7843_ (
);

FILL FILL_1__7423_ (
);

FILL FILL_2__14613_ (
);

FILL FILL_3__7349_ (
);

FILL FILL_5__12193_ (
);

FILL FILL_1__13606_ (
);

FILL FILL_4__11186_ (
);

FILL FILL_3__8710_ (
);

FILL FILL_1__16078_ (
);

FILL FILL_5__8636_ (
);

FILL FILL_5__8216_ (
);

FILL FILL_3__10179_ (
);

NOR2X1 _15776_ (
    .A(_6236_),
    .B(_6237_),
    .Y(_6238_)
);

AOI22X1 _15356_ (
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .B(_5567_),
    .C(_5486_),
    .D(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_5829_)
);

FILL FILL_3__16405_ (
);

OAI21X1 _10491_ (
    .A(_1824_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1825_),
    .Y(_1823_[1])
);

FILL FILL_5__10926_ (
);

DFFSR _10071_ (
    .Q(\datapath_1.regfile_1.regOut[25] [1]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_1563_[1])
);

FILL FILL_3__11960_ (
);

FILL FILL_5__10506_ (
);

FILL FILL_1__8628_ (
);

FILL FILL_1__8208_ (
);

FILL FILL_3__11540_ (
);

FILL FILL_3__11120_ (
);

FILL FILL_2__15818_ (
);

FILL SFILL63880x80050 (
);

FILL FILL_0__16012_ (
);

FILL FILL_2__10953_ (
);

FILL FILL_2__10533_ (
);

FILL FILL_5__13398_ (
);

FILL FILL_2__10113_ (
);

NAND2X1 _7698_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_411_)
);

DFFSR _7278_ (
    .Q(\datapath_1.regfile_1.regOut[3] [24]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_133_[24])
);

FILL FILL_3__9915_ (
);

FILL SFILL18840x40050 (
);

FILL FILL_0__6953_ (
);

FILL FILL_4__13752_ (
);

FILL FILL_4__13332_ (
);

FILL SFILL110280x82050 (
);

AOI21X1 _11696_ (
    .A(_2165_),
    .B(_2757_),
    .C(_2458_),
    .Y(_2796_)
);

OAI21X1 _11276_ (
    .A(_2381_),
    .B(_2390_),
    .C(_2394_),
    .Y(_2395_)
);

FILL FILL_3__12745_ (
);

FILL FILL_3__12325_ (
);

FILL FILL_4__7838_ (
);

FILL FILL_4__7418_ (
);

FILL SFILL69960x70050 (
);

FILL FILL_2__11738_ (
);

FILL FILL_0__12772_ (
);

FILL FILL_2__11318_ (
);

FILL SFILL109240x77050 (
);

FILL FILL_0__12352_ (
);

FILL SFILL74120x9050 (
);

FILL FILL_5__15964_ (
);

FILL FILL_5__15544_ (
);

FILL FILL_0__7738_ (
);

FILL FILL_5__15124_ (
);

DFFSR _9844_ (
    .Q(\datapath_1.regfile_1.regOut[23] [30]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1433_[30])
);

FILL FILL_0__7318_ (
);

INVX1 _9424_ (
    .A(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_1297_)
);

INVX1 _9004_ (
    .A(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_1078_)
);

FILL FILL_1__8381_ (
);

FILL FILL_4__14957_ (
);

FILL SFILL48920x79050 (
);

FILL FILL_2__15991_ (
);

FILL FILL_4__14537_ (
);

FILL FILL_2__15571_ (
);

FILL FILL_4__14117_ (
);

FILL FILL_2__15151_ (
);

FILL FILL_1__14984_ (
);

FILL FILL_1__14564_ (
);

FILL FILL_1__14144_ (
);

FILL FILL_0__13977_ (
);

INVX1 _13842_ (
    .A(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_4346_)
);

FILL FILL_0__13557_ (
);

INVX1 _13422_ (
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_3934_)
);

FILL FILL_0__13137_ (
);

INVX1 _13002_ (
    .A(_2_[17]),
    .Y(_3653_)
);

FILL FILL_5__9594_ (
);

FILL FILL_5__16329_ (
);

FILL FILL_5__11884_ (
);

FILL FILL_5__11464_ (
);

FILL FILL_1__9166_ (
);

FILL FILL_5__11044_ (
);

FILL FILL_2__16356_ (
);

FILL FILL_4__7591_ (
);

FILL FILL_4__7171_ (
);

FILL FILL_4__10877_ (
);

FILL SFILL48920x34050 (
);

FILL FILL_4__10037_ (
);

FILL FILL_2__11491_ (
);

FILL FILL_2__11071_ (
);

FILL FILL_1__15769_ (
);

FILL FILL_1__15349_ (
);

FILL FILL_1__10064_ (
);

INVX1 _14627_ (
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_5115_)
);

INVX1 _14207_ (
    .A(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_4704_)
);

FILL FILL_0__7491_ (
);

FILL FILL_2__7089_ (
);

FILL FILL_0__7071_ (
);

FILL SFILL48520x20050 (
);

FILL FILL_3__10811_ (
);

FILL FILL_4__14290_ (
);

FILL FILL_0__15703_ (
);

FILL SFILL13720x28050 (
);

FILL FILL_2__8870_ (
);

FILL FILL_2__8450_ (
);

FILL FILL_5__12249_ (
);

FILL FILL_3__13283_ (
);

NAND2X1 _6969_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_47_)
);

FILL FILL_4__8376_ (
);

FILL FILL_2__12696_ (
);

FILL FILL_2__12276_ (
);

FILL FILL_5__13610_ (
);

DFFSR _7910_ (
    .Q(\datapath_1.regfile_1.regOut[8] [16]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_458_[16])
);

FILL FILL_1__11689_ (
);

FILL FILL_1__11269_ (
);

FILL FILL_4__12603_ (
);

FILL FILL_0__8696_ (
);

FILL FILL_5__16082_ (
);

INVX1 _10967_ (
    .A(\control_1.op [0]),
    .Y(_2042_)
);

FILL FILL_6__9663_ (
);

FILL FILL_0__8276_ (
);

NAND2X1 _10547_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1863_)
);

NAND2X1 _10127_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1644_)
);

FILL FILL_1__12630_ (
);

FILL FILL_4__15495_ (
);

FILL FILL_4__15075_ (
);

FILL FILL_1__12210_ (
);

FILL FILL_2__9655_ (
);

FILL FILL_3__14488_ (
);

FILL FILL_0__11623_ (
);

FILL FILL_2__9235_ (
);

FILL FILL_3__14068_ (
);

FILL FILL_0__11203_ (
);

FILL SFILL83960x72050 (
);

FILL FILL_5__7240_ (
);

FILL SFILL3560x76050 (
);

NOR2X1 _14380_ (
    .A(_4860_),
    .B(_4872_),
    .Y(_4873_)
);

FILL FILL_0__14095_ (
);

FILL FILL_5__14815_ (
);

FILL FILL_1__7232_ (
);

FILL FILL_4__13808_ (
);

FILL SFILL99160x43050 (
);

FILL FILL_2__14842_ (
);

FILL FILL_3__7998_ (
);

FILL FILL_2__14422_ (
);

FILL FILL_2__14002_ (
);

FILL FILL_3__7578_ (
);

FILL FILL_3__7158_ (
);

FILL FILL_1__13835_ (
);

FILL FILL_1__13415_ (
);

FILL FILL_0__12828_ (
);

FILL FILL_0__12408_ (
);

FILL SFILL38840x39050 (
);

FILL FILL_5__8865_ (
);

FILL FILL_5__8445_ (
);

NAND3X1 _15585_ (
    .A(_6050_),
    .B(_6051_),
    .C(_6049_),
    .Y(_6052_)
);

NAND2X1 _15165_ (
    .A(_5642_),
    .B(_5638_),
    .Y(_5643_)
);

FILL FILL_3__16214_ (
);

FILL SFILL28920x75050 (
);

FILL SFILL3560x31050 (
);

FILL FILL_1__8857_ (
);

FILL FILL_5__10315_ (
);

FILL FILL_1__8017_ (
);

FILL FILL_2__15627_ (
);

FILL FILL_2__15207_ (
);

FILL FILL_4__6862_ (
);

FILL FILL_0__16241_ (
);

FILL FILL_2__10762_ (
);

INVX1 _7087_ (
    .A(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_105_)
);

FILL FILL112200x26050 (
);

FILL SFILL99480x19050 (
);

FILL FILL_3__9724_ (
);

FILL SFILL3480x38050 (
);

FILL FILL_4__13981_ (
);

FILL FILL_4__13561_ (
);

FILL FILL_4__13141_ (
);

AOI21X1 _11085_ (
    .A(_2201_),
    .B(_2188_),
    .C(_2203_),
    .Y(_2204_)
);

FILL FILL_3__12974_ (
);

FILL FILL_2__7721_ (
);

FILL FILL_2__7301_ (
);

FILL FILL_3__12134_ (
);

FILL SFILL28920x30050 (
);

FILL FILL_4__7227_ (
);

FILL FILL_2__11967_ (
);

FILL FILL_2__11547_ (
);

FILL FILL_0__12581_ (
);

FILL FILL_2__11127_ (
);

FILL FILL_0__12161_ (
);

FILL FILL_6__16360_ (
);

FILL SFILL89960x24050 (
);

FILL FILL_5__15773_ (
);

FILL FILL_5__15353_ (
);

FILL FILL_0__7967_ (
);

FILL FILL_0__7547_ (
);

INVX1 _9653_ (
    .A(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_1409_)
);

INVX1 _9233_ (
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_1190_)
);

FILL FILL_1__8190_ (
);

FILL SFILL28840x37050 (
);

FILL FILL_1__11901_ (
);

FILL FILL_4__14766_ (
);

FILL FILL_4__14346_ (
);

FILL FILL_2__15380_ (
);

FILL FILL_2__8506_ (
);

FILL FILL_3__13759_ (
);

FILL FILL_3__13339_ (
);

FILL FILL_1__14793_ (
);

FILL FILL_1__14373_ (
);

FILL FILL_5__6931_ (
);

FILL FILL_0__13786_ (
);

OAI22X1 _13651_ (
    .A(_3916_),
    .B(_4157_),
    .C(_3971__bF$buf1),
    .D(_4158_),
    .Y(_4159_)
);

FILL FILL_0__13366_ (
);

NAND2X1 _13231_ (
    .A(_3770_),
    .B(_3758_),
    .Y(_3774_)
);

FILL FILL_3__14700_ (
);

FILL FILL_1__6923_ (
);

FILL FILL_6__12280_ (
);

FILL SFILL115000x14050 (
);

FILL FILL_3__6849_ (
);

FILL FILL_5__16138_ (
);

FILL FILL_5__11693_ (
);

FILL FILL_1__9395_ (
);

FILL FILL_5__11273_ (
);

FILL FILL_2__16165_ (
);

FILL FILL_4__10686_ (
);

FILL FILL_4__10266_ (
);

FILL FILL_1__15998_ (
);

FILL FILL_1__15578_ (
);

FILL FILL_1__15158_ (
);

FILL FILL_5__7716_ (
);

FILL FILL_2_BUFX2_insert500 (
);

FILL FILL_2_BUFX2_insert501 (
);

FILL FILL_1__10293_ (
);

FILL FILL_2_BUFX2_insert502 (
);

FILL FILL_2_BUFX2_insert503 (
);

OAI22X1 _14856_ (
    .A(_3905__bF$buf1),
    .B(_5338_),
    .C(_3930__bF$buf3),
    .D(_5337_),
    .Y(_5339_)
);

OAI22X1 _14436_ (
    .A(_3960_),
    .B(_4927_),
    .C(_3944__bF$buf1),
    .D(_4926_),
    .Y(_4928_)
);

FILL FILL_2_BUFX2_insert504 (
);

FILL FILL_2_BUFX2_insert505 (
);

INVX1 _14016_ (
    .A(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_4517_)
);

FILL FILL_2_BUFX2_insert506 (
);

FILL FILL_3__15905_ (
);

FILL FILL_2_BUFX2_insert507 (
);

FILL FILL_2_BUFX2_insert508 (
);

FILL FILL_2_BUFX2_insert509 (
);

FILL FILL_1__7708_ (
);

FILL FILL_6__13485_ (
);

FILL FILL_3__10620_ (
);

FILL FILL_0_CLKBUF1_insert200 (
);

FILL FILL_0_CLKBUF1_insert201 (
);

FILL FILL_0__15932_ (
);

FILL FILL_0_CLKBUF1_insert202 (
);

FILL FILL_0_CLKBUF1_insert203 (
);

FILL FILL_0__15512_ (
);

FILL FILL_0_CLKBUF1_insert204 (
);

FILL FILL_0_CLKBUF1_insert205 (
);

FILL FILL_5__12898_ (
);

FILL FILL_0_CLKBUF1_insert206 (
);

FILL FILL_5__12478_ (
);

FILL FILL_0_CLKBUF1_insert207 (
);

FILL FILL_5__12058_ (
);

FILL FILL_0_CLKBUF1_insert208 (
);

FILL FILL_3__13092_ (
);

FILL FILL_0_CLKBUF1_insert209 (
);

FILL FILL_4__8185_ (
);

FILL SFILL18840x35050 (
);

FILL FILL_2__12085_ (
);

FILL FILL_1__11498_ (
);

FILL FILL_1__11078_ (
);

FILL FILL_4__12832_ (
);

FILL FILL_4__12412_ (
);

FILL FILL_6__9472_ (
);

NAND2X1 _10776_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1975_)
);

FILL FILL_0__8085_ (
);

DFFSR _10356_ (
    .Q(\datapath_1.regfile_1.regOut[27] [30]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_1693_[30])
);

FILL FILL_3__11825_ (
);

FILL FILL_3__11405_ (
);

FILL FILL_4__6918_ (
);

FILL FILL_2__9884_ (
);

FILL FILL_2__10818_ (
);

FILL FILL_2__9464_ (
);

FILL FILL_0__11852_ (
);

FILL FILL_3__14297_ (
);

FILL FILL_2__9044_ (
);

FILL FILL_0__11432_ (
);

FILL FILL_0__11012_ (
);

FILL FILL_5__14624_ (
);

FILL FILL_5__14204_ (
);

DFFSR _8924_ (
    .Q(\datapath_1.regfile_1.regOut[16] [6]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_978_[6])
);

INVX1 _8504_ (
    .A(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_826_)
);

FILL FILL_1__7881_ (
);

FILL FILL_1__7461_ (
);

FILL FILL_1__7041_ (
);

FILL FILL_4__13617_ (
);

FILL FILL_2__14651_ (
);

FILL FILL_2__14231_ (
);

FILL FILL_1__13644_ (
);

FILL FILL_1__13224_ (
);

FILL FILL_4__16089_ (
);

FILL FILL_1_BUFX2_insert520 (
);

FILL FILL_1_BUFX2_insert521 (
);

FILL FILL_0__12637_ (
);

DFFSR _12922_ (
    .Q(\datapath_1.a [3]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3555_[3])
);

FILL FILL_1_BUFX2_insert522 (
);

FILL SFILL114520x83050 (
);

FILL FILL_1_BUFX2_insert523 (
);

INVX1 _12502_ (
    .A(ALUOut[21]),
    .Y(_3401_)
);

FILL FILL_0__12217_ (
);

FILL FILL_1_BUFX2_insert524 (
);

FILL FILL_1_BUFX2_insert525 (
);

FILL FILL_6__16416_ (
);

FILL FILL_1_BUFX2_insert526 (
);

FILL FILL_5__8254_ (
);

FILL FILL_1_BUFX2_insert527 (
);

FILL FILL_1_BUFX2_insert528 (
);

FILL FILL_1_BUFX2_insert529 (
);

OAI22X1 _15394_ (
    .A(_5865_),
    .B(_5544__bF$buf2),
    .C(_5480__bF$buf0),
    .D(_4373_),
    .Y(_5866_)
);

FILL FILL_5__15829_ (
);

FILL FILL_5__15409_ (
);

DFFSR _9709_ (
    .Q(\datapath_1.regfile_1.regOut[22] [23]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1368_[23])
);

FILL FILL_3__16023_ (
);

FILL FILL_5__10964_ (
);

FILL FILL_5__10544_ (
);

FILL FILL_5__10124_ (
);

FILL FILL_1__8246_ (
);

FILL FILL_2__15856_ (
);

FILL FILL_2__15436_ (
);

FILL FILL_2__15016_ (
);

FILL FILL_0__16050_ (
);

FILL SFILL48920x29050 (
);

FILL FILL_2__10991_ (
);

FILL FILL_2__10571_ (
);

FILL FILL_2__10151_ (
);

FILL FILL_1__14849_ (
);

FILL FILL_1__14429_ (
);

FILL FILL_1__14009_ (
);

FILL FILL_3__9533_ (
);

FILL FILL_3__9113_ (
);

INVX1 _13707_ (
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_4214_)
);

FILL FILL_0__6991_ (
);

FILL FILL_5__9879_ (
);

FILL FILL_5__9039_ (
);

FILL FILL_4__13790_ (
);

FILL FILL_6__12336_ (
);

NOR2X1 _16179_ (
    .A(_6630_),
    .B(_6624_),
    .Y(_6631_)
);

FILL FILL_4__13370_ (
);

FILL FILL_2__7950_ (
);

FILL FILL_5__11749_ (
);

FILL FILL_3__12783_ (
);

FILL FILL_5__11329_ (
);

FILL SFILL38600x51050 (
);

FILL FILL_3__12363_ (
);

FILL FILL_2__7110_ (
);

FILL FILL_4__7876_ (
);

FILL FILL_4__7456_ (
);

FILL FILL_4__7036_ (
);

FILL FILL_2__11776_ (
);

FILL FILL_2__11356_ (
);

FILL FILL_0__12390_ (
);

FILL FILL_1__10769_ (
);

FILL SFILL3640x64050 (
);

FILL FILL_5__15582_ (
);

FILL FILL_5__15162_ (
);

FILL FILL_0__7356_ (
);

FILL FILL_6__8743_ (
);

INVX1 _9882_ (
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_1521_)
);

INVX1 _9462_ (
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_1366_)
);

OAI21X1 _9042_ (
    .A(_1102_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .C(_1103_),
    .Y(_1043_[30])
);

FILL SFILL104520x81050 (
);

FILL SFILL43880x71050 (
);

FILL FILL_4__14995_ (
);

FILL FILL_4__14575_ (
);

FILL FILL_1__11710_ (
);

FILL FILL_4__14155_ (
);

NAND3X1 _12099_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[28]),
    .C(_3032__bF$buf4),
    .Y(_3120_)
);

FILL FILL_3__13988_ (
);

FILL FILL_2__8735_ (
);

FILL SFILL7960x72050 (
);

FILL FILL_0__10703_ (
);

FILL FILL_2__8315_ (
);

FILL FILL_3__13568_ (
);

FILL SFILL3560x2050 (
);

FILL FILL_3__13148_ (
);

FILL FILL_1__14182_ (
);

FILL FILL_6__14902_ (
);

FILL SFILL59080x42050 (
);

FILL FILL_0__13595_ (
);

NOR2X1 _13880_ (
    .A(_4383_),
    .B(_4380_),
    .Y(_4384_)
);

NAND3X1 _13460_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3904_),
    .C(_3883_),
    .Y(_3972_)
);

OAI21X1 _13040_ (
    .A(_3677_),
    .B(vdd),
    .C(_3678_),
    .Y(_3620_[29])
);

FILL FILL_4__9602_ (
);

FILL FILL_2__13922_ (
);

FILL FILL_5__16367_ (
);

FILL FILL_2__13502_ (
);

FILL SFILL3160x57050 (
);

FILL FILL_5__11082_ (
);

FILL SFILL99320x50 (
);

FILL FILL_1__12915_ (
);

FILL FILL_2__16394_ (
);

FILL FILL_4__10495_ (
);

FILL FILL_0__9922_ (
);

FILL FILL_0__11908_ (
);

FILL FILL_0__9502_ (
);

FILL FILL_1__15387_ (
);

FILL FILL_5__7945_ (
);

FILL FILL_4__16301_ (
);

FILL FILL_5__7105_ (
);

FILL SFILL59000x40050 (
);

FILL FILL_6__10822_ (
);

OAI22X1 _14665_ (
    .A(_3902__bF$buf3),
    .B(_5150_),
    .C(_5151_),
    .D(_3935__bF$buf0),
    .Y(_5152_)
);

INVX1 _14245_ (
    .A(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_4741_)
);

FILL FILL_3__15714_ (
);

FILL SFILL3560x26050 (
);

FILL FILL_1__7937_ (
);

FILL SFILL104440x43050 (
);

FILL FILL_2__14707_ (
);

FILL FILL_0__15741_ (
);

FILL FILL_0__15321_ (
);

FILL FILL_5__12287_ (
);

FILL SFILL49000x83050 (
);

FILL FILL_4__12641_ (
);

FILL FILL_4__12221_ (
);

DFFSR _10585_ (
    .Q(\datapath_1.regfile_1.regOut[29] [3]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_1823_[3])
);

FILL FILL_6__9281_ (
);

INVX1 _10165_ (
    .A(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_1669_)
);

FILL FILL_3__11634_ (
);

FILL FILL_3__11214_ (
);

FILL FILL_0__16106_ (
);

FILL FILL_2__10627_ (
);

FILL FILL_2__9273_ (
);

FILL FILL_0__11661_ (
);

FILL FILL_0__11241_ (
);

FILL FILL_6__15020_ (
);

FILL FILL_2__13099_ (
);

FILL FILL_5__14853_ (
);

FILL FILL_5__14433_ (
);

FILL FILL_5__14013_ (
);

INVX1 _8733_ (
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_938_)
);

INVX1 _8313_ (
    .A(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_719_)
);

FILL FILL_1__7690_ (
);

FILL FILL_4__13846_ (
);

FILL FILL_2__14880_ (
);

FILL FILL_4__13426_ (
);

FILL FILL_2__14460_ (
);

FILL FILL_4__13006_ (
);

FILL FILL_2__14040_ (
);

FILL FILL_0__9099_ (
);

FILL FILL_3__7196_ (
);

FILL FILL_3__12839_ (
);

FILL FILL_1__13873_ (
);

FILL FILL_3__12419_ (
);

FILL FILL_1__13453_ (
);

FILL FILL_1__13033_ (
);

FILL FILL_0__12866_ (
);

INVX1 _12731_ (
    .A(\datapath_1.PCJump [14]),
    .Y(_3513_)
);

FILL FILL_0__12446_ (
);

FILL SFILL59000x50 (
);

FILL FILL_0__12026_ (
);

NAND3X1 _12311_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3272_)
);

FILL FILL_5__8483_ (
);

FILL FILL_5__8063_ (
);

FILL FILL_5__15638_ (
);

FILL FILL_5__15218_ (
);

OAI21X1 _9938_ (
    .A(_1557_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .C(_1558_),
    .Y(_1498_[30])
);

FILL FILL_3__16252_ (
);

OAI21X1 _9518_ (
    .A(_1338_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1339_),
    .Y(_1303_[18])
);

FILL FILL_1__8895_ (
);

FILL FILL_5__10773_ (
);

FILL FILL_1__8475_ (
);

FILL FILL_1__8055_ (
);

FILL FILL_2__15665_ (
);

FILL FILL_2__15245_ (
);

FILL SFILL94360x54050 (
);

FILL FILL_2__10380_ (
);

FILL FILL_1__14658_ (
);

FILL FILL_1__14238_ (
);

FILL FILL_3__9762_ (
);

INVX1 _13936_ (
    .A(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_4438_)
);

FILL FILL_3__9342_ (
);

INVX1 _13516_ (
    .A(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_4027_)
);

FILL SFILL79160x34050 (
);

FILL FILL_5__9268_ (
);

FILL FILL_5__11978_ (
);

FILL FILL_5__11558_ (
);

FILL FILL_3__12592_ (
);

FILL FILL_5__11138_ (
);

FILL FILL_3__12172_ (
);

FILL FILL_4__7685_ (
);

FILL FILL_2__11585_ (
);

FILL FILL_2__11165_ (
);

FILL FILL_1__10998_ (
);

FILL FILL_1__10578_ (
);

FILL FILL_1__10158_ (
);

FILL FILL_4__11912_ (
);

FILL FILL_5__15391_ (
);

FILL FILL_0__7585_ (
);

FILL FILL_0__7165_ (
);

DFFSR _9691_ (
    .Q(\datapath_1.regfile_1.regOut[22] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_1368_[5])
);

OAI21X1 _9271_ (
    .A(_1214_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .C(_1215_),
    .Y(_1173_[21])
);

FILL FILL_3__10905_ (
);

FILL FILL_4__14384_ (
);

FILL SFILL8760x71050 (
);

FILL FILL_2__8964_ (
);

FILL FILL_0__10932_ (
);

FILL FILL_3__13797_ (
);

FILL FILL_0__10512_ (
);

FILL FILL_2__8124_ (
);

FILL FILL_3__13377_ (
);

FILL FILL_5__13704_ (
);

FILL SFILL53960x61050 (
);

FILL SFILL84360x52050 (
);

FILL FILL_1__6961_ (
);

FILL FILL_4__9411_ (
);

FILL FILL_2__13731_ (
);

FILL FILL_2__13311_ (
);

FILL FILL_5__16176_ (
);

FILL FILL_3__6887_ (
);

FILL FILL_1__12724_ (
);

FILL FILL_4__15589_ (
);

FILL FILL_4__15169_ (
);

FILL FILL_1__12304_ (
);

FILL FILL_0__9731_ (
);

FILL FILL_2__9749_ (
);

FILL SFILL114520x78050 (
);

FILL FILL_0__11717_ (
);

FILL FILL_1__15196_ (
);

FILL FILL_5__7754_ (
);

FILL FILL_5__7334_ (
);

FILL FILL_4__16110_ (
);

OAI22X1 _14894_ (
    .A(_5374_),
    .B(_3966__bF$buf1),
    .C(_3924__bF$buf2),
    .D(_5375_),
    .Y(_5376_)
);

FILL FILL_6__10631_ (
);

INVX1 _14474_ (
    .A(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_4965_)
);

FILL FILL_0__14189_ (
);

OAI22X1 _14054_ (
    .A(_3916_),
    .B(_4552_),
    .C(_3935__bF$buf3),
    .D(_4553_),
    .Y(_4554_)
);

FILL FILL_5__14909_ (
);

FILL FILL_3__15943_ (
);

FILL FILL_3__15523_ (
);

FILL FILL_3__15103_ (
);

FILL FILL_1__7746_ (
);

FILL FILL_1__7326_ (
);

FILL SFILL69080x39050 (
);

FILL FILL_2__14936_ (
);

FILL FILL_0__15970_ (
);

FILL FILL_2__14516_ (
);

FILL FILL_0__15550_ (
);

FILL FILL_0__15130_ (
);

FILL FILL_5__12096_ (
);

FILL FILL_1__13929_ (
);

FILL SFILL38200x77050 (
);

FILL FILL_1__13509_ (
);

FILL FILL_4__11089_ (
);

FILL FILL_3__8613_ (
);

FILL FILL_5__8959_ (
);

FILL SFILL114520x33050 (
);

FILL FILL_5__8119_ (
);

NAND3X1 _15679_ (
    .A(_6134_),
    .B(_6140_),
    .C(_6143_),
    .Y(_6144_)
);

FILL FILL_4__12870_ (
);

FILL FILL_4__12450_ (
);

AOI21X1 _15259_ (
    .A(_5734_),
    .B(_5706_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [4])
);

FILL FILL_4__12030_ (
);

FILL SFILL3720x52050 (
);

FILL FILL_3__16308_ (
);

FILL FILL_6__9090_ (
);

INVX1 _10394_ (
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_1781_)
);

FILL FILL_5__10829_ (
);

FILL FILL_5__10409_ (
);

FILL FILL_3__11863_ (
);

FILL FILL_5__9900_ (
);

FILL FILL_3__11443_ (
);

FILL FILL_3__11023_ (
);

FILL FILL_4__6956_ (
);

FILL FILL_0__16335_ (
);

NOR2X1 _16200_ (
    .A(_6648_),
    .B(_6651_),
    .Y(_6652_)
);

FILL FILL_2__10436_ (
);

FILL FILL_0__11890_ (
);

FILL FILL_2__10016_ (
);

FILL FILL_2__9082_ (
);

FILL FILL_0__11470_ (
);

FILL FILL_0__11050_ (
);

FILL SFILL38200x32050 (
);

FILL FILL_5__14662_ (
);

FILL FILL_5__14242_ (
);

FILL FILL_0__6856_ (
);

INVX1 _8962_ (
    .A(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_1050_)
);

DFFSR _8542_ (
    .Q(\datapath_1.regfile_1.regOut[13] [8]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_783_[8])
);

FILL SFILL104520x76050 (
);

OAI21X1 _8122_ (
    .A(_631_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .C(_632_),
    .Y(_588_[22])
);

FILL SFILL43880x66050 (
);

FILL FILL_4__13655_ (
);

FILL FILL_4__13235_ (
);

NAND3X1 _11599_ (
    .A(_2470__bF$buf0),
    .B(_2705_),
    .C(_2702_),
    .Y(_2706_)
);

INVX1 _11179_ (
    .A(\datapath_1.alu_1.ALUInA [24]),
    .Y(_2298_)
);

FILL FILL_2__7815_ (
);

FILL FILL_3__12648_ (
);

FILL FILL_1__13682_ (
);

FILL FILL_3__12228_ (
);

FILL FILL_1__13262_ (
);

FILL FILL_1_BUFX2_insert900 (
);

FILL SFILL59080x37050 (
);

FILL FILL_1_BUFX2_insert901 (
);

INVX1 _12960_ (
    .A(_2_[3]),
    .Y(_3625_)
);

FILL FILL_1_BUFX2_insert902 (
);

FILL FILL_1_BUFX2_insert903 (
);

DFFSR _12540_ (
    .Q(ALUOut[5]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[5])
);

FILL FILL_0__12255_ (
);

FILL FILL_1_BUFX2_insert904 (
);

OAI21X1 _12120_ (
    .A(_3132_),
    .B(ALUSrcA_bF$buf3),
    .C(_3133_),
    .Y(\datapath_1.alu_1.ALUInA [1])
);

FILL FILL_1_BUFX2_insert905 (
);

FILL FILL_1_BUFX2_insert906 (
);

FILL FILL_1_BUFX2_insert907 (
);

FILL FILL_1_BUFX2_insert908 (
);

FILL FILL_1_BUFX2_insert909 (
);

FILL FILL_5__15867_ (
);

FILL FILL_5__15447_ (
);

FILL FILL_5__15027_ (
);

OAI21X1 _9747_ (
    .A(_1450_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1451_),
    .Y(_1433_[9])
);

FILL FILL_3__16061_ (
);

DFFSR _9327_ (
    .Q(\datapath_1.regfile_1.regOut[19] [25]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_1173_[25])
);

FILL SFILL3640x14050 (
);

FILL FILL_5__10162_ (
);

FILL SFILL64760x62050 (
);

FILL FILL_2__15894_ (
);

FILL FILL_2__15474_ (
);

FILL SFILL104520x31050 (
);

FILL FILL_2__15054_ (
);

FILL SFILL43880x21050 (
);

FILL FILL_1__14887_ (
);

FILL FILL_1__14467_ (
);

FILL FILL_1__14047_ (
);

FILL FILL_4__15801_ (
);

FILL FILL_3__9991_ (
);

FILL FILL_3__9151_ (
);

OAI22X1 _13745_ (
    .A(_3960_),
    .B(_4250_),
    .C(_3944__bF$buf0),
    .D(_4249_),
    .Y(_4251_)
);

NAND2X1 _13325_ (
    .A(_3750_),
    .B(_3782_),
    .Y(_3854_)
);

FILL FILL_5__9497_ (
);

FILL SFILL104440x38050 (
);

FILL FILL_0__14821_ (
);

FILL FILL_0__14401_ (
);

FILL FILL_5__11787_ (
);

FILL FILL_5__11367_ (
);

FILL FILL_1__9489_ (
);

FILL FILL_2__16259_ (
);

FILL FILL_4__7494_ (
);

FILL SFILL33880x64050 (
);

FILL FILL_4__7074_ (
);

FILL FILL_2__11394_ (
);

FILL FILL_1__10387_ (
);

FILL SFILL49000x78050 (
);

FILL FILL_4__11721_ (
);

FILL FILL_4__11301_ (
);

FILL FILL_6__8361_ (
);

OAI21X1 _9080_ (
    .A(_1171_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .C(_1172_),
    .Y(_1108_[0])
);

FILL FILL_4__14193_ (
);

FILL FILL_0__15606_ (
);

FILL FILL_2__8773_ (
);

FILL FILL_2__8353_ (
);

FILL FILL_0__10321_ (
);

FILL FILL_4__8699_ (
);

FILL FILL_2__12599_ (
);

FILL FILL_2__12179_ (
);

FILL FILL_5__13933_ (
);

FILL FILL_5__13513_ (
);

INVX1 _7813_ (
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_467_)
);

FILL FILL_4_BUFX2_insert410 (
);

FILL FILL_4__9640_ (
);

FILL FILL_4_BUFX2_insert411 (
);

FILL FILL_4__9220_ (
);

FILL FILL_4_BUFX2_insert412 (
);

FILL FILL_4__12506_ (
);

FILL FILL_4_BUFX2_insert413 (
);

FILL FILL_2__13960_ (
);

FILL FILL_4_BUFX2_insert414 (
);

FILL FILL_2__13540_ (
);

FILL FILL_4_BUFX2_insert415 (
);

FILL FILL_0__8599_ (
);

FILL FILL_2__13120_ (
);

FILL SFILL49000x33050 (
);

FILL FILL_4_BUFX2_insert416 (
);

FILL FILL_6__9146_ (
);

FILL FILL_4_BUFX2_insert417 (
);

FILL FILL_4_BUFX2_insert418 (
);

FILL FILL_4_BUFX2_insert419 (
);

FILL FILL_3__11919_ (
);

FILL FILL_1__12953_ (
);

FILL FILL_4__15398_ (
);

FILL FILL_1__12533_ (
);

FILL FILL_1__12113_ (
);

FILL FILL_2__9978_ (
);

FILL SFILL94440x42050 (
);

FILL FILL_0__11946_ (
);

FILL FILL_0__9540_ (
);

FILL FILL_0__9120_ (
);

FILL FILL_2__9138_ (
);

AND2X2 _11811_ (
    .A(_2901_),
    .B(_2124_),
    .Y(_2902_)
);

FILL FILL_0__11526_ (
);

FILL FILL_0__11106_ (
);

FILL FILL_6__15725_ (
);

FILL FILL_5__7983_ (
);

FILL FILL_5__7563_ (
);

AOI22X1 _14283_ (
    .A(\datapath_1.regfile_1.regOut[18] [17]),
    .B(_4135_),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_4778_)
);

FILL FILL_5__14718_ (
);

FILL FILL_3__15752_ (
);

FILL SFILL54280x53050 (
);

FILL FILL_3__15332_ (
);

FILL FILL_1__7975_ (
);

FILL FILL_1__7555_ (
);

FILL FILL_2__14745_ (
);

FILL FILL_2__14325_ (
);

FILL SFILL39000x76050 (
);

FILL SFILL94360x49050 (
);

FILL FILL_1__13738_ (
);

FILL FILL_1__13318_ (
);

FILL FILL_3__8842_ (
);

FILL FILL_3__8002_ (
);

FILL SFILL79160x29050 (
);

FILL FILL_5__8768_ (
);

FILL FILL_5__8348_ (
);

FILL FILL_6__11645_ (
);

INVX1 _15488_ (
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_5958_)
);

NAND2X1 _15068_ (
    .A(_5500__bF$buf2),
    .B(_5465_),
    .Y(_5548_)
);

FILL FILL_3__16117_ (
);

FILL FILL_5__10638_ (
);

FILL FILL_3__11672_ (
);

FILL FILL_3__11252_ (
);

FILL FILL_0__16144_ (
);

FILL FILL_2__10665_ (
);

FILL FILL_2__10245_ (
);

FILL SFILL39000x31050 (
);

FILL FILL_3__9627_ (
);

FILL FILL_3_BUFX2_insert430 (
);

FILL FILL_3_BUFX2_insert431 (
);

FILL FILL_3__9207_ (
);

FILL FILL_5__14891_ (
);

FILL FILL_3_BUFX2_insert432 (
);

FILL FILL_3_BUFX2_insert433 (
);

FILL FILL_5__14471_ (
);

FILL FILL_3_BUFX2_insert434 (
);

FILL FILL_5__14051_ (
);

FILL FILL_3_BUFX2_insert435 (
);

FILL FILL_6__7632_ (
);

OAI21X1 _8771_ (
    .A(_962_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_963_),
    .Y(_913_[25])
);

FILL FILL_3_BUFX2_insert436 (
);

OAI21X1 _8351_ (
    .A(_743_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .C(_744_),
    .Y(_718_[13])
);

FILL FILL_3_BUFX2_insert437 (
);

FILL FILL_3_BUFX2_insert438 (
);

FILL FILL_4__13884_ (
);

FILL FILL_3_BUFX2_insert439 (
);

FILL FILL_4__13464_ (
);

FILL FILL_4__13044_ (
);

FILL SFILL4040x44050 (
);

FILL FILL_3__12877_ (
);

FILL FILL_2__7624_ (
);

FILL FILL_2__7204_ (
);

FILL FILL_3__12457_ (
);

FILL FILL_3__12037_ (
);

FILL FILL_1__13491_ (
);

FILL FILL_0__12484_ (
);

FILL SFILL114600x66050 (
);

FILL FILL_0__12064_ (
);

FILL SFILL53960x56050 (
);

FILL SFILL84360x47050 (
);

FILL FILL_6__16263_ (
);

FILL FILL_4__8911_ (
);

FILL FILL_5__15676_ (
);

FILL FILL_5__15256_ (
);

OAI21X1 _9976_ (
    .A(_1626_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .C(_1627_),
    .Y(_1563_[0])
);

FILL FILL_3__16290_ (
);

FILL FILL_6__8837_ (
);

NAND2X1 _9556_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1365_)
);

NAND2X1 _9136_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1146_)
);

FILL FILL_5__10391_ (
);

FILL FILL_1__8093_ (
);

FILL FILL_1__11804_ (
);

FILL FILL_4__14669_ (
);

FILL FILL_4__14249_ (
);

FILL FILL_2__15283_ (
);

FILL FILL_2__8829_ (
);

FILL SFILL8760x21050 (
);

FILL FILL_1__14696_ (
);

FILL FILL_1__14276_ (
);

FILL FILL_0_BUFX2_insert560 (
);

FILL FILL_4__15610_ (
);

FILL FILL_0_BUFX2_insert561 (
);

FILL FILL_0_BUFX2_insert562 (
);

FILL FILL_0_BUFX2_insert563 (
);

FILL FILL_3__9380_ (
);

FILL FILL_0_BUFX2_insert564 (
);

FILL FILL_0__13689_ (
);

NOR2X1 _13974_ (
    .A(_4475_),
    .B(_4465_),
    .Y(_4476_)
);

FILL FILL_0__13269_ (
);

FILL FILL_0_BUFX2_insert565 (
);

OAI22X1 _13554_ (
    .A(_3881_),
    .B(_4062_),
    .C(_3966__bF$buf2),
    .D(_4063_),
    .Y(_4064_)
);

FILL FILL_0_BUFX2_insert566 (
);

NAND2X1 _13134_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [18]),
    .Y(_3721_)
);

FILL FILL_0_BUFX2_insert567 (
);

FILL FILL_3__14603_ (
);

FILL FILL_0_BUFX2_insert568 (
);

FILL FILL_0_BUFX2_insert569 (
);

FILL SFILL114120x59050 (
);

FILL SFILL53960x11050 (
);

FILL FILL_6__12183_ (
);

FILL FILL_0__14630_ (
);

FILL FILL_0__14210_ (
);

FILL FILL_5__11596_ (
);

FILL FILL_5__11176_ (
);

FILL FILL_1__9298_ (
);

FILL FILL_2__16068_ (
);

FILL FILL_4__10169_ (
);

FILL SFILL114520x28050 (
);

FILL FILL_5__7619_ (
);

FILL FILL_1__10196_ (
);

FILL FILL_4__11950_ (
);

INVX1 _14759_ (
    .A(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_5244_)
);

OAI22X1 _14339_ (
    .A(_3983__bF$buf3),
    .B(_4831_),
    .C(_3971__bF$buf3),
    .D(_4832_),
    .Y(_4833_)
);

FILL FILL_4__11530_ (
);

FILL SFILL3720x47050 (
);

FILL FILL_4__11110_ (
);

FILL FILL_3__15808_ (
);

FILL FILL_1__16002_ (
);

FILL SFILL104600x64050 (
);

FILL FILL_3__10943_ (
);

FILL FILL_6__13388_ (
);

FILL FILL_3__10523_ (
);

FILL FILL_3__10103_ (
);

FILL FILL_0__15835_ (
);

NOR2X1 _15700_ (
    .A(_4753_),
    .B(_5534__bF$buf2),
    .Y(_6164_)
);

FILL FILL_0__15415_ (
);

FILL FILL_0__10970_ (
);

FILL FILL_2__8582_ (
);

FILL FILL_0__10550_ (
);

FILL FILL_0__10130_ (
);

FILL FILL_4__8088_ (
);

FILL FILL_5__13742_ (
);

FILL FILL_5__13322_ (
);

OAI21X1 _7622_ (
    .A(_379_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .C(_380_),
    .Y(_328_[26])
);

OAI21X1 _7202_ (
    .A(_160_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_161_),
    .Y(_133_[14])
);

FILL FILL_4__12735_ (
);

FILL FILL_4__12315_ (
);

OAI21X1 _10679_ (
    .A(_1929_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1930_),
    .Y(_1888_[21])
);

OAI21X1 _10259_ (
    .A(_1710_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .C(_1711_),
    .Y(_1693_[9])
);

FILL FILL_3__11728_ (
);

FILL FILL_1__12762_ (
);

FILL FILL_3__11308_ (
);

FILL FILL_1__12342_ (
);

FILL FILL112280x65050 (
);

FILL FILL_2__9787_ (
);

FILL FILL_2__9367_ (
);

FILL FILL_0__11755_ (
);

FILL FILL_0__11335_ (
);

OAI22X1 _11620_ (
    .A(_2480_),
    .B(_2418_),
    .C(_2419_),
    .D(_2344__bF$buf3),
    .Y(_2725_)
);

NOR2X1 _11200_ (
    .A(_2317_),
    .B(_2318_),
    .Y(_2319_)
);

FILL FILL_5__7372_ (
);

FILL FILL_5__14947_ (
);

NOR2X1 _14092_ (
    .A(_4587_),
    .B(_4590_),
    .Y(_4591_)
);

FILL FILL_3__15981_ (
);

FILL FILL_5__14527_ (
);

FILL FILL_3__15561_ (
);

FILL FILL_5__14107_ (
);

FILL FILL_3__15141_ (
);

OAI21X1 _8827_ (
    .A(_979_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .C(_980_),
    .Y(_978_[1])
);

DFFSR _8407_ (
    .Q(\datapath_1.regfile_1.regOut[12] [1]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_718_[1])
);

FILL FILL_1__7364_ (
);

FILL FILL_2__14974_ (
);

FILL SFILL104520x26050 (
);

FILL FILL_2__14554_ (
);

FILL SFILL43880x16050 (
);

FILL FILL_2__14134_ (
);

FILL FILL_1__13967_ (
);

FILL FILL_1__13547_ (
);

FILL FILL_1__13127_ (
);

FILL FILL_1_CLKBUF1_insert1074 (
);

FILL FILL_3__8651_ (
);

FILL FILL_3__8231_ (
);

OAI21X1 _12825_ (
    .A(_3618_),
    .B(vdd),
    .C(_3619_),
    .Y(_3555_[0])
);

FILL FILL_1_CLKBUF1_insert1075 (
);

OAI21X1 _12405_ (
    .A(_3334_),
    .B(MemToReg_bF$buf0),
    .C(_3335_),
    .Y(\datapath_1.mux_wd3.dout [20])
);

FILL FILL_1_CLKBUF1_insert1076 (
);

FILL FILL_1_CLKBUF1_insert1077 (
);

FILL FILL112280x20050 (
);

FILL FILL_1_CLKBUF1_insert1078 (
);

FILL FILL_5__8997_ (
);

FILL SFILL84280x3050 (
);

FILL FILL_5__8577_ (
);

FILL FILL_6__16319_ (
);

FILL FILL_1_CLKBUF1_insert1079 (
);

NAND2X1 _15297_ (
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .B(_5481_),
    .Y(_5771_)
);

FILL FILL_0__13901_ (
);

FILL SFILL28200x25050 (
);

FILL FILL_3__16346_ (
);

FILL FILL_1__8989_ (
);

FILL FILL_5__10447_ (
);

FILL FILL_1__8569_ (
);

FILL FILL_1__8149_ (
);

FILL FILL_5__10027_ (
);

FILL FILL_3__11481_ (
);

FILL FILL_3__11061_ (
);

FILL FILL_2__15759_ (
);

FILL FILL_2__15339_ (
);

FILL FILL_4__6994_ (
);

FILL SFILL33880x59050 (
);

FILL FILL_0__16373_ (
);

FILL FILL_2__10894_ (
);

FILL FILL_2__10054_ (
);

FILL FILL_1__9930_ (
);

FILL FILL_1__9510_ (
);

FILL FILL_3__9856_ (
);

FILL FILL_3__9016_ (
);

FILL FILL_4__10801_ (
);

FILL FILL_0__6894_ (
);

FILL FILL_5__14280_ (
);

OAI21X1 _8580_ (
    .A(_855_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .C(_856_),
    .Y(_848_[4])
);

FILL FILL_6__7441_ (
);

DFFSR _8160_ (
    .Q(\datapath_1.regfile_1.regOut[10] [10]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_588_[10])
);

FILL FILL_6__12239_ (
);

FILL FILL_4__13693_ (
);

FILL FILL_4__13273_ (
);

FILL FILL_2__7853_ (
);

FILL FILL_2__7433_ (
);

FILL FILL_3__12266_ (
);

FILL FILL_4__7359_ (
);

FILL FILL_2__11679_ (
);

FILL FILL_2__11259_ (
);

FILL FILL_0__12293_ (
);

FILL FILL_4__8720_ (
);

FILL FILL_2__12620_ (
);

FILL FILL_5__15485_ (
);

FILL FILL_0__7679_ (
);

FILL FILL_5__15065_ (
);

FILL FILL_2__12200_ (
);

NAND2X1 _9785_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1477_)
);

FILL FILL_6__8226_ (
);

NAND2X1 _9365_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1258_)
);

FILL FILL_4__14898_ (
);

FILL FILL_4__14478_ (
);

FILL FILL_1__11613_ (
);

FILL FILL_4__14058_ (
);

FILL FILL_2__15092_ (
);

FILL FILL_2__8638_ (
);

FILL FILL_0__8620_ (
);

FILL FILL_0__8200_ (
);

FILL FILL_2__8218_ (
);

FILL FILL_1__14085_ (
);

FILL FILL_6__14805_ (
);

INVX1 _13783_ (
    .A(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_4289_)
);

FILL FILL_0__13498_ (
);

NAND2X1 _13363_ (
    .A(\datapath_1.a3 [1]),
    .B(_3875_),
    .Y(_3877_)
);

FILL SFILL23880x57050 (
);

FILL FILL_3__14832_ (
);

FILL FILL_3__14412_ (
);

FILL FILL_4__9925_ (
);

FILL FILL_4__9505_ (
);

FILL FILL_2__13825_ (
);

FILL FILL_2__13405_ (
);

FILL FILL_2__16297_ (
);

CLKBUF1 CLKBUF1_insert111 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf113)
);

CLKBUF1 CLKBUF1_insert112 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf112)
);

FILL FILL_4__10398_ (
);

CLKBUF1 CLKBUF1_insert113 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf111)
);

FILL FILL_3__7502_ (
);

CLKBUF1 CLKBUF1_insert114 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf110)
);

FILL FILL_0__9405_ (
);

CLKBUF1 CLKBUF1_insert115 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf109)
);

CLKBUF1 CLKBUF1_insert116 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf108)
);

CLKBUF1 CLKBUF1_insert117 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf107)
);

FILL FILL_5__7848_ (
);

CLKBUF1 CLKBUF1_insert118 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf106)
);

CLKBUF1 CLKBUF1_insert119 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf105)
);

FILL FILL_5__7428_ (
);

FILL FILL_4__16204_ (
);

AND2X2 _14988_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5468_)
);

NOR2X1 _14568_ (
    .A(_5053_),
    .B(_5056_),
    .Y(_5057_)
);

FILL FILL_6__10305_ (
);

FILL SFILL23800x55050 (
);

INVX1 _14148_ (
    .A(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_4646_)
);

FILL FILL_3__15617_ (
);

FILL FILL_1__16231_ (
);

FILL SFILL79320x4050 (
);

FILL SFILL23880x12050 (
);

FILL FILL_3__10752_ (
);

FILL SFILL79240x9050 (
);

FILL FILL_0__15644_ (
);

FILL FILL_0__15224_ (
);

FILL FILL_2__8391_ (
);

FILL SFILL39000x26050 (
);

FILL FILL_3__8707_ (
);

FILL FILL_5__13971_ (
);

FILL FILL_5__13551_ (
);

FILL FILL_5__13131_ (
);

OAI21X1 _7851_ (
    .A(_491_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .C(_492_),
    .Y(_458_[17])
);

OAI21X1 _7431_ (
    .A(_272_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .C(_273_),
    .Y(_263_[5])
);

DFFSR _7011_ (
    .Q(\datapath_1.regfile_1.regOut[1] [13]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_3_[13])
);

FILL FILL_4__12964_ (
);

FILL FILL_4__12124_ (
);

OAI21X1 _10488_ (
    .A(_1886_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1887_),
    .Y(_1823_[0])
);

NAND2X1 _10068_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1625_)
);

FILL SFILL23800x10050 (
);

FILL FILL_3__11957_ (
);

FILL FILL_1__12991_ (
);

FILL FILL_3__11537_ (
);

FILL FILL_1__12571_ (
);

FILL FILL_3__11117_ (
);

FILL FILL_1__12151_ (
);

FILL SFILL84040x21050 (
);

FILL FILL_0__16009_ (
);

FILL FILL_0__11984_ (
);

FILL FILL_2__9596_ (
);

FILL FILL_0__11564_ (
);

FILL FILL_0__11144_ (
);

FILL FILL_5__7181_ (
);

FILL FILL_5__14756_ (
);

FILL FILL_3__15790_ (
);

FILL FILL_5__14336_ (
);

FILL FILL_3__15370_ (
);

NAND2X1 _8636_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_894_)
);

NAND2X1 _8216_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_675_)
);

FILL FILL_1__7593_ (
);

FILL FILL_1__7173_ (
);

FILL FILL_4__13749_ (
);

FILL FILL_4__13329_ (
);

FILL FILL_2__14783_ (
);

FILL FILL_2__14363_ (
);

FILL FILL_3__7099_ (
);

FILL SFILL8760x16050 (
);

FILL SFILL13800x53050 (
);

FILL FILL_1__13776_ (
);

FILL FILL_1__13356_ (
);

FILL SFILL13880x10050 (
);

FILL FILL_3__8880_ (
);

FILL FILL_0__12769_ (
);

FILL FILL_3__8460_ (
);

NAND2X1 _12634_ (
    .A(vdd),
    .B(memoryOutData[22]),
    .Y(_3469_)
);

FILL FILL_0__12349_ (
);

NAND3X1 _12214_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\aluControl_1.inst [0]),
    .C(_3198__bF$buf1),
    .Y(_3199_)
);

FILL FILL_5__8386_ (
);

FILL SFILL114600x16050 (
);

FILL FILL_0__13710_ (
);

FILL FILL_3__16155_ (
);

FILL FILL_5__10676_ (
);

FILL FILL_5__10256_ (
);

FILL FILL_1__8378_ (
);

FILL FILL_3__11290_ (
);

FILL FILL_2__15988_ (
);

FILL FILL_2__15568_ (
);

FILL FILL_2__15148_ (
);

FILL FILL_0__16182_ (
);

FILL FILL_2__10283_ (
);

FILL FILL_3_BUFX2_insert810 (
);

FILL FILL_3__9665_ (
);

NOR2X1 _13839_ (
    .A(_4331_),
    .B(_4343_),
    .Y(_4344_)
);

FILL FILL_3_BUFX2_insert811 (
);

FILL FILL_3__9245_ (
);

NAND2X1 _13419_ (
    .A(_3889_),
    .B(_3919_),
    .Y(_3931_)
);

FILL FILL_3_BUFX2_insert812 (
);

FILL FILL_3_BUFX2_insert813 (
);

FILL FILL_3_BUFX2_insert814 (
);

FILL FILL_1__15922_ (
);

FILL FILL_3_BUFX2_insert815 (
);

FILL FILL_3_BUFX2_insert816 (
);

FILL FILL_1__15502_ (
);

FILL FILL_3_BUFX2_insert817 (
);

FILL SFILL43960x49050 (
);

FILL FILL_3_BUFX2_insert818 (
);

FILL FILL_3_BUFX2_insert819 (
);

FILL FILL_4__13082_ (
);

FILL FILL_0__14915_ (
);

FILL SFILL49640x9050 (
);

FILL FILL_2__7242_ (
);

FILL FILL_3__12495_ (
);

FILL FILL_3__12075_ (
);

FILL FILL_4__7588_ (
);

FILL FILL_4__7168_ (
);

FILL FILL112360x53050 (
);

FILL FILL_2__11488_ (
);

FILL FILL_2__11068_ (
);

FILL FILL_5__12402_ (
);

FILL SFILL23960x4050 (
);

FILL FILL_4__11815_ (
);

FILL SFILL23880x9050 (
);

FILL FILL_5__15294_ (
);

FILL FILL_0__7488_ (
);

FILL FILL_0__7068_ (
);

NAND2X1 _9594_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1370_)
);

DFFSR _9174_ (
    .Q(\datapath_1.regfile_1.regOut[18] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_1108_[0])
);

FILL FILL_3__10808_ (
);

FILL FILL_1__11842_ (
);

FILL FILL_4__14287_ (
);

FILL FILL_1__11422_ (
);

FILL FILL_1__11002_ (
);

FILL FILL_2__8867_ (
);

FILL FILL_2__8447_ (
);

FILL FILL_0__10835_ (
);

OAI21X1 _10700_ (
    .A(_1943_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1944_),
    .Y(_1888_[28])
);

FILL FILL_0__10415_ (
);

FILL FILL_0_BUFX2_insert940 (
);

FILL FILL_5__6872_ (
);

FILL FILL_0_BUFX2_insert941 (
);

FILL FILL_0_BUFX2_insert942 (
);

FILL FILL_0_BUFX2_insert943 (
);

FILL FILL_0_BUFX2_insert944 (
);

AOI22X1 _13592_ (
    .A(_3950__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[11] [3]),
    .C(\datapath_1.regfile_1.regOut[2] [3]),
    .D(_3998__bF$buf2),
    .Y(_4101_)
);

FILL FILL_0_BUFX2_insert945 (
);

FILL SFILL108920x22050 (
);

FILL FILL_0_BUFX2_insert946 (
);

INVX1 _13172_ (
    .A(\datapath_1.PCJump [31]),
    .Y(_3746_)
);

FILL FILL_5__13607_ (
);

FILL FILL_0_BUFX2_insert947 (
);

FILL FILL_3__14641_ (
);

FILL FILL_0_BUFX2_insert948 (
);

FILL FILL_3__14221_ (
);

FILL FILL_0_BUFX2_insert949 (
);

DFFSR _7907_ (
    .Q(\datapath_1.regfile_1.regOut[8] [13]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_458_[13])
);

FILL FILL_1__6864_ (
);

FILL FILL_4__9734_ (
);

FILL FILL_2__13634_ (
);

FILL FILL_2__13214_ (
);

FILL FILL_5__16079_ (
);

FILL FILL_1__12627_ (
);

FILL FILL_1__12207_ (
);

FILL FILL_0__9634_ (
);

FILL FILL_3__7731_ (
);

FILL FILL_3__7311_ (
);

INVX1 _11905_ (
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_2978_)
);

FILL FILL_0__9214_ (
);

FILL FILL112280x15050 (
);

FILL FILL_1__15099_ (
);

FILL FILL_5__7237_ (
);

FILL FILL_4__16013_ (
);

INVX1 _14797_ (
    .A(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_5281_)
);

FILL FILL_6__10114_ (
);

NOR2X1 _14377_ (
    .A(_4869_),
    .B(_3944__bF$buf1),
    .Y(_4870_)
);

FILL FILL_3__15846_ (
);

FILL FILL_3__15426_ (
);

FILL FILL_3__15006_ (
);

FILL FILL_1__16040_ (
);

FILL FILL_3__10981_ (
);

FILL FILL_1__7229_ (
);

FILL FILL_3__10561_ (
);

FILL FILL_6_BUFX2_insert321 (
);

FILL FILL_3__10141_ (
);

FILL FILL_2__14839_ (
);

FILL FILL_2__14419_ (
);

FILL FILL_0__15873_ (
);

FILL FILL_0__15453_ (
);

FILL FILL_0__15033_ (
);

FILL FILL_6_BUFX2_insert326 (
);

FILL FILL_3__8516_ (
);

FILL FILL_5__13780_ (
);

FILL FILL_5__13360_ (
);

DFFSR _7660_ (
    .Q(\datapath_1.regfile_1.regOut[6] [22]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_328_[22])
);

NAND2X1 _7240_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_187_)
);

FILL FILL_4__12773_ (
);

FILL FILL_4__12353_ (
);

NAND2X1 _10297_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1737_)
);

FILL FILL_2__6933_ (
);

FILL FILL_5__9803_ (
);

FILL FILL_3__11766_ (
);

FILL FILL_3__11346_ (
);

FILL FILL_1__12380_ (
);

FILL FILL_4__6859_ (
);

FILL FILL_0__16238_ (
);

NAND2X1 _16103_ (
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .B(_5649_),
    .Y(_6557_)
);

FILL FILL_2__10759_ (
);

FILL FILL_0__11793_ (
);

FILL FILL_0__11373_ (
);

FILL FILL_6__15992_ (
);

FILL FILL_6__15572_ (
);

FILL FILL_4__7800_ (
);

FILL FILL_5__14985_ (
);

FILL FILL_5__14565_ (
);

FILL FILL_2__11700_ (
);

FILL FILL_5__14145_ (
);

NAND2X1 _8865_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1006_)
);

NAND2X1 _8445_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_787_)
);

DFFSR _8025_ (
    .Q(\datapath_1.regfile_1.regOut[9] [3]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_523_[3])
);

FILL FILL_4__13978_ (
);

FILL FILL_4__13558_ (
);

FILL FILL_2__14592_ (
);

FILL FILL_4__13138_ (
);

FILL FILL_2__14172_ (
);

FILL FILL_2__7718_ (
);

FILL FILL_0__7700_ (
);

FILL FILL_1__13585_ (
);

FILL FILL_1__13165_ (
);

FILL FILL_0__12998_ (
);

FILL FILL_0__12578_ (
);

NAND2X1 _12863_ (
    .A(vdd),
    .B(\datapath_1.rd1 [13]),
    .Y(_3581_)
);

FILL FILL_0__12158_ (
);

NAND2X1 _12443_ (
    .A(vdd),
    .B(\datapath_1.ALUResult [1]),
    .Y(_3362_)
);

NAND3X1 _12023_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[9]),
    .C(_3032__bF$buf3),
    .Y(_3063_)
);

FILL FILL_3__13912_ (
);

FILL FILL_5__8195_ (
);

FILL SFILL79160x71050 (
);

FILL SFILL59080x4050 (
);

FILL FILL_6__11492_ (
);

FILL FILL_5_BUFX2_insert340 (
);

FILL FILL_6__11072_ (
);

FILL FILL_5_BUFX2_insert341 (
);

FILL FILL_2__12905_ (
);

FILL FILL_5_BUFX2_insert342 (
);

FILL FILL_3__16384_ (
);

FILL FILL_5_BUFX2_insert343 (
);

FILL FILL_5_BUFX2_insert344 (
);

FILL FILL_5_BUFX2_insert345 (
);

FILL FILL_5_BUFX2_insert346 (
);

FILL FILL_5_BUFX2_insert347 (
);

FILL FILL_1__8187_ (
);

FILL FILL_5__10065_ (
);

FILL FILL_5_BUFX2_insert348 (
);

FILL FILL_2__15797_ (
);

FILL FILL_5_BUFX2_insert349 (
);

FILL FILL_2__15377_ (
);

FILL FILL_0__8905_ (
);

FILL FILL_5__6928_ (
);

FILL FILL_4__15704_ (
);

FILL FILL_3__9894_ (
);

FILL FILL_3__9474_ (
);

NAND3X1 _13648_ (
    .A(_4153_),
    .B(_4155_),
    .C(_4152_),
    .Y(_4156_)
);

INVX1 _13228_ (
    .A(\datapath_1.a3 [2]),
    .Y(_3771_)
);

FILL SFILL109480x5050 (
);

FILL SFILL8040x66050 (
);

FILL FILL_1__15731_ (
);

FILL SFILL84520x23050 (
);

FILL FILL_1__15311_ (
);

FILL FILL_6__12697_ (
);

FILL FILL_0__14724_ (
);

FILL FILL_0__14304_ (
);

FILL FILL_2__7891_ (
);

FILL FILL_2__7471_ (
);

FILL FILL_2__7051_ (
);

FILL FILL_2__11297_ (
);

FILL FILL_5__12631_ (
);

FILL FILL_5__12211_ (
);

OAI21X1 _6931_ (
    .A(_20_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_21_),
    .Y(_3_[9])
);

FILL FILL_2_BUFX2_insert470 (
);

FILL FILL_2_BUFX2_insert471 (
);

FILL FILL_2_BUFX2_insert472 (
);

FILL FILL_2_BUFX2_insert473 (
);

FILL FILL_2_BUFX2_insert474 (
);

FILL FILL_4__11624_ (
);

FILL FILL_2_BUFX2_insert475 (
);

FILL FILL_4__11204_ (
);

FILL FILL_2_BUFX2_insert476 (
);

FILL FILL_0__7297_ (
);

FILL FILL_2_BUFX2_insert477 (
);

FILL FILL_2_BUFX2_insert478 (
);

FILL FILL_2_BUFX2_insert479 (
);

FILL FILL_3__10617_ (
);

FILL FILL_0_CLKBUF1_insert170 (
);

FILL FILL_1__11651_ (
);

FILL FILL_1__11231_ (
);

FILL FILL_4__14096_ (
);

FILL FILL_0_CLKBUF1_insert171 (
);

FILL FILL_0__15929_ (
);

FILL FILL_0_CLKBUF1_insert172 (
);

FILL FILL_0_CLKBUF1_insert173 (
);

FILL FILL_0__15509_ (
);

FILL FILL_0_CLKBUF1_insert174 (
);

FILL FILL_0_CLKBUF1_insert175 (
);

FILL FILL_0_CLKBUF1_insert176 (
);

FILL FILL_2__8256_ (
);

FILL FILL_0_CLKBUF1_insert177 (
);

FILL FILL_0__10644_ (
);

FILL FILL_3__13089_ (
);

FILL FILL_0_CLKBUF1_insert178 (
);

FILL FILL_0_CLKBUF1_insert179 (
);

FILL SFILL109720x21050 (
);

FILL SFILL13480x36050 (
);

FILL FILL_5__13836_ (
);

FILL FILL_3__14870_ (
);

FILL FILL_5__13416_ (
);

FILL FILL_3__14450_ (
);

NAND2X1 _7716_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_423_)
);

FILL FILL_3__14030_ (
);

FILL FILL_4__9543_ (
);

FILL SFILL13000x65050 (
);

FILL FILL_4__9123_ (
);

FILL FILL_4__12829_ (
);

FILL FILL_2__13863_ (
);

FILL FILL_4__12409_ (
);

FILL FILL_2__13443_ (
);

FILL FILL_2__13023_ (
);

FILL SFILL13800x48050 (
);

FILL FILL_1__12856_ (
);

FILL FILL_1__12436_ (
);

FILL FILL_1__12016_ (
);

FILL FILL_3__7960_ (
);

FILL FILL_0__9863_ (
);

FILL FILL_0__11849_ (
);

FILL FILL_0__9023_ (
);

FILL FILL_3__7120_ (
);

FILL FILL_0__11429_ (
);

AND2X2 _11714_ (
    .A(_2812_),
    .B(_2188_),
    .Y(_2813_)
);

FILL FILL_0__11009_ (
);

FILL FILL_5__7886_ (
);

FILL FILL_6__15628_ (
);

FILL FILL_5__7466_ (
);

FILL FILL_4__16242_ (
);

FILL FILL_5__7046_ (
);

AOI22X1 _14186_ (
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .B(_4005__bF$buf3),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_4683_)
);

FILL FILL_3__15655_ (
);

FILL FILL_3__15235_ (
);

FILL FILL_1__7878_ (
);

FILL FILL_3__10790_ (
);

FILL FILL_1__7458_ (
);

FILL FILL_3__10370_ (
);

FILL FILL_1__7038_ (
);

FILL SFILL28840x1050 (
);

FILL FILL_2__14648_ (
);

FILL FILL_0__15682_ (
);

FILL FILL_2__14228_ (
);

FILL FILL_0__15262_ (
);

FILL SFILL28760x6050 (
);

FILL FILL_1_BUFX2_insert490 (
);

FILL SFILL78760x36050 (
);

FILL FILL_3__8745_ (
);

FILL FILL_1_BUFX2_insert491 (
);

DFFSR _12919_ (
    .Q(\datapath_1.a [0]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3555_[0])
);

FILL FILL_1_BUFX2_insert492 (
);

FILL FILL_3__8325_ (
);

FILL FILL_1_BUFX2_insert493 (
);

FILL FILL_1_BUFX2_insert494 (
);

FILL FILL_1_BUFX2_insert495 (
);

FILL FILL_1_BUFX2_insert496 (
);

FILL FILL_1_BUFX2_insert497 (
);

FILL SFILL8680x2050 (
);

FILL FILL_1_BUFX2_insert498 (
);

FILL FILL_6__11968_ (
);

FILL FILL_1_BUFX2_insert499 (
);

FILL FILL_6__11548_ (
);

FILL FILL_4__12582_ (
);

FILL FILL_4__12162_ (
);

FILL SFILL64120x50050 (
);

FILL FILL_3__11995_ (
);

FILL FILL_5__9612_ (
);

FILL FILL_3__11575_ (
);

FILL FILL_3__11155_ (
);

OAI21X1 _16332_ (
    .A(_6774_),
    .B(gnd),
    .C(_6775_),
    .Y(_6769_[3])
);

FILL FILL_0__16047_ (
);

FILL FILL112360x48050 (
);

FILL FILL_2__10988_ (
);

FILL FILL_2__10568_ (
);

FILL FILL_2__10148_ (
);

FILL FILL_0__11182_ (
);

FILL FILL_5__11902_ (
);

FILL FILL_1__9604_ (
);

FILL SFILL68760x79050 (
);

FILL SFILL64040x57050 (
);

FILL FILL_5__14794_ (
);

FILL FILL_0__6988_ (
);

FILL FILL_5__14374_ (
);

DFFSR _8674_ (
    .Q(\datapath_1.regfile_1.regOut[14] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_848_[12])
);

INVX1 _8254_ (
    .A(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_700_)
);

FILL FILL_6__7115_ (
);

FILL FILL_1__10922_ (
);

FILL FILL_4__13787_ (
);

FILL FILL_4__13367_ (
);

FILL FILL_1__10502_ (
);

FILL FILL_2__7947_ (
);

FILL FILL_2__7107_ (
);

FILL FILL_1__13394_ (
);

DFFSR _12672_ (
    .Q(\datapath_1.Data [9]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_3425_[9])
);

FILL FILL_0__12387_ (
);

NAND3X1 _12252_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [11]),
    .C(_3198__bF$buf3),
    .Y(_3228_)
);

FILL FILL_3__13721_ (
);

FILL FILL_3__13301_ (
);

FILL FILL_5__15999_ (
);

FILL FILL_2__12714_ (
);

FILL FILL_5__15579_ (
);

FILL FILL_5__15159_ (
);

FILL FILL_3__16193_ (
);

INVX1 _9879_ (
    .A(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_1519_)
);

DFFSR _9459_ (
    .Q(\datapath_1.regfile_1.regOut[20] [29]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_1238_[29])
);

OAI21X1 _9039_ (
    .A(_1100_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1101_),
    .Y(_1043_[29])
);

FILL SFILL64040x12050 (
);

FILL FILL_5__10294_ (
);

FILL FILL_1__11707_ (
);

FILL FILL_2__15186_ (
);

FILL FILL_0__8714_ (
);

FILL FILL_5__16100_ (
);

FILL SFILL89240x61050 (
);

FILL FILL_1__14599_ (
);

FILL FILL_1__14179_ (
);

FILL FILL_4__15933_ (
);

FILL FILL_4__15513_ (
);

FILL FILL_6_BUFX2_insert1093 (
);

INVX1 _13877_ (
    .A(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_4381_)
);

FILL FILL_3__9283_ (
);

INVX1 _13457_ (
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_3969_)
);

OAI21X1 _13037_ (
    .A(_3675_),
    .B(vdd),
    .C(_3676_),
    .Y(_3620_[28])
);

FILL FILL_3__14926_ (
);

FILL FILL_1__15960_ (
);

FILL FILL_3__14506_ (
);

FILL SFILL18680x81050 (
);

FILL FILL_1__15540_ (
);

FILL FILL_1__15120_ (
);

FILL FILL_2__13919_ (
);

FILL FILL_0__14953_ (
);

FILL FILL_0__14533_ (
);

FILL FILL_0__14113_ (
);

FILL FILL_5__11499_ (
);

FILL SFILL54040x55050 (
);

FILL FILL_5__11079_ (
);

FILL FILL_0__9919_ (
);

FILL FILL_5__12860_ (
);

FILL FILL_5__12440_ (
);

FILL FILL_5__12020_ (
);

FILL FILL_4__11853_ (
);

FILL FILL_4__11433_ (
);

FILL FILL_4__11013_ (
);

FILL FILL_1__16325_ (
);

FILL FILL_1__11880_ (
);

FILL FILL_3__10426_ (
);

FILL FILL_1__11460_ (
);

FILL FILL_3__10006_ (
);

FILL FILL_1__11040_ (
);

FILL FILL_0__15738_ (
);

FILL FILL_0__15318_ (
);

OAI22X1 _15603_ (
    .A(_5495__bF$buf0),
    .B(_4589_),
    .C(_4616_),
    .D(_5534__bF$buf3),
    .Y(_6070_)
);

FILL FILL_2__8485_ (
);

FILL FILL_0__10873_ (
);

FILL FILL_2__8065_ (
);

FILL FILL_0__10453_ (
);

FILL FILL_0__10033_ (
);

FILL FILL_6__14232_ (
);

FILL SFILL54040x10050 (
);

FILL FILL_5__13645_ (
);

FILL FILL_5__13225_ (
);

NAND2X1 _7945_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_535_)
);

DFFSR _7525_ (
    .Q(\datapath_1.regfile_1.regOut[5] [15]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_263_[15])
);

INVX1 _7105_ (
    .A(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_117_)
);

FILL FILL_4__9772_ (
);

FILL FILL_4__9352_ (
);

FILL FILL_4__12638_ (
);

FILL FILL_2__13672_ (
);

FILL FILL_4__12218_ (
);

FILL FILL_2__13252_ (
);

FILL FILL_1__12245_ (
);

FILL FILL_0__9672_ (
);

FILL FILL_0__9252_ (
);

OAI21X1 _11943_ (
    .A(_3002_),
    .B(IorD_bF$buf6),
    .C(_3003_),
    .Y(_1_[18])
);

FILL FILL_0__11658_ (
);

FILL FILL_0__11238_ (
);

INVX1 _11523_ (
    .A(_2278_),
    .Y(_2634_)
);

INVX1 _11103_ (
    .A(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2222_)
);

FILL FILL_5__7695_ (
);

FILL SFILL44040x53050 (
);

FILL FILL_4__16051_ (
);

FILL FILL_3__15884_ (
);

FILL FILL_3__15464_ (
);

FILL FILL_3__15044_ (
);

FILL FILL_1__7687_ (
);

FILL FILL_6_BUFX2_insert700 (
);

FILL FILL_2__14877_ (
);

FILL FILL_2__14457_ (
);

FILL FILL_2__14037_ (
);

FILL FILL_0__15491_ (
);

FILL FILL_0__15071_ (
);

FILL FILL_6_BUFX2_insert705 (
);

FILL FILL_3__8974_ (
);

INVX1 _12728_ (
    .A(\datapath_1.PCJump [13]),
    .Y(_3511_)
);

FILL FILL_3__8134_ (
);

NAND3X1 _12308_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf4),
    .Y(_3270_)
);

FILL FILL_1__14811_ (
);

FILL SFILL109400x40050 (
);

FILL FILL_4__12391_ (
);

FILL FILL_0__13804_ (
);

FILL FILL_3__16249_ (
);

FILL FILL_2__6971_ (
);

FILL FILL_5__9421_ (
);

FILL FILL_3__11384_ (
);

FILL FILL_5__9001_ (
);

FILL FILL_4__6897_ (
);

FILL FILL_0__16276_ (
);

NOR3X1 _16141_ (
    .A(_5515__bF$buf2),
    .B(_5261_),
    .C(_5521__bF$buf1),
    .Y(_6594_)
);

FILL FILL_2__10797_ (
);

FILL FILL_2__10377_ (
);

FILL FILL_5__11711_ (
);

FILL FILL_1__9413_ (
);

FILL FILL_3__9759_ (
);

FILL FILL_3__9339_ (
);

FILL FILL_4__10704_ (
);

FILL FILL_5__14183_ (
);

INVX1 _8483_ (
    .A(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_812_)
);

INVX1 _8063_ (
    .A(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_593_)
);

FILL FILL_4__13596_ (
);

FILL FILL_1__10311_ (
);

FILL SFILL69160x64050 (
);

FILL FILL_2__7756_ (
);

FILL FILL_3__12589_ (
);

FILL FILL_2__7336_ (
);

FILL FILL_3__12169_ (
);

FILL SFILL74120x47050 (
);

INVX1 _12481_ (
    .A(ALUOut[14]),
    .Y(_3387_)
);

FILL FILL_0__12196_ (
);

AOI22X1 _12061_ (
    .A(\datapath_1.ALUResult [18]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3092_)
);

FILL FILL_5__12916_ (
);

FILL FILL_3__13950_ (
);

FILL FILL_3__13530_ (
);

FILL FILL_3__13110_ (
);

FILL FILL_4__8623_ (
);

FILL FILL_4__8203_ (
);

FILL FILL_4__11909_ (
);

FILL FILL_5_BUFX2_insert720 (
);

FILL SFILL34440x20050 (
);

FILL FILL_5_BUFX2_insert721 (
);

FILL FILL_5__15388_ (
);

FILL FILL_2__12523_ (
);

FILL FILL_5_BUFX2_insert722 (
);

FILL FILL_2__12103_ (
);

FILL FILL_5_BUFX2_insert723 (
);

FILL FILL_5_BUFX2_insert724 (
);

DFFSR _9688_ (
    .Q(\datapath_1.regfile_1.regOut[22] [2]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_1368_[2])
);

FILL FILL_5_BUFX2_insert725 (
);

OAI21X1 _9268_ (
    .A(_1212_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1213_),
    .Y(_1173_[20])
);

FILL FILL_5_BUFX2_insert726 (
);

FILL FILL_5_BUFX2_insert727 (
);

FILL FILL_1__11936_ (
);

FILL FILL_5_BUFX2_insert728 (
);

FILL FILL_1__11516_ (
);

FILL FILL_5_BUFX2_insert729 (
);

FILL FILL_0__10929_ (
);

FILL FILL_0__8523_ (
);

FILL FILL_0__10509_ (
);

FILL FILL_0__8103_ (
);

FILL FILL_5__6966_ (
);

FILL FILL_4__15742_ (
);

FILL FILL_4__15322_ (
);

FILL FILL_3__9092_ (
);

AOI21X1 _13686_ (
    .A(_4172_),
    .B(_4193_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [4])
);

AOI22X1 _13266_ (
    .A(_3763_),
    .B(_3804_),
    .C(_3775_),
    .D(_3750_),
    .Y(_3808_)
);

FILL FILL_2__9902_ (
);

FILL FILL_3__14735_ (
);

FILL FILL_3__14315_ (
);

FILL FILL_1__6958_ (
);

FILL FILL_4__9408_ (
);

FILL FILL_2__13728_ (
);

FILL FILL_2__13308_ (
);

FILL FILL_0__14762_ (
);

FILL SFILL99320x51050 (
);

FILL FILL_0__14342_ (
);

FILL FILL_0__9728_ (
);

FILL FILL_3__7825_ (
);

FILL SFILL28760x71050 (
);

FILL FILL_2_BUFX2_insert850 (
);

FILL FILL_2_BUFX2_insert851 (
);

FILL FILL_4__16107_ (
);

FILL FILL_2_BUFX2_insert852 (
);

FILL FILL_2_BUFX2_insert853 (
);

FILL FILL_2_BUFX2_insert854 (
);

FILL FILL_4__11662_ (
);

FILL FILL_2_BUFX2_insert855 (
);

FILL FILL_4__11242_ (
);

FILL SFILL64120x45050 (
);

FILL FILL_2_BUFX2_insert856 (
);

FILL FILL_2_BUFX2_insert857 (
);

FILL FILL_2_BUFX2_insert858 (
);

FILL FILL_2_BUFX2_insert859 (
);

FILL FILL_1__16134_ (
);

FILL FILL_3__10655_ (
);

FILL FILL_3__10235_ (
);

FILL FILL_0__15967_ (
);

FILL FILL_0__15547_ (
);

OAI22X1 _15832_ (
    .A(_5480__bF$buf2),
    .B(_6291_),
    .C(_6292_),
    .D(_5499__bF$buf3),
    .Y(_6293_)
);

NAND3X1 _15412_ (
    .A(_5877_),
    .B(_5883_),
    .C(_5871_),
    .Y(_5884_)
);

FILL FILL_0__15127_ (
);

FILL FILL_0__10682_ (
);

FILL FILL_0__10262_ (
);

FILL FILL_6__14881_ (
);

FILL FILL_5__13874_ (
);

FILL FILL_5__13454_ (
);

FILL FILL_5__13034_ (
);

INVX1 _7754_ (
    .A(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_448_)
);

INVX1 _7334_ (
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_229_)
);

FILL FILL_4__12867_ (
);

FILL FILL_4__9161_ (
);

FILL FILL_4__12447_ (
);

FILL FILL_4__12027_ (
);

FILL FILL_2__13481_ (
);

FILL FILL_1__12894_ (
);

FILL FILL_1__12474_ (
);

FILL FILL_1__12054_ (
);

FILL SFILL49560x74050 (
);

FILL FILL_0__11887_ (
);

FILL FILL_0__9481_ (
);

FILL FILL_2__9499_ (
);

FILL FILL_2__9079_ (
);

FILL FILL_0__11467_ (
);

OAI21X1 _11752_ (
    .A(_2846_),
    .B(_2847_),
    .C(_2845_),
    .Y(_2848_)
);

NOR2X1 _11332_ (
    .A(_2320_),
    .B(_2319_),
    .Y(_2451_)
);

FILL FILL_0__11047_ (
);

FILL FILL_5__7084_ (
);

FILL FILL_4__16280_ (
);

FILL SFILL54520x57050 (
);

FILL FILL_5__14659_ (
);

FILL FILL_5__14239_ (
);

FILL FILL_3__15693_ (
);

INVX1 _8959_ (
    .A(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_1048_)
);

FILL FILL_3__15273_ (
);

DFFSR _8539_ (
    .Q(\datapath_1.regfile_1.regOut[13] [5]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_783_[5])
);

OAI21X1 _8119_ (
    .A(_629_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .C(_630_),
    .Y(_588_[21])
);

FILL FILL_1__7496_ (
);

FILL FILL_1__7076_ (
);

FILL FILL_2__14686_ (
);

FILL FILL_2__14266_ (
);

FILL FILL_5__15600_ (
);

FILL SFILL89240x56050 (
);

INVX1 _9900_ (
    .A(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_1533_)
);

FILL SFILL54120x43050 (
);

FILL FILL_1__13679_ (
);

FILL FILL_1__13259_ (
);

FILL FILL_1_BUFX2_insert870 (
);

FILL FILL_3__8783_ (
);

FILL FILL_1_BUFX2_insert871 (
);

FILL FILL_1_BUFX2_insert872 (
);

FILL FILL_3__8363_ (
);

INVX1 _12957_ (
    .A(_2_[2]),
    .Y(_3623_)
);

DFFSR _12537_ (
    .Q(ALUOut[2]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3360_[2])
);

FILL FILL_1_BUFX2_insert873 (
);

FILL FILL_1_BUFX2_insert874 (
);

OAI21X1 _12117_ (
    .A(_3194_),
    .B(ALUSrcA_bF$buf1),
    .C(_3195_),
    .Y(\datapath_1.alu_1.ALUInA [0])
);

FILL FILL_1_BUFX2_insert875 (
);

FILL SFILL18680x76050 (
);

FILL FILL_1_BUFX2_insert876 (
);

FILL FILL_1__14620_ (
);

FILL FILL_1_BUFX2_insert877 (
);

FILL FILL_1__14200_ (
);

FILL FILL_1_BUFX2_insert878 (
);

FILL FILL_1_BUFX2_insert879 (
);

FILL FILL_0__13613_ (
);

FILL FILL_3__16058_ (
);

FILL FILL_5__10999_ (
);

FILL FILL_5__10579_ (
);

FILL FILL_5__10159_ (
);

FILL FILL_5__9650_ (
);

FILL FILL_5__9230_ (
);

FILL FILL_3__11193_ (
);

NAND2X1 _16370_ (
    .A(gnd),
    .B(gnd),
    .Y(_6801_)
);

FILL FILL_0__16085_ (
);

FILL FILL_2__10186_ (
);

FILL FILL_5__11940_ (
);

FILL FILL_1__9642_ (
);

FILL FILL_5__11520_ (
);

FILL FILL_1__9222_ (
);

FILL FILL_5__11100_ (
);

FILL SFILL89240x11050 (
);

FILL FILL_3__9988_ (
);

FILL FILL_2__16412_ (
);

FILL FILL_3__9148_ (
);

FILL FILL_4__10933_ (
);

FILL FILL_4__10513_ (
);

FILL FILL_1__15825_ (
);

FILL FILL_1__15405_ (
);

DFFSR _8292_ (
    .Q(\datapath_1.regfile_1.regOut[11] [14]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_653_[14])
);

FILL FILL_1__10960_ (
);

FILL FILL_1__10540_ (
);

FILL FILL_1__10120_ (
);

FILL FILL_0__14818_ (
);

FILL FILL_2__7985_ (
);

FILL FILL_2__7565_ (
);

BUFX2 BUFX2_insert540 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf67)
);

FILL FILL_3__12398_ (
);

BUFX2 BUFX2_insert541 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf66)
);

BUFX2 BUFX2_insert542 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf65)
);

BUFX2 BUFX2_insert543 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf64)
);

BUFX2 BUFX2_insert544 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf63)
);

BUFX2 BUFX2_insert545 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf62)
);

BUFX2 BUFX2_insert546 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf61)
);

BUFX2 BUFX2_insert547 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf60)
);

BUFX2 BUFX2_insert548 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf59)
);

BUFX2 BUFX2_insert549 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf58)
);

NAND3X1 _12290_ (
    .A(_3254_),
    .B(_3255_),
    .C(_3256_),
    .Y(\datapath_1.alu_1.ALUInB [18])
);

FILL FILL_5__12725_ (
);

FILL FILL_5__12305_ (
);

FILL SFILL79240x54050 (
);

FILL FILL_4__8852_ (
);

FILL FILL_4__8012_ (
);

FILL FILL_4__11718_ (
);

FILL FILL_2__12752_ (
);

FILL FILL_5__15197_ (
);

FILL FILL_2__12332_ (
);

OAI21X1 _9497_ (
    .A(_1324_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1325_),
    .Y(_1303_[11])
);

DFFSR _9077_ (
    .Q(\datapath_1.regfile_1.regOut[17] [31]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_1043_[31])
);

FILL FILL_1__11745_ (
);

FILL FILL_1__11325_ (
);

FILL FILL_0__8752_ (
);

FILL FILL_0__8332_ (
);

DFFSR _10603_ (
    .Q(\datapath_1.regfile_1.regOut[29] [21]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1823_[21])
);

FILL FILL_0__10318_ (
);

FILL FILL_0_BUFX2_insert60 (
);

FILL FILL_0_BUFX2_insert61 (
);

FILL FILL_4__15971_ (
);

FILL FILL_0_BUFX2_insert62 (
);

FILL SFILL44040x48050 (
);

FILL FILL_4__15551_ (
);

FILL FILL_0_BUFX2_insert63 (
);

FILL FILL_0_BUFX2_insert64 (
);

FILL FILL_4__15131_ (
);

FILL FILL_0_BUFX2_insert65 (
);

FILL FILL_0_BUFX2_insert66 (
);

FILL FILL_0_BUFX2_insert67 (
);

AOI22X1 _13495_ (
    .A(_3942__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[3] [1]),
    .C(\datapath_1.regfile_1.regOut[12] [1]),
    .D(_4005__bF$buf1),
    .Y(_4006_)
);

DFFSR _13075_ (
    .Q(_2_[28]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_3620_[28])
);

FILL FILL_0_BUFX2_insert68 (
);

FILL FILL_0_BUFX2_insert69 (
);

FILL FILL_3__14964_ (
);

FILL FILL_3__14544_ (
);

FILL FILL_3__14124_ (
);

FILL FILL_4_BUFX2_insert380 (
);

FILL FILL_4__9637_ (
);

FILL FILL_4_BUFX2_insert381 (
);

FILL FILL_4__9217_ (
);

FILL FILL_4_BUFX2_insert382 (
);

FILL FILL_4_BUFX2_insert383 (
);

FILL FILL_2__13957_ (
);

FILL FILL_0__14991_ (
);

FILL FILL_4_BUFX2_insert384 (
);

FILL FILL_2__13537_ (
);

FILL FILL_0__14571_ (
);

FILL FILL_4_BUFX2_insert385 (
);

FILL FILL_2__13117_ (
);

FILL FILL_0__14151_ (
);

FILL FILL_4_BUFX2_insert386 (
);

FILL FILL_4_BUFX2_insert387 (
);

FILL FILL_4_BUFX2_insert388 (
);

FILL FILL_4_BUFX2_insert389 (
);

FILL FILL111880x22050 (
);

FILL FILL_3__7634_ (
);

FILL FILL_0__9537_ (
);

FILL FILL_3__7214_ (
);

NAND3X1 _11808_ (
    .A(_2897_),
    .B(_2899_),
    .C(_2894_),
    .Y(\datapath_1.ALUResult [4])
);

FILL FILL_0__9117_ (
);

FILL SFILL8520x18050 (
);

FILL FILL_4__16336_ (
);

FILL FILL_4__11891_ (
);

FILL FILL_4__11471_ (
);

FILL FILL_4__11051_ (
);

FILL FILL_3__15749_ (
);

FILL FILL_3__15329_ (
);

FILL FILL_1__16363_ (
);

FILL FILL_3__10884_ (
);

FILL FILL_5__8501_ (
);

FILL FILL_3__10044_ (
);

FILL FILL_0__15776_ (
);

FILL SFILL69240x52050 (
);

FILL FILL_0__15356_ (
);

NAND2X1 _15641_ (
    .A(_6100_),
    .B(_6106_),
    .Y(_6107_)
);

NOR3X1 _15221_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5493_),
    .C(_5696_),
    .Y(_5697_)
);

FILL FILL_0__10491_ (
);

FILL FILL_1__8913_ (
);

FILL FILL_3__8839_ (
);

FILL FILL_5__13683_ (
);

FILL FILL_5__13263_ (
);

INVX1 _7983_ (
    .A(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_560_)
);

INVX1 _7563_ (
    .A(\datapath_1.regfile_1.regOut[6] [7]),
    .Y(_341_)
);

DFFSR _7143_ (
    .Q(\datapath_1.regfile_1.regOut[2] [17]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_68_[17])
);

FILL FILL_4__9390_ (
);

FILL FILL_4__12256_ (
);

FILL FILL_2__13290_ (
);

FILL FILL_2__6836_ (
);

FILL FILL_3__11669_ (
);

FILL FILL_3__11249_ (
);

FILL FILL_1__12283_ (
);

DFFSR _16426_ (
    .Q(\datapath_1.regfile_1.regOut[0] [9]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_6769_[9])
);

AOI21X1 _16006_ (
    .A(_6441_),
    .B(_6462_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [23])
);

NAND2X1 _11981_ (
    .A(IorD_bF$buf6),
    .B(ALUOut[31]),
    .Y(_3029_)
);

FILL FILL_0__9290_ (
);

FILL FILL_0__11696_ (
);

NAND2X1 _11561_ (
    .A(_2669_),
    .B(_2430_),
    .Y(_2670_)
);

FILL FILL_0__11276_ (
);

NAND2X1 _11141_ (
    .A(_2238_),
    .B(_2259_),
    .Y(_2260_)
);

FILL FILL_3__12610_ (
);

FILL FILL_6__15475_ (
);

FILL FILL_6__15055_ (
);

FILL FILL_4__7703_ (
);

FILL FILL_5__14888_ (
);

FILL FILL_5__14468_ (
);

FILL FILL_2__11603_ (
);

FILL FILL_5__14048_ (
);

OAI21X1 _8768_ (
    .A(_960_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_961_),
    .Y(_913_[24])
);

FILL FILL_3__15082_ (
);

OAI21X1 _8348_ (
    .A(_741_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_742_),
    .Y(_718_[12])
);

FILL FILL_2__14495_ (
);

FILL FILL_2__14075_ (
);

FILL SFILL69160x14050 (
);

FILL FILL_0__7603_ (
);

FILL FILL_1__13488_ (
);

FILL FILL_4__14822_ (
);

FILL FILL_4__14402_ (
);

FILL FILL_3__8592_ (
);

OAI21X1 _12766_ (
    .A(_3535_),
    .B(IRWrite_bF$buf7),
    .C(_3536_),
    .Y(_3490_[23])
);

INVX1 _12346_ (
    .A(ALUOut[1]),
    .Y(_3296_)
);

FILL FILL_3__13815_ (
);

FILL FILL_5__8098_ (
);

FILL FILL_4__8908_ (
);

FILL FILL_6__11395_ (
);

FILL SFILL99320x46050 (
);

FILL FILL_0__13842_ (
);

FILL FILL_0__13422_ (
);

FILL FILL_3__16287_ (
);

FILL FILL_0__13002_ (
);

FILL FILL_5__10388_ (
);

FILL SFILL89400x82050 (
);

FILL SFILL28760x66050 (
);

FILL FILL_3__6905_ (
);

FILL FILL_1__9871_ (
);

FILL FILL_1__9031_ (
);

FILL FILL_4__15607_ (
);

FILL FILL_2__16221_ (
);

FILL FILL_3__9797_ (
);

FILL FILL_3__9377_ (
);

FILL FILL_4__10742_ (
);

FILL FILL_4__10322_ (
);

FILL FILL_1__15634_ (
);

FILL FILL_1__15214_ (
);

FILL FILL_0__14627_ (
);

OAI22X1 _14912_ (
    .A(_5392_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf0),
    .D(_5393_),
    .Y(_5394_)
);

FILL FILL_0__14207_ (
);

FILL FILL_2__7374_ (
);

FILL FILL_6__13961_ (
);

FILL FILL_6__13541_ (
);

FILL FILL_5__12954_ (
);

FILL FILL_5__12534_ (
);

FILL FILL_5__12114_ (
);

FILL SFILL28760x21050 (
);

FILL SFILL59160x12050 (
);

FILL FILL_4__8661_ (
);

FILL FILL_4__11947_ (
);

FILL FILL_4__8241_ (
);

FILL FILL_2__12981_ (
);

FILL FILL_4__11527_ (
);

FILL FILL_4__11107_ (
);

FILL FILL_2__12141_ (
);

FILL FILL_1__11974_ (
);

FILL FILL_1__11554_ (
);

FILL FILL_1__11134_ (
);

FILL FILL_2__8999_ (
);

FILL FILL_0__8981_ (
);

FILL FILL_0__10967_ (
);

FILL FILL_2__8579_ (
);

FILL FILL_0__8141_ (
);

INVX1 _10832_ (
    .A(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_2012_)
);

FILL FILL_0__10547_ (
);

FILL SFILL89320x44050 (
);

FILL FILL_0__10127_ (
);

INVX1 _10412_ (
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_1793_)
);

FILL FILL_4__15780_ (
);

FILL FILL_4__15360_ (
);

FILL FILL_2__9940_ (
);

FILL FILL_5__13739_ (
);

FILL FILL_5__13319_ (
);

FILL FILL_3__14773_ (
);

FILL FILL_2__9520_ (
);

FILL FILL_2__9100_ (
);

FILL FILL_3__14353_ (
);

FILL SFILL18760x64050 (
);

OAI21X1 _7619_ (
    .A(_377_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_378_),
    .Y(_328_[25])
);

FILL FILL_1__6996_ (
);

FILL FILL_4__9866_ (
);

FILL FILL_4__9026_ (
);

FILL FILL_2__13766_ (
);

FILL FILL_2__13346_ (
);

FILL FILL_0__14380_ (
);

FILL FILL_1__12759_ (
);

FILL FILL_1__12339_ (
);

FILL FILL_3__7863_ (
);

FILL FILL_0__9766_ (
);

FILL FILL_0__9346_ (
);

FILL FILL_3__7443_ (
);

OAI21X1 _11617_ (
    .A(_2254_),
    .B(_2255_),
    .C(_2721_),
    .Y(_2722_)
);

FILL FILL_5__7369_ (
);

FILL FILL_1__13700_ (
);

FILL FILL_4__16145_ (
);

INVX1 _14089_ (
    .A(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_4588_)
);

FILL FILL_4__11280_ (
);

FILL FILL_3__15978_ (
);

FILL FILL_3__15558_ (
);

FILL FILL_3__15138_ (
);

FILL FILL_1__16172_ (
);

FILL FILL_3__10693_ (
);

FILL FILL_5__8730_ (
);

FILL FILL_3__10273_ (
);

FILL FILL_5__8310_ (
);

OAI22X1 _15870_ (
    .A(_4931_),
    .B(_5544__bF$buf1),
    .C(_5499__bF$buf3),
    .D(_4932_),
    .Y(_6330_)
);

FILL FILL_0__15585_ (
);

INVX1 _15450_ (
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_5921_)
);

FILL FILL_0__15165_ (
);

NAND2X1 _15030_ (
    .A(\datapath_1.PCJump [24]),
    .B(_5460_),
    .Y(_5510_)
);

FILL FILL_1__8722_ (
);

FILL FILL_2__15912_ (
);

FILL FILL_3__8648_ (
);

FILL FILL_3__8228_ (
);

FILL FILL_5__13492_ (
);

FILL SFILL23960x82050 (
);

DFFSR _7792_ (
    .Q(\datapath_1.regfile_1.regOut[7] [26]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_393_[26])
);

FILL FILL_1__14905_ (
);

OAI21X1 _7372_ (
    .A(_253_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .C(_254_),
    .Y(_198_[28])
);

FILL SFILL79320x42050 (
);

FILL FILL_4__12485_ (
);

FILL FILL_4__12065_ (
);

FILL FILL_5__9935_ (
);

FILL FILL_3__11898_ (
);

FILL FILL_5__9515_ (
);

FILL FILL_3__11478_ (
);

FILL FILL_3__11058_ (
);

FILL FILL_1__12092_ (
);

OAI22X1 _16235_ (
    .A(_5480__bF$buf3),
    .B(_6685_),
    .C(_5326_),
    .D(_5499__bF$buf2),
    .Y(_6686_)
);

NOR3X1 _11790_ (
    .A(_2337_),
    .B(_2880_),
    .C(_2882_),
    .Y(_2883_)
);

OAI21X1 _11370_ (
    .A(_2354_),
    .B(_2355_),
    .C(_2121_),
    .Y(_2487_)
);

FILL FILL_0__11085_ (
);

FILL FILL_1__9927_ (
);

FILL FILL_5__11805_ (
);

FILL FILL_1__9507_ (
);

FILL FILL_4__7932_ (
);

FILL FILL_5__14697_ (
);

FILL FILL_2__11832_ (
);

FILL FILL_5__14277_ (
);

FILL FILL_2__11412_ (
);

OAI21X1 _8997_ (
    .A(_1072_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .C(_1073_),
    .Y(_1043_[15])
);

OAI21X1 _8577_ (
    .A(_853_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_854_),
    .Y(_848_[3])
);

DFFSR _8157_ (
    .Q(\datapath_1.regfile_1.regOut[10] [7]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_588_[7])
);

FILL FILL_1__10825_ (
);

FILL FILL_1__10405_ (
);

FILL FILL_0__7832_ (
);

FILL FILL_1__13297_ (
);

FILL FILL_4__14631_ (
);

FILL SFILL94360x9050 (
);

FILL FILL_4__14211_ (
);

FILL FILL111960x10050 (
);

OAI21X1 _12995_ (
    .A(_3647_),
    .B(vdd),
    .C(_3648_),
    .Y(_3620_[14])
);

OAI21X1 _12575_ (
    .A(_3428_),
    .B(vdd),
    .C(_3429_),
    .Y(_3425_[2])
);

NAND2X1 _12155_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [13]),
    .Y(_3157_)
);

FILL FILL_3__13624_ (
);

FILL FILL_4__8717_ (
);

FILL FILL_2__12617_ (
);

FILL FILL_0__13651_ (
);

FILL FILL_0__13231_ (
);

FILL FILL_3__16096_ (
);

FILL FILL_5__10197_ (
);

FILL SFILL13960x80050 (
);

FILL SFILL29560x65050 (
);

FILL FILL_2__15089_ (
);

FILL FILL_0__8617_ (
);

FILL FILL_5__16003_ (
);

FILL FILL_1__9680_ (
);

FILL FILL_1__9260_ (
);

FILL FILL_4__15836_ (
);

FILL FILL_4__15416_ (
);

FILL FILL_2__16450_ (
);

FILL FILL_2__16030_ (
);

FILL FILL_4__10971_ (
);

FILL FILL_4__10551_ (
);

FILL FILL_4__10131_ (
);

FILL FILL_3__14829_ (
);

FILL FILL_3__14409_ (
);

FILL FILL_1__15863_ (
);

FILL FILL_1__15443_ (
);

FILL FILL_1__15023_ (
);

FILL SFILL69240x47050 (
);

FILL FILL_0__14856_ (
);

OAI22X1 _14721_ (
    .A(_3983__bF$buf1),
    .B(_5205_),
    .C(_3971__bF$buf0),
    .D(_5206_),
    .Y(_5207_)
);

FILL FILL_0__14436_ (
);

FILL FILL_0__14016_ (
);

OAI22X1 _14301_ (
    .A(_4795_),
    .B(_3936__bF$buf3),
    .C(_3967__bF$buf2),
    .D(_4794_),
    .Y(_4796_)
);

BUFX2 BUFX2_insert920 (
    .A(_5549_),
    .Y(_5549__bF$buf0)
);

FILL FILL_2__7183_ (
);

BUFX2 BUFX2_insert921 (
    .A(_3882_),
    .Y(_3882__bF$buf3)
);

BUFX2 BUFX2_insert922 (
    .A(_3882_),
    .Y(_3882__bF$buf2)
);

BUFX2 BUFX2_insert923 (
    .A(_3882_),
    .Y(_3882__bF$buf1)
);

BUFX2 BUFX2_insert924 (
    .A(_3882_),
    .Y(_3882__bF$buf0)
);

BUFX2 BUFX2_insert925 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf4 )
);

BUFX2 BUFX2_insert926 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf3 )
);

BUFX2 BUFX2_insert927 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf2 )
);

BUFX2 BUFX2_insert928 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf1 )
);

BUFX2 BUFX2_insert929 (
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf0 )
);

FILL FILL_5__12763_ (
);

FILL FILL_5__12343_ (
);

FILL FILL_4__8890_ (
);

FILL FILL_4__8470_ (
);

FILL FILL_4__11756_ (
);

FILL FILL_2__12790_ (
);

FILL FILL_4__11336_ (
);

FILL FILL_2__12370_ (
);

FILL FILL_1__16228_ (
);

FILL FILL_3__10749_ (
);

FILL FILL_1__11783_ (
);

FILL FILL_1__11363_ (
);

NOR2X1 _15926_ (
    .A(_6383_),
    .B(_6384_),
    .Y(_6385_)
);

OAI22X1 _15506_ (
    .A(_5974_),
    .B(_5469__bF$buf0),
    .C(_5472__bF$buf3),
    .D(_4509_),
    .Y(_5975_)
);

FILL FILL_0__10776_ (
);

FILL FILL_2__8388_ (
);

FILL FILL_0__8370_ (
);

FILL SFILL104360x72050 (
);

INVX1 _10641_ (
    .A(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_1905_)
);

DFFSR _10221_ (
    .Q(\datapath_1.regfile_1.regOut[26] [23]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1628_[23])
);

FILL FILL_5__13968_ (
);

FILL FILL_5__13548_ (
);

FILL FILL_3__14582_ (
);

FILL FILL_5__13128_ (
);

OAI21X1 _7848_ (
    .A(_489_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .C(_490_),
    .Y(_458_[16])
);

FILL FILL_3__14162_ (
);

OAI21X1 _7428_ (
    .A(_270_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_271_),
    .Y(_263_[4])
);

FILL FILL_4_BUFX2_insert760 (
);

DFFSR _7008_ (
    .Q(\datapath_1.regfile_1.regOut[1] [10]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_3_[10])
);

FILL FILL_4__9675_ (
);

FILL FILL_4_BUFX2_insert761 (
);

FILL FILL_4__9255_ (
);

FILL FILL_4_BUFX2_insert762 (
);

FILL FILL_4_BUFX2_insert763 (
);

FILL FILL_2__13995_ (
);

FILL FILL_4_BUFX2_insert764 (
);

FILL FILL_2__13575_ (
);

FILL FILL_4_BUFX2_insert765 (
);

FILL FILL_2__13155_ (
);

FILL SFILL99400x34050 (
);

FILL FILL_4_BUFX2_insert766 (
);

FILL FILL_4_BUFX2_insert767 (
);

FILL FILL_4_BUFX2_insert768 (
);

FILL FILL_4_BUFX2_insert769 (
);

FILL FILL_1__12988_ (
);

FILL FILL_1__12568_ (
);

FILL FILL_1__12148_ (
);

FILL FILL_4__13902_ (
);

FILL FILL_0__9995_ (
);

FILL FILL_3__7672_ (
);

FILL FILL_3__7252_ (
);

OAI21X1 _11846_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .C(_2620_),
    .Y(_2934_)
);

FILL FILL_0__9155_ (
);

AND2X2 _11426_ (
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2542_)
);

AOI21X1 _11006_ (
    .A(_2121_),
    .B(_2124_),
    .C(_2119_),
    .Y(_2125_)
);

FILL FILL_5__7598_ (
);

FILL FILL_5__7178_ (
);

FILL FILL_4__16374_ (
);

FILL FILL_3__15787_ (
);

FILL FILL_3__15367_ (
);

FILL FILL_0__12502_ (
);

FILL FILL_0__15394_ (
);

FILL SFILL64040x2050 (
);

FILL FILL_1__8951_ (
);

FILL FILL_1__8531_ (
);

FILL SFILL3720x9050 (
);

FILL FILL_1__8111_ (
);

FILL FILL_2__15721_ (
);

FILL FILL_2__15301_ (
);

FILL FILL_3__8877_ (
);

FILL FILL_3__8457_ (
);

FILL FILL_1__14714_ (
);

OAI21X1 _7181_ (
    .A(_146_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_147_),
    .Y(_133_[7])
);

FILL FILL_4__12294_ (
);

FILL FILL_0__13707_ (
);

FILL FILL_2__6874_ (
);

FILL FILL_5__9744_ (
);

FILL FILL_3__11287_ (
);

FILL FILL_0__16179_ (
);

FILL SFILL114440x3050 (
);

NAND2X1 _16044_ (
    .A(_6495_),
    .B(_6499_),
    .Y(_6500_)
);

FILL SFILL89400x32050 (
);

FILL FILL_1__9736_ (
);

FILL FILL_5__11614_ (
);

FILL FILL_4__7741_ (
);

FILL FILL_3_BUFX2_insert780 (
);

FILL FILL_4__7321_ (
);

FILL FILL_3_BUFX2_insert781 (
);

FILL FILL_3_BUFX2_insert782 (
);

FILL FILL_3_BUFX2_insert783 (
);

FILL FILL_2__11641_ (
);

FILL FILL_2__11221_ (
);

FILL FILL_3_BUFX2_insert784 (
);

FILL FILL_5__14086_ (
);

FILL FILL_1__15919_ (
);

FILL FILL_3_BUFX2_insert785 (
);

FILL FILL_3_BUFX2_insert786 (
);

NAND2X1 _8386_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_768_)
);

FILL FILL_3_BUFX2_insert787 (
);

FILL FILL_3_BUFX2_insert788 (
);

FILL FILL_3_BUFX2_insert789 (
);

FILL FILL_1__10634_ (
);

FILL FILL_4__13499_ (
);

FILL FILL_4__13079_ (
);

FILL SFILL33960x79050 (
);

FILL FILL_0__7221_ (
);

FILL FILL_2__7239_ (
);

FILL FILL_4__14860_ (
);

FILL FILL_4__14440_ (
);

FILL FILL_4__14020_ (
);

FILL FILL_0__12099_ (
);

OAI21X1 _12384_ (
    .A(_3320_),
    .B(MemToReg_bF$buf4),
    .C(_3321_),
    .Y(\datapath_1.mux_wd3.dout [13])
);

FILL FILL_3__13853_ (
);

FILL FILL_2__8600_ (
);

FILL SFILL18760x59050 (
);

FILL FILL_3__13433_ (
);

FILL FILL_6__16298_ (
);

FILL FILL_3__13013_ (
);

FILL FILL_4__8526_ (
);

FILL SFILL8600x50 (
);

FILL FILL_4__8106_ (
);

FILL FILL_2__12846_ (
);

FILL FILL_0__13880_ (
);

FILL FILL_2__12426_ (
);

FILL FILL_0__13460_ (
);

FILL FILL_2__12006_ (
);

FILL FILL_0__13040_ (
);

FILL FILL_1__11839_ (
);

FILL FILL_1__11419_ (
);

FILL FILL_0__8846_ (
);

FILL FILL_5__16232_ (
);

FILL FILL_3__6943_ (
);

FILL FILL_6__9813_ (
);

FILL FILL_0__8006_ (
);

FILL SFILL33960x34050 (
);

FILL FILL_5__6869_ (
);

FILL FILL_4__15645_ (
);

FILL FILL_4__15225_ (
);

INVX1 _13589_ (
    .A(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_4098_)
);

FILL FILL_4__10780_ (
);

FILL FILL_4__10360_ (
);

INVX1 _13169_ (
    .A(\datapath_1.PCJump [30]),
    .Y(_3744_)
);

FILL FILL_2__9805_ (
);

FILL FILL_4_BUFX2_insert10 (
);

FILL FILL_4_BUFX2_insert11 (
);

FILL FILL_3__14638_ (
);

FILL FILL_3__14218_ (
);

FILL FILL_1__15672_ (
);

FILL FILL_4_BUFX2_insert12 (
);

FILL FILL_1__15252_ (
);

FILL FILL_4_BUFX2_insert13 (
);

FILL FILL_4_BUFX2_insert14 (
);

FILL FILL_5__7810_ (
);

FILL FILL_4_BUFX2_insert15 (
);

FILL FILL_4_BUFX2_insert16 (
);

FILL SFILL18760x14050 (
);

FILL FILL_4_BUFX2_insert17 (
);

FILL SFILL84280x81050 (
);

FILL FILL_4_BUFX2_insert18 (
);

NOR2X1 _14950_ (
    .A(_5427_),
    .B(_5430_),
    .Y(_5431_)
);

FILL FILL_4_BUFX2_insert19 (
);

FILL FILL_0__14665_ (
);

FILL FILL_0__14245_ (
);

INVX1 _14530_ (
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_5020_)
);

INVX1 _14110_ (
    .A(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_4609_)
);

FILL FILL_1__7802_ (
);

FILL FILL_3__7728_ (
);

FILL FILL_3__7308_ (
);

FILL FILL_5__12992_ (
);

FILL FILL_5__12572_ (
);

FILL FILL_5__12152_ (
);

BUFX2 _6872_ (
    .A(_2_[2]),
    .Y(memoryWriteData[2])
);

FILL SFILL79320x37050 (
);

FILL SFILL59000x8050 (
);

FILL FILL_4__11985_ (
);

FILL FILL_4__11565_ (
);

FILL FILL_4__11145_ (
);

FILL FILL_1__16037_ (
);

FILL FILL_3__10978_ (
);

FILL FILL_3__10558_ (
);

FILL FILL_6_BUFX2_insert290 (
);

FILL FILL_3__10138_ (
);

FILL FILL_1__11592_ (
);

FILL FILL_1__11172_ (
);

FILL SFILL39640x10050 (
);

NAND2X1 _15735_ (
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .B(_5562_),
    .Y(_6198_)
);

FILL FILL_6_BUFX2_insert295 (
);

NOR2X1 _15315_ (
    .A(_5788_),
    .B(_5549__bF$buf2),
    .Y(_5789_)
);

INVX1 _10870_ (
    .A(\aluControl_1.inst [4]),
    .Y(_2018_)
);

FILL FILL_2__8197_ (
);

FILL FILL_0__10165_ (
);

OAI21X1 _10450_ (
    .A(_1817_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1818_),
    .Y(_1758_[30])
);

FILL SFILL33320x3050 (
);

OAI21X1 _10030_ (
    .A(_1598_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .C(_1599_),
    .Y(_1563_[18])
);

BUFX2 BUFX2_insert70 (
    .A(_3905_),
    .Y(_3905__bF$buf1)
);

FILL FILL_6__14784_ (
);

BUFX2 BUFX2_insert71 (
    .A(_3905_),
    .Y(_3905__bF$buf0)
);

BUFX2 BUFX2_insert72 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf4 )
);

BUFX2 BUFX2_insert73 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf3 )
);

BUFX2 BUFX2_insert74 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf2 )
);

BUFX2 BUFX2_insert75 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf1 )
);

BUFX2 BUFX2_insert76 (
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf0 )
);

FILL FILL_2__10912_ (
);

FILL FILL_5__13777_ (
);

BUFX2 BUFX2_insert77 (
    .A(_5495_),
    .Y(_5495__bF$buf3)
);

FILL FILL_5__13357_ (
);

BUFX2 BUFX2_insert78 (
    .A(_5495_),
    .Y(_5495__bF$buf2)
);

BUFX2 BUFX2_insert79 (
    .A(_5495_),
    .Y(_5495__bF$buf1)
);

FILL FILL_3__14391_ (
);

DFFSR _7657_ (
    .Q(\datapath_1.regfile_1.regOut[6] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_328_[19])
);

NAND2X1 _7237_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_185_)
);

FILL FILL_4__9484_ (
);

FILL FILL_2__13384_ (
);

FILL SFILL114440x62050 (
);

FILL FILL_0__6912_ (
);

FILL FILL_1__12377_ (
);

FILL FILL_4__13711_ (
);

FILL FILL_0__9384_ (
);

FILL FILL_3__7481_ (
);

FILL FILL_3__7061_ (
);

AOI21X1 _11655_ (
    .A(_2753_),
    .B(_2757_),
    .C(_2754_),
    .Y(_2758_)
);

AND2X2 _11235_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2354_)
);

FILL FILL_3__12704_ (
);

FILL FILL_4__16183_ (
);

FILL FILL_6__10284_ (
);

FILL FILL_0__12731_ (
);

FILL FILL_3__15596_ (
);

FILL FILL_3__15176_ (
);

FILL FILL_0__12311_ (
);

FILL FILL_2__14589_ (
);

FILL FILL_2__14169_ (
);

FILL FILL_5__15923_ (
);

FILL FILL_5__15503_ (
);

NAND2X1 _9803_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1489_)
);

FILL FILL_1__8760_ (
);

FILL FILL_1__8340_ (
);

FILL FILL_4__14916_ (
);

FILL FILL_2__15950_ (
);

FILL FILL_2__15530_ (
);

FILL FILL_2__15110_ (
);

FILL FILL_3__8266_ (
);

FILL FILL_3__13909_ (
);

FILL FILL_1__14943_ (
);

FILL FILL_1__14523_ (
);

FILL FILL_1__14103_ (
);

FILL FILL_0__13936_ (
);

INVX1 _13801_ (
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_4306_)
);

FILL FILL_0__13516_ (
);

FILL FILL_5__9553_ (
);

FILL FILL_5__9133_ (
);

FILL FILL_3__11096_ (
);

NOR2X1 _16273_ (
    .A(_6722_),
    .B(_6721_),
    .Y(_6723_)
);

FILL FILL_5__11843_ (
);

FILL FILL_1__9545_ (
);

FILL FILL_5__11423_ (
);

FILL FILL_1__9125_ (
);

FILL FILL_5__11003_ (
);

FILL FILL_4__7970_ (
);

FILL FILL_2__16315_ (
);

FILL FILL_4__7550_ (
);

FILL FILL_4__10836_ (
);

FILL FILL_2__11870_ (
);

FILL FILL_4__10416_ (
);

FILL FILL_2__11450_ (
);

FILL FILL_2__11030_ (
);

FILL FILL_1__15728_ (
);

NAND2X1 _8195_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_661_)
);

FILL FILL_1__15308_ (
);

FILL FILL_1__10443_ (
);

FILL FILL_1__10023_ (
);

FILL FILL_0__7870_ (
);

FILL FILL_2__7888_ (
);

FILL SFILL104360x67050 (
);

FILL FILL_0__7450_ (
);

FILL FILL_2__7468_ (
);

FILL FILL_2__7048_ (
);

FILL FILL_0__7030_ (
);

FILL SFILL43880x6050 (
);

INVX1 _12193_ (
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3182_)
);

FILL FILL_5__12628_ (
);

FILL FILL_3__13662_ (
);

FILL FILL_5__12208_ (
);

FILL FILL_3__13242_ (
);

OAI21X1 _6928_ (
    .A(_18_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_19_),
    .Y(_3_[8])
);

FILL FILL_4__8755_ (
);

FILL SFILL8600x6050 (
);

FILL FILL_4__8335_ (
);

FILL FILL_2__12655_ (
);

FILL SFILL99400x29050 (
);

FILL FILL_2__12235_ (
);

FILL FILL_1__11648_ (
);

FILL FILL_1__11228_ (
);

FILL FILL_0__8655_ (
);

FILL FILL_5__16041_ (
);

FILL FILL112440x73050 (
);

NOR2X1 _10926_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2047_),
    .Y(ALUOp[0])
);

FILL FILL_0__8235_ (
);

FILL FILL_6__9622_ (
);

OAI21X1 _10506_ (
    .A(_1834_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1835_),
    .Y(_1823_[6])
);

FILL FILL_4__15874_ (
);

FILL SFILL104360x22050 (
);

FILL FILL_4__15454_ (
);

FILL FILL_4__15034_ (
);

NAND2X1 _13398_ (
    .A(_3880_),
    .B(_3889_),
    .Y(_3910_)
);

FILL FILL_2__9614_ (
);

FILL FILL_3__14867_ (
);

FILL FILL_3__14447_ (
);

FILL FILL_3__14027_ (
);

FILL FILL_1__15481_ (
);

FILL FILL_1__15061_ (
);

FILL SFILL108680x30050 (
);

FILL FILL_0__14894_ (
);

FILL FILL_0__14474_ (
);

FILL FILL_0__14054_ (
);

FILL FILL_1__7611_ (
);

FILL FILL_2__14801_ (
);

FILL FILL_3__7957_ (
);

FILL FILL_3__7117_ (
);

FILL FILL_5__12381_ (
);

FILL FILL_4__16239_ (
);

FILL FILL_4__11794_ (
);

FILL FILL_4__11374_ (
);

FILL FILL_1__16266_ (
);

FILL FILL_3__10787_ (
);

FILL FILL_5__8824_ (
);

FILL FILL_3__10367_ (
);

FILL FILL_5__8404_ (
);

FILL FILL_0__15679_ (
);

OAI22X1 _15964_ (
    .A(_5549__bF$buf3),
    .B(_6421_),
    .C(_5466__bF$buf2),
    .D(_6420_),
    .Y(_6422_)
);

FILL FILL_0__15259_ (
);

OAI22X1 _15544_ (
    .A(_5489__bF$buf3),
    .B(_6011_),
    .C(_5527__bF$buf4),
    .D(_4553_),
    .Y(_6012_)
);

NOR2X1 _15124_ (
    .A(_5600_),
    .B(_5602_),
    .Y(_5603_)
);

FILL FILL_0__10394_ (
);

FILL SFILL89400x27050 (
);

FILL FILL_0__16200_ (
);

FILL FILL_5__13586_ (
);

FILL FILL_2__10301_ (
);

FILL FILL_5__13166_ (
);

NAND2X1 _7886_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_516_)
);

NAND2X1 _7466_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_297_)
);

NAND2X1 _7046_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_78_)
);

FILL FILL_4__9293_ (
);

FILL FILL_4__12999_ (
);

FILL FILL_4__12579_ (
);

FILL FILL_4__12159_ (
);

FILL FILL_5__9609_ (
);

FILL FILL_1__12186_ (
);

FILL FILL_4__13940_ (
);

FILL FILL_4__13520_ (
);

OAI21X1 _16329_ (
    .A(_6772_),
    .B(gnd),
    .C(_6773_),
    .Y(_6769_[2])
);

FILL FILL_4__13100_ (
);

INVX1 _11884_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_2966_)
);

FILL FILL_3__7290_ (
);

FILL FILL_0__11599_ (
);

FILL FILL_0__11179_ (
);

AOI21X1 _11464_ (
    .A(_2309_),
    .B(_2578_),
    .C(_2288_),
    .Y(_2579_)
);

NOR2X1 _11044_ (
    .A(_2161_),
    .B(_2162_),
    .Y(_2163_)
);

FILL FILL_6__15378_ (
);

FILL FILL_3__12513_ (
);

FILL FILL_4__7606_ (
);

FILL SFILL94280x33050 (
);

FILL FILL_2__11926_ (
);

FILL FILL_0__12960_ (
);

FILL FILL_2__11506_ (
);

FILL FILL_0__12120_ (
);

FILL FILL_1__10919_ (
);

FILL FILL_2__14398_ (
);

FILL FILL_5__15732_ (
);

FILL FILL_5__15312_ (
);

FILL FILL_0__7926_ (
);

FILL SFILL79800x39050 (
);

FILL FILL_0__7506_ (
);

NAND2X1 _9612_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1382_)
);

FILL SFILL33960x29050 (
);

FILL FILL_4__14725_ (
);

FILL FILL_4__14305_ (
);

FILL FILL_3__8495_ (
);

DFFSR _12669_ (
    .Q(\datapath_1.Data [6]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3425_[6])
);

FILL FILL_3__8075_ (
);

AOI22X1 _12249_ (
    .A(_2_[8]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [8]),
    .Y(_3226_)
);

FILL FILL_3__13718_ (
);

FILL FILL_1__14752_ (
);

FILL FILL_1__14332_ (
);

FILL FILL_6__11298_ (
);

FILL SFILL84280x76050 (
);

FILL FILL_0__13745_ (
);

FILL FILL_0__13325_ (
);

NAND3X1 _13610_ (
    .A(_4114_),
    .B(_4118_),
    .C(_4111_),
    .Y(_4119_)
);

FILL FILL_5__9782_ (
);

FILL FILL_5__9362_ (
);

FILL SFILL23640x51050 (
);

OAI22X1 _16082_ (
    .A(_6536_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf0),
    .D(_5169_),
    .Y(_6537_)
);

FILL FILL_5__11652_ (
);

FILL FILL_1__9774_ (
);

FILL FILL_1__9354_ (
);

FILL FILL_5__11232_ (
);

FILL FILL_2__16124_ (
);

FILL FILL_4__10645_ (
);

FILL FILL_1__15957_ (
);

FILL FILL_1__15537_ (
);

FILL FILL_1__15117_ (
);

FILL FILL_1__10672_ (
);

FILL FILL_1__10252_ (
);

OAI22X1 _14815_ (
    .A(_5298_),
    .B(_3902__bF$buf1),
    .C(_3954__bF$buf4),
    .D(_5297_),
    .Y(_5299_)
);

FILL SFILL84280x31050 (
);

FILL FILL_2__7697_ (
);

FILL FILL_6__13444_ (
);

FILL SFILL109480x74050 (
);

FILL SFILL23160x44050 (
);

FILL FILL_5__12857_ (
);

FILL FILL_5__12437_ (
);

FILL FILL_3__13891_ (
);

FILL FILL_5__12017_ (
);

FILL FILL_3__13471_ (
);

FILL FILL_4__8984_ (
);

FILL FILL_4__8144_ (
);

FILL FILL_2__12884_ (
);

FILL SFILL114440x57050 (
);

FILL FILL_2__12464_ (
);

FILL FILL_2__12044_ (
);

FILL FILL_1__11877_ (
);

FILL FILL_1__11457_ (
);

FILL FILL_1__11037_ (
);

FILL FILL_3__6981_ (
);

FILL FILL_5__16270_ (
);

FILL FILL_0__8884_ (
);

FILL FILL_0__8464_ (
);

DFFSR _10735_ (
    .Q(\datapath_1.regfile_1.regOut[30] [25]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_1888_[25])
);

NAND2X1 _10315_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1749_)
);

FILL FILL_4__15683_ (
);

FILL FILL_4__15263_ (
);

FILL FILL_2__9423_ (
);

FILL FILL_0__11811_ (
);

FILL FILL_3__14676_ (
);

FILL FILL_3__14256_ (
);

FILL FILL_2__9003_ (
);

FILL FILL_1__15290_ (
);

FILL FILL_1__6899_ (
);

FILL FILL_4__9769_ (
);

FILL FILL_4__9349_ (
);

FILL FILL_2__13669_ (
);

FILL FILL_2__13249_ (
);

FILL FILL_0__14283_ (
);

FILL SFILL114440x12050 (
);

FILL FILL_1__7840_ (
);

FILL FILL_1__7420_ (
);

FILL FILL_2__14610_ (
);

FILL SFILL74200x72050 (
);

FILL FILL_0__9669_ (
);

FILL FILL_0__9249_ (
);

FILL FILL_3__7346_ (
);

FILL FILL_5__12190_ (
);

FILL FILL_1__13603_ (
);

FILL FILL_4__16048_ (
);

FILL FILL_1_BUFX2_insert110 (
);

FILL FILL_4__11183_ (
);

FILL FILL_1__16075_ (
);

FILL FILL_5__8633_ (
);

FILL FILL_3__10176_ (
);

FILL FILL_5__8213_ (
);

FILL SFILL59800x35050 (
);

FILL FILL_6_BUFX2_insert674 (
);

INVX1 _15773_ (
    .A(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_6235_)
);

FILL FILL_0__15488_ (
);

NOR2X1 _15353_ (
    .A(_5825_),
    .B(_5824_),
    .Y(_5826_)
);

FILL FILL_0__15068_ (
);

FILL FILL_3__16402_ (
);

FILL FILL_6_BUFX2_insert679 (
);

FILL FILL_5__10923_ (
);

FILL FILL_1__8625_ (
);

FILL FILL_5__10503_ (
);

FILL FILL_1__8205_ (
);

FILL FILL_2__15815_ (
);

FILL FILL_2__10950_ (
);

FILL FILL_2__10530_ (
);

FILL FILL_5__13395_ (
);

FILL FILL_2__10110_ (
);

NAND2X1 _7695_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_409_)
);

FILL FILL_1__14808_ (
);

DFFSR _7275_ (
    .Q(\datapath_1.regfile_1.regOut[3] [21]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_133_[21])
);

FILL FILL_4__12388_ (
);

FILL FILL_3__9912_ (
);

FILL FILL_0__6950_ (
);

FILL FILL_2__6968_ (
);

FILL FILL_5__9418_ (
);

NOR2X1 _16138_ (
    .A(_6590_),
    .B(_6587_),
    .Y(_6591_)
);

NAND2X1 _11693_ (
    .A(_2185_),
    .B(_2480_),
    .Y(_2793_)
);

NOR2X1 _11273_ (
    .A(_2391_),
    .B(_2202_),
    .Y(_2392_)
);

FILL FILL_5__11708_ (
);

FILL FILL_3__12742_ (
);

FILL FILL_3__12322_ (
);

FILL SFILL104440x10050 (
);

FILL FILL_4__7835_ (
);

FILL FILL_4__7415_ (
);

FILL FILL_2__11735_ (
);

FILL FILL_2__11315_ (
);

FILL SFILL64200x70050 (
);

FILL FILL_1__10308_ (
);

FILL FILL_5__15961_ (
);

FILL FILL_5__15541_ (
);

FILL FILL112440x68050 (
);

FILL FILL_0__7735_ (
);

FILL FILL_5__15121_ (
);

DFFSR _9841_ (
    .Q(\datapath_1.regfile_1.regOut[23] [27]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1433_[27])
);

FILL FILL_0__7315_ (
);

FILL FILL_6__8702_ (
);

INVX1 _9421_ (
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_1295_)
);

INVX1 _9001_ (
    .A(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_1076_)
);

FILL FILL_4__14954_ (
);

FILL FILL_4__14534_ (
);

FILL FILL_4__14114_ (
);

INVX1 _12898_ (
    .A(\datapath_1.a [25]),
    .Y(_3604_)
);

INVX1 _12478_ (
    .A(ALUOut[13]),
    .Y(_3385_)
);

NAND3X1 _12058_ (
    .A(_3087_),
    .B(_3088_),
    .C(_3089_),
    .Y(\datapath_1.mux_pcsrc.dout [17])
);

FILL FILL_3__13947_ (
);

FILL FILL_3__13527_ (
);

FILL FILL_1__14981_ (
);

FILL FILL_1__14561_ (
);

FILL FILL_3__13107_ (
);

FILL FILL_1__14141_ (
);

FILL FILL112040x54050 (
);

FILL FILL_5_BUFX2_insert690 (
);

FILL FILL_5_BUFX2_insert691 (
);

FILL FILL_5_BUFX2_insert692 (
);

FILL FILL_0__13974_ (
);

FILL FILL_5_BUFX2_insert693 (
);

FILL FILL_0__13554_ (
);

FILL FILL_5_BUFX2_insert694 (
);

FILL FILL_0__13134_ (
);

FILL FILL_5_BUFX2_insert695 (
);

FILL FILL_5_BUFX2_insert696 (
);

FILL FILL_5__9591_ (
);

FILL FILL_5_BUFX2_insert697 (
);

FILL FILL_5__9171_ (
);

FILL FILL_5_BUFX2_insert698 (
);

FILL FILL_5_BUFX2_insert699 (
);

FILL FILL_5__16326_ (
);

FILL FILL_5__11881_ (
);

FILL FILL_5__11461_ (
);

FILL FILL_1__9163_ (
);

FILL FILL_5__11041_ (
);

FILL FILL112440x23050 (
);

FILL FILL_4__15739_ (
);

FILL FILL_4__15319_ (
);

FILL FILL_2__16353_ (
);

FILL FILL_3__9089_ (
);

FILL FILL_4__10874_ (
);

FILL FILL_4__10034_ (
);

FILL SFILL48840x50 (
);

FILL FILL_1__15766_ (
);

FILL FILL_6__7094_ (
);

FILL FILL_1__15346_ (
);

FILL FILL_1__10061_ (
);

FILL FILL_0__14759_ (
);

OAI22X1 _14624_ (
    .A(_5111_),
    .B(_3971__bF$buf4),
    .C(_3924__bF$buf3),
    .D(_5110_),
    .Y(_5112_)
);

FILL FILL_0__14339_ (
);

NOR2X1 _14204_ (
    .A(_4697_),
    .B(_4700_),
    .Y(_4701_)
);

FILL FILL_2__7086_ (
);

FILL FILL_0__15700_ (
);

FILL FILL_5__12246_ (
);

FILL FILL_3__13280_ (
);

NAND2X1 _6966_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_45_)
);

FILL FILL_4__8373_ (
);

FILL FILL_4__11659_ (
);

FILL FILL_4__11239_ (
);

FILL FILL_2__12273_ (
);

FILL FILL_1__11686_ (
);

FILL FILL_1__11266_ (
);

OAI21X1 _15829_ (
    .A(_5524__bF$buf1),
    .B(_4865_),
    .C(_6289_),
    .Y(_6290_)
);

FILL FILL_4__12600_ (
);

INVX1 _15409_ (
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_5881_)
);

FILL FILL_0__10679_ (
);

NAND3X1 _10964_ (
    .A(_2091_),
    .B(_2095_),
    .C(_2094_),
    .Y(\control_1.next [2])
);

FILL FILL_0__8273_ (
);

FILL FILL_6__9240_ (
);

NAND2X1 _10544_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1861_)
);

FILL FILL_0__10259_ (
);

NAND2X1 _10124_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1642_)
);

FILL FILL_4__15492_ (
);

FILL FILL_4__15072_ (
);

FILL SFILL94280x28050 (
);

FILL FILL_2__9652_ (
);

FILL FILL_2__9232_ (
);

FILL FILL_3__14485_ (
);

FILL FILL_0__11620_ (
);

FILL FILL_3__14065_ (
);

FILL FILL_0__11200_ (
);

FILL FILL_4__9998_ (
);

FILL FILL_4__9158_ (
);

FILL FILL_2__13898_ (
);

FILL FILL_2__13478_ (
);

FILL FILL_0__14092_ (
);

FILL FILL_5__14812_ (
);

FILL FILL_4__13805_ (
);

FILL FILL_3__7995_ (
);

FILL FILL_0__9898_ (
);

FILL FILL_3__7575_ (
);

FILL FILL_0__9478_ (
);

AOI21X1 _11749_ (
    .A(_2841_),
    .B(_2844_),
    .C(_2843_),
    .Y(_2845_)
);

OAI21X1 _11329_ (
    .A(_2292_),
    .B(_2286_),
    .C(_2290_),
    .Y(_2448_)
);

FILL FILL_1__13832_ (
);

FILL FILL_1__13412_ (
);

FILL FILL_4__16277_ (
);

FILL FILL_6__10378_ (
);

FILL FILL_0__12825_ (
);

FILL FILL_0__12405_ (
);

FILL FILL_5__8862_ (
);

FILL FILL_5__8442_ (
);

FILL SFILL23640x46050 (
);

FILL FILL_0__15297_ (
);

AOI21X1 _15582_ (
    .A(\datapath_1.regfile_1.regOut[7] [13]),
    .B(_5490_),
    .C(_6048_),
    .Y(_6049_)
);

OAI22X1 _15162_ (
    .A(_5495__bF$buf0),
    .B(_5639_),
    .C(_4085_),
    .D(_5534__bF$buf3),
    .Y(_5640_)
);

FILL FILL_3__16211_ (
);

FILL FILL_1__8854_ (
);

FILL FILL_5__10312_ (
);

FILL FILL_1__8014_ (
);

FILL SFILL13720x82050 (
);

FILL FILL_2__15624_ (
);

FILL FILL_2__15204_ (
);

FILL SFILL23240x32050 (
);

FILL FILL_1__14617_ (
);

INVX1 _7084_ (
    .A(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_103_)
);

FILL SFILL84200x69050 (
);

FILL FILL_4__12197_ (
);

FILL FILL_3__9721_ (
);

FILL FILL_3__9301_ (
);

FILL SFILL84280x26050 (
);

FILL FILL_5__9647_ (
);

FILL FILL_5__9227_ (
);

NAND2X1 _16367_ (
    .A(gnd),
    .B(gnd),
    .Y(_6799_)
);

FILL SFILL109480x69050 (
);

FILL FILL_5__11937_ (
);

NOR2X1 _11082_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2190_),
    .Y(_2201_)
);

FILL FILL_1__9639_ (
);

FILL FILL_3__12971_ (
);

FILL FILL_5__11517_ (
);

FILL FILL_1__9219_ (
);

FILL SFILL8600x43050 (
);

FILL FILL_3__12131_ (
);

FILL FILL_2__16409_ (
);

FILL FILL_4__7224_ (
);

FILL FILL_2__11964_ (
);

FILL FILL_2__11544_ (
);

FILL FILL_3_CLKBUF1_insert220 (
);

FILL FILL_2__11124_ (
);

FILL FILL_3_CLKBUF1_insert221 (
);

DFFSR _8289_ (
    .Q(\datapath_1.regfile_1.regOut[11] [11]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_653_[11])
);

FILL FILL_3_CLKBUF1_insert222 (
);

FILL FILL_3_CLKBUF1_insert223 (
);

FILL FILL_3_CLKBUF1_insert224 (
);

FILL FILL_1__10957_ (
);

FILL FILL_1__10537_ (
);

FILL FILL_1__10117_ (
);

FILL SFILL84200x24050 (
);

FILL FILL_5__15770_ (
);

FILL SFILL74280x69050 (
);

FILL FILL_5__15350_ (
);

FILL FILL_0__7964_ (
);

FILL FILL_0__7544_ (
);

FILL FILL_0__7124_ (
);

INVX1 _9650_ (
    .A(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_1407_)
);

FILL SFILL114040x38050 (
);

INVX1 _9230_ (
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_1188_)
);

FILL FILL_4__14763_ (
);

FILL FILL_4__14343_ (
);

FILL SFILL13640x44050 (
);

NAND3X1 _12287_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3254_)
);

FILL FILL_2__8503_ (
);

FILL FILL_3__13756_ (
);

FILL FILL_3__13336_ (
);

FILL FILL_1__14790_ (
);

FILL FILL_1__14370_ (
);

FILL FILL_4__8849_ (
);

FILL FILL_4__8009_ (
);

FILL FILL_2__12749_ (
);

FILL FILL_0__13783_ (
);

FILL FILL_2__12329_ (
);

FILL FILL_0__13363_ (
);

FILL FILL_1__6920_ (
);

FILL SFILL74200x67050 (
);

FILL FILL_3__6846_ (
);

FILL FILL_0__8749_ (
);

FILL FILL_5__16135_ (
);

FILL FILL_0__8329_ (
);

FILL FILL_5__11690_ (
);

FILL FILL_1__9392_ (
);

FILL FILL_5__11270_ (
);

FILL SFILL74280x24050 (
);

FILL FILL_4__15968_ (
);

FILL FILL_4__15548_ (
);

FILL FILL_4__15128_ (
);

FILL FILL_2__16162_ (
);

FILL FILL_4__10683_ (
);

FILL FILL_4__10263_ (
);

FILL FILL_1__15995_ (
);

FILL FILL112200x80050 (
);

FILL FILL_1__15575_ (
);

FILL SFILL99480x73050 (
);

FILL FILL_1__15155_ (
);

FILL FILL_5__7713_ (
);

FILL FILL_1__10290_ (
);

FILL FILL_0__14988_ (
);

FILL FILL_0__14568_ (
);

OAI22X1 _14853_ (
    .A(_5335_),
    .B(_3936__bF$buf2),
    .C(_3955__bF$buf3),
    .D(_5334_),
    .Y(_5336_)
);

FILL FILL_0__14148_ (
);

OAI22X1 _14433_ (
    .A(_4924_),
    .B(_3902__bF$buf3),
    .C(_3954__bF$buf4),
    .D(_4923_),
    .Y(_4925_)
);

INVX1 _14013_ (
    .A(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_4514_)
);

FILL FILL_3__15902_ (
);

FILL FILL_1__7705_ (
);

FILL FILL_5__12895_ (
);

FILL SFILL43800x31050 (
);

FILL FILL_5__12475_ (
);

FILL SFILL74200x22050 (
);

FILL FILL_5__12055_ (
);

FILL FILL_4__11888_ (
);

FILL FILL_4__8182_ (
);

FILL FILL_4__11468_ (
);

FILL FILL_4__11048_ (
);

FILL FILL_2__12082_ (
);

FILL FILL_1__11495_ (
);

FILL FILL_1__11075_ (
);

INVX1 _15638_ (
    .A(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_6104_)
);

AOI22X1 _15218_ (
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .B(_5693_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_5694_)
);

FILL FILL_0__10488_ (
);

NAND2X1 _10773_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1973_)
);

FILL FILL_0__8082_ (
);

FILL FILL_0__10068_ (
);

DFFSR _10353_ (
    .Q(\datapath_1.regfile_1.regOut[27] [27]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_1693_[27])
);

FILL FILL_3__11822_ (
);

FILL FILL_6__14687_ (
);

FILL FILL_6__14267_ (
);

FILL FILL_3__11402_ (
);

FILL FILL_4__6915_ (
);

FILL FILL_2__10815_ (
);

FILL FILL_2__9881_ (
);

FILL SFILL33800x74050 (
);

FILL SFILL64200x65050 (
);

FILL FILL_2__9041_ (
);

FILL FILL_3__14294_ (
);

FILL FILL112120x42050 (
);

FILL FILL_4__9387_ (
);

FILL FILL_2__13287_ (
);

FILL FILL_5__14621_ (
);

FILL FILL_5__14201_ (
);

DFFSR _8921_ (
    .Q(\datapath_1.regfile_1.regOut[16] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_978_[3])
);

INVX1 _8501_ (
    .A(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_824_)
);

FILL FILL_4__13614_ (
);

NAND2X1 _11978_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[30]),
    .Y(_3027_)
);

FILL FILL_0__9287_ (
);

INVX1 _11558_ (
    .A(_2666_),
    .Y(_2667_)
);

NAND2X1 _11138_ (
    .A(_2253_),
    .B(_2256_),
    .Y(_2257_)
);

FILL SFILL89720x8050 (
);

FILL FILL_3__12607_ (
);

FILL FILL_1__13641_ (
);

FILL FILL112040x49050 (
);

FILL FILL_1__13221_ (
);

FILL FILL_4__16086_ (
);

FILL FILL_0__12634_ (
);

FILL FILL_3__15499_ (
);

FILL FILL_0__12214_ (
);

FILL FILL_3__15079_ (
);

FILL SFILL89400x2050 (
);

FILL FILL_5__8251_ (
);

FILL SFILL64200x20050 (
);

INVX1 _15391_ (
    .A(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_5863_)
);

FILL FILL_5__15826_ (
);

FILL FILL_5__15406_ (
);

FILL FILL_3__16020_ (
);

DFFSR _9706_ (
    .Q(\datapath_1.regfile_1.regOut[22] [20]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1368_[20])
);

FILL FILL_5__10961_ (
);

FILL FILL_5__10541_ (
);

FILL FILL112440x18050 (
);

FILL FILL_5__10121_ (
);

FILL FILL_1__8243_ (
);

FILL FILL_4__14819_ (
);

FILL FILL_2__15853_ (
);

FILL FILL_2__15433_ (
);

FILL FILL_3__8589_ (
);

FILL FILL_2__15013_ (
);

FILL FILL_1__14846_ (
);

FILL FILL_1__14426_ (
);

FILL FILL_1__14006_ (
);

FILL FILL_0__13839_ (
);

FILL FILL_3__9530_ (
);

FILL FILL_0__13419_ (
);

OAI22X1 _13704_ (
    .A(_3884__bF$buf3),
    .B(_4209_),
    .C(_3955__bF$buf2),
    .D(_4210_),
    .Y(_4211_)
);

FILL FILL_3__9110_ (
);

FILL FILL_5__9876_ (
);

FILL FILL_5__9036_ (
);

FILL FILL_6__12753_ (
);

AOI22X1 _16176_ (
    .A(_5567_),
    .B(\datapath_1.regfile_1.regOut[28] [28]),
    .C(\datapath_1.regfile_1.regOut[31] [28]),
    .D(_5571_),
    .Y(_6628_)
);

FILL FILL_1__9868_ (
);

FILL FILL_5__11746_ (
);

FILL FILL_3__12780_ (
);

FILL FILL_5__11326_ (
);

FILL FILL_1__9028_ (
);

FILL FILL_3__12360_ (
);

FILL FILL_2__16218_ (
);

FILL FILL_4__7873_ (
);

FILL FILL_4__7453_ (
);

FILL FILL_4__7033_ (
);

FILL FILL_4__10319_ (
);

FILL FILL_2__11773_ (
);

FILL FILL_2__11353_ (
);

OAI21X1 _8098_ (
    .A(_615_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_616_),
    .Y(_588_[14])
);

FILL SFILL23720x79050 (
);

FILL FILL_1__10766_ (
);

FILL FILL_2_CLKBUF1_insert210 (
);

FILL FILL_2_CLKBUF1_insert211 (
);

AOI22X1 _14909_ (
    .A(\datapath_1.regfile_1.regOut[4] [30]),
    .B(_3891__bF$buf1),
    .C(_3998__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_5391_)
);

FILL FILL_2_CLKBUF1_insert212 (
);

FILL FILL_2_CLKBUF1_insert213 (
);

FILL FILL_2_CLKBUF1_insert214 (
);

FILL FILL_2_CLKBUF1_insert215 (
);

FILL FILL_0__7353_ (
);

FILL FILL_2_CLKBUF1_insert216 (
);

FILL FILL_6__8320_ (
);

FILL FILL_2_CLKBUF1_insert217 (
);

FILL FILL_2_CLKBUF1_insert218 (
);

FILL FILL_4__14992_ (
);

FILL FILL_2_CLKBUF1_insert219 (
);

FILL FILL_4__14572_ (
);

FILL FILL_4__14152_ (
);

NAND3X1 _12096_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_27_bF$buf3 ),
    .C(_3034__bF$buf1),
    .Y(_3118_)
);

FILL FILL_3__13985_ (
);

FILL FILL_2__8732_ (
);

FILL FILL_0__10700_ (
);

FILL FILL_2__8312_ (
);

FILL FILL_3__13565_ (
);

FILL FILL_3__13145_ (
);

FILL FILL_4__8658_ (
);

FILL FILL_4__8238_ (
);

FILL FILL_2__12978_ (
);

FILL FILL_0__13592_ (
);

FILL FILL_2__12138_ (
);

FILL FILL_0__13172_ (
);

FILL FILL_5__16364_ (
);

FILL FILL_0__8978_ (
);

INVX1 _10829_ (
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_2010_)
);

FILL FILL_0__8138_ (
);

INVX1 _10409_ (
    .A(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_1791_)
);

FILL FILL_6__9105_ (
);

FILL FILL_1__12912_ (
);

FILL FILL_4__15777_ (
);

FILL FILL_4__15357_ (
);

FILL SFILL48920x83050 (
);

FILL FILL_2__16391_ (
);

FILL FILL_4__10492_ (
);

FILL FILL_2__9937_ (
);

FILL FILL_0__11905_ (
);

FILL FILL_2__9517_ (
);

FILL FILL_1__15384_ (
);

FILL FILL_5__7942_ (
);

FILL FILL_5__7102_ (
);

FILL FILL_0__14797_ (
);

FILL FILL_0__14377_ (
);

OAI22X1 _14662_ (
    .A(_5148_),
    .B(_3931__bF$buf1),
    .C(_3966__bF$buf1),
    .D(_5147_),
    .Y(_5149_)
);

NAND2X1 _14242_ (
    .A(_4730_),
    .B(_4737_),
    .Y(_4738_)
);

FILL FILL_3__15711_ (
);

FILL FILL_1__7934_ (
);

FILL SFILL13720x77050 (
);

FILL FILL_2__14704_ (
);

FILL SFILL109560x57050 (
);

FILL FILL_5__12284_ (
);

FILL FILL_4__11697_ (
);

FILL FILL_4__11277_ (
);

FILL SFILL99480x9050 (
);

FILL FILL_1__16169_ (
);

FILL FILL_5__8727_ (
);

NOR3X1 _15867_ (
    .A(_5515__bF$buf0),
    .B(_4910_),
    .C(_5521__bF$buf2),
    .Y(_6327_)
);

FILL FILL_6__11604_ (
);

INVX1 _15447_ (
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_5918_)
);

NAND3X1 _15027_ (
    .A(_5491_),
    .B(_5497_),
    .C(_5506_),
    .Y(_5507_)
);

DFFSR _10582_ (
    .Q(\datapath_1.regfile_1.regOut[29] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_1823_[0])
);

FILL FILL_0__10297_ (
);

INVX1 _10162_ (
    .A(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_1667_)
);

FILL FILL_1__8719_ (
);

FILL SFILL8600x38050 (
);

FILL FILL_3__11631_ (
);

FILL FILL_3__11211_ (
);

FILL FILL_2__15909_ (
);

FILL FILL_0__16103_ (
);

FILL SFILL13720x32050 (
);

FILL SFILL29320x17050 (
);

FILL FILL_2__10624_ (
);

FILL FILL_5__13489_ (
);

FILL FILL_2__9270_ (
);

DFFSR _7789_ (
    .Q(\datapath_1.regfile_1.regOut[7] [23]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_393_[23])
);

OAI21X1 _7369_ (
    .A(_251_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .C(_252_),
    .Y(_198_[27])
);

FILL FILL_2__13096_ (
);

FILL SFILL38920x81050 (
);

FILL SFILL84200x19050 (
);

FILL FILL_5__14850_ (
);

FILL FILL_5_BUFX2_insert80 (
);

FILL FILL_5__14430_ (
);

FILL FILL_5__14010_ (
);

FILL FILL_5_BUFX2_insert81 (
);

INVX1 _8730_ (
    .A(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_936_)
);

FILL FILL_5_BUFX2_insert82 (
);

FILL FILL_5_BUFX2_insert83 (
);

INVX1 _8310_ (
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_781_)
);

FILL FILL_5_BUFX2_insert84 (
);

FILL FILL_1__12089_ (
);

FILL FILL_5_BUFX2_insert85 (
);

FILL FILL_4__13843_ (
);

FILL FILL_5_BUFX2_insert86 (
);

FILL FILL_5_BUFX2_insert87 (
);

FILL FILL_4__13423_ (
);

FILL FILL_5_BUFX2_insert88 (
);

FILL FILL_4__13003_ (
);

FILL FILL_5_BUFX2_insert89 (
);

FILL SFILL13640x39050 (
);

FILL FILL_0__9096_ (
);

FILL FILL_3__7193_ (
);

AOI21X1 _11787_ (
    .A(_2878_),
    .B(_2879_),
    .C(_2367_),
    .Y(_2880_)
);

AOI21X1 _11367_ (
    .A(_2451_),
    .B(_2478_),
    .C(_2483_),
    .Y(_2484_)
);

FILL FILL_3__12836_ (
);

FILL SFILL109480x19050 (
);

FILL FILL_3__12416_ (
);

FILL FILL_1__13870_ (
);

FILL FILL_1__13450_ (
);

FILL FILL_1__13030_ (
);

FILL FILL_4__7929_ (
);

FILL FILL_4__7509_ (
);

FILL FILL_2__11829_ (
);

FILL FILL_0__12863_ (
);

FILL FILL_2__11409_ (
);

FILL FILL_0__12443_ (
);

FILL FILL_0__12023_ (
);

FILL FILL_6__16222_ (
);

FILL FILL_5__8480_ (
);

FILL FILL_5__8060_ (
);

FILL SFILL3560x80050 (
);

FILL FILL_5__15635_ (
);

FILL FILL_5__15215_ (
);

FILL FILL_0__7829_ (
);

OAI21X1 _9935_ (
    .A(_1555_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1556_),
    .Y(_1498_[29])
);

OAI21X1 _9515_ (
    .A(_1336_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .C(_1337_),
    .Y(_1303_[17])
);

FILL FILL_1__8892_ (
);

FILL FILL_5__10770_ (
);

FILL SFILL74280x19050 (
);

FILL FILL_1__8472_ (
);

FILL FILL_4__14628_ (
);

FILL FILL_2__15662_ (
);

FILL FILL_4__14208_ (
);

FILL FILL_2__15242_ (
);

FILL FILL_3__8398_ (
);

FILL FILL112200x75050 (
);

FILL SFILL99480x68050 (
);

FILL FILL_1__14655_ (
);

FILL FILL_1__14235_ (
);

FILL FILL_0__13648_ (
);

NOR2X1 _13933_ (
    .A(_4434_),
    .B(_3944__bF$buf1),
    .Y(_4435_)
);

FILL FILL_0__13228_ (
);

INVX1 _13513_ (
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_4024_)
);

FILL FILL_5__9685_ (
);

FILL FILL_5__9265_ (
);

FILL FILL_6__12142_ (
);

FILL SFILL43800x26050 (
);

FILL FILL_5__11975_ (
);

FILL SFILL74200x17050 (
);

FILL FILL_1__9677_ (
);

FILL FILL_5__11555_ (
);

FILL FILL_1__9257_ (
);

FILL FILL_5__11135_ (
);

BUFX2 BUFX2_insert1070 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf3 )
);

BUFX2 BUFX2_insert1071 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf2 )
);

BUFX2 BUFX2_insert1072 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf1 )
);

FILL FILL_2__16027_ (
);

FILL FILL_4__7682_ (
);

FILL FILL_4__10968_ (
);

BUFX2 BUFX2_insert1073 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf0 )
);

FILL FILL_4__10548_ (
);

FILL FILL_4__10128_ (
);

FILL FILL_2__11582_ (
);

FILL FILL_2__11162_ (
);

FILL FILL_6__7188_ (
);

FILL FILL_1__10995_ (
);

FILL FILL112200x30050 (
);

FILL FILL_1__10575_ (
);

FILL SFILL99480x23050 (
);

FILL FILL_1__10155_ (
);

OAI22X1 _14718_ (
    .A(_5203_),
    .B(_3954__bF$buf0),
    .C(_3924__bF$buf2),
    .D(_5202_),
    .Y(_5204_)
);

BUFX2 BUFX2_insert890 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf4 )
);

FILL FILL_0__7582_ (
);

BUFX2 BUFX2_insert891 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf3 )
);

FILL FILL_0__7162_ (
);

BUFX2 BUFX2_insert892 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf2 )
);

BUFX2 BUFX2_insert893 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf1 )
);

FILL FILL_1_CLKBUF1_insert200 (
);

BUFX2 BUFX2_insert894 (
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf0 )
);

FILL FILL_3__10902_ (
);

FILL FILL_1_CLKBUF1_insert201 (
);

FILL FILL_6__13347_ (
);

BUFX2 BUFX2_insert895 (
    .A(_3982_),
    .Y(_3982__bF$buf3)
);

FILL FILL_1_CLKBUF1_insert202 (
);

FILL FILL_1_CLKBUF1_insert203 (
);

BUFX2 BUFX2_insert896 (
    .A(_3982_),
    .Y(_3982__bF$buf2)
);

FILL FILL_4__14381_ (
);

BUFX2 BUFX2_insert897 (
    .A(_3982_),
    .Y(_3982__bF$buf1)
);

FILL FILL_1_CLKBUF1_insert204 (
);

FILL FILL_1_CLKBUF1_insert205 (
);

BUFX2 BUFX2_insert898 (
    .A(_3982_),
    .Y(_3982__bF$buf0)
);

FILL FILL_1_CLKBUF1_insert206 (
);

BUFX2 BUFX2_insert899 (
    .A(_5552_),
    .Y(_5552__bF$buf3)
);

FILL FILL_1_CLKBUF1_insert207 (
);

FILL SFILL33800x69050 (
);

FILL FILL_1_CLKBUF1_insert208 (
);

FILL FILL_2__8961_ (
);

FILL FILL_3__13794_ (
);

FILL FILL_1_CLKBUF1_insert209 (
);

FILL FILL_2__8121_ (
);

FILL FILL_3__13374_ (
);

FILL FILL112120x37050 (
);

FILL FILL_4__8887_ (
);

FILL FILL_4__8467_ (
);

FILL FILL_2__12787_ (
);

FILL FILL_2__12367_ (
);

FILL FILL_5__13701_ (
);

FILL FILL_5__16173_ (
);

FILL FILL_3__6884_ (
);

FILL FILL_0__8787_ (
);

FILL FILL_0__8367_ (
);

INVX1 _10638_ (
    .A(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_1903_)
);

DFFSR _10218_ (
    .Q(\datapath_1.regfile_1.regOut[26] [20]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1628_[20])
);

FILL FILL_1__12721_ (
);

FILL FILL_4__15586_ (
);

FILL SFILL28840x41050 (
);

FILL FILL_1__12301_ (
);

FILL FILL_4__15166_ (
);

FILL FILL_3__14999_ (
);

FILL FILL_2__9746_ (
);

FILL FILL_3__14579_ (
);

FILL FILL_0__11714_ (
);

FILL FILL_3__14159_ (
);

FILL FILL_1__15193_ (
);

FILL SFILL33800x24050 (
);

FILL FILL_5__7751_ (
);

FILL SFILL64200x15050 (
);

FILL FILL_5__7331_ (
);

NAND3X1 _14891_ (
    .A(_5371_),
    .B(_5372_),
    .C(_5370_),
    .Y(_5373_)
);

AOI22X1 _14471_ (
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .B(_3894_),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_4962_)
);

FILL FILL_0__14186_ (
);

OAI22X1 _14051_ (
    .A(_4550_),
    .B(_3954__bF$buf4),
    .C(_3924__bF$buf1),
    .D(_4549_),
    .Y(_4551_)
);

FILL FILL_5__14906_ (
);

FILL FILL_3__15940_ (
);

FILL FILL_3__15520_ (
);

FILL FILL_3__15100_ (
);

FILL FILL_1__7743_ (
);

FILL FILL_1__7323_ (
);

FILL FILL_2__14933_ (
);

FILL FILL_2__14513_ (
);

FILL FILL_3__7249_ (
);

FILL FILL_5__12093_ (
);

FILL FILL_1__13926_ (
);

FILL FILL_1__13506_ (
);

FILL FILL_4__11086_ (
);

FILL FILL_3__8610_ (
);

FILL FILL_1__16398_ (
);

FILL FILL_5__8956_ (
);

FILL FILL_3__10499_ (
);

FILL FILL_5__8116_ (
);

INVX1 _15676_ (
    .A(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_6141_)
);

NOR2X1 _15256_ (
    .A(_5729_),
    .B(_5731_),
    .Y(_5732_)
);

FILL FILL_3__16305_ (
);

INVX1 _10391_ (
    .A(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_1779_)
);

FILL FILL_5__10826_ (
);

FILL FILL_5__10406_ (
);

FILL FILL_3__11860_ (
);

FILL FILL_1__8528_ (
);

FILL FILL_3__11440_ (
);

FILL FILL_1__8108_ (
);

FILL FILL_3__11020_ (
);

FILL FILL_2__15718_ (
);

FILL FILL_4__6953_ (
);

FILL FILL_0__16332_ (
);

FILL SFILL44040x50 (
);

FILL FILL_5__13298_ (
);

FILL FILL_2__10433_ (
);

FILL FILL_2__10013_ (
);

OAI21X1 _7598_ (
    .A(_363_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_364_),
    .Y(_328_[18])
);

OAI21X1 _7178_ (
    .A(_144_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .C(_145_),
    .Y(_133_[6])
);

FILL FILL_0__6853_ (
);

FILL FILL_4__13652_ (
);

FILL FILL_4__13232_ (
);

OAI21X1 _11596_ (
    .A(_2547_),
    .B(_2548_),
    .C(_2420_),
    .Y(_2703_)
);

NOR2X1 _11176_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2295_)
);

FILL FILL_2__7812_ (
);

FILL FILL_3__12645_ (
);

FILL FILL_3__12225_ (
);

FILL FILL_4__7738_ (
);

FILL FILL_4__7318_ (
);

FILL FILL_2__11638_ (
);

FILL FILL_2__11218_ (
);

FILL FILL_0__12252_ (
);

FILL SFILL74120x8050 (
);

FILL FILL_5__15864_ (
);

FILL FILL_5__15444_ (
);

FILL SFILL38840x4050 (
);

FILL FILL_5__15024_ (
);

OAI21X1 _9744_ (
    .A(_1448_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .C(_1449_),
    .Y(_1433_[8])
);

FILL FILL_0__7218_ (
);

DFFSR _9324_ (
    .Q(\datapath_1.regfile_1.regOut[19] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1173_[22])
);

FILL FILL_4__14857_ (
);

FILL SFILL48920x78050 (
);

FILL FILL_4__14437_ (
);

FILL FILL_2__15891_ (
);

FILL FILL_4__14017_ (
);

FILL FILL_2__15471_ (
);

FILL SFILL44200x56050 (
);

FILL FILL_2__15051_ (
);

FILL FILL_1__14884_ (
);

FILL FILL_1__14464_ (
);

FILL FILL_1__14044_ (
);

FILL FILL_0__13877_ (
);

AOI22X1 _13742_ (
    .A(_4154_),
    .B(\datapath_1.regfile_1.regOut[14] [6]),
    .C(\datapath_1.regfile_1.regOut[31] [6]),
    .D(_3995__bF$buf4),
    .Y(_4248_)
);

FILL FILL_0__13457_ (
);

INVX1 _13322_ (
    .A(_3851_),
    .Y(_3852_)
);

FILL FILL_0__13037_ (
);

FILL FILL_5__9494_ (
);

FILL SFILL109240x31050 (
);

FILL FILL_5__16229_ (
);

FILL FILL_5__11784_ (
);

FILL FILL_1__9486_ (
);

FILL FILL_5__11364_ (
);

FILL FILL_2__16256_ (
);

FILL FILL_4__7491_ (
);

FILL FILL_4__10777_ (
);

FILL FILL_4__7071_ (
);

FILL FILL_2__11391_ (
);

FILL FILL_1__15669_ (
);

FILL FILL_1__15249_ (
);

FILL SFILL109160x38050 (
);

FILL FILL_5__7807_ (
);

FILL FILL_1__10384_ (
);

INVX1 _14947_ (
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_5428_)
);

NOR2X1 _14527_ (
    .A(_5002_),
    .B(_5016_),
    .Y(_5017_)
);

INVX1 _14107_ (
    .A(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_4606_)
);

FILL FILL_6__13996_ (
);

FILL FILL_6__13156_ (
);

FILL FILL_4__14190_ (
);

FILL FILL_0__15603_ (
);

FILL FILL_5__12989_ (
);

FILL FILL_5__12569_ (
);

FILL FILL_2__8770_ (
);

FILL FILL_5__12149_ (
);

FILL FILL_2__8350_ (
);

BUFX2 _6869_ (
    .A(_1_[31]),
    .Y(memoryAddress[31])
);

FILL FILL_4__8696_ (
);

FILL FILL_4__8276_ (
);

FILL FILL_2__12596_ (
);

FILL SFILL38920x76050 (
);

FILL FILL_2__12176_ (
);

FILL FILL_5__13930_ (
);

FILL FILL_5__13510_ (
);

INVX1 _7810_ (
    .A(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_465_)
);

FILL FILL_1__11589_ (
);

FILL FILL_1__11169_ (
);

FILL FILL_4__12503_ (
);

FILL FILL_0__8596_ (
);

DFFSR _10867_ (
    .Q(\datapath_1.regfile_1.regOut[31] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_1953_[29])
);

OAI21X1 _10447_ (
    .A(_1815_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1816_),
    .Y(_1758_[29])
);

OAI21X1 _10027_ (
    .A(_1596_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1597_),
    .Y(_1563_[17])
);

FILL FILL_3__11916_ (
);

FILL FILL_4__15395_ (
);

FILL FILL_1__12530_ (
);

FILL FILL_1__12110_ (
);

FILL FILL_2__10909_ (
);

FILL FILL_2__9975_ (
);

FILL FILL_0__11943_ (
);

FILL FILL_2__9555_ (
);

FILL FILL_3__14388_ (
);

FILL FILL_2__9135_ (
);

FILL FILL_0__11523_ (
);

FILL FILL_0__11103_ (
);

FILL SFILL83960x71050 (
);

FILL FILL_5__7980_ (
);

FILL FILL_5__7560_ (
);

FILL SFILL3560x75050 (
);

INVX1 _14280_ (
    .A(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_4775_)
);

FILL FILL_5__14715_ (
);

FILL FILL_0__6909_ (
);

FILL FILL_1__7972_ (
);

FILL FILL_1__7552_ (
);

FILL FILL_4__13708_ (
);

FILL FILL_2__14742_ (
);

FILL FILL_2__14322_ (
);

FILL FILL_3__7478_ (
);

FILL FILL_3__7058_ (
);

FILL SFILL44120x7050 (
);

FILL FILL_1__13735_ (
);

FILL FILL_1__13315_ (
);

FILL SFILL3960x44050 (
);

FILL FILL_0__12728_ (
);

FILL FILL_0__12308_ (
);

FILL SFILL38840x38050 (
);

FILL FILL_5__8765_ (
);

FILL FILL_5__8345_ (
);

OAI22X1 _15485_ (
    .A(_5954_),
    .B(_5518__bF$buf0),
    .C(_5478__bF$buf3),
    .D(_5953_),
    .Y(_5955_)
);

NAND3X1 _15065_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5462_),
    .C(_5468_),
    .Y(_5545_)
);

FILL FILL_3__16114_ (
);

FILL SFILL28920x74050 (
);

FILL SFILL3560x30050 (
);

FILL FILL_5__10635_ (
);

FILL FILL_1__8757_ (
);

FILL FILL_1__8337_ (
);

FILL FILL_2__15947_ (
);

FILL FILL_2__15527_ (
);

FILL FILL_2__15107_ (
);

FILL FILL_0__16141_ (
);

FILL FILL_2__10662_ (
);

FILL FILL_2__10242_ (
);

FILL FILL112200x25050 (
);

FILL FILL_3__9624_ (
);

FILL FILL_3_BUFX2_insert400 (
);

FILL FILL_3_BUFX2_insert401 (
);

FILL FILL_3_BUFX2_insert402 (
);

FILL FILL_3_BUFX2_insert403 (
);

FILL FILL_3_BUFX2_insert404 (
);

FILL SFILL3480x37050 (
);

FILL FILL_3_BUFX2_insert405 (
);

FILL FILL_3_BUFX2_insert406 (
);

FILL FILL_3_BUFX2_insert407 (
);

FILL FILL_3_BUFX2_insert408 (
);

FILL FILL_4__13881_ (
);

FILL FILL_3_BUFX2_insert409 (
);

FILL FILL_4__13461_ (
);

FILL FILL_4__13041_ (
);

FILL FILL_2__7621_ (
);

FILL FILL_3__12874_ (
);

FILL FILL_2__7201_ (
);

FILL FILL_3__12454_ (
);

FILL FILL_3__12034_ (
);

FILL FILL_4__7967_ (
);

FILL FILL_4__7547_ (
);

FILL FILL_2__11867_ (
);

FILL FILL_2__11447_ (
);

FILL FILL_0__12481_ (
);

FILL FILL_2__11027_ (
);

FILL FILL_0__12061_ (
);

FILL FILL_5__15673_ (
);

FILL FILL_0__7867_ (
);

FILL FILL_5__15253_ (
);

FILL FILL_0__7447_ (
);

DFFSR _9973_ (
    .Q(\datapath_1.regfile_1.regOut[24] [31]),
    .CLK(clk_bF$buf15),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_1498_[31])
);

NAND2X1 _9553_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1363_)
);

NAND2X1 _9133_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1144_)
);

FILL FILL_1__8090_ (
);

FILL SFILL28840x36050 (
);

FILL FILL_1__11801_ (
);

FILL FILL_4__14666_ (
);

FILL FILL_4__14246_ (
);

FILL FILL_2__15280_ (
);

FILL FILL_2__8826_ (
);

FILL FILL_3__13659_ (
);

FILL FILL_3__13239_ (
);

FILL FILL_1__14693_ (
);

FILL FILL_1__14273_ (
);

FILL SFILL33800x19050 (
);

FILL SFILL18920x72050 (
);

FILL FILL_0_BUFX2_insert530 (
);

FILL FILL_0_BUFX2_insert531 (
);

FILL FILL_0_BUFX2_insert532 (
);

FILL FILL_0_BUFX2_insert533 (
);

FILL FILL_0_BUFX2_insert534 (
);

FILL FILL_0__13686_ (
);

AOI22X1 _13971_ (
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .B(_4154_),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_4473_)
);

FILL FILL_0_BUFX2_insert535 (
);

FILL FILL_0__13266_ (
);

NOR2X1 _13551_ (
    .A(_4057_),
    .B(_4060_),
    .Y(_4061_)
);

FILL FILL_0_BUFX2_insert536 (
);

NAND2X1 _13131_ (
    .A(PCEn_bF$buf0),
    .B(\datapath_1.mux_pcsrc.dout [17]),
    .Y(_3719_)
);

FILL FILL_0_BUFX2_insert537 (
);

FILL FILL_3__14600_ (
);

FILL FILL_0_BUFX2_insert538 (
);

FILL FILL_0_BUFX2_insert539 (
);

FILL SFILL73880x31050 (
);

FILL SFILL89480x16050 (
);

FILL FILL_5__16038_ (
);

FILL FILL_5__11593_ (
);

FILL FILL_1__9295_ (
);

FILL FILL_5__11173_ (
);

FILL FILL_2__16065_ (
);

FILL FILL_4__10166_ (
);

FILL FILL_1__15898_ (
);

FILL FILL_1__15478_ (
);

FILL FILL_1__15058_ (
);

FILL FILL_5__7616_ (
);

FILL FILL_1__10193_ (
);

FILL SFILL13800x9050 (
);

INVX1 _14756_ (
    .A(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_5241_)
);

OAI22X1 _14336_ (
    .A(_4828_),
    .B(_3955__bF$buf1),
    .C(_3924__bF$buf1),
    .D(_4829_),
    .Y(_4830_)
);

FILL FILL_3__15805_ (
);

FILL FILL_3__10940_ (
);

FILL FILL_1__7608_ (
);

FILL FILL_3__10520_ (
);

FILL FILL_0__15832_ (
);

FILL SFILL79480x59050 (
);

FILL FILL_0__15412_ (
);

FILL FILL_5__12378_ (
);

FILL FILL_4__8085_ (
);

FILL SFILL18840x34050 (
);

FILL FILL_1__11398_ (
);

FILL FILL_4__12732_ (
);

FILL FILL_4__12312_ (
);

FILL FILL_6__9792_ (
);

OAI21X1 _10676_ (
    .A(_1927_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .C(_1928_),
    .Y(_1888_[20])
);

OAI21X1 _10256_ (
    .A(_1708_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1709_),
    .Y(_1693_[8])
);

FILL FILL_3__11725_ (
);

FILL FILL_3__11305_ (
);

FILL FILL_2__9784_ (
);

FILL FILL_0__11752_ (
);

FILL FILL_2__9364_ (
);

FILL FILL_3__14197_ (
);

FILL FILL_0__11332_ (
);

FILL FILL_6__15951_ (
);

FILL FILL_6__15531_ (
);

FILL FILL_5__14944_ (
);

FILL FILL_5__14524_ (
);

FILL FILL_5__14104_ (
);

OAI21X1 _8824_ (
    .A(_1041_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1042_),
    .Y(_978_[0])
);

NAND2X1 _8404_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_780_)
);

FILL FILL_1__7361_ (
);

FILL FILL_4__13937_ (
);

FILL FILL_2__14971_ (
);

FILL FILL_4__13517_ (
);

FILL FILL_2__14551_ (
);

FILL FILL_2__14131_ (
);

FILL FILL_3__7287_ (
);

FILL FILL_1__13964_ (
);

FILL FILL_1__13544_ (
);

FILL FILL_1__13124_ (
);

FILL FILL_0__12957_ (
);

DFFSR _12822_ (
    .Q(\control_1.op [5]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3490_[31])
);

FILL SFILL114520x82050 (
);

OAI21X1 _12402_ (
    .A(_3332_),
    .B(MemToReg_bF$buf6),
    .C(_3333_),
    .Y(\datapath_1.mux_wd3.dout [19])
);

FILL FILL_0__12117_ (
);

FILL FILL_5__8994_ (
);

FILL FILL_5__8574_ (
);

FILL FILL_6__11871_ (
);

FILL FILL_6__11451_ (
);

FILL FILL_6__11031_ (
);

NAND2X1 _15294_ (
    .A(_5768_),
    .B(_5764_),
    .Y(_5769_)
);

FILL FILL_5__15729_ (
);

FILL FILL_5__15309_ (
);

FILL FILL_3__16343_ (
);

NAND2X1 _9609_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1380_)
);

FILL FILL_1__8986_ (
);

FILL FILL_5__10444_ (
);

FILL FILL_1__8566_ (
);

FILL FILL_5__10024_ (
);

FILL FILL_1__8146_ (
);

FILL SFILL69080x43050 (
);

FILL FILL_2__15756_ (
);

FILL FILL_4__6991_ (
);

FILL FILL_2__15336_ (
);

FILL FILL_0__16370_ (
);

FILL FILL_2__10891_ (
);

FILL FILL_2__10051_ (
);

FILL FILL_1__14749_ (
);

FILL FILL_1__14329_ (
);

FILL FILL_3__9853_ (
);

INVX1 _13607_ (
    .A(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_4116_)
);

FILL FILL_3__9013_ (
);

FILL FILL_0__6891_ (
);

FILL FILL_5__9779_ (
);

FILL FILL_5__9359_ (
);

FILL FILL_4__13690_ (
);

FILL FILL_4__13270_ (
);

OAI22X1 _16079_ (
    .A(_5148_),
    .B(_5548__bF$buf4),
    .C(_5489__bF$buf3),
    .D(_5163_),
    .Y(_6534_)
);

FILL FILL_2__7850_ (
);

FILL FILL_5__11649_ (
);

FILL FILL_5__11229_ (
);

FILL FILL_2__7430_ (
);

FILL FILL_3__12263_ (
);

FILL FILL_4__7356_ (
);

FILL SFILL85000x50 (
);

FILL FILL_2__11676_ (
);

FILL FILL_2__11256_ (
);

FILL FILL_0__12290_ (
);

FILL FILL_1__10669_ (
);

FILL FILL_1__10249_ (
);

FILL SFILL3640x63050 (
);

FILL FILL_5__15482_ (
);

FILL FILL_5__15062_ (
);

FILL FILL_0__7676_ (
);

NAND2X1 _9782_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1475_)
);

NAND2X1 _9362_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1256_)
);

FILL SFILL43880x70050 (
);

FILL FILL_4__14895_ (
);

FILL FILL_4__14475_ (
);

FILL FILL_1__11610_ (
);

FILL FILL_4__14055_ (
);

FILL FILL_2__8635_ (
);

FILL FILL_3__13888_ (
);

FILL FILL_3__13468_ (
);

FILL FILL_2__8215_ (
);

FILL SFILL3560x1050 (
);

FILL FILL_1__14082_ (
);

FILL SFILL59080x41050 (
);

INVX1 _13780_ (
    .A(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_4286_)
);

FILL FILL_0__13495_ (
);

OAI21X1 _13360_ (
    .A(_3765_),
    .B(_3753_),
    .C(_3875_),
    .Y(_3876_)
);

FILL SFILL38920x26050 (
);

FILL FILL_4__9922_ (
);

FILL FILL_4__9502_ (
);

FILL FILL_2__13822_ (
);

FILL FILL_2__13402_ (
);

FILL FILL_5__16267_ (
);

FILL FILL_3__6978_ (
);

FILL FILL_2__16294_ (
);

FILL FILL_4__10395_ (
);

FILL FILL_0__9402_ (
);

FILL FILL_0__11808_ (
);

FILL FILL_1__15287_ (
);

FILL FILL_5__7845_ (
);

FILL FILL_5__7425_ (
);

FILL FILL_4__16201_ (
);

NOR2X1 _14985_ (
    .A(\datapath_1.PCJump [25]),
    .B(_5464_),
    .Y(_5465_)
);

INVX1 _14565_ (
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_5054_)
);

AOI22X1 _14145_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [14]),
    .C(\datapath_1.regfile_1.regOut[6] [14]),
    .D(_4001__bF$buf3),
    .Y(_4643_)
);

FILL FILL_3__15614_ (
);

FILL SFILL28920x69050 (
);

FILL SFILL3560x25050 (
);

FILL FILL_1__7837_ (
);

FILL FILL_1__7417_ (
);

FILL FILL_2__14607_ (
);

FILL FILL_0__15641_ (
);

FILL FILL_0__15221_ (
);

FILL FILL_5__12187_ (
);

FILL FILL_3__8704_ (
);

FILL FILL_6__11927_ (
);

FILL FILL_4__12961_ (
);

FILL FILL_6__11507_ (
);

FILL FILL_4__12121_ (
);

DFFSR _10485_ (
    .Q(\datapath_1.regfile_1.regOut[28] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1758_[31])
);

NAND2X1 _10065_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1623_)
);

FILL FILL_3__11954_ (
);

FILL FILL_3__11534_ (
);

FILL FILL_3__11114_ (
);

FILL FILL_0__16006_ (
);

FILL FILL_2__10947_ (
);

FILL FILL_0__11981_ (
);

FILL FILL_2__9593_ (
);

FILL FILL_2__10527_ (
);

FILL FILL_2__9173_ (
);

FILL FILL_0__11561_ (
);

FILL FILL_2__10107_ (
);

FILL FILL_0__11141_ (
);

FILL FILL_4__9099_ (
);

FILL FILL_3__9909_ (
);

FILL FILL_5__14753_ (
);

FILL FILL_0__6947_ (
);

FILL FILL_5__14333_ (
);

NAND2X1 _8633_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_892_)
);

NAND2X1 _8213_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_673_)
);

FILL FILL_1__7590_ (
);

FILL FILL_1__7170_ (
);

FILL FILL_4__13746_ (
);

FILL FILL_4__13326_ (
);

FILL FILL_2__14780_ (
);

FILL FILL_2__14360_ (
);

FILL FILL_3__7096_ (
);

FILL FILL_3__12739_ (
);

FILL FILL_1__13773_ (
);

FILL FILL_3__12319_ (
);

FILL FILL_1__13353_ (
);

FILL SFILL18920x67050 (
);

FILL FILL_0__12766_ (
);

NAND2X1 _12631_ (
    .A(vdd),
    .B(memoryOutData[21]),
    .Y(_3467_)
);

FILL FILL_0__12346_ (
);

INVX8 _12211_ (
    .A(ALUSrcB_1_bF$buf2),
    .Y(_3196_)
);

FILL FILL_5__8383_ (
);

FILL FILL_6__16125_ (
);

FILL FILL_5__15958_ (
);

FILL FILL_5__15538_ (
);

FILL FILL_5__15118_ (
);

DFFSR _9838_ (
    .Q(\datapath_1.regfile_1.regOut[23] [24]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_1433_[24])
);

FILL FILL_3__16152_ (
);

INVX1 _9418_ (
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_1293_)
);

FILL FILL_5__10673_ (
);

FILL FILL_1__8375_ (
);

FILL FILL_5__10253_ (
);

FILL FILL_2__15985_ (
);

FILL FILL_2__15565_ (
);

FILL FILL_2__15145_ (
);

FILL FILL_2__10280_ (
);

FILL FILL_1__14978_ (
);

FILL FILL_1__14558_ (
);

FILL FILL_1__14138_ (
);

FILL FILL_3__9662_ (
);

OAI22X1 _13836_ (
    .A(_4340_),
    .B(_3982__bF$buf1),
    .C(_3983__bF$buf4),
    .D(_4339_),
    .Y(_4341_)
);

FILL FILL_3__9242_ (
);

INVX1 _13416_ (
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_3928_)
);

FILL SFILL79160x33050 (
);

FILL FILL_5__9168_ (
);

FILL FILL_0__14912_ (
);

FILL FILL_5__11878_ (
);

FILL FILL_5__11458_ (
);

FILL FILL_3__12492_ (
);

FILL FILL_5__11038_ (
);

FILL FILL_3__12072_ (
);

FILL FILL_4__7585_ (
);

FILL FILL_4__7165_ (
);

FILL SFILL18840x29050 (
);

FILL FILL_2__11485_ (
);

FILL FILL_2__11065_ (
);

FILL FILL_1__10898_ (
);

FILL FILL_1__10058_ (
);

FILL FILL_4__11812_ (
);

FILL FILL_5__15291_ (
);

FILL FILL_6__8872_ (
);

FILL FILL_0__7485_ (
);

NAND2X1 _9591_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .Y(_1432_)
);

FILL FILL_0__7065_ (
);

INVX1 _9171_ (
    .A(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_1169_)
);

FILL FILL_3__10805_ (
);

FILL FILL_4__14284_ (
);

FILL FILL111720x44050 (
);

FILL FILL_2__8864_ (
);

FILL FILL_0__10832_ (
);

FILL FILL_2__8444_ (
);

FILL FILL_3__13697_ (
);

FILL FILL_3__13277_ (
);

FILL FILL_0__10412_ (
);

FILL FILL_0_BUFX2_insert910 (
);

FILL FILL_0_BUFX2_insert911 (
);

FILL FILL_0_BUFX2_insert912 (
);

FILL FILL_0_BUFX2_insert913 (
);

FILL FILL_0_BUFX2_insert914 (
);

FILL FILL_0_BUFX2_insert915 (
);

FILL FILL_0_BUFX2_insert916 (
);

FILL SFILL114600x70050 (
);

FILL FILL_5__13604_ (
);

FILL FILL_0_BUFX2_insert917 (
);

FILL FILL_0_BUFX2_insert918 (
);

FILL SFILL84360x51050 (
);

FILL FILL_0_BUFX2_insert919 (
);

DFFSR _7904_ (
    .Q(\datapath_1.regfile_1.regOut[8] [10]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_458_[10])
);

FILL FILL_1__6861_ (
);

FILL FILL_4__9731_ (
);

FILL FILL_2__13631_ (
);

FILL FILL_2__13211_ (
);

FILL FILL_5__16076_ (
);

FILL FILL_1__12624_ (
);

FILL FILL_4__15489_ (
);

FILL FILL_1__12204_ (
);

FILL FILL_4__15069_ (
);

FILL FILL_6_CLKBUF1_insert1083 (
);

FILL FILL_2__9649_ (
);

FILL FILL_0__9631_ (
);

FILL FILL_2__9229_ (
);

INVX1 _11902_ (
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_2976_)
);

FILL FILL_0__9211_ (
);

FILL FILL_0__11617_ (
);

FILL FILL_1__15096_ (
);

FILL FILL_5__7234_ (
);

FILL FILL_4__16010_ (
);

FILL FILL_6__10951_ (
);

INVX1 _14794_ (
    .A(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_5278_)
);

NOR2X1 _14374_ (
    .A(_4863_),
    .B(_4866_),
    .Y(_4867_)
);

FILL FILL_0__14089_ (
);

FILL FILL_5__14809_ (
);

FILL FILL_3__15843_ (
);

FILL FILL_3__15423_ (
);

FILL FILL_3__15003_ (
);

FILL FILL_1__7226_ (
);

FILL SFILL69080x38050 (
);

FILL FILL_2__14836_ (
);

FILL FILL_0__15870_ (
);

FILL FILL_2__14416_ (
);

FILL FILL_0__15450_ (
);

FILL FILL_0__15030_ (
);

FILL SFILL114920x46050 (
);

FILL FILL_1__13829_ (
);

FILL FILL_1__13409_ (
);

FILL FILL_3__8513_ (
);

FILL FILL_5__8859_ (
);

FILL FILL_5__8439_ (
);

FILL SFILL114520x32050 (
);

FILL FILL_5__8019_ (
);

INVX1 _15999_ (
    .A(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_6456_)
);

FILL FILL_4__12770_ (
);

NOR2X1 _15579_ (
    .A(_6045_),
    .B(_6043_),
    .Y(_6046_)
);

FILL FILL_4__12350_ (
);

OAI22X1 _15159_ (
    .A(_5527__bF$buf3),
    .B(_4045_),
    .C(_5636_),
    .D(_5532__bF$buf1),
    .Y(_5637_)
);

FILL FILL_3__16208_ (
);

NAND2X1 _10294_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1735_)
);

FILL FILL_2__6930_ (
);

FILL FILL_5__10309_ (
);

FILL FILL_3__11763_ (
);

FILL FILL_5__9800_ (
);

FILL FILL_3__11343_ (
);

FILL FILL_4__6856_ (
);

FILL FILL_0__16235_ (
);

NOR2X1 _16100_ (
    .A(_6553_),
    .B(_6552_),
    .Y(_6554_)
);

FILL FILL_2__10756_ (
);

FILL FILL_0__11790_ (
);

FILL FILL_0__11370_ (
);

FILL FILL_3__9718_ (
);

FILL FILL_5__14982_ (
);

FILL FILL_5__14562_ (
);

FILL FILL_5__14142_ (
);

NAND2X1 _8862_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1004_)
);

NAND2X1 _8442_ (
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_785_)
);

FILL SFILL104520x75050 (
);

DFFSR _8022_ (
    .Q(\datapath_1.regfile_1.regOut[9] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_523_[0])
);

FILL FILL_4__13975_ (
);

FILL FILL_4__13555_ (
);

FILL FILL_4__13135_ (
);

OAI21X1 _11499_ (
    .A(_2261_),
    .B(_2284_),
    .C(_2611_),
    .Y(_2612_)
);

NAND2X1 _11079_ (
    .A(\datapath_1.alu_1.ALUInA [8]),
    .B(_2197_),
    .Y(_2198_)
);

FILL SFILL7960x66050 (
);

FILL FILL_2__7715_ (
);

FILL FILL_3__12968_ (
);

FILL FILL_3__12128_ (
);

FILL FILL_1__13582_ (
);

FILL FILL_1__13162_ (
);

FILL SFILL59080x36050 (
);

FILL FILL_0__12995_ (
);

FILL FILL_3_CLKBUF1_insert190 (
);

FILL FILL_0__12575_ (
);

NAND2X1 _12860_ (
    .A(vdd),
    .B(\datapath_1.rd1 [12]),
    .Y(_3579_)
);

FILL FILL_3_CLKBUF1_insert191 (
);

NAND2X1 _12440_ (
    .A(\datapath_1.ALUResult [0]),
    .B(vdd),
    .Y(_3424_)
);

FILL FILL_0__12155_ (
);

FILL FILL_3_CLKBUF1_insert192 (
);

NAND3X1 _12020_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [8]),
    .C(_3034__bF$buf0),
    .Y(_3061_)
);

FILL FILL_3_CLKBUF1_insert193 (
);

FILL FILL_3_CLKBUF1_insert194 (
);

FILL FILL_5__8192_ (
);

FILL FILL_3_CLKBUF1_insert195 (
);

FILL FILL_3_CLKBUF1_insert196 (
);

FILL FILL_3_CLKBUF1_insert197 (
);

FILL FILL_3_CLKBUF1_insert198 (
);

FILL FILL_3_CLKBUF1_insert199 (
);

FILL FILL_5_BUFX2_insert310 (
);

FILL FILL_2__12902_ (
);

FILL FILL_5__15767_ (
);

FILL FILL_5_BUFX2_insert311 (
);

FILL FILL_5__15347_ (
);

FILL FILL_5_BUFX2_insert312 (
);

FILL FILL_5_BUFX2_insert313 (
);

FILL FILL_3__16381_ (
);

FILL FILL_5_BUFX2_insert314 (
);

INVX1 _9647_ (
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_1405_)
);

INVX1 _9227_ (
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_1186_)
);

FILL FILL_5_BUFX2_insert315 (
);

FILL SFILL3640x13050 (
);

FILL FILL_5_BUFX2_insert316 (
);

FILL FILL_5__10062_ (
);

FILL FILL_5_BUFX2_insert317 (
);

FILL FILL_1__8184_ (
);

FILL FILL_5_BUFX2_insert318 (
);

FILL FILL_5_BUFX2_insert319 (
);

FILL FILL_2__15794_ (
);

FILL FILL_2__15374_ (
);

FILL SFILL104520x30050 (
);

FILL SFILL43880x20050 (
);

FILL FILL_0__8902_ (
);

FILL FILL_1__14787_ (
);

FILL FILL_1__14367_ (
);

FILL FILL_5__6925_ (
);

FILL FILL_4__15701_ (
);

FILL FILL_3__9891_ (
);

FILL FILL_3__9471_ (
);

AOI22X1 _13645_ (
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .B(_3950__bF$buf1),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_4153_)
);

OAI22X1 _13225_ (
    .A(_3752_),
    .B(_3767_),
    .C(_3765_),
    .D(_3766_),
    .Y(_3768_)
);

FILL FILL_5__9397_ (
);

FILL FILL_1__6917_ (
);

FILL SFILL104440x37050 (
);

FILL FILL_0__14721_ (
);

FILL FILL_0__14301_ (
);

FILL FILL_5__11687_ (
);

FILL FILL_1__9389_ (
);

FILL FILL_5__11267_ (
);

FILL FILL_2__16159_ (
);

FILL FILL_2__11294_ (
);

FILL FILL_2_BUFX2_insert440 (
);

FILL FILL_1__10287_ (
);

FILL FILL_2_BUFX2_insert441 (
);

FILL FILL_2_BUFX2_insert442 (
);

FILL FILL_2_BUFX2_insert443 (
);

FILL FILL_2_BUFX2_insert444 (
);

FILL FILL_4__11621_ (
);

FILL FILL_2_BUFX2_insert445 (
);

FILL FILL_4__11201_ (
);

FILL FILL_2_BUFX2_insert446 (
);

FILL FILL_2_BUFX2_insert447 (
);

FILL FILL_0__7294_ (
);

FILL SFILL49080x34050 (
);

FILL FILL_2_BUFX2_insert448 (
);

FILL FILL_2_BUFX2_insert449 (
);

FILL FILL_6__13899_ (
);

FILL FILL_3__10614_ (
);

FILL FILL_0_CLKBUF1_insert140 (
);

FILL FILL_0_CLKBUF1_insert141 (
);

FILL FILL_4__14093_ (
);

FILL FILL_0_CLKBUF1_insert142 (
);

FILL FILL_0__15926_ (
);

FILL FILL_0__15506_ (
);

FILL FILL_0_CLKBUF1_insert143 (
);

FILL FILL_0_CLKBUF1_insert144 (
);

FILL FILL_0_CLKBUF1_insert145 (
);

FILL FILL_0_CLKBUF1_insert146 (
);

FILL FILL_2__8253_ (
);

FILL FILL_0__10641_ (
);

FILL FILL_0_CLKBUF1_insert147 (
);

FILL FILL_3__13086_ (
);

FILL FILL_0_CLKBUF1_insert148 (
);

FILL FILL_0_CLKBUF1_insert149 (
);

FILL FILL_6__14840_ (
);

FILL FILL_4__8599_ (
);

FILL FILL_2__12499_ (
);

FILL FILL_2__12079_ (
);

FILL FILL_5__13833_ (
);

FILL FILL_5__13413_ (
);

NAND2X1 _7713_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_421_)
);

FILL FILL_4__9540_ (
);

FILL FILL_4__9120_ (
);

FILL FILL_4__12826_ (
);

FILL FILL_4__12406_ (
);

FILL FILL_2__13860_ (
);

FILL FILL_2__13440_ (
);

FILL FILL_2__13020_ (
);

FILL FILL_0__8499_ (
);

FILL FILL_6__9886_ (
);

FILL SFILL49000x32050 (
);

FILL FILL_0__8079_ (
);

FILL FILL_3__11819_ (
);

FILL FILL_1__12853_ (
);

FILL FILL_4__15298_ (
);

FILL FILL_1__12433_ (
);

FILL FILL_1__12013_ (
);

FILL FILL_0__9860_ (
);

FILL FILL_2__9878_ (
);

FILL FILL_0__11846_ (
);

FILL FILL_2__9038_ (
);

FILL FILL_0__9020_ (
);

FILL FILL_0__11426_ (
);

INVX1 _11711_ (
    .A(_2192_),
    .Y(_2810_)
);

FILL FILL_0__11006_ (
);

FILL FILL_5__7883_ (
);

FILL FILL_5__7463_ (
);

FILL FILL_5__7043_ (
);

FILL FILL_6__10760_ (
);

FILL SFILL18520x48050 (
);

INVX1 _14183_ (
    .A(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_4680_)
);

FILL FILL_5__14618_ (
);

FILL SFILL23880x61050 (
);

FILL FILL_3__15652_ (
);

DFFSR _8918_ (
    .Q(\datapath_1.regfile_1.regOut[16] [0]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_978_[0])
);

FILL FILL_3__15232_ (
);

FILL FILL_1__7875_ (
);

FILL FILL_1__7455_ (
);

FILL FILL_1__7035_ (
);

FILL FILL_2__14645_ (
);

FILL FILL_2__14225_ (
);

FILL SFILL39000x75050 (
);

FILL SFILL94360x48050 (
);

FILL FILL_1__13638_ (
);

FILL FILL_1__13218_ (
);

FILL FILL_1_BUFX2_insert460 (
);

FILL FILL_3__8742_ (
);

FILL FILL_1_BUFX2_insert461 (
);

FILL FILL_3__8322_ (
);

FILL FILL_1_BUFX2_insert462 (
);

INVX1 _12916_ (
    .A(\datapath_1.a [31]),
    .Y(_3616_)
);

FILL FILL_1_BUFX2_insert463 (
);

FILL FILL_1_BUFX2_insert464 (
);

FILL FILL_1_BUFX2_insert465 (
);

FILL SFILL79160x28050 (
);

FILL FILL_1_BUFX2_insert466 (
);

FILL FILL_5__8248_ (
);

FILL FILL_1_BUFX2_insert467 (
);

FILL FILL_1_BUFX2_insert468 (
);

FILL FILL_1_BUFX2_insert469 (
);

NAND3X1 _15388_ (
    .A(_5854_),
    .B(_5855_),
    .C(_5859_),
    .Y(_5860_)
);

FILL FILL_3__16017_ (
);

FILL FILL_5__10958_ (
);

FILL FILL_3__11992_ (
);

FILL FILL_5__10538_ (
);

FILL FILL_3__11572_ (
);

FILL FILL_5__10118_ (
);

FILL FILL_3__11152_ (
);

FILL FILL_0__16044_ (
);

FILL FILL_2__10565_ (
);

FILL FILL_2__10145_ (
);

FILL SFILL63960x12050 (
);

FILL SFILL39000x30050 (
);

FILL FILL_1__9601_ (
);

FILL FILL_3__9527_ (
);

FILL FILL_3__9107_ (
);

FILL FILL_5__14791_ (
);

FILL FILL_5__14371_ (
);

FILL FILL_0__6985_ (
);

FILL FILL112280x3050 (
);

DFFSR _8671_ (
    .Q(\datapath_1.regfile_1.regOut[14] [9]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_848_[9])
);

FILL FILL111960x6050 (
);

INVX1 _8251_ (
    .A(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_698_)
);

FILL FILL_4__13784_ (
);

FILL FILL_4__13364_ (
);

FILL FILL_2__7944_ (
);

FILL FILL_3__12777_ (
);

FILL FILL_2__7104_ (
);

FILL FILL_3__12357_ (
);

FILL FILL_1__13391_ (
);

FILL FILL_0__12384_ (
);

FILL SFILL53960x55050 (
);

FILL SFILL29000x73050 (
);

FILL FILL_2_CLKBUF1_insert180 (
);

FILL FILL_2_CLKBUF1_insert181 (
);

FILL FILL_5__15996_ (
);

FILL FILL_2_CLKBUF1_insert182 (
);

FILL FILL_2__12711_ (
);

FILL FILL_2_CLKBUF1_insert183 (
);

FILL FILL_5__15576_ (
);

FILL FILL_2_CLKBUF1_insert184 (
);

FILL FILL_5__15156_ (
);

FILL FILL_2_CLKBUF1_insert185 (
);

FILL FILL_3__16190_ (
);

INVX1 _9876_ (
    .A(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_1517_)
);

FILL FILL_2_CLKBUF1_insert186 (
);

DFFSR _9456_ (
    .Q(\datapath_1.regfile_1.regOut[20] [26]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_1238_[26])
);

FILL FILL_2_CLKBUF1_insert187 (
);

OAI21X1 _9036_ (
    .A(_1098_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .C(_1099_),
    .Y(_1043_[28])
);

FILL FILL_2_CLKBUF1_insert188 (
);

FILL FILL_5__10291_ (
);

FILL FILL_4__14989_ (
);

FILL FILL_2_CLKBUF1_insert189 (
);

FILL FILL_4__14569_ (
);

FILL FILL_1__11704_ (
);

FILL FILL_4__14149_ (
);

FILL FILL_2__15183_ (
);

FILL FILL_2__8729_ (
);

FILL FILL_0__8711_ (
);

FILL SFILL8760x20050 (
);

FILL FILL_1__14596_ (
);

FILL FILL_1__14176_ (
);

FILL FILL_4__15930_ (
);

FILL FILL_4__15510_ (
);

FILL FILL_6_BUFX2_insert1063 (
);

FILL FILL_3__9280_ (
);

FILL FILL_0__13589_ (
);

INVX1 _13874_ (
    .A(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_4378_)
);

NAND3X1 _13454_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3919_),
    .C(_3879_),
    .Y(_3966_)
);

FILL FILL_0__13169_ (
);

OAI21X1 _13034_ (
    .A(_3673_),
    .B(vdd),
    .C(_3674_),
    .Y(_3620_[27])
);

FILL FILL_6_BUFX2_insert1068 (
);

FILL FILL_3__14923_ (
);

FILL FILL_3__14503_ (
);

FILL SFILL114120x58050 (
);

FILL SFILL114600x20050 (
);

FILL SFILL53960x10050 (
);

FILL FILL_2__13916_ (
);

FILL FILL_0__14950_ (
);

FILL FILL_0__14530_ (
);

FILL FILL_0__14110_ (
);

FILL FILL_5__11496_ (
);

FILL FILL_5__11076_ (
);

FILL FILL_1__12909_ (
);

FILL FILL_2__16388_ (
);

FILL FILL_4__10489_ (
);

FILL FILL_0__9916_ (
);

FILL FILL_4__10069_ (
);

FILL FILL_5__7939_ (
);

FILL SFILL114520x27050 (
);

FILL SFILL53880x17050 (
);

FILL FILL_6__10816_ (
);

FILL FILL_4__11850_ (
);

AOI22X1 _14659_ (
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .B(_3942__bF$buf3),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_5146_)
);

INVX1 _14239_ (
    .A(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_4735_)
);

FILL FILL_4__11430_ (
);

FILL FILL_4__11010_ (
);

FILL FILL_3__15708_ (
);

FILL FILL_6__8490_ (
);

FILL FILL_1__16322_ (
);

FILL SFILL104600x63050 (
);

FILL SFILL43960x53050 (
);

FILL FILL_3__10423_ (
);

FILL FILL_3__10003_ (
);

FILL FILL_0__15735_ (
);

FILL FILL_0__15315_ (
);

INVX1 _15600_ (
    .A(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_6067_)
);

FILL FILL_2__8482_ (
);

FILL FILL_0__10870_ (
);

FILL FILL_2__8062_ (
);

FILL FILL_0__10450_ (
);

FILL FILL_0__10030_ (
);

FILL FILL_5__13642_ (
);

FILL FILL_5__13222_ (
);

NAND2X1 _7942_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_533_)
);

DFFSR _7522_ (
    .Q(\datapath_1.regfile_1.regOut[5] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_263_[12])
);

INVX1 _7102_ (
    .A(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_115_)
);

FILL FILL_4__12635_ (
);

FILL FILL_4__12215_ (
);

INVX1 _10999_ (
    .A(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2118_)
);

FILL FILL_6__9275_ (
);

INVX1 _10579_ (
    .A(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_1884_)
);

INVX1 _10159_ (
    .A(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_1665_)
);

FILL FILL_3__11628_ (
);

FILL FILL_1__12662_ (
);

FILL FILL_3__11208_ (
);

FILL FILL_1__12242_ (
);

FILL FILL112280x64050 (
);

OAI21X1 _11940_ (
    .A(_3000_),
    .B(IorD_bF$buf1),
    .C(_3001_),
    .Y(_1_[17])
);

FILL FILL_2__9267_ (
);

FILL FILL_0__11655_ (
);

FILL FILL_0__11235_ (
);

AOI21X1 _11520_ (
    .A(_2275_),
    .B(_2630_),
    .C(_2629_),
    .Y(_2631_)
);

INVX2 _11100_ (
    .A(_2218_),
    .Y(_2219_)
);

FILL FILL_5__7692_ (
);

FILL FILL_6__15434_ (
);

FILL FILL_6__15014_ (
);

FILL FILL_5__14847_ (
);

FILL FILL_3__15881_ (
);

FILL FILL_5__14427_ (
);

FILL FILL_5__14007_ (
);

FILL FILL_3__15461_ (
);

INVX1 _8727_ (
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_934_)
);

FILL FILL_3__15041_ (
);

DFFSR _8307_ (
    .Q(\datapath_1.regfile_1.regOut[11] [29]),
    .CLK(clk_bF$buf7),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_653_[29])
);

FILL FILL_1__7684_ (
);

FILL FILL_2__14874_ (
);

FILL FILL_2__14454_ (
);

FILL SFILL43880x15050 (
);

FILL FILL_2__14034_ (
);

FILL SFILL68280x81050 (
);

FILL FILL_1__13867_ (
);

FILL FILL_1__13447_ (
);

FILL FILL_1__13027_ (
);

FILL SFILL59000x29050 (
);

FILL FILL_3__8971_ (
);

INVX1 _12725_ (
    .A(\datapath_1.PCJump [12]),
    .Y(_3509_)
);

FILL FILL_3__8131_ (
);

AOI22X1 _12305_ (
    .A(_2_[22]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3268_)
);

FILL FILL_5__8897_ (
);

FILL SFILL84280x2050 (
);

FILL FILL_5__8477_ (
);

FILL FILL_5__8057_ (
);

FILL FILL_6__11354_ (
);

OAI22X1 _15197_ (
    .A(_4125_),
    .B(_5501_),
    .C(_5524__bF$buf3),
    .D(_4109_),
    .Y(_5674_)
);

FILL FILL_0__13801_ (
);

FILL FILL_3__16246_ (
);

FILL FILL_5__10767_ (
);

FILL FILL_1__8889_ (
);

FILL FILL_1__8469_ (
);

FILL FILL_3__11381_ (
);

FILL FILL_2__15659_ (
);

FILL FILL_2__15239_ (
);

FILL FILL_4__6894_ (
);

FILL SFILL33880x58050 (
);

FILL FILL_0__16273_ (
);

FILL FILL_2__10794_ (
);

FILL FILL_2__10374_ (
);

FILL FILL_1__9410_ (
);

FILL FILL_3__9756_ (
);

FILL FILL_3__9336_ (
);

FILL FILL_4__10701_ (
);

FILL FILL_5__14180_ (
);

FILL SFILL33480x44050 (
);

FILL FILL_6__7761_ (
);

INVX1 _8480_ (
    .A(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_810_)
);

INVX1 _8060_ (
    .A(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_591_)
);

FILL FILL_4__13593_ (
);

FILL FILL_4__13173_ (
);

FILL FILL_2__7753_ (
);

FILL FILL_3__12586_ (
);

FILL FILL_2__7333_ (
);

FILL FILL_3__12166_ (
);

FILL FILL_6__13920_ (
);

FILL FILL_4__7679_ (
);

FILL FILL_6__13500_ (
);

FILL FILL_2__11999_ (
);

FILL FILL_2__11579_ (
);

FILL FILL_2__11159_ (
);

FILL FILL_0__12193_ (
);

FILL FILL_5__12913_ (
);

FILL FILL_4__8620_ (
);

FILL FILL_4__8200_ (
);

FILL FILL_4__11906_ (
);

FILL FILL_0__7999_ (
);

FILL FILL_5__15385_ (
);

FILL FILL_2__12520_ (
);

FILL FILL_2__12100_ (
);

FILL FILL_0__7579_ (
);

FILL FILL_6__8966_ (
);

FILL FILL_0__7159_ (
);

OAI21X1 _9685_ (
    .A(_1429_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1430_),
    .Y(_1368_[31])
);

OAI21X1 _9265_ (
    .A(_1210_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1211_),
    .Y(_1173_[19])
);

FILL FILL_1_CLKBUF1_insert170 (
);

FILL FILL_1_CLKBUF1_insert171 (
);

FILL FILL_1__11933_ (
);

FILL FILL_4__14798_ (
);

FILL FILL_1_CLKBUF1_insert172 (
);

FILL FILL_1_CLKBUF1_insert173 (
);

FILL FILL_4__14378_ (
);

FILL FILL_1__11513_ (
);

FILL FILL_1_CLKBUF1_insert174 (
);

FILL FILL_1_CLKBUF1_insert175 (
);

FILL FILL_1_CLKBUF1_insert176 (
);

FILL FILL_1_CLKBUF1_insert177 (
);

FILL SFILL94440x36050 (
);

FILL FILL_1_CLKBUF1_insert178 (
);

FILL FILL_2__8958_ (
);

FILL FILL_0__10926_ (
);

FILL FILL_1_CLKBUF1_insert179 (
);

FILL FILL_0__8520_ (
);

FILL FILL_0__8100_ (
);

FILL FILL_2__8118_ (
);

FILL FILL_0__10506_ (
);

FILL FILL_5__6963_ (
);

FILL FILL_0__13398_ (
);

AOI22X1 _13683_ (
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .B(_4102_),
    .C(_3891__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_4191_)
);

NAND3X1 _13263_ (
    .A(_3803_),
    .B(_3805_),
    .C(_3802_),
    .Y(_3806_)
);

FILL FILL_3__14732_ (
);

FILL SFILL98760x44050 (
);

FILL FILL_3__14312_ (
);

FILL FILL_1__6955_ (
);

FILL FILL_4__9405_ (
);

FILL FILL_2__13725_ (
);

FILL FILL_2__13305_ (
);

FILL FILL_1__12718_ (
);

FILL FILL_2__16197_ (
);

FILL FILL_4__10298_ (
);

FILL FILL_3__7822_ (
);

FILL FILL_0__9725_ (
);

FILL FILL_5__7748_ (
);

FILL FILL_5__7328_ (
);

FILL FILL_2_BUFX2_insert820 (
);

FILL FILL_4__16104_ (
);

FILL FILL_2_BUFX2_insert821 (
);

FILL FILL_2_BUFX2_insert822 (
);

FILL FILL_2_BUFX2_insert823 (
);

NOR2X1 _14888_ (
    .A(_5366_),
    .B(_5369_),
    .Y(_5370_)
);

INVX1 _14468_ (
    .A(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_4959_)
);

FILL FILL_2_BUFX2_insert824 (
);

FILL FILL_2_BUFX2_insert825 (
);

NOR2X1 _14048_ (
    .A(_4547_),
    .B(_4536_),
    .Y(_4548_)
);

FILL FILL_3__15937_ (
);

FILL FILL_2_BUFX2_insert826 (
);

FILL FILL_2_BUFX2_insert827 (
);

FILL FILL_3__15517_ (
);

FILL FILL_2_BUFX2_insert828 (
);

FILL FILL_2_BUFX2_insert829 (
);

FILL FILL_1__16131_ (
);

FILL SFILL23880x11050 (
);

FILL FILL_3__10652_ (
);

FILL FILL_3__10232_ (
);

FILL FILL_0__15964_ (
);

FILL FILL_0__15544_ (
);

FILL FILL_0__15124_ (
);

FILL SFILL53960x4050 (
);

FILL FILL111800x27050 (
);

FILL SFILL39000x25050 (
);

FILL FILL_3__8607_ (
);

FILL FILL_5__13871_ (
);

FILL FILL_5__13451_ (
);

FILL FILL_5__13031_ (
);

INVX1 _7751_ (
    .A(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_446_)
);

INVX1 _7331_ (
    .A(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_227_)
);

FILL FILL_4__12864_ (
);

FILL FILL_4__12444_ (
);

FILL FILL_4__12024_ (
);

INVX1 _10388_ (
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_1777_)
);

FILL FILL_3__11857_ (
);

FILL FILL_1__12891_ (
);

FILL FILL_3__11437_ (
);

FILL FILL_1__12471_ (
);

FILL FILL_3__11017_ (
);

FILL FILL_1__12051_ (
);

FILL FILL_0__16329_ (
);

FILL FILL_0__11884_ (
);

FILL FILL_2__9496_ (
);

FILL FILL_0__11464_ (
);

FILL FILL_0__11044_ (
);

FILL FILL_5__7081_ (
);

FILL FILL_5__14656_ (
);

FILL FILL_3__15690_ (
);

FILL FILL_5__14236_ (
);

FILL FILL_3__15270_ (
);

INVX1 _8956_ (
    .A(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_1046_)
);

DFFSR _8536_ (
    .Q(\datapath_1.regfile_1.regOut[13] [2]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_783_[2])
);

OAI21X1 _8116_ (
    .A(_627_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_628_),
    .Y(_588_[20])
);

FILL FILL_1__7493_ (
);

FILL FILL_1__7073_ (
);

FILL FILL_4__13649_ (
);

FILL FILL_4__13229_ (
);

FILL FILL_2__14683_ (
);

FILL FILL_2__14263_ (
);

FILL SFILL8760x15050 (
);

FILL FILL_2__7809_ (
);

FILL SFILL13800x52050 (
);

FILL FILL_1__13676_ (
);

FILL FILL_1__13256_ (
);

FILL FILL_1_BUFX2_insert840 (
);

FILL FILL_3__8780_ (
);

FILL FILL_1_BUFX2_insert841 (
);

FILL FILL_3__8360_ (
);

FILL FILL_1_BUFX2_insert842 (
);

INVX1 _12954_ (
    .A(_2_[1]),
    .Y(_3621_)
);

OAI21X1 _12534_ (
    .A(_3421_),
    .B(vdd),
    .C(_3422_),
    .Y(_3360_[31])
);

FILL FILL_0__12249_ (
);

FILL FILL_1_BUFX2_insert843 (
);

NAND3X1 _12114_ (
    .A(_3129_),
    .B(_3130_),
    .C(_3131_),
    .Y(\datapath_1.mux_pcsrc.dout [31])
);

FILL FILL_1_BUFX2_insert844 (
);

FILL FILL_1_BUFX2_insert845 (
);

FILL FILL_1_BUFX2_insert846 (
);

FILL FILL_1_BUFX2_insert847 (
);

FILL FILL_1_BUFX2_insert848 (
);

FILL FILL_1_BUFX2_insert849 (
);

FILL FILL_0__13610_ (
);

FILL FILL_3__16055_ (
);

FILL FILL_5__10996_ (
);

FILL FILL_5__10576_ (
);

FILL FILL_1__8698_ (
);

FILL FILL_5__10156_ (
);

FILL FILL_3__11190_ (
);

FILL FILL_2__15888_ (
);

FILL FILL_2__15468_ (
);

FILL FILL_2__15048_ (
);

FILL FILL_0__16082_ (
);

FILL FILL_2__10183_ (
);

FILL FILL_3__9985_ (
);

FILL FILL_4__10930_ (
);

FILL FILL_3__9145_ (
);

AOI21X1 _13739_ (
    .A(_4221_),
    .B(_4245_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [5])
);

FILL FILL_4__10510_ (
);

OAI21X1 _13319_ (
    .A(\datapath_1.a3 [0]),
    .B(_3786_),
    .C(_3848_),
    .Y(_3850_)
);

FILL FILL_1__15822_ (
);

FILL FILL_6__7570_ (
);

FILL FILL_1__15402_ (
);

FILL SFILL43960x48050 (
);

FILL FILL_0__14815_ (
);

FILL FILL_2__7982_ (
);

BUFX2 BUFX2_insert510 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf97)
);

FILL FILL_2__7562_ (
);

BUFX2 BUFX2_insert511 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf96)
);

FILL FILL_3__12395_ (
);

BUFX2 BUFX2_insert512 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf95)
);

BUFX2 BUFX2_insert513 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf94)
);

BUFX2 BUFX2_insert514 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf93)
);

BUFX2 BUFX2_insert515 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf92)
);

FILL FILL_4__7488_ (
);

BUFX2 BUFX2_insert516 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf91)
);

FILL FILL_4__7068_ (
);

BUFX2 BUFX2_insert517 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf90)
);

FILL FILL112360x52050 (
);

BUFX2 BUFX2_insert518 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf89)
);

FILL FILL_2__11388_ (
);

BUFX2 BUFX2_insert519 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf88)
);

FILL FILL_5__12722_ (
);

FILL FILL_5__12302_ (
);

FILL FILL_4__11715_ (
);

FILL SFILL64040x61050 (
);

FILL SFILL23880x8050 (
);

FILL FILL_5__15194_ (
);

OAI21X1 _9494_ (
    .A(_1322_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1323_),
    .Y(_1303_[10])
);

DFFSR _9074_ (
    .Q(\datapath_1.regfile_1.regOut[17] [28]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_1043_[28])
);

FILL FILL_3__10708_ (
);

FILL FILL_1__11742_ (
);

FILL FILL_4__14187_ (
);

FILL FILL_1__11322_ (
);

FILL FILL112280x59050 (
);

FILL FILL_2__8767_ (
);

FILL FILL_2__8347_ (
);

FILL FILL_0__10315_ (
);

DFFSR _10600_ (
    .Q(\datapath_1.regfile_1.regOut[29] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_1823_[18])
);

FILL FILL_0_BUFX2_insert30 (
);

FILL FILL_0_BUFX2_insert31 (
);

FILL FILL_0_BUFX2_insert32 (
);

FILL FILL_0_BUFX2_insert33 (
);

FILL FILL_0_BUFX2_insert34 (
);

FILL FILL_0_BUFX2_insert35 (
);

FILL FILL_0_BUFX2_insert36 (
);

FILL FILL_0_BUFX2_insert37 (
);

NOR2X1 _13492_ (
    .A(_4002_),
    .B(_3977__bF$buf2),
    .Y(_4003_)
);

FILL FILL_0_BUFX2_insert38 (
);

FILL FILL_5__13927_ (
);

DFFSR _13072_ (
    .Q(_2_[25]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_3620_[25])
);

FILL FILL_3__14961_ (
);

FILL FILL_5__13507_ (
);

FILL FILL_0_BUFX2_insert39 (
);

FILL FILL_3__14541_ (
);

INVX1 _7807_ (
    .A(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_463_)
);

FILL FILL_3__14121_ (
);

FILL FILL_4_BUFX2_insert350 (
);

FILL FILL_4__9634_ (
);

FILL FILL_4_BUFX2_insert351 (
);

FILL FILL_4__9214_ (
);

FILL FILL_4_BUFX2_insert352 (
);

FILL FILL_4_BUFX2_insert353 (
);

FILL FILL_2__13954_ (
);

FILL FILL_4_BUFX2_insert354 (
);

FILL FILL_5__16399_ (
);

FILL FILL_2__13534_ (
);

FILL FILL_4_BUFX2_insert355 (
);

FILL FILL_2__13114_ (
);

FILL FILL_4_BUFX2_insert356 (
);

FILL FILL_4_BUFX2_insert357 (
);

FILL FILL_4_BUFX2_insert358 (
);

FILL FILL_4_BUFX2_insert359 (
);

FILL FILL_1__12527_ (
);

FILL FILL_1__12107_ (
);

FILL FILL_3__7631_ (
);

FILL FILL_0__9534_ (
);

FILL FILL_0__9114_ (
);

FILL FILL_3__7211_ (
);

AOI21X1 _11805_ (
    .A(_2887_),
    .B(_2620_),
    .C(_2896_),
    .Y(_2897_)
);

FILL FILL112280x14050 (
);

FILL FILL_5__7977_ (
);

FILL FILL_5__7557_ (
);

FILL FILL_4__16333_ (
);

OAI22X1 _14697_ (
    .A(_5182_),
    .B(_3936__bF$buf1),
    .C(_3905__bF$buf0),
    .D(_5181_),
    .Y(_5183_)
);

FILL FILL_6__10434_ (
);

INVX1 _14277_ (
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_4772_)
);

FILL FILL_3__15746_ (
);

FILL FILL_3__15326_ (
);

FILL FILL_1__16360_ (
);

FILL FILL_1__7969_ (
);

FILL FILL_3__10881_ (
);

FILL FILL_1__7549_ (
);

FILL FILL_3__10041_ (
);

FILL SFILL94520x69050 (
);

FILL FILL_2__14739_ (
);

FILL FILL_2__14319_ (
);

FILL FILL_0__15773_ (
);

FILL FILL_0__15353_ (
);

FILL FILL_1__8910_ (
);

FILL FILL_3__8836_ (
);

FILL SFILL98840x77050 (
);

FILL FILL_5__13680_ (
);

FILL FILL_5__13260_ (
);

INVX1 _7980_ (
    .A(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_558_)
);

INVX1 _7560_ (
    .A(\datapath_1.regfile_1.regOut[6] [6]),
    .Y(_339_)
);

DFFSR _7140_ (
    .Q(\datapath_1.regfile_1.regOut[2] [14]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_68_[14])
);

FILL FILL_4__12253_ (
);

OAI21X1 _10197_ (
    .A(_1689_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1690_),
    .Y(_1628_[31])
);

FILL FILL_3__11666_ (
);

FILL FILL_3__11246_ (
);

FILL FILL_1__12280_ (
);

DFFSR _16423_ (
    .Q(\datapath_1.regfile_1.regOut[0] [6]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_6769_[6])
);

FILL FILL_0__16138_ (
);

NOR2X1 _16003_ (
    .A(_6457_),
    .B(_6459_),
    .Y(_6460_)
);

FILL FILL_2__10659_ (
);

FILL FILL_2__10239_ (
);

FILL FILL_0__11693_ (
);

FILL FILL_0__11273_ (
);

FILL SFILL58280x74050 (
);

FILL FILL_3_BUFX2_insert370 (
);

FILL FILL_4__7700_ (
);

FILL FILL_3_BUFX2_insert371 (
);

FILL FILL_3_BUFX2_insert372 (
);

FILL FILL_5__14885_ (
);

FILL FILL_5__14465_ (
);

FILL FILL_3_BUFX2_insert373 (
);

FILL FILL_2__11600_ (
);

FILL FILL_5__14045_ (
);

FILL FILL_3_BUFX2_insert374 (
);

OAI21X1 _8765_ (
    .A(_958_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .C(_959_),
    .Y(_913_[23])
);

FILL FILL_3_BUFX2_insert375 (
);

OAI21X1 _8345_ (
    .A(_739_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .C(_740_),
    .Y(_718_[11])
);

FILL FILL_3_BUFX2_insert376 (
);

FILL FILL_3_BUFX2_insert377 (
);

FILL FILL_3_BUFX2_insert378 (
);

FILL FILL_4__13878_ (
);

FILL FILL_3_BUFX2_insert379 (
);

FILL FILL_4__13458_ (
);

FILL FILL_2__14492_ (
);

FILL FILL_4__13038_ (
);

FILL FILL_2__14072_ (
);

FILL SFILL18920x9050 (
);

FILL FILL_0__7600_ (
);

FILL FILL_2__7618_ (
);

FILL FILL_1__13485_ (
);

FILL SFILL58680x43050 (
);

FILL FILL_0__12898_ (
);

OAI21X1 _12763_ (
    .A(_3533_),
    .B(IRWrite_bF$buf5),
    .C(_3534_),
    .Y(_3490_[22])
);

FILL FILL_0__12478_ (
);

INVX1 _12343_ (
    .A(ALUOut[0]),
    .Y(_3358_)
);

FILL FILL_0__12058_ (
);

FILL SFILL58840x1050 (
);

FILL FILL_3__13812_ (
);

FILL FILL_5__8095_ (
);

FILL SFILL79160x70050 (
);

FILL SFILL59080x3050 (
);

FILL FILL_4__8905_ (
);

FILL FILL_3__16284_ (
);

FILL SFILL88840x75050 (
);

FILL FILL_5__10385_ (
);

FILL FILL_1__8087_ (
);

FILL FILL_2__15697_ (
);

FILL FILL_2__15277_ (
);

FILL FILL_3__6902_ (
);

FILL FILL_4__15604_ (
);

FILL FILL_3__9794_ (
);

INVX1 _13968_ (
    .A(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_4470_)
);

FILL FILL_3__9374_ (
);

FILL SFILL23800x49050 (
);

INVX1 _13548_ (
    .A(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_4058_)
);

NAND2X1 _13128_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [16]),
    .Y(_3717_)
);

FILL SFILL8040x65050 (
);

FILL FILL_1__15631_ (
);

FILL FILL_1__15211_ (
);

FILL FILL_6__12177_ (
);

FILL FILL_0__14624_ (
);

FILL FILL_0__14204_ (
);

FILL FILL_2__7371_ (
);

FILL SFILL44360x33050 (
);

FILL FILL_4__7297_ (
);

FILL FILL_2__11197_ (
);

FILL FILL_5__12951_ (
);

FILL FILL_5__12531_ (
);

FILL FILL_5__12111_ (
);

FILL FILL_4__11944_ (
);

FILL FILL_4__11524_ (
);

FILL FILL_4__11104_ (
);

FILL FILL_0__7197_ (
);

FILL FILL_1__16416_ (
);

FILL FILL_3__10937_ (
);

FILL FILL_1__11971_ (
);

FILL FILL_3__10517_ (
);

FILL FILL_1__11551_ (
);

FILL FILL_1__11131_ (
);

FILL FILL_0__15829_ (
);

FILL FILL_0__15409_ (
);

FILL FILL_2__8996_ (
);

FILL FILL_2__8576_ (
);

FILL FILL_0__10964_ (
);

FILL FILL_0__10544_ (
);

FILL FILL_0__10124_ (
);

FILL FILL_6__14743_ (
);

FILL SFILL74120x51050 (
);

FILL FILL_5__13736_ (
);

FILL FILL_5__13316_ (
);

FILL FILL_3__14770_ (
);

FILL FILL_3__14350_ (
);

OAI21X1 _7616_ (
    .A(_375_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .C(_376_),
    .Y(_328_[24])
);

FILL FILL_1__6993_ (
);

FILL FILL_4__9863_ (
);

FILL FILL_4__12729_ (
);

FILL FILL_4__9023_ (
);

FILL FILL_2__13763_ (
);

FILL FILL_4__12309_ (
);

FILL FILL_2__13343_ (
);

FILL FILL_6__9369_ (
);

FILL SFILL13800x47050 (
);

FILL FILL_1__12756_ (
);

FILL FILL_1__12336_ (
);

FILL FILL_0__9763_ (
);

FILL FILL_3__7860_ (
);

FILL FILL_3__7440_ (
);

FILL FILL_0__9343_ (
);

FILL FILL_0__11749_ (
);

FILL FILL_0__11329_ (
);

INVX1 _11614_ (
    .A(_2419_),
    .Y(_2719_)
);

FILL FILL_5__7366_ (
);

FILL FILL_4__16142_ (
);

FILL FILL_6__10243_ (
);

INVX1 _14086_ (
    .A(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_4585_)
);

FILL FILL_3__15975_ (
);

FILL FILL_3__15555_ (
);

FILL FILL_3__15135_ (
);

FILL FILL_1__7358_ (
);

FILL FILL_3__10690_ (
);

FILL FILL_3__10270_ (
);

FILL FILL_2__14968_ (
);

FILL FILL_2__14548_ (
);

FILL FILL_2__14128_ (
);

FILL FILL_0__15582_ (
);

FILL FILL_0__15162_ (
);

FILL SFILL28760x5050 (
);

FILL SFILL78760x35050 (
);

FILL FILL_3__8645_ (
);

DFFSR _12819_ (
    .Q(\control_1.op [2]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3490_[28])
);

FILL FILL_3__8225_ (
);

FILL FILL_1__14902_ (
);

FILL SFILL8680x1050 (
);

FILL FILL_4__12482_ (
);

FILL FILL_4__12062_ (
);

FILL FILL_5__9932_ (
);

FILL FILL_3__11895_ (
);

FILL FILL_5__9512_ (
);

FILL FILL_3__11475_ (
);

FILL FILL_3__11055_ (
);

FILL FILL_4__6988_ (
);

FILL FILL_0__16367_ (
);

NAND3X1 _16232_ (
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .B(_5500__bF$buf2),
    .C(_5471__bF$buf0),
    .Y(_6683_)
);

FILL FILL112360x47050 (
);

FILL FILL_2__10888_ (
);

FILL FILL_2__10048_ (
);

FILL FILL_0__11082_ (
);

FILL FILL_1__9924_ (
);

FILL FILL_5__11802_ (
);

FILL FILL_1__9504_ (
);

FILL SFILL64040x56050 (
);

FILL FILL_5__14694_ (
);

FILL FILL_0__6888_ (
);

FILL FILL_5__14274_ (
);

OAI21X1 _8994_ (
    .A(_1070_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1071_),
    .Y(_1043_[14])
);

OAI21X1 _8574_ (
    .A(_851_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .C(_852_),
    .Y(_848_[2])
);

DFFSR _8154_ (
    .Q(\datapath_1.regfile_1.regOut[10] [4]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_588_[4])
);

FILL FILL_1__10822_ (
);

FILL FILL_4__13687_ (
);

FILL FILL_4__13267_ (
);

FILL FILL_1__10402_ (
);

FILL FILL_2__7847_ (
);

FILL FILL_2__7427_ (
);

FILL FILL_1__13294_ (
);

OAI21X1 _12992_ (
    .A(_3645_),
    .B(vdd),
    .C(_3646_),
    .Y(_3620_[13])
);

OAI21X1 _12572_ (
    .A(_3426_),
    .B(vdd),
    .C(_3427_),
    .Y(_3425_[1])
);

FILL FILL_0__12287_ (
);

NAND2X1 _12152_ (
    .A(ALUSrcA_bF$buf2),
    .B(\datapath_1.a [12]),
    .Y(_3155_)
);

FILL FILL_3__13621_ (
);

FILL FILL_4__8714_ (
);

FILL FILL_5__15899_ (
);

FILL FILL_2__12614_ (
);

FILL FILL_5__15479_ (
);

FILL FILL_5__15059_ (
);

FILL FILL_3__16093_ (
);

NAND2X1 _9779_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1473_)
);

NAND2X1 _9359_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1254_)
);

FILL SFILL64040x11050 (
);

FILL FILL_5__10194_ (
);

FILL FILL_1__11607_ (
);

FILL FILL_2__15086_ (
);

FILL FILL_5__16000_ (
);

FILL FILL_0__8614_ (
);

FILL SFILL89240x60050 (
);

FILL FILL_1__14499_ (
);

FILL FILL_1__14079_ (
);

FILL FILL_4__15833_ (
);

FILL FILL_4__15413_ (
);

INVX1 _13777_ (
    .A(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_4283_)
);

NAND2X1 _13357_ (
    .A(\datapath_1.a3 [4]),
    .B(_3782_),
    .Y(_3873_)
);

FILL FILL_3__14826_ (
);

FILL FILL_1__15860_ (
);

FILL FILL_3__14406_ (
);

FILL SFILL18680x80050 (
);

FILL FILL_1__15440_ (
);

FILL FILL_1__15020_ (
);

FILL FILL_4__9919_ (
);

FILL FILL_2__13819_ (
);

CLKBUF1 CLKBUF1_insert1080 (
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1081 (
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

FILL FILL_0__14853_ (
);

FILL FILL_0__14433_ (
);

CLKBUF1 CLKBUF1_insert1082 (
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert1083 (
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

FILL FILL_0__14013_ (
);

FILL FILL_5__11399_ (
);

FILL SFILL54040x54050 (
);

FILL FILL_2__7180_ (
);

FILL FILL_5__12760_ (
);

FILL FILL_5__12340_ (
);

FILL FILL_4__11753_ (
);

FILL FILL_4__11333_ (
);

FILL FILL_1__16225_ (
);

FILL FILL_3__10746_ (
);

FILL FILL_1__11780_ (
);

FILL FILL_1__11360_ (
);

NOR2X1 _15923_ (
    .A(_6381_),
    .B(_6379_),
    .Y(_6382_)
);

FILL FILL_0__15638_ (
);

FILL FILL_0__15218_ (
);

AOI22X1 _15503_ (
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .B(_5579_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_5972_)
);

FILL FILL_0__10773_ (
);

FILL FILL_2__8385_ (
);

FILL FILL_5__13965_ (
);

FILL FILL_5__13545_ (
);

FILL FILL_5__13125_ (
);

OAI21X1 _7845_ (
    .A(_487_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_488_),
    .Y(_458_[15])
);

OAI21X1 _7425_ (
    .A(_268_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_269_),
    .Y(_263_[3])
);

DFFSR _7005_ (
    .Q(\datapath_1.regfile_1.regOut[1] [7]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf29),
    .S(vdd),
    .D(_3_[7])
);

FILL FILL_4_BUFX2_insert730 (
);

FILL FILL_4_BUFX2_insert731 (
);

FILL FILL_4__9672_ (
);

FILL FILL_4__9252_ (
);

FILL FILL_4_BUFX2_insert732 (
);

FILL FILL_4__12958_ (
);

FILL FILL_2__13992_ (
);

FILL FILL_4_BUFX2_insert733 (
);

FILL FILL_4_BUFX2_insert734 (
);

FILL FILL_4__12118_ (
);

FILL FILL_2__13572_ (
);

FILL FILL_2__13152_ (
);

FILL FILL_4_BUFX2_insert735 (
);

FILL FILL_4_BUFX2_insert736 (
);

FILL FILL_4_BUFX2_insert737 (
);

FILL FILL_4_BUFX2_insert738 (
);

FILL FILL_4_BUFX2_insert739 (
);

FILL FILL_1__12985_ (
);

FILL FILL111880x71050 (
);

FILL FILL_1__12145_ (
);

FILL FILL_0__9992_ (
);

FILL FILL_0__11978_ (
);

FILL FILL_0__9152_ (
);

OR2X2 _11843_ (
    .A(_2333_),
    .B(ALUControl[0]),
    .Y(_2931_)
);

FILL FILL_0__11558_ (
);

OAI21X1 _11423_ (
    .A(_2322_),
    .B(_2347__bF$buf0),
    .C(_2538_),
    .Y(_2539_)
);

FILL FILL_0__11138_ (
);

NAND2X1 _11003_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2122_)
);

FILL FILL_6__15337_ (
);

FILL FILL_5__7595_ (
);

FILL FILL_4__16371_ (
);

FILL FILL_5__7175_ (
);

FILL SFILL44040x52050 (
);

FILL FILL_3__15784_ (
);

FILL FILL_3__15364_ (
);

FILL FILL_1__7587_ (
);

FILL FILL_1__7167_ (
);

FILL FILL_2__14777_ (
);

FILL SFILL109000x70050 (
);

FILL FILL_2__14357_ (
);

FILL FILL_0__15391_ (
);

FILL SFILL109800x53050 (
);

FILL FILL_3__8874_ (
);

FILL FILL_3__8454_ (
);

NAND2X1 _12628_ (
    .A(vdd),
    .B(memoryOutData[20]),
    .Y(_3465_)
);

INVX1 _12208_ (
    .A(\datapath_1.PCJump [31]),
    .Y(_3192_)
);

FILL FILL_1__14711_ (
);

FILL FILL_6__11257_ (
);

FILL FILL_4__12291_ (
);

FILL FILL_0__13704_ (
);

FILL FILL_3__16149_ (
);

FILL FILL_2__6871_ (
);

FILL FILL_5__9741_ (
);

FILL FILL_3__11284_ (
);

FILL FILL_0__16176_ (
);

OAI22X1 _16041_ (
    .A(_6496_),
    .B(_5548__bF$buf0),
    .C(_5534__bF$buf4),
    .D(_5129_),
    .Y(_6497_)
);

FILL FILL_2__10697_ (
);

FILL FILL_2__10277_ (
);

FILL SFILL8440x29050 (
);

FILL FILL_1__9733_ (
);

FILL FILL_5__11611_ (
);

FILL FILL_3__9659_ (
);

FILL FILL_3_BUFX2_insert750 (
);

FILL FILL_3_BUFX2_insert751 (
);

FILL FILL_3__9239_ (
);

FILL FILL_3_BUFX2_insert752 (
);

FILL FILL_3_BUFX2_insert753 (
);

FILL FILL_3_BUFX2_insert754 (
);

FILL FILL_5__14083_ (
);

FILL FILL_1__15916_ (
);

FILL FILL_3_BUFX2_insert755 (
);

FILL FILL_6__7244_ (
);

NAND2X1 _8383_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_766_)
);

FILL FILL_3_BUFX2_insert756 (
);

FILL FILL_3_BUFX2_insert757 (
);

FILL FILL_3_BUFX2_insert758 (
);

FILL FILL_3_BUFX2_insert759 (
);

FILL FILL_4__13496_ (
);

FILL FILL_1__10631_ (
);

FILL SFILL69160x63050 (
);

FILL FILL_0__14909_ (
);

FILL FILL_2__7236_ (
);

FILL FILL_3__12489_ (
);

FILL FILL_3__12069_ (
);

FILL FILL_6__13403_ (
);

FILL SFILL74120x46050 (
);

OAI21X1 _12381_ (
    .A(_3318_),
    .B(MemToReg_bF$buf0),
    .C(_3319_),
    .Y(\datapath_1.mux_wd3.dout [12])
);

FILL FILL_0__12096_ (
);

FILL FILL_3__13850_ (
);

FILL FILL_3__13430_ (
);

FILL FILL_3__13010_ (
);

FILL SFILL38680x79050 (
);

FILL FILL_4__8523_ (
);

FILL FILL_4__8103_ (
);

FILL FILL_4__11809_ (
);

FILL FILL_2__12843_ (
);

FILL FILL_2__12423_ (
);

FILL FILL_5__15288_ (
);

FILL FILL_2__12003_ (
);

FILL FILL_6__8449_ (
);

DFFSR _9588_ (
    .Q(\datapath_1.regfile_1.regOut[21] [30]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_1303_[30])
);

INVX1 _9168_ (
    .A(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_1167_)
);

FILL FILL_1__11836_ (
);

FILL FILL_1__11416_ (
);

FILL FILL_0__8843_ (
);

FILL FILL_3__6940_ (
);

FILL FILL_0__10829_ (
);

FILL FILL_0__10409_ (
);

FILL FILL_0__8003_ (
);

FILL FILL_5__6866_ (
);

FILL FILL_0_BUFX2_insert880 (
);

FILL FILL_4__15642_ (
);

FILL FILL_0_BUFX2_insert881 (
);

FILL FILL_4__15222_ (
);

FILL FILL_0_BUFX2_insert882 (
);

FILL FILL_0_BUFX2_insert883 (
);

FILL FILL_0_BUFX2_insert884 (
);

INVX1 _13586_ (
    .A(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_4095_)
);

FILL FILL_0_BUFX2_insert885 (
);

INVX1 _13166_ (
    .A(\datapath_1.PCJump [29]),
    .Y(_3742_)
);

FILL FILL_0_BUFX2_insert886 (
);

FILL FILL_0_BUFX2_insert887 (
);

FILL FILL_2__9802_ (
);

FILL FILL_3__14635_ (
);

FILL FILL_0_BUFX2_insert888 (
);

FILL FILL_3__14215_ (
);

FILL FILL_0_BUFX2_insert889 (
);

FILL FILL_1__6858_ (
);

FILL FILL_4__9728_ (
);

FILL FILL_2__13628_ (
);

FILL FILL_2__13208_ (
);

FILL FILL_0__14662_ (
);

FILL SFILL99320x50050 (
);

FILL FILL_0__14242_ (
);

FILL FILL_0__9628_ (
);

FILL FILL_3__7725_ (
);

FILL SFILL28760x70050 (
);

FILL FILL_3__7305_ (
);

FILL FILL_0__9208_ (
);

FILL FILL_4__16007_ (
);

FILL FILL_4__11982_ (
);

FILL FILL_4__11562_ (
);

FILL FILL_4__11142_ (
);

FILL SFILL64120x44050 (
);

FILL FILL_1__16034_ (
);

FILL FILL_3__10975_ (
);

FILL FILL_3__10555_ (
);

FILL FILL_6_BUFX2_insert260 (
);

FILL FILL_3__10135_ (
);

FILL FILL_0__15867_ (
);

AOI21X1 _15732_ (
    .A(_6170_),
    .B(_6195_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [16])
);

FILL FILL_0__15447_ (
);

NAND2X1 _15312_ (
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .B(_5785_),
    .Y(_5786_)
);

FILL FILL_0__15027_ (
);

FILL FILL_6_BUFX2_insert265 (
);

FILL FILL_2__8194_ (
);

FILL FILL_0__10162_ (
);

BUFX2 BUFX2_insert40 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf1 )
);

BUFX2 BUFX2_insert41 (
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf0 )
);

BUFX2 BUFX2_insert42 (
    .A(_5466_),
    .Y(_5466__bF$buf4)
);

BUFX2 BUFX2_insert43 (
    .A(_5466_),
    .Y(_5466__bF$buf3)
);

BUFX2 BUFX2_insert44 (
    .A(_5466_),
    .Y(_5466__bF$buf2)
);

BUFX2 BUFX2_insert45 (
    .A(_5466_),
    .Y(_5466__bF$buf1)
);

BUFX2 BUFX2_insert46 (
    .A(_5466_),
    .Y(_5466__bF$buf0)
);

FILL FILL_5__13774_ (
);

BUFX2 BUFX2_insert47 (
    .A(_3893_),
    .Y(_3893__bF$buf3)
);

FILL FILL_5__13354_ (
);

BUFX2 BUFX2_insert48 (
    .A(_3893_),
    .Y(_3893__bF$buf2)
);

BUFX2 BUFX2_insert49 (
    .A(_3893_),
    .Y(_3893__bF$buf1)
);

DFFSR _7654_ (
    .Q(\datapath_1.regfile_1.regOut[6] [16]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_328_[16])
);

NAND2X1 _7234_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_183_)
);

FILL FILL_4__9481_ (
);

FILL FILL_4__12767_ (
);

FILL FILL_4__12347_ (
);

FILL FILL_2__13381_ (
);

FILL FILL_2__6927_ (
);

FILL FILL_1__12374_ (
);

FILL FILL_0__9381_ (
);

FILL FILL_2__9399_ (
);

FILL FILL_0__11787_ (
);

FILL FILL_0__11367_ (
);

INVX1 _11652_ (
    .A(_2382_),
    .Y(_2755_)
);

AND2X2 _11232_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2351_)
);

FILL FILL_6__15986_ (
);

FILL FILL_3__12701_ (
);

FILL FILL_4__16180_ (
);

FILL FILL_5__14979_ (
);

FILL FILL_5__14559_ (
);

FILL FILL_5__14139_ (
);

FILL FILL_3__15593_ (
);

FILL FILL_3__15173_ (
);

NAND2X1 _8859_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1002_)
);

NAND2X1 _8439_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .Y(_847_)
);

INVX1 _8019_ (
    .A(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_584_)
);

FILL FILL_2__14586_ (
);

FILL FILL_2__14166_ (
);

FILL FILL_5__15920_ (
);

FILL FILL_5__15500_ (
);

FILL FILL_1__13999_ (
);

NAND2X1 _9800_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1487_)
);

FILL SFILL54120x42050 (
);

FILL FILL_1__13579_ (
);

FILL FILL_1__13159_ (
);

FILL FILL_4__14913_ (
);

NAND2X1 _12857_ (
    .A(vdd),
    .B(\datapath_1.rd1 [11]),
    .Y(_3577_)
);

FILL FILL_3__8263_ (
);

NAND2X1 _12437_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [31]),
    .Y(_3357_)
);

AOI22X1 _12017_ (
    .A(\datapath_1.ALUResult [7]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3059_)
);

FILL FILL_3__13906_ (
);

FILL SFILL18680x75050 (
);

FILL FILL_1__14940_ (
);

FILL FILL_1__14520_ (
);

FILL FILL_5__8189_ (
);

FILL FILL_1__14100_ (
);

FILL FILL_5_BUFX2_insert280 (
);

FILL FILL_5_BUFX2_insert281 (
);

FILL FILL_5_BUFX2_insert282 (
);

FILL FILL_0__13933_ (
);

FILL FILL_5_BUFX2_insert283 (
);

FILL FILL_3__16378_ (
);

FILL FILL_0__13513_ (
);

FILL FILL_5_BUFX2_insert284 (
);

FILL FILL_5__10899_ (
);

FILL FILL_5_BUFX2_insert285 (
);

FILL SFILL54040x49050 (
);

FILL FILL_5_BUFX2_insert286 (
);

FILL FILL_5__9550_ (
);

FILL FILL_5__10059_ (
);

FILL FILL_5_BUFX2_insert287 (
);

FILL FILL_5_BUFX2_insert1070 (
);

FILL FILL_5_BUFX2_insert1071 (
);

FILL FILL_5_BUFX2_insert288 (
);

FILL FILL_5__9130_ (
);

FILL FILL_3__11093_ (
);

FILL FILL_5_BUFX2_insert1072 (
);

FILL FILL_5_BUFX2_insert289 (
);

FILL FILL_5_BUFX2_insert1073 (
);

INVX1 _16270_ (
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_6720_)
);

FILL FILL_5__11840_ (
);

FILL FILL_1__9542_ (
);

FILL FILL_5__11420_ (
);

FILL FILL_1__9122_ (
);

FILL FILL_5__11000_ (
);

FILL FILL_3__9888_ (
);

FILL FILL_2__16312_ (
);

FILL FILL_3__9468_ (
);

FILL FILL_4__10833_ (
);

FILL FILL_4__10413_ (
);

FILL FILL_1__15725_ (
);

NAND2X1 _8192_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_659_)
);

FILL FILL_6__7053_ (
);

FILL FILL_1__15305_ (
);

FILL SFILL18680x30050 (
);

FILL FILL_1__10440_ (
);

FILL FILL_1__10020_ (
);

FILL FILL_0__14718_ (
);

FILL FILL_2__7885_ (
);

FILL FILL_2__7465_ (
);

FILL FILL_3__12298_ (
);

FILL FILL_2__7045_ (
);

INVX1 _12190_ (
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3180_)
);

FILL FILL_5__12625_ (
);

FILL FILL_5__12205_ (
);

OAI21X1 _6925_ (
    .A(_16_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .C(_17_),
    .Y(_3_[7])
);

FILL SFILL79240x53050 (
);

FILL FILL_4__8752_ (
);

FILL FILL_4__8332_ (
);

FILL FILL_4__11618_ (
);

FILL FILL_2__12652_ (
);

FILL FILL_5__15097_ (
);

FILL FILL_2__12232_ (
);

INVX1 _9397_ (
    .A(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_1279_)
);

FILL FILL111880x66050 (
);

FILL FILL_1__11645_ (
);

FILL FILL_1__11225_ (
);

FILL FILL_0__8652_ (
);

FILL FILL_0__10638_ (
);

NOR2X1 _10923_ (
    .A(_2049_),
    .B(_2053_),
    .Y(_0_)
);

FILL FILL_0__8232_ (
);

OAI21X1 _10503_ (
    .A(_1832_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1833_),
    .Y(_1823_[5])
);

FILL SFILL109400x79050 (
);

FILL FILL_4__15871_ (
);

FILL FILL_4__15451_ (
);

FILL FILL_4__15031_ (
);

INVX1 _13395_ (
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_3907_)
);

FILL FILL_3__14864_ (
);

FILL FILL_2__9611_ (
);

FILL FILL_3__14444_ (
);

FILL FILL_3__14024_ (
);

FILL FILL112200x7050 (
);

FILL FILL_4__9537_ (
);

FILL FILL_4__9117_ (
);

FILL FILL_2__13857_ (
);

FILL FILL_2__13437_ (
);

FILL FILL_0__14891_ (
);

FILL FILL_0__14471_ (
);

FILL FILL_2__13017_ (
);

FILL FILL_0__14051_ (
);

FILL FILL111880x21050 (
);

FILL FILL_0__9857_ (
);

FILL FILL_3__7954_ (
);

FILL FILL_3__7114_ (
);

FILL FILL_0__9017_ (
);

OAI21X1 _11708_ (
    .A(_2341__bF$buf1),
    .B(_2393_),
    .C(_2806_),
    .Y(_2807_)
);

FILL FILL_4__16236_ (
);

FILL SFILL109400x34050 (
);

FILL SFILL48760x24050 (
);

FILL FILL_4__11791_ (
);

FILL FILL_4__11371_ (
);

FILL FILL_3__15649_ (
);

FILL FILL_3__15229_ (
);

FILL FILL_1__16263_ (
);

FILL FILL_3__10784_ (
);

FILL FILL_5__8401_ (
);

FILL FILL_3__10364_ (
);

FILL FILL_0__15676_ (
);

OAI22X1 _15961_ (
    .A(_5534__bF$buf0),
    .B(_5021_),
    .C(_5532__bF$buf3),
    .D(_6418_),
    .Y(_6419_)
);

FILL SFILL69240x51050 (
);

FILL FILL_0__15256_ (
);

NOR2X1 _15541_ (
    .A(_6007_),
    .B(_6008_),
    .Y(_6009_)
);

OAI21X1 _15121_ (
    .A(_4027_),
    .B(_5535__bF$buf1),
    .C(_5599_),
    .Y(_5600_)
);

FILL FILL_0__10391_ (
);

FILL FILL_6__14590_ (
);

FILL FILL_6__14170_ (
);

FILL FILL_3__8739_ (
);

FILL FILL_3__8319_ (
);

FILL FILL_5__13583_ (
);

FILL FILL_5__13163_ (
);

NAND2X1 _7883_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_514_)
);

NAND2X1 _7463_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_295_)
);

NAND2X1 _7043_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_76_)
);

FILL SFILL99400x83050 (
);

FILL FILL_4__12996_ (
);

FILL FILL_4__9290_ (
);

FILL FILL_4__12576_ (
);

FILL SFILL69160x58050 (
);

FILL SFILL69640x20050 (
);

FILL FILL_4__12156_ (
);

FILL FILL_3__11989_ (
);

FILL FILL_3__11569_ (
);

FILL FILL_5__9606_ (
);

FILL FILL_3__11149_ (
);

FILL FILL_1__12183_ (
);

FILL FILL_6__12903_ (
);

OAI21X1 _16326_ (
    .A(_6770_),
    .B(gnd),
    .C(_6771_),
    .Y(_6769_[1])
);

INVX1 _11881_ (
    .A(\datapath_1.PCJump [21]),
    .Y(_2964_)
);

FILL FILL_0__11596_ (
);

FILL FILL_0__11176_ (
);

NAND3X1 _11461_ (
    .A(_2438_),
    .B(_2573_),
    .C(_2575_),
    .Y(_2576_)
);

OAI21X1 _11041_ (
    .A(_2153_),
    .B(_2140_),
    .C(_2159_),
    .Y(_2160_)
);

FILL FILL_3__12510_ (
);

FILL FILL_4__7603_ (
);

FILL FILL_2__11923_ (
);

FILL FILL_5__14788_ (
);

FILL FILL_5__14368_ (
);

FILL FILL_2__11503_ (
);

DFFSR _8668_ (
    .Q(\datapath_1.regfile_1.regOut[14] [6]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_848_[6])
);

INVX1 _8248_ (
    .A(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_696_)
);

FILL FILL_1__10916_ (
);

FILL FILL_2__14395_ (
);

FILL SFILL69160x13050 (
);

FILL FILL_0__7503_ (
);

FILL FILL_1__13388_ (
);

FILL FILL_4__14722_ (
);

FILL FILL_4__14302_ (
);

FILL FILL_3__8492_ (
);

FILL SFILL93640x24050 (
);

DFFSR _12666_ (
    .Q(\datapath_1.Data [3]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3425_[3])
);

FILL FILL_3__8072_ (
);

NAND3X1 _12246_ (
    .A(_3221_),
    .B(_3222_),
    .C(_3223_),
    .Y(\datapath_1.alu_1.ALUInB [7])
);

FILL FILL_3__13715_ (
);

FILL FILL_2__12708_ (
);

FILL FILL_0__13742_ (
);

FILL FILL_0__13322_ (
);

FILL FILL_3__16187_ (
);

FILL FILL_5__10288_ (
);

FILL SFILL89400x81050 (
);

FILL FILL_0__8708_ (
);

FILL SFILL59160x56050 (
);

FILL FILL_1__9771_ (
);

FILL FILL_1__9351_ (
);

FILL SFILL38280x15050 (
);

FILL FILL_4__15927_ (
);

FILL FILL_4__15507_ (
);

FILL FILL_2__16121_ (
);

FILL FILL_3__9277_ (
);

FILL FILL_4__10642_ (
);

FILL SFILL64120x39050 (
);

FILL FILL_1__15954_ (
);

FILL FILL_1__15534_ (
);

FILL FILL_1__15114_ (
);

FILL FILL_0__14947_ (
);

NOR2X1 _14812_ (
    .A(_5285_),
    .B(_5295_),
    .Y(_5296_)
);

FILL FILL_0__14527_ (
);

FILL FILL_0__14107_ (
);

FILL FILL_2__7694_ (
);

FILL FILL_5__12854_ (
);

FILL FILL_5__12434_ (
);

FILL FILL_5__12014_ (
);

FILL SFILL59160x11050 (
);

FILL SFILL84200x6050 (
);

FILL FILL_4__8981_ (
);

FILL FILL_4__8141_ (
);

FILL FILL_4__11847_ (
);

FILL FILL_2__12881_ (
);

FILL FILL_4__11427_ (
);

FILL FILL_2__12461_ (
);

FILL FILL_4__11007_ (
);

FILL FILL_2__12041_ (
);

FILL FILL_6__8067_ (
);

FILL FILL_1__16319_ (
);

FILL FILL_1__11874_ (
);

FILL FILL_1__11454_ (
);

FILL FILL_1__11034_ (
);

FILL SFILL33960x83050 (
);

FILL SFILL49560x68050 (
);

FILL FILL_0__8881_ (
);

FILL FILL_2__8899_ (
);

FILL FILL_0__8461_ (
);

FILL FILL_2__8479_ (
);

FILL FILL_0__10447_ (
);

DFFSR _10732_ (
    .Q(\datapath_1.regfile_1.regOut[30] [22]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1888_[22])
);

FILL FILL_2__8059_ (
);

FILL SFILL89320x43050 (
);

NAND2X1 _10312_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1747_)
);

FILL FILL_0__10027_ (
);

FILL FILL_6__14646_ (
);

FILL FILL_4__15680_ (
);

FILL FILL_4__15260_ (
);

FILL FILL_5__13639_ (
);

FILL FILL_5__13219_ (
);

FILL FILL_2__9420_ (
);

FILL FILL_3__14673_ (
);

FILL FILL_2__9000_ (
);

FILL FILL_3__14253_ (
);

NAND2X1 _7939_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_531_)
);

FILL SFILL18760x63050 (
);

DFFSR _7519_ (
    .Q(\datapath_1.regfile_1.regOut[5] [9]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_263_[9])
);

FILL FILL_1__6896_ (
);

FILL FILL_4__9766_ (
);

FILL FILL_4__9346_ (
);

FILL FILL_2__13666_ (
);

FILL FILL_2__13246_ (
);

FILL FILL_0__14280_ (
);

FILL FILL_1__12659_ (
);

FILL FILL_1__12239_ (
);

FILL FILL_3__7763_ (
);

FILL FILL_0__9666_ (
);

OAI21X1 _11937_ (
    .A(_2998_),
    .B(IorD_bF$buf0),
    .C(_2999_),
    .Y(_1_[16])
);

FILL FILL_3__7343_ (
);

FILL FILL_0__9246_ (
);

INVX1 _11517_ (
    .A(_2280_),
    .Y(_2628_)
);

FILL FILL_5__7689_ (
);

FILL FILL_1__13600_ (
);

FILL FILL_4__16045_ (
);

FILL FILL_4__11180_ (
);

FILL FILL_3__15878_ (
);

FILL FILL_3__15458_ (
);

FILL FILL_3__15038_ (
);

FILL FILL_1__16072_ (
);

FILL FILL_5__8630_ (
);

FILL FILL_3__10173_ (
);

FILL FILL_5__8210_ (
);

FILL FILL_6_BUFX2_insert643 (
);

AOI21X1 _15770_ (
    .A(_6209_),
    .B(_6232_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [17])
);

FILL FILL_0__15485_ (
);

AOI22X1 _15350_ (
    .A(_5565__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [7]),
    .C(\datapath_1.regfile_1.regOut[5] [7]),
    .D(_5700_),
    .Y(_5823_)
);

FILL FILL_0__15065_ (
);

FILL FILL_6_BUFX2_insert648 (
);

FILL FILL_5__10920_ (
);

FILL FILL_5__10500_ (
);

FILL FILL_1__8622_ (
);

FILL FILL_1__8202_ (
);

FILL FILL_2__15812_ (
);

FILL FILL_3__8968_ (
);

FILL FILL_3__8128_ (
);

FILL FILL_5__13392_ (
);

NAND2X1 _7692_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_407_)
);

FILL FILL_1__14805_ (
);

DFFSR _7272_ (
    .Q(\datapath_1.regfile_1.regOut[3] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_133_[18])
);

FILL SFILL79320x41050 (
);

FILL SFILL18680x25050 (
);

FILL FILL_4__12385_ (
);

FILL FILL_2__6965_ (
);

FILL FILL_3__11798_ (
);

FILL FILL_5__9415_ (
);

FILL FILL_3__11378_ (
);

FILL FILL_6__12712_ (
);

FILL SFILL39160x52050 (
);

INVX1 _16135_ (
    .A(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_6588_)
);

INVX1 _11690_ (
    .A(_2790_),
    .Y(\datapath_1.ALUResult [13])
);

NOR2X1 _11270_ (
    .A(_2197_),
    .B(_2388_),
    .Y(_2389_)
);

FILL FILL_5__11705_ (
);

FILL FILL_1__9407_ (
);

FILL SFILL79240x48050 (
);

FILL FILL_4__7832_ (
);

FILL FILL_5__14597_ (
);

FILL FILL_2__11732_ (
);

FILL FILL_5__14177_ (
);

FILL FILL_2__11312_ (
);

INVX1 _8897_ (
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_1027_)
);

INVX1 _8477_ (
    .A(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_808_)
);

INVX1 _8057_ (
    .A(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_589_)
);

FILL FILL_1__10305_ (
);

FILL SFILL54200x5050 (
);

FILL FILL_0__7732_ (
);

FILL FILL_0__7312_ (
);

FILL SFILL94440x3050 (
);

FILL FILL_4__14951_ (
);

FILL FILL_4__14531_ (
);

FILL SFILL94360x8050 (
);

FILL FILL_4__14111_ (
);

INVX1 _12895_ (
    .A(\datapath_1.a [24]),
    .Y(_3602_)
);

INVX1 _12475_ (
    .A(ALUOut[12]),
    .Y(_3383_)
);

NAND3X1 _12055_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[17]),
    .C(_3032__bF$buf1),
    .Y(_3087_)
);

FILL FILL_3__13944_ (
);

FILL FILL_3__13524_ (
);

FILL FILL_3__13104_ (
);

FILL FILL_4__8617_ (
);

FILL FILL_5_BUFX2_insert660 (
);

FILL FILL_5_BUFX2_insert661 (
);

FILL FILL_2__12517_ (
);

FILL FILL_0__13971_ (
);

FILL FILL_5_BUFX2_insert662 (
);

FILL FILL_5_BUFX2_insert663 (
);

FILL FILL_0__13551_ (
);

FILL FILL_0__13131_ (
);

FILL FILL_5_BUFX2_insert664 (
);

FILL FILL_5_BUFX2_insert665 (
);

FILL FILL_5_BUFX2_insert666 (
);

FILL FILL_5_BUFX2_insert667 (
);

FILL FILL_5_BUFX2_insert668 (
);

FILL FILL_5_BUFX2_insert669 (
);

FILL SFILL104600x6050 (
);

FILL FILL_5__16323_ (
);

FILL FILL_0__8517_ (
);

FILL FILL_1__9160_ (
);

FILL FILL_4__15736_ (
);

FILL FILL_4__15316_ (
);

FILL SFILL109400x29050 (
);

FILL FILL_2__16350_ (
);

FILL FILL_4__10871_ (
);

FILL FILL_3__9086_ (
);

FILL FILL_4__10451_ (
);

FILL FILL_4__10031_ (
);

FILL FILL_3__14729_ (
);

FILL FILL_1__15763_ (
);

FILL FILL_3__14309_ (
);

FILL FILL_1__15343_ (
);

FILL SFILL69240x46050 (
);

FILL FILL_0__14756_ (
);

OAI22X1 _14621_ (
    .A(_3947__bF$buf3),
    .B(_5108_),
    .C(_3909_),
    .D(_5107_),
    .Y(_5109_)
);

FILL FILL_0__14336_ (
);

INVX1 _14201_ (
    .A(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_4698_)
);

FILL FILL_2__7083_ (
);

FILL FILL_3__7819_ (
);

FILL FILL_5__12243_ (
);

NAND2X1 _6963_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_43_)
);

FILL FILL_2_BUFX2_insert790 (
);

FILL FILL_2_BUFX2_insert791 (
);

FILL SFILL99400x78050 (
);

FILL FILL_2_BUFX2_insert792 (
);

FILL FILL_2_BUFX2_insert793 (
);

FILL FILL_4__8370_ (
);

FILL FILL_2_BUFX2_insert794 (
);

FILL FILL_4__11656_ (
);

FILL FILL_2_BUFX2_insert795 (
);

FILL FILL_4__11236_ (
);

FILL FILL_2__12270_ (
);

FILL FILL_2_BUFX2_insert796 (
);

FILL FILL_2_BUFX2_insert797 (
);

FILL FILL_2_BUFX2_insert798 (
);

FILL FILL_2_BUFX2_insert799 (
);

FILL FILL_1__16128_ (
);

FILL FILL_3__10649_ (
);

FILL FILL_1__11683_ (
);

FILL FILL_1__11263_ (
);

INVX1 _15826_ (
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_6287_)
);

INVX1 _15406_ (
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_5878_)
);

NOR2X1 _10961_ (
    .A(\control_1.op [0]),
    .B(_2092_),
    .Y(_2093_)
);

FILL FILL_0__8270_ (
);

FILL FILL_0__10676_ (
);

FILL SFILL104360x71050 (
);

FILL FILL_0__10256_ (
);

NAND2X1 _10541_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1859_)
);

NAND2X1 _10121_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1640_)
);

FILL FILL_5__13868_ (
);

FILL FILL_5__13448_ (
);

FILL SFILL3800x66050 (
);

FILL FILL_3__14482_ (
);

FILL FILL_5__13028_ (
);

FILL FILL_3__14062_ (
);

INVX1 _7748_ (
    .A(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_444_)
);

INVX1 _7328_ (
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_225_)
);

FILL FILL_4__9995_ (
);

FILL FILL_4__9155_ (
);

FILL FILL_2__13895_ (
);

FILL FILL_2__13475_ (
);

FILL SFILL99400x33050 (
);

FILL FILL_1__12888_ (
);

FILL FILL_1__12468_ (
);

FILL FILL_1__12048_ (
);

FILL FILL_4__13802_ (
);

FILL FILL_0__9895_ (
);

FILL FILL_3__7992_ (
);

FILL FILL_0__9475_ (
);

FILL FILL_3__7572_ (
);

NAND2X1 _11746_ (
    .A(_2389_),
    .B(_2481__bF$buf0),
    .Y(_2842_)
);

INVX1 _11326_ (
    .A(_2444_),
    .Y(_2445_)
);

FILL FILL_5__7498_ (
);

FILL FILL_5__7078_ (
);

FILL FILL_4__16274_ (
);

FILL FILL_3__15687_ (
);

FILL FILL_0__12402_ (
);

FILL FILL_3__15267_ (
);

FILL FILL_0__15294_ (
);

FILL SFILL89400x76050 (
);

FILL SFILL64040x1050 (
);

FILL FILL_1__8851_ (
);

FILL FILL_1__8011_ (
);

FILL FILL_2__15621_ (
);

FILL FILL_2__15201_ (
);

FILL FILL_3__8777_ (
);

FILL FILL_3__8357_ (
);

FILL FILL_1__14614_ (
);

INVX1 _7081_ (
    .A(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_101_)
);

FILL SFILL115080x5050 (
);

FILL FILL_4__12194_ (
);

FILL FILL_0__13607_ (
);

FILL FILL_5__9644_ (
);

FILL FILL_5__9224_ (
);

FILL FILL_3__11187_ (
);

FILL FILL_6__12101_ (
);

NAND2X1 _16364_ (
    .A(gnd),
    .B(gnd),
    .Y(_6797_)
);

FILL FILL_0__16079_ (
);

FILL FILL_5__11934_ (
);

FILL SFILL89400x31050 (
);

FILL FILL_1__9636_ (
);

FILL FILL_5__11514_ (
);

FILL SFILL28760x15050 (
);

FILL FILL_1__9216_ (
);

FILL SFILL94280x82050 (
);

FILL FILL_2__16406_ (
);

FILL FILL_4__7221_ (
);

FILL FILL_4__10927_ (
);

FILL FILL_4__10507_ (
);

FILL FILL_2__11961_ (
);

FILL FILL_2__11541_ (
);

FILL FILL_2__11121_ (
);

FILL FILL_1__15819_ (
);

DFFSR _8286_ (
    .Q(\datapath_1.regfile_1.regOut[11] [8]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_653_[8])
);

FILL SFILL113720x4050 (
);

FILL SFILL49240x42050 (
);

FILL FILL_1__10954_ (
);

FILL FILL_1__10534_ (
);

FILL FILL_4__13399_ (
);

FILL FILL_1__10114_ (
);

FILL SFILL33960x78050 (
);

FILL FILL_0__7961_ (
);

FILL FILL_2__7979_ (
);

BUFX2 BUFX2_insert480 (
    .A(_5459_),
    .Y(_5459__bF$buf3)
);

FILL FILL_2__7559_ (
);

FILL SFILL89320x38050 (
);

BUFX2 BUFX2_insert481 (
    .A(_5459_),
    .Y(_5459__bF$buf2)
);

FILL FILL_0__7121_ (
);

BUFX2 BUFX2_insert482 (
    .A(_5459_),
    .Y(_5459__bF$buf1)
);

BUFX2 BUFX2_insert483 (
    .A(_5459_),
    .Y(_5459__bF$buf0)
);

BUFX2 BUFX2_insert484 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf4 )
);

FILL FILL_6__13306_ (
);

FILL FILL_4__14760_ (
);

BUFX2 BUFX2_insert485 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf3 )
);

FILL FILL_4__14340_ (
);

BUFX2 BUFX2_insert486 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf2 )
);

BUFX2 BUFX2_insert487 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf1 )
);

BUFX2 BUFX2_insert488 (
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf0 )
);

BUFX2 BUFX2_insert489 (
    .A(_3983_),
    .Y(_3983__bF$buf4)
);

FILL SFILL33880x50 (
);

NAND3X1 _12284_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf4),
    .Y(_3252_)
);

FILL FILL_5__12719_ (
);

FILL FILL_3__13753_ (
);

FILL FILL_2__8500_ (
);

FILL SFILL94200x80050 (
);

FILL SFILL18760x58050 (
);

FILL FILL_3__13333_ (
);

FILL FILL_4__8846_ (
);

FILL FILL_4__8006_ (
);

FILL FILL_2__12746_ (
);

FILL FILL_0__13780_ (
);

FILL FILL_2__12326_ (
);

FILL FILL_0__13360_ (
);

FILL FILL_1__11739_ (
);

FILL FILL_1__11319_ (
);

FILL SFILL33160x50050 (
);

FILL FILL_3__6843_ (
);

FILL FILL_0__8746_ (
);

FILL FILL_5__16132_ (
);

FILL FILL_0__8326_ (
);

FILL SFILL33960x33050 (
);

FILL FILL_4__15965_ (
);

FILL FILL_4__15545_ (
);

FILL FILL_4__15125_ (
);

FILL FILL_4__10680_ (
);

NAND3X1 _13489_ (
    .A(_3996_),
    .B(_3999_),
    .C(_3994_),
    .Y(_4000_)
);

DFFSR _13069_ (
    .Q(_2_[22]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3620_[22])
);

FILL FILL_4__10260_ (
);

FILL FILL_3__14958_ (
);

FILL FILL_1__15992_ (
);

FILL FILL_3__14538_ (
);

FILL FILL_1__15572_ (
);

FILL FILL_3__14118_ (
);

FILL FILL_1__15152_ (
);

FILL FILL_5__7710_ (
);

FILL SFILL18760x13050 (
);

FILL SFILL84280x80050 (
);

FILL FILL_0__14985_ (
);

FILL FILL_0__14565_ (
);

AOI21X1 _14850_ (
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .B(_4225_),
    .C(_5332_),
    .Y(_5333_)
);

FILL FILL_0__14145_ (
);

NOR2X1 _14430_ (
    .A(_4921_),
    .B(_4918_),
    .Y(_4922_)
);

OAI22X1 _14010_ (
    .A(_4510_),
    .B(_3905__bF$buf2),
    .C(_3954__bF$buf3),
    .D(_4509_),
    .Y(_4511_)
);

FILL FILL_1__7702_ (
);

FILL FILL_3__7628_ (
);

FILL FILL_3__7208_ (
);

FILL FILL_5__12892_ (
);

FILL FILL_5__12472_ (
);

FILL FILL_5__12052_ (
);

FILL SFILL59000x7050 (
);

FILL FILL_4__11885_ (
);

FILL FILL_4__11465_ (
);

FILL FILL_4__11045_ (
);

FILL FILL_1__16357_ (
);

FILL FILL_3__10878_ (
);

FILL FILL_5__8915_ (
);

FILL FILL111960x49050 (
);

FILL FILL_3__10038_ (
);

FILL FILL_1__11492_ (
);

FILL FILL_1__11072_ (
);

INVX1 _15635_ (
    .A(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_6101_)
);

NOR3X1 _15215_ (
    .A(_5687_),
    .B(_5689_),
    .C(_5690_),
    .Y(_5691_)
);

FILL FILL_2__8097_ (
);

NAND2X1 _10770_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1971_)
);

DFFSR _10350_ (
    .Q(\datapath_1.regfile_1.regOut[27] [24]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_1693_[24])
);

FILL FILL_0__10065_ (
);

FILL FILL_1__8907_ (
);

FILL FILL_4__6912_ (
);

FILL FILL_2__10812_ (
);

FILL FILL_5__13677_ (
);

FILL FILL_5__13257_ (
);

FILL FILL_3__14291_ (
);

INVX1 _7977_ (
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_556_)
);

INVX1 _7557_ (
    .A(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_337_)
);

DFFSR _7137_ (
    .Q(\datapath_1.regfile_1.regOut[2] [11]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_68_[11])
);

FILL FILL_4__9384_ (
);

FILL FILL_2__13284_ (
);

FILL SFILL114440x61050 (
);

FILL FILL_1__12697_ (
);

FILL FILL_1__12277_ (
);

FILL FILL_4__13611_ (
);

NAND2X1 _11975_ (
    .A(IorD_bF$buf2),
    .B(ALUOut[29]),
    .Y(_3025_)
);

FILL FILL_0__9284_ (
);

FILL FILL_3__7381_ (
);

NOR2X1 _11555_ (
    .A(_2230_),
    .B(_2347__bF$buf0),
    .Y(_2664_)
);

INVX2 _11135_ (
    .A(\datapath_1.alu_1.ALUInA [16]),
    .Y(_2254_)
);

FILL FILL_6__15889_ (
);

FILL FILL_3__12604_ (
);

FILL FILL_4__16083_ (
);

FILL FILL_0__12631_ (
);

FILL FILL_3__15496_ (
);

FILL FILL_3__15076_ (
);

FILL FILL_0__12211_ (
);

FILL FILL_1__7299_ (
);

FILL FILL_2__14489_ (
);

FILL FILL_2__14069_ (
);

FILL FILL_5__15823_ (
);

FILL FILL_5__15403_ (
);

DFFSR _9703_ (
    .Q(\datapath_1.regfile_1.regOut[22] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_1368_[17])
);

FILL FILL_1__8660_ (
);

FILL FILL_1__8240_ (
);

FILL FILL_4__14816_ (
);

FILL SFILL93800x45050 (
);

FILL FILL_2__15850_ (
);

FILL FILL_2__15430_ (
);

FILL FILL_3__8586_ (
);

FILL FILL_2__15010_ (
);

FILL FILL_3__13809_ (
);

FILL FILL_1__14843_ (
);

FILL FILL_1__14423_ (
);

FILL FILL_1__14003_ (
);

FILL FILL_0__13836_ (
);

FILL FILL_0__13416_ (
);

OAI22X1 _13701_ (
    .A(_3967__bF$buf1),
    .B(_4207_),
    .C(_3944__bF$buf4),
    .D(_4206_),
    .Y(_4208_)
);

FILL FILL_5__9873_ (
);

FILL FILL_5__9033_ (
);

INVX1 _16173_ (
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_6625_)
);

FILL FILL_1__9865_ (
);

FILL FILL_5__11743_ (
);

FILL FILL_5__11323_ (
);

FILL FILL_1__9025_ (
);

FILL FILL_4__7870_ (
);

FILL FILL_2__16215_ (
);

FILL FILL_4__7450_ (
);

FILL FILL_4__7030_ (
);

FILL FILL_4__10316_ (
);

FILL FILL_2__11770_ (
);

FILL FILL_2__11350_ (
);

FILL FILL_1__15628_ (
);

FILL FILL_1__15208_ (
);

OAI21X1 _8095_ (
    .A(_613_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_614_),
    .Y(_588_[13])
);

FILL FILL_1__10763_ (
);

FILL SFILL59720x46050 (
);

NAND2X1 _14906_ (
    .A(_5380_),
    .B(_5387_),
    .Y(_5388_)
);

FILL SFILL104360x66050 (
);

FILL FILL_0__7350_ (
);

FILL FILL_2__7368_ (
);

FILL FILL_6__13955_ (
);

FILL FILL_6__13115_ (
);

FILL SFILL69160x9050 (
);

FILL SFILL43880x5050 (
);

AOI22X1 _12093_ (
    .A(\datapath_1.ALUResult [26]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3116_)
);

FILL FILL_5__12528_ (
);

FILL FILL_3__13982_ (
);

FILL FILL_5__12108_ (
);

FILL FILL_3__13562_ (
);

FILL FILL_3__13142_ (
);

FILL FILL_4__8655_ (
);

FILL SFILL8600x5050 (
);

FILL FILL_4__8235_ (
);

FILL FILL_2__12975_ (
);

FILL SFILL99400x28050 (
);

FILL FILL_2__12135_ (
);

FILL FILL_1__11968_ (
);

FILL FILL_1__11548_ (
);

FILL FILL_1__11128_ (
);

FILL FILL_0__8975_ (
);

FILL FILL_5__16361_ (
);

FILL FILL112440x72050 (
);

INVX1 _10826_ (
    .A(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_2008_)
);

FILL FILL_0__8135_ (
);

INVX1 _10406_ (
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_1789_)
);

FILL FILL_4__15774_ (
);

FILL SFILL104360x21050 (
);

FILL FILL_4__15354_ (
);

OAI21X1 _13298_ (
    .A(_3757_),
    .B(_3797_),
    .C(_3798_),
    .Y(_3834_)
);

FILL FILL_2__9934_ (
);

FILL FILL_0__11902_ (
);

FILL FILL_3__14767_ (
);

FILL FILL_2__9514_ (
);

FILL FILL_3__14347_ (
);

FILL FILL_1__15381_ (
);

FILL FILL_0__14794_ (
);

FILL FILL_0__14374_ (
);

FILL FILL_1__7931_ (
);

FILL FILL_2__14701_ (
);

FILL FILL_3__7857_ (
);

FILL FILL_3__7437_ (
);

FILL FILL_5__12281_ (
);

FILL FILL_4__16139_ (
);

FILL FILL_4__11694_ (
);

FILL FILL_4__11274_ (
);

FILL FILL_1__16166_ (
);

FILL FILL_3__10687_ (
);

FILL FILL_5__8724_ (
);

FILL FILL_3__10267_ (
);

FILL FILL_0__15999_ (
);

AOI22X1 _15864_ (
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [20]),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_6324_)
);

FILL FILL_0__15579_ (
);

OAI22X1 _15444_ (
    .A(_5914_),
    .B(_5518__bF$buf3),
    .C(_5478__bF$buf3),
    .D(_5913_),
    .Y(_5915_)
);

FILL FILL_0__15159_ (
);

NAND3X1 _15024_ (
    .A(_5459__bF$buf2),
    .B(_5462_),
    .C(_5476_),
    .Y(_5504_)
);

FILL FILL_0__10294_ (
);

FILL FILL_1__8716_ (
);

FILL SFILL94280x77050 (
);

FILL FILL_6__14493_ (
);

FILL FILL_6__14073_ (
);

FILL FILL_2__15906_ (
);

FILL FILL_0__16100_ (
);

FILL FILL_5__13486_ (
);

FILL FILL_2__10621_ (
);

DFFSR _7786_ (
    .Q(\datapath_1.regfile_1.regOut[7] [20]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_393_[20])
);

OAI21X1 _7366_ (
    .A(_249_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .C(_250_),
    .Y(_198_[26])
);

FILL FILL_4__12899_ (
);

FILL FILL_4__12479_ (
);

FILL FILL_4__12059_ (
);

FILL FILL_2__13093_ (
);

FILL FILL_5_BUFX2_insert50 (
);

FILL FILL_5_BUFX2_insert51 (
);

FILL FILL_5__9929_ (
);

FILL FILL_5__9509_ (
);

FILL FILL_5_BUFX2_insert52 (
);

FILL FILL_5_BUFX2_insert53 (
);

FILL FILL_1__12086_ (
);

FILL FILL_5_BUFX2_insert54 (
);

FILL FILL_5_BUFX2_insert55 (
);

FILL FILL_4__13840_ (
);

FILL FILL_5_BUFX2_insert56 (
);

FILL FILL_5_BUFX2_insert57 (
);

OAI22X1 _16229_ (
    .A(_5466__bF$buf3),
    .B(_5353_),
    .C(_5331_),
    .D(_5526__bF$buf2),
    .Y(_6680_)
);

FILL FILL_4__13420_ (
);

FILL FILL_4__13000_ (
);

FILL FILL_5_BUFX2_insert58 (
);

FILL FILL_5_BUFX2_insert59 (
);

NAND3X1 _11784_ (
    .A(_2874_),
    .B(_2877_),
    .C(_2870_),
    .Y(\datapath_1.ALUResult [6])
);

FILL FILL_3__7190_ (
);

FILL FILL_0__11499_ (
);

FILL FILL_0__9093_ (
);

INVX8 _11364_ (
    .A(_2346_),
    .Y(_2481_)
);

FILL FILL_0__11079_ (
);

FILL FILL_3__12833_ (
);

FILL FILL_3__12413_ (
);

FILL FILL_4__7926_ (
);

FILL FILL_4__7506_ (
);

FILL SFILL94280x32050 (
);

FILL FILL_4_CLKBUF1_insert220 (
);

FILL FILL_2__11826_ (
);

FILL FILL_4_CLKBUF1_insert221 (
);

FILL FILL_0__12860_ (
);

FILL FILL_4_CLKBUF1_insert222 (
);

FILL FILL_2__11406_ (
);

FILL FILL_4_CLKBUF1_insert223 (
);

FILL FILL_0__12440_ (
);

FILL FILL_4_CLKBUF1_insert224 (
);

FILL FILL_0__12020_ (
);

FILL FILL_1__10819_ (
);

FILL SFILL79000x55050 (
);

FILL FILL_2__14298_ (
);

FILL FILL_5__15632_ (
);

FILL FILL_5__15212_ (
);

FILL FILL_0__7826_ (
);

OAI21X1 _9932_ (
    .A(_1553_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .C(_1554_),
    .Y(_1498_[28])
);

OAI21X1 _9512_ (
    .A(_1334_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1335_),
    .Y(_1303_[16])
);

FILL FILL_4__14625_ (
);

FILL FILL_4__14205_ (
);

FILL FILL_3__8395_ (
);

OAI21X1 _12989_ (
    .A(_3643_),
    .B(vdd),
    .C(_3644_),
    .Y(_3620_[12])
);

OAI21X1 _12569_ (
    .A(_3488_),
    .B(vdd),
    .C(_3489_),
    .Y(_3425_[0])
);

NAND2X1 _12149_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.a [11]),
    .Y(_3153_)
);

FILL FILL_3__13618_ (
);

FILL FILL_1__14652_ (
);

FILL FILL_1__14232_ (
);

FILL SFILL84280x75050 (
);

FILL FILL_0__13645_ (
);

AOI21X1 _13930_ (
    .A(_4432_),
    .B(_4411_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [9])
);

FILL FILL_0__13225_ (
);

OAI22X1 _13510_ (
    .A(_4020_),
    .B(_3972__bF$buf2),
    .C(_3920_),
    .D(_4019_),
    .Y(_4021_)
);

FILL FILL_5__9682_ (
);

FILL FILL_5__9262_ (
);

FILL SFILL79000x10050 (
);

FILL FILL_5__11972_ (
);

FILL FILL_1__9674_ (
);

FILL FILL_5__11552_ (
);

FILL FILL_1__9254_ (
);

FILL FILL_5__11132_ (
);

BUFX2 BUFX2_insert1040 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf7 )
);

BUFX2 BUFX2_insert1041 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf6 )
);

BUFX2 BUFX2_insert1042 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf5 )
);

FILL FILL_2__16024_ (
);

BUFX2 BUFX2_insert1043 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf4 )
);

FILL FILL_4__10965_ (
);

BUFX2 BUFX2_insert1044 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf3 )
);

FILL FILL_4__10545_ (
);

FILL FILL_4__10125_ (
);

BUFX2 BUFX2_insert1045 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf2 )
);

BUFX2 BUFX2_insert1046 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf1 )
);

BUFX2 BUFX2_insert1047 (
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf0 )
);

FILL FILL_1__15857_ (
);

BUFX2 BUFX2_insert1048 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf4 )
);

FILL FILL_1__15437_ (
);

FILL SFILL4280x48050 (
);

FILL FILL_1__15017_ (
);

BUFX2 BUFX2_insert1049 (
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf3 )
);

FILL FILL_1__10992_ (
);

FILL SFILL84200x73050 (
);

FILL FILL_1__10572_ (
);

FILL FILL_1__10152_ (
);

NOR2X1 _14715_ (
    .A(_5200_),
    .B(_5188_),
    .Y(_5201_)
);

FILL SFILL84280x30050 (
);

BUFX2 BUFX2_insert860 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf3 )
);

FILL FILL_2__7597_ (
);

FILL FILL_2__7177_ (
);

BUFX2 BUFX2_insert861 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf2 )
);

BUFX2 BUFX2_insert862 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf1 )
);

BUFX2 BUFX2_insert863 (
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf0 )
);

BUFX2 BUFX2_insert864 (
    .A(_3950_),
    .Y(_3950__bF$buf3)
);

BUFX2 BUFX2_insert865 (
    .A(_3950_),
    .Y(_3950__bF$buf2)
);

BUFX2 BUFX2_insert866 (
    .A(_3950_),
    .Y(_3950__bF$buf1)
);

BUFX2 BUFX2_insert867 (
    .A(_3950_),
    .Y(_3950__bF$buf0)
);

BUFX2 BUFX2_insert868 (
    .A(_3891_),
    .Y(_3891__bF$buf3)
);

BUFX2 BUFX2_insert869 (
    .A(_3891_),
    .Y(_3891__bF$buf2)
);

FILL SFILL109480x73050 (
);

FILL FILL_5__12757_ (
);

FILL FILL_3__13791_ (
);

FILL FILL_5__12337_ (
);

FILL FILL_3__13371_ (
);

FILL FILL_4__8884_ (
);

FILL FILL_4__8464_ (
);

FILL FILL_2__12784_ (
);

FILL FILL_2__12364_ (
);

FILL FILL_1__11777_ (
);

FILL FILL_1__11357_ (
);

FILL FILL_5__16170_ (
);

FILL FILL_3__6881_ (
);

FILL FILL_0__8784_ (
);

FILL FILL_6__9751_ (
);

FILL FILL_0__8364_ (
);

INVX1 _10635_ (
    .A(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_1901_)
);

DFFSR _10215_ (
    .Q(\datapath_1.regfile_1.regOut[26] [17]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_1628_[17])
);

FILL FILL_6__14549_ (
);

FILL FILL_6__14129_ (
);

FILL FILL_4__15583_ (
);

FILL FILL_4__15163_ (
);

FILL FILL_2__9743_ (
);

FILL FILL_3__14996_ (
);

FILL FILL_3__14576_ (
);

FILL FILL_0__11711_ (
);

FILL FILL_3__14156_ (
);

FILL FILL_1__15190_ (
);

FILL FILL_6__15910_ (
);

FILL FILL_4__9669_ (
);

FILL FILL_4__9249_ (
);

FILL FILL_2__13989_ (
);

FILL FILL_2__13569_ (
);

FILL FILL_2__13149_ (
);

FILL FILL_0__14183_ (
);

FILL FILL_5__14903_ (
);

FILL SFILL114440x11050 (
);

FILL FILL_1__7740_ (
);

FILL FILL_1__7320_ (
);

FILL FILL_2__14930_ (
);

FILL FILL_2__14510_ (
);

FILL FILL_0__9989_ (
);

FILL FILL_0__9149_ (
);

FILL FILL_3__7246_ (
);

FILL FILL_5__12090_ (
);

FILL FILL_1__13923_ (
);

FILL FILL_4__16368_ (
);

FILL FILL_1__13503_ (
);

FILL FILL_6__10889_ (
);

FILL FILL_4__11083_ (
);

FILL FILL_0__12916_ (
);

FILL FILL_1__16395_ (
);

FILL FILL_5__8953_ (
);

FILL SFILL13160x41050 (
);

FILL FILL_3__10496_ (
);

FILL FILL_5__8533_ (
);

FILL FILL_5__8113_ (
);

FILL FILL_6__11830_ (
);

FILL FILL_0__15388_ (
);

INVX1 _15673_ (
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_6138_)
);

FILL FILL_6__11410_ (
);

OAI22X1 _15253_ (
    .A(_5727_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf2),
    .D(_5728_),
    .Y(_5729_)
);

FILL FILL_3__16302_ (
);

FILL FILL_5__10823_ (
);

FILL FILL_1__8525_ (
);

FILL FILL_5__10403_ (
);

FILL FILL_1__8105_ (
);

FILL FILL_2__15715_ (
);

FILL FILL_4__6950_ (
);

FILL FILL_5__13295_ (
);

FILL FILL_2__10430_ (
);

FILL FILL_2__10010_ (
);

FILL FILL_1__14708_ (
);

OAI21X1 _7595_ (
    .A(_361_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_362_),
    .Y(_328_[17])
);

OAI21X1 _7175_ (
    .A(_142_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_143_),
    .Y(_133_[5])
);

FILL FILL_4_BUFX2_insert1084 (
);

FILL FILL_4_BUFX2_insert1085 (
);

FILL FILL_4__12288_ (
);

FILL FILL_4_BUFX2_insert1086 (
);

FILL FILL_3__9812_ (
);

FILL FILL_4_BUFX2_insert1087 (
);

FILL FILL_4_BUFX2_insert1088 (
);

FILL FILL_4_BUFX2_insert1089 (
);

FILL FILL_0__6850_ (
);

FILL FILL_2__6868_ (
);

FILL FILL_5__9738_ (
);

OAI21X1 _16038_ (
    .A(_5526__bF$buf3),
    .B(_5111_),
    .C(_6493_),
    .Y(_6494_)
);

AOI21X1 _11593_ (
    .A(_2407_),
    .B(_2565_),
    .C(_2566_),
    .Y(_2700_)
);

NOR2X1 _11173_ (
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2292_)
);

FILL FILL_5__11608_ (
);

FILL FILL_3__12642_ (
);

FILL FILL_3__12222_ (
);

FILL FILL_4__7735_ (
);

FILL FILL_4__7315_ (
);

FILL FILL_2__11635_ (
);

FILL FILL_2__11215_ (
);

FILL FILL_1__10628_ (
);

FILL FILL_5__15861_ (
);

FILL FILL_5__15441_ (
);

FILL FILL112440x67050 (
);

FILL FILL_5__15021_ (
);

FILL FILL_0__7635_ (
);

OAI21X1 _9741_ (
    .A(_1446_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1447_),
    .Y(_1433_[7])
);

FILL FILL_0__7215_ (
);

DFFSR _9321_ (
    .Q(\datapath_1.regfile_1.regOut[19] [19]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_1173_[19])
);

FILL SFILL104360x16050 (
);

FILL FILL_4__14854_ (
);

FILL FILL_4__14434_ (
);

FILL FILL_4__14014_ (
);

DFFSR _12798_ (
    .Q(\datapath_1.PCJump [9]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[7])
);

OAI21X1 _12378_ (
    .A(_3316_),
    .B(MemToReg_bF$buf0),
    .C(_3317_),
    .Y(\datapath_1.mux_wd3.dout [11])
);

FILL FILL_3__13847_ (
);

FILL FILL_1__14881_ (
);

FILL FILL_3__13427_ (
);

FILL FILL_1__14461_ (
);

FILL FILL_3__13007_ (
);

FILL FILL_1__14041_ (
);

FILL FILL112040x53050 (
);

FILL FILL_0__13874_ (
);

FILL FILL_0__13454_ (
);

FILL FILL_0__13034_ (
);

FILL FILL_5__9491_ (
);

FILL FILL_5__16226_ (
);

FILL FILL_3__6937_ (
);

FILL FILL_5__11781_ (
);

FILL FILL_1__9483_ (
);

FILL FILL_5__11361_ (
);

FILL FILL112440x22050 (
);

FILL FILL_4__15639_ (
);

FILL FILL_4__15219_ (
);

FILL FILL_2__16253_ (
);

FILL FILL_4__10774_ (
);

FILL FILL_1__15666_ (
);

FILL FILL_1__15246_ (
);

FILL SFILL33720x40050 (
);

FILL FILL_5__7804_ (
);

FILL FILL_1__10381_ (
);

INVX1 _14944_ (
    .A(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_5425_)
);

FILL FILL_0__14659_ (
);

FILL FILL_0__14239_ (
);

NOR2X1 _14524_ (
    .A(_5013_),
    .B(_3954__bF$buf4),
    .Y(_5014_)
);

OAI22X1 _14104_ (
    .A(_4602_),
    .B(_3936__bF$buf4),
    .C(_3905__bF$buf3),
    .D(_4601_),
    .Y(_4603_)
);

FILL FILL_0__15600_ (
);

FILL FILL_5__12986_ (
);

FILL FILL_5__12146_ (
);

BUFX2 _6866_ (
    .A(_1_[28]),
    .Y(memoryAddress[28])
);

FILL FILL_4__11979_ (
);

FILL FILL_4__8273_ (
);

FILL FILL_4__11559_ (
);

FILL FILL_2__12593_ (
);

FILL FILL_4__11139_ (
);

FILL FILL_2__12173_ (
);

FILL SFILL23720x83050 (
);

FILL FILL_1__11586_ (
);

FILL FILL_1__11166_ (
);

NOR2X1 _15729_ (
    .A(_6192_),
    .B(_6190_),
    .Y(_6193_)
);

NAND3X1 _15309_ (
    .A(_5778_),
    .B(_5779_),
    .C(_5782_),
    .Y(_5783_)
);

FILL FILL_4__12500_ (
);

FILL FILL_0__10999_ (
);

FILL FILL_0__8593_ (
);

DFFSR _10864_ (
    .Q(\datapath_1.regfile_1.regOut[31] [26]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_1953_[26])
);

FILL FILL_0__10579_ (
);

OAI21X1 _10444_ (
    .A(_1813_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1814_),
    .Y(_1758_[28])
);

FILL FILL_0__10159_ (
);

OAI21X1 _10024_ (
    .A(_1594_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1595_),
    .Y(_1563_[16])
);

FILL FILL_3__11913_ (
);

FILL FILL_4__15392_ (
);

FILL SFILL94280x27050 (
);

FILL FILL_2__10906_ (
);

FILL FILL_0__11940_ (
);

FILL FILL_2__9552_ (
);

FILL FILL_2__9132_ (
);

FILL FILL_3__14385_ (
);

FILL FILL_0__11520_ (
);

FILL FILL_0__11100_ (
);

FILL FILL_4__9898_ (
);

FILL FILL_4__9478_ (
);

FILL FILL_2__13798_ (
);

FILL FILL_2__13378_ (
);

FILL FILL_5__14712_ (
);

FILL FILL_0__6906_ (
);

FILL FILL_4__13705_ (
);

FILL FILL_0__9798_ (
);

FILL FILL_0__9378_ (
);

FILL FILL_3__7475_ (
);

FILL FILL_3__7055_ (
);

INVX2 _11649_ (
    .A(_2162_),
    .Y(_2752_)
);

OAI22X1 _11229_ (
    .A(_2108_),
    .B(_2346_),
    .C(_2347__bF$buf2),
    .D(_2107_),
    .Y(_2348_)
);

FILL FILL_1__13732_ (
);

FILL FILL_1__13312_ (
);

FILL FILL_4__16177_ (
);

FILL FILL_0__12725_ (
);

FILL FILL_0__12305_ (
);

FILL FILL_5__8762_ (
);

FILL FILL_5__8342_ (
);

FILL FILL_0__15197_ (
);

NAND3X1 _15482_ (
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5952_)
);

FILL FILL_5__15917_ (
);

NOR3X1 _15062_ (
    .A(_3964_),
    .B(_5459__bF$buf0),
    .C(_5541_),
    .Y(_5542_)
);

FILL FILL_3__16111_ (
);

FILL FILL_5__10632_ (
);

FILL FILL_1__8754_ (
);

FILL FILL_1__8334_ (
);

FILL SFILL8680x44050 (
);

FILL FILL_2__15944_ (
);

FILL SFILL13720x81050 (
);

FILL FILL_2__15524_ (
);

FILL FILL_2__15104_ (
);

FILL SFILL109560x61050 (
);

FILL FILL_1__14937_ (
);

FILL FILL_1__14517_ (
);

FILL SFILL84200x68050 (
);

FILL FILL_4__12097_ (
);

FILL FILL_3__9621_ (
);

FILL SFILL84280x25050 (
);

FILL FILL_5__9547_ (
);

FILL FILL_5__9127_ (
);

FILL FILL_6__12004_ (
);

NAND3X1 _16267_ (
    .A(_6710_),
    .B(_6716_),
    .C(_6712_),
    .Y(_6717_)
);

FILL FILL_5__11837_ (
);

FILL FILL_3__12871_ (
);

FILL FILL_5__11417_ (
);

FILL FILL_1__9539_ (
);

FILL FILL_3__12451_ (
);

FILL FILL_1__9119_ (
);

FILL FILL_3__12031_ (
);

FILL FILL_4__7964_ (
);

FILL FILL_2__16309_ (
);

FILL FILL_4__7544_ (
);

FILL FILL_4__7124_ (
);

FILL FILL_2__11864_ (
);

FILL FILL_2__11444_ (
);

FILL FILL_2__11024_ (
);

NAND2X1 _8189_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_657_)
);

FILL FILL_1__10437_ (
);

FILL FILL_1__10017_ (
);

FILL FILL_5__15670_ (
);

FILL SFILL74280x68050 (
);

FILL FILL_5__15250_ (
);

FILL FILL_0__7864_ (
);

DFFSR _9970_ (
    .Q(\datapath_1.regfile_1.regOut[24] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_1498_[28])
);

FILL FILL_0__7444_ (
);

NAND2X1 _9550_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1361_)
);

NAND2X1 _9130_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1142_)
);

FILL FILL_4__14663_ (
);

FILL FILL_4__14243_ (
);

FILL SFILL13640x43050 (
);

INVX1 _12187_ (
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3178_)
);

FILL FILL_2__8823_ (
);

FILL FILL_3__13656_ (
);

FILL FILL_2__8403_ (
);

FILL FILL_3__13236_ (
);

FILL FILL_1__14690_ (
);

FILL SFILL109480x23050 (
);

FILL FILL_1__14270_ (
);

FILL FILL_0_BUFX2_insert500 (
);

FILL FILL_4__8749_ (
);

FILL FILL_0_BUFX2_insert501 (
);

FILL FILL_4__8329_ (
);

FILL FILL_0_BUFX2_insert502 (
);

FILL FILL_2__12649_ (
);

FILL FILL_0_BUFX2_insert503 (
);

FILL FILL_0__13683_ (
);

FILL FILL_2__12229_ (
);

FILL FILL_0_BUFX2_insert504 (
);

FILL FILL_0__13263_ (
);

FILL FILL_0_BUFX2_insert505 (
);

FILL FILL_0_BUFX2_insert506 (
);

FILL FILL_0_BUFX2_insert507 (
);

FILL SFILL104920x4050 (
);

FILL FILL_0_BUFX2_insert508 (
);

FILL FILL_0_BUFX2_insert509 (
);

FILL SFILL74200x66050 (
);

FILL FILL_5__16035_ (
);

FILL FILL_0__8649_ (
);

FILL FILL_0__8229_ (
);

FILL FILL_5__11590_ (
);

FILL FILL_1__9292_ (
);

FILL FILL_5__11170_ (
);

FILL SFILL74280x23050 (
);

FILL FILL_4__15868_ (
);

FILL FILL_4__15448_ (
);

FILL FILL_4__15028_ (
);

FILL FILL_2__16062_ (
);

FILL FILL_4__10163_ (
);

FILL FILL_2__9608_ (
);

FILL FILL_1__15895_ (
);

FILL FILL_1__15475_ (
);

FILL FILL_1__15055_ (
);

FILL FILL_5__7613_ (
);

FILL FILL_1__10190_ (
);

FILL FILL_6__10910_ (
);

FILL FILL_0__14888_ (
);

FILL FILL_0__14468_ (
);

NOR2X1 _14753_ (
    .A(_5234_),
    .B(_5237_),
    .Y(_5238_)
);

FILL FILL_0__14048_ (
);

NOR2X1 _14333_ (
    .A(_4816_),
    .B(_4826_),
    .Y(_4827_)
);

FILL FILL_3__15802_ (
);

FILL FILL_1__7605_ (
);

FILL FILL_6__13382_ (
);

FILL FILL_5__12375_ (
);

FILL SFILL74200x21050 (
);

FILL FILL_4__11788_ (
);

FILL FILL_4__8082_ (
);

FILL FILL_4__11368_ (
);

FILL FILL_1__11395_ (
);

OAI22X1 _15958_ (
    .A(_6415_),
    .B(_5548__bF$buf1),
    .C(_5463__bF$buf1),
    .D(_5031_),
    .Y(_6416_)
);

AOI22X1 _15538_ (
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [12]),
    .C(\datapath_1.regfile_1.regOut[6] [12]),
    .D(_5565__bF$buf2),
    .Y(_6006_)
);

OAI22X1 _15118_ (
    .A(_5480__bF$buf1),
    .B(_5595_),
    .C(_5596_),
    .D(_5499__bF$buf0),
    .Y(_5597_)
);

OAI21X1 _10673_ (
    .A(_1925_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .C(_1926_),
    .Y(_1888_[19])
);

FILL FILL_0__10388_ (
);

OAI21X1 _10253_ (
    .A(_1706_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .C(_1707_),
    .Y(_1693_[7])
);

FILL FILL_3__11722_ (
);

FILL FILL_3__11302_ (
);

FILL FILL_2__9781_ (
);

FILL SFILL33800x73050 (
);

FILL FILL_2__9361_ (
);

FILL SFILL64200x64050 (
);

FILL FILL_3__14194_ (
);

FILL FILL_4__9287_ (
);

FILL FILL_5__14941_ (
);

FILL FILL_5__14521_ (
);

FILL FILL_5__14101_ (
);

DFFSR _8821_ (
    .Q(\datapath_1.regfile_1.regOut[15] [31]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_913_[31])
);

NAND2X1 _8401_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_778_)
);

FILL SFILL68520x72050 (
);

FILL FILL_4__13934_ (
);

FILL FILL_4__13514_ (
);

INVX1 _11878_ (
    .A(\datapath_1.PCJump [20]),
    .Y(_2962_)
);

INVX1 _11458_ (
    .A(_2313_),
    .Y(_2573_)
);

INVX1 _11038_ (
    .A(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2157_)
);

FILL FILL_3__12507_ (
);

FILL FILL_1__13961_ (
);

FILL FILL_1__13541_ (
);

FILL FILL112040x48050 (
);

FILL FILL_1__13121_ (
);

FILL FILL_0__12954_ (
);

FILL FILL_3__15399_ (
);

FILL FILL_0__12534_ (
);

FILL FILL_0__12114_ (
);

FILL SFILL89400x1050 (
);

FILL FILL_5__8991_ (
);

FILL SFILL68920x41050 (
);

FILL FILL_5__8571_ (
);

OAI22X1 _15291_ (
    .A(_5765_),
    .B(_5548__bF$buf4),
    .C(_5534__bF$buf3),
    .D(_4216_),
    .Y(_5766_)
);

FILL FILL_5__15726_ (
);

FILL FILL_5__15306_ (
);

FILL FILL_3__16340_ (
);

NAND2X1 _9606_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1378_)
);

FILL FILL_1__8983_ (
);

FILL FILL_5__10441_ (
);

FILL FILL112440x17050 (
);

FILL FILL_1__8143_ (
);

FILL FILL_5__10021_ (
);

FILL FILL_4__14719_ (
);

FILL FILL_2__15753_ (
);

FILL FILL_2__15333_ (
);

FILL FILL_3__8489_ (
);

FILL FILL_3__8069_ (
);

FILL FILL_1__14746_ (
);

FILL FILL_1__14326_ (
);

FILL FILL_3__9850_ (
);

FILL FILL_0__13739_ (
);

FILL FILL_0__13319_ (
);

NOR2X1 _13604_ (
    .A(_4112_),
    .B(_3935__bF$buf3),
    .Y(_4113_)
);

FILL FILL_3__9010_ (
);

FILL FILL_5__9776_ (
);

FILL FILL_5__9356_ (
);

NAND3X1 _16076_ (
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6531_)
);

FILL FILL_1__9768_ (
);

FILL FILL_5__11646_ (
);

FILL FILL_1__9348_ (
);

FILL FILL_5__11226_ (
);

FILL FILL_3__12260_ (
);

FILL FILL_2__16118_ (
);

FILL FILL_4__7353_ (
);

FILL FILL_4__10639_ (
);

FILL FILL_2__11673_ (
);

FILL FILL_2__11253_ (
);

FILL FILL_6__7699_ (
);

FILL SFILL23720x78050 (
);

FILL FILL_1__10666_ (
);

FILL FILL_1__10246_ (
);

OAI22X1 _14809_ (
    .A(_3884__bF$buf1),
    .B(_5291_),
    .C(_3977__bF$buf1),
    .D(_5292_),
    .Y(_5293_)
);

FILL FILL_0__7673_ (
);

FILL FILL_6__8640_ (
);

FILL FILL_0__7253_ (
);

FILL FILL_6__13858_ (
);

FILL FILL_4__14892_ (
);

FILL FILL_4__14472_ (
);

FILL FILL_4__14052_ (
);

FILL FILL_3__13885_ (
);

FILL FILL_2__8632_ (
);

FILL FILL_3__13465_ (
);

FILL FILL_2__8212_ (
);

FILL FILL_3__13045_ (
);

FILL FILL_4__8978_ (
);

FILL FILL_4__8138_ (
);

FILL FILL_2__12878_ (
);

FILL FILL_2__12458_ (
);

FILL FILL_2__12038_ (
);

FILL FILL_0__13492_ (
);

FILL FILL_3__6975_ (
);

FILL FILL_0__8878_ (
);

FILL FILL_5__16264_ (
);

FILL FILL_0__8458_ (
);

DFFSR _10729_ (
    .Q(\datapath_1.regfile_1.regOut[30] [19]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1888_[19])
);

FILL FILL_6__9425_ (
);

NAND2X1 _10309_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1745_)
);

FILL FILL_4__15677_ (
);

FILL FILL_4__15257_ (
);

FILL FILL_2__16291_ (
);

FILL FILL_4__10392_ (
);

FILL FILL_2__9417_ (
);

FILL FILL_0__11805_ (
);

FILL FILL_1__15284_ (
);

FILL FILL_5__7842_ (
);

FILL FILL_5__7422_ (
);

AND2X2 _14982_ (
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5462_)
);

FILL FILL_0__14697_ (
);

INVX1 _14562_ (
    .A(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_5051_)
);

FILL FILL_0__14277_ (
);

NOR2X1 _14142_ (
    .A(_4639_),
    .B(_4636_),
    .Y(_4640_)
);

FILL FILL_3__15611_ (
);

FILL FILL_1__7834_ (
);

FILL FILL_1__7414_ (
);

FILL SFILL13720x76050 (
);

FILL SFILL44120x67050 (
);

FILL FILL_2__14604_ (
);

FILL SFILL109560x56050 (
);

FILL SFILL23240x26050 (
);

FILL FILL_5__12184_ (
);

FILL SFILL99560x3050 (
);

FILL FILL_4__11597_ (
);

FILL FILL_4__11177_ (
);

FILL FILL_3__8701_ (
);

FILL FILL_1__16069_ (
);

FILL FILL_5__8627_ (
);

FILL FILL_5__8207_ (
);

NOR2X1 _15767_ (
    .A(_6228_),
    .B(_6229_),
    .Y(_6230_)
);

NOR2X1 _15347_ (
    .A(_5818_),
    .B(_5819_),
    .Y(_5820_)
);

DFFSR _10482_ (
    .Q(\datapath_1.regfile_1.regOut[28] [28]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_1758_[28])
);

FILL FILL_0__10197_ (
);

NAND2X1 _10062_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1621_)
);

FILL FILL_5__10917_ (
);

FILL FILL_3__11951_ (
);

FILL FILL_1__8619_ (
);

FILL FILL_3__11531_ (
);

FILL FILL_3__11111_ (
);

FILL FILL_2__15809_ (
);

FILL FILL_0__16003_ (
);

FILL FILL_2__10944_ (
);

FILL SFILL13720x31050 (
);

FILL FILL_5__13389_ (
);

FILL FILL_2__9590_ (
);

FILL FILL_2__10524_ (
);

FILL FILL_2__10104_ (
);

FILL FILL_2__9170_ (
);

NAND2X1 _7689_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_405_)
);

DFFSR _7269_ (
    .Q(\datapath_1.regfile_1.regOut[3] [15]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_133_[15])
);

FILL FILL_4__9096_ (
);

FILL FILL_3__9906_ (
);

FILL SFILL38920x80050 (
);

FILL SFILL84200x18050 (
);

FILL FILL_5__14750_ (
);

FILL FILL_0__6944_ (
);

FILL FILL_5__14330_ (
);

NAND2X1 _8630_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_890_)
);

NAND2X1 _8210_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_671_)
);

FILL FILL_4__13743_ (
);

FILL FILL_4__13323_ (
);

FILL SFILL13640x38050 (
);

FILL FILL_3__7093_ (
);

NAND3X1 _11687_ (
    .A(_2514_),
    .B(_2462__bF$buf3),
    .C(_2743_),
    .Y(_2788_)
);

NOR2X1 _11267_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2386_)
);

FILL FILL_3__12736_ (
);

FILL SFILL109480x18050 (
);

FILL FILL_1__13770_ (
);

FILL FILL_3__12316_ (
);

FILL FILL_1__13350_ (
);

FILL FILL_4__7829_ (
);

FILL FILL_2__11729_ (
);

FILL FILL_0__12763_ (
);

FILL FILL_2__11309_ (
);

FILL FILL_0__12343_ (
);

FILL FILL_5__8380_ (
);

FILL FILL_5__15955_ (
);

FILL FILL_5__15535_ (
);

FILL FILL_0__7729_ (
);

FILL FILL_5__15115_ (
);

DFFSR _9835_ (
    .Q(\datapath_1.regfile_1.regOut[23] [21]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1433_[21])
);

FILL FILL_0__7309_ (
);

INVX1 _9415_ (
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_1291_)
);

FILL FILL_5__10670_ (
);

FILL FILL_5__10250_ (
);

FILL FILL_1__8372_ (
);

FILL FILL_4__14948_ (
);

FILL FILL_2__15982_ (
);

FILL FILL_4__14528_ (
);

FILL FILL_2__15562_ (
);

FILL FILL_4__14108_ (
);

FILL FILL_2__15142_ (
);

FILL FILL_1__14975_ (
);

FILL SFILL99480x67050 (
);

FILL FILL_1__14555_ (
);

FILL FILL_1__14135_ (
);

FILL FILL_0__13968_ (
);

OAI22X1 _13833_ (
    .A(_3978_),
    .B(_4336_),
    .C(_3977__bF$buf3),
    .D(_4337_),
    .Y(_4338_)
);

FILL FILL_0__13548_ (
);

NAND2X1 _13413_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3901_),
    .Y(_3925_)
);

FILL FILL_0__13128_ (
);

FILL FILL_5__9165_ (
);

FILL FILL_6__12882_ (
);

FILL FILL_1__9997_ (
);

FILL FILL_5__11875_ (
);

FILL SFILL74200x16050 (
);

FILL FILL_5__11455_ (
);

FILL FILL_1__9157_ (
);

FILL FILL_5__11035_ (
);

FILL FILL_2__16347_ (
);

FILL FILL_4__7582_ (
);

FILL FILL_4__7162_ (
);

FILL FILL_4__10448_ (
);

FILL FILL_4__10028_ (
);

FILL FILL_2__11482_ (
);

FILL FILL_2__11062_ (
);

FILL FILL_1__10895_ (
);

FILL SFILL99480x22050 (
);

FILL FILL_1__10055_ (
);

NOR2X1 _14618_ (
    .A(_5095_),
    .B(_5105_),
    .Y(_5106_)
);

FILL FILL_0__7482_ (
);

FILL FILL_0__7062_ (
);

FILL SFILL24120x63050 (
);

FILL FILL_3__10802_ (
);

FILL FILL_4__14281_ (
);

FILL SFILL33800x68050 (
);

FILL FILL_2__8861_ (
);

FILL FILL_2__8441_ (
);

FILL FILL_3__13694_ (
);

FILL FILL_3__13274_ (
);

FILL FILL_2__8021_ (
);

FILL FILL112120x36050 (
);

FILL FILL_4__8787_ (
);

FILL FILL_4__8367_ (
);

FILL FILL_2__12267_ (
);

FILL FILL_5__13601_ (
);

DFFSR _7901_ (
    .Q(\datapath_1.regfile_1.regOut[8] [7]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_458_[7])
);

FILL SFILL73880x80050 (
);

FILL FILL_5__16073_ (
);

NOR2X1 _10958_ (
    .A(_2075_),
    .B(_2089_),
    .Y(_2090_)
);

FILL FILL_0__8267_ (
);

NAND2X1 _10538_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1857_)
);

NAND2X1 _10118_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1638_)
);

FILL FILL_1__12621_ (
);

FILL FILL_4__15486_ (
);

FILL SFILL28840x40050 (
);

FILL FILL_4__15066_ (
);

FILL FILL_1__12201_ (
);

FILL FILL_2__9646_ (
);

FILL FILL_3__14899_ (
);

FILL FILL_3__14479_ (
);

FILL FILL_2__9226_ (
);

FILL FILL_0__11614_ (
);

FILL FILL_3__14059_ (
);

FILL FILL_1__15093_ (
);

FILL SFILL33800x23050 (
);

FILL SFILL64200x14050 (
);

FILL FILL_5__7231_ (
);

AOI21X1 _14791_ (
    .A(_5250_),
    .B(_5275_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [27])
);

INVX1 _14371_ (
    .A(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_4864_)
);

FILL FILL_0__14086_ (
);

FILL FILL_5__14806_ (
);

FILL FILL_3__15840_ (
);

FILL FILL_3__15420_ (
);

FILL FILL_3__15000_ (
);

FILL FILL_1__7223_ (
);

FILL FILL_2__14833_ (
);

FILL SFILL68520x22050 (
);

FILL FILL_3__7989_ (
);

FILL FILL_2__14413_ (
);

FILL FILL_3__7569_ (
);

FILL FILL_1__13826_ (
);

FILL FILL_1__13406_ (
);

FILL SFILL18840x83050 (
);

FILL FILL_3__8510_ (
);

FILL FILL_1__16298_ (
);

FILL FILL_5__8856_ (
);

FILL FILL_3__10399_ (
);

FILL FILL_5__8016_ (
);

OAI21X1 _15996_ (
    .A(_5526__bF$buf2),
    .B(_5074_),
    .C(_6452_),
    .Y(_6453_)
);

OAI22X1 _15576_ (
    .A(_5472__bF$buf0),
    .B(_4613_),
    .C(_4612_),
    .D(_5552__bF$buf1),
    .Y(_6043_)
);

FILL FILL_6__11313_ (
);

NAND2X1 _15156_ (
    .A(_5628_),
    .B(_5633_),
    .Y(_5634_)
);

FILL FILL_3__16205_ (
);

NAND2X1 _10291_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1733_)
);

FILL FILL_1__8848_ (
);

FILL FILL_3__11760_ (
);

FILL FILL_5__10306_ (
);

FILL FILL_3__11340_ (
);

FILL FILL_1__8008_ (
);

FILL FILL_2__15618_ (
);

FILL FILL_4__6853_ (
);

FILL FILL_0__16232_ (
);

FILL FILL_2__10753_ (
);

FILL SFILL79240x50 (
);

INVX1 _7498_ (
    .A(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_318_)
);

INVX1 _7078_ (
    .A(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_99_)
);

FILL FILL_6__7720_ (
);

FILL FILL_4__13972_ (
);

FILL FILL_4__13552_ (
);

FILL FILL_4__13132_ (
);

AND2X2 _11496_ (
    .A(_2608_),
    .B(_2607_),
    .Y(_2609_)
);

FILL SFILL103560x54050 (
);

INVX1 _11076_ (
    .A(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2195_)
);

FILL FILL_2__7712_ (
);

FILL FILL_3__12965_ (
);

FILL FILL_3__12125_ (
);

FILL FILL_4__7218_ (
);

FILL FILL_2__11958_ (
);

FILL FILL_0__12992_ (
);

FILL FILL_2__11538_ (
);

FILL FILL_3_CLKBUF1_insert160 (
);

FILL FILL_0__12572_ (
);

FILL FILL_2__11118_ (
);

FILL FILL_0__12152_ (
);

FILL FILL_3_CLKBUF1_insert161 (
);

FILL FILL_3_CLKBUF1_insert162 (
);

FILL FILL_3_CLKBUF1_insert163 (
);

FILL FILL_3_CLKBUF1_insert164 (
);

FILL FILL_3_CLKBUF1_insert165 (
);

FILL FILL_3_CLKBUF1_insert166 (
);

FILL SFILL74120x7050 (
);

FILL FILL_3_CLKBUF1_insert167 (
);

FILL SFILL23720x28050 (
);

FILL FILL_3_CLKBUF1_insert168 (
);

FILL FILL_3_CLKBUF1_insert169 (
);

FILL FILL_5__15764_ (
);

FILL FILL_5__15344_ (
);

FILL FILL_0__7958_ (
);

FILL FILL_0__7118_ (
);

FILL FILL_6__8505_ (
);

INVX1 _9644_ (
    .A(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_1403_)
);

INVX1 _9224_ (
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_1184_)
);

FILL FILL_4__14757_ (
);

FILL FILL_2__15791_ (
);

FILL FILL_4__14337_ (
);

FILL FILL_2__15371_ (
);

FILL FILL_2__8917_ (
);

FILL FILL_1__14784_ (
);

FILL FILL_1__14364_ (
);

FILL FILL_5__6922_ (
);

FILL FILL_0__13777_ (
);

FILL FILL_0__13357_ (
);

INVX1 _13642_ (
    .A(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_4150_)
);

NOR2X1 _13222_ (
    .A(_3752_),
    .B(_3764_),
    .Y(_3765_)
);

FILL FILL_5__9394_ (
);

FILL FILL_1__6914_ (
);

FILL FILL_5__16129_ (
);

FILL FILL_5__11684_ (
);

FILL FILL_1__9386_ (
);

FILL FILL_5__11264_ (
);

FILL FILL_2__16156_ (
);

FILL FILL_4__10677_ (
);

FILL FILL_4__10257_ (
);

FILL SFILL48920x32050 (
);

FILL FILL_2__11291_ (
);

FILL FILL_1__15989_ (
);

FILL FILL_1__15569_ (
);

FILL FILL_1__15149_ (
);

FILL FILL_5__7707_ (
);

FILL FILL_2_BUFX2_insert410 (
);

FILL FILL_2_BUFX2_insert411 (
);

FILL FILL_1__10284_ (
);

FILL FILL_2_BUFX2_insert412 (
);

AOI22X1 _14847_ (
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .B(_4090_),
    .C(_3998__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_5330_)
);

FILL FILL_2_BUFX2_insert413 (
);

FILL FILL_2_BUFX2_insert414 (
);

INVX1 _14427_ (
    .A(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_4919_)
);

OAI22X1 _14007_ (
    .A(_4506_),
    .B(_3931__bF$buf2),
    .C(_3947__bF$buf1),
    .D(_4507_),
    .Y(_4508_)
);

FILL FILL_2_BUFX2_insert415 (
);

FILL FILL_2_BUFX2_insert416 (
);

FILL FILL_2_BUFX2_insert417 (
);

FILL FILL_0__7291_ (
);

FILL FILL_2_BUFX2_insert418 (
);

FILL FILL_2_BUFX2_insert419 (
);

FILL FILL_0_CLKBUF1_insert111 (
);

FILL FILL_4__14090_ (
);

FILL FILL_0__15923_ (
);

FILL FILL_0_CLKBUF1_insert112 (
);

FILL FILL_0__15503_ (
);

FILL FILL_0_CLKBUF1_insert113 (
);

FILL SFILL48840x39050 (
);

FILL FILL_0_CLKBUF1_insert114 (
);

FILL SFILL13720x26050 (
);

FILL FILL_5__12889_ (
);

FILL FILL_0_CLKBUF1_insert115 (
);

FILL FILL_5__12469_ (
);

FILL FILL_0_CLKBUF1_insert116 (
);

FILL FILL_2__8250_ (
);

FILL FILL_5__12049_ (
);

FILL FILL_0_CLKBUF1_insert117 (
);

FILL FILL_3__13083_ (
);

FILL FILL_0_CLKBUF1_insert118 (
);

FILL FILL_0_CLKBUF1_insert119 (
);

FILL FILL_4__8596_ (
);

FILL FILL_2__12496_ (
);

FILL SFILL38920x75050 (
);

FILL FILL_2__12076_ (
);

FILL FILL_5__13830_ (
);

FILL FILL_5__13410_ (
);

NAND2X1 _7710_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_419_)
);

FILL FILL_1__11489_ (
);

FILL FILL_1__11069_ (
);

FILL FILL_4__12823_ (
);

FILL FILL_4__12403_ (
);

FILL FILL_0__8496_ (
);

NAND2X1 _10767_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1969_)
);

FILL FILL_0__8076_ (
);

DFFSR _10347_ (
    .Q(\datapath_1.regfile_1.regOut[27] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_1693_[21])
);

FILL FILL_6__9043_ (
);

FILL SFILL93880x34050 (
);

FILL FILL_3__11816_ (
);

FILL FILL_1__12850_ (
);

FILL FILL_1__12430_ (
);

FILL FILL_4__15295_ (
);

FILL FILL_1__12010_ (
);

FILL FILL_4__6909_ (
);

FILL FILL_2__10809_ (
);

FILL FILL_2__9875_ (
);

FILL FILL_0__11843_ (
);

FILL FILL_2__9035_ (
);

FILL FILL_3__14288_ (
);

FILL FILL_0__11423_ (
);

FILL FILL_0__11003_ (
);

FILL FILL_5__7880_ (
);

FILL FILL_5__7460_ (
);

FILL FILL_5__7040_ (
);

FILL SFILL3560x74050 (
);

AOI22X1 _14180_ (
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .B(_3995__bF$buf4),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_4677_)
);

FILL FILL_5__14615_ (
);

INVX1 _8915_ (
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_1039_)
);

FILL SFILL38920x30050 (
);

FILL FILL_1__7872_ (
);

FILL FILL_1__7452_ (
);

FILL FILL_1__7032_ (
);

FILL FILL_4__13608_ (
);

FILL FILL_2__14642_ (
);

FILL FILL_2__14222_ (
);

FILL FILL_3__7798_ (
);

FILL FILL_3__7378_ (
);

FILL FILL112200x69050 (
);

FILL FILL_1__13635_ (
);

FILL FILL_1__13215_ (
);

FILL FILL_1_BUFX2_insert430 (
);

FILL FILL_1_BUFX2_insert431 (
);

FILL FILL_0__12628_ (
);

INVX1 _12913_ (
    .A(\datapath_1.a [30]),
    .Y(_3614_)
);

FILL FILL_1_BUFX2_insert432 (
);

FILL FILL_1_BUFX2_insert433 (
);

FILL FILL_0__12208_ (
);

FILL FILL_1_BUFX2_insert434 (
);

FILL SFILL38840x37050 (
);

FILL FILL_1_BUFX2_insert435 (
);

FILL FILL_1_BUFX2_insert436 (
);

FILL FILL_6_BUFX2_insert991 (
);

FILL FILL_5__8245_ (
);

FILL FILL_1_BUFX2_insert437 (
);

FILL FILL_1_BUFX2_insert438 (
);

FILL FILL_1_BUFX2_insert439 (
);

INVX1 _15385_ (
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_5857_)
);

FILL FILL_6_BUFX2_insert996 (
);

FILL FILL_3__16014_ (
);

FILL SFILL28920x73050 (
);

FILL FILL_5__10955_ (
);

FILL FILL_5__10535_ (
);

FILL FILL_1__8657_ (
);

FILL FILL_5__10115_ (
);

FILL FILL_1__8237_ (
);

FILL FILL_2__15847_ (
);

FILL FILL_2__15427_ (
);

FILL FILL_2__15007_ (
);

FILL FILL_0__16041_ (
);

FILL FILL_2__10982_ (
);

FILL FILL_2__10562_ (
);

FILL FILL_2__10142_ (
);

FILL SFILL9240x50050 (
);

FILL SFILL99480x17050 (
);

FILL FILL_3__9524_ (
);

FILL FILL_3__9104_ (
);

FILL FILL_0__6982_ (
);

FILL FILL_4__13781_ (
);

FILL FILL_4__13361_ (
);

FILL FILL_2__7941_ (
);

FILL SFILL9160x57050 (
);

FILL FILL_3__12774_ (
);

BUFX2 BUFX2_insert100 (
    .A(_5489_),
    .Y(_5489__bF$buf2)
);

FILL FILL_2__7101_ (
);

FILL FILL_3__12354_ (
);

BUFX2 BUFX2_insert101 (
    .A(_5489_),
    .Y(_5489__bF$buf1)
);

BUFX2 BUFX2_insert102 (
    .A(_5489_),
    .Y(_5489__bF$buf0)
);

BUFX2 BUFX2_insert103 (
    .A(IorD),
    .Y(IorD_bF$buf7)
);

FILL FILL_4__7867_ (
);

BUFX2 BUFX2_insert104 (
    .A(IorD),
    .Y(IorD_bF$buf6)
);

BUFX2 BUFX2_insert105 (
    .A(IorD),
    .Y(IorD_bF$buf5)
);

FILL FILL_4__7447_ (
);

BUFX2 BUFX2_insert106 (
    .A(IorD),
    .Y(IorD_bF$buf4)
);

BUFX2 BUFX2_insert107 (
    .A(IorD),
    .Y(IorD_bF$buf3)
);

FILL FILL_2__11767_ (
);

BUFX2 BUFX2_insert108 (
    .A(IorD),
    .Y(IorD_bF$buf2)
);

FILL FILL_2__11347_ (
);

FILL FILL_0__12381_ (
);

BUFX2 BUFX2_insert109 (
    .A(IorD),
    .Y(IorD_bF$buf1)
);

FILL FILL_6__16160_ (
);

FILL FILL_2_CLKBUF1_insert150 (
);

FILL FILL_2_CLKBUF1_insert151 (
);

FILL FILL_5__15993_ (
);

FILL FILL_2_CLKBUF1_insert152 (
);

FILL FILL_2_CLKBUF1_insert153 (
);

FILL FILL_5__15573_ (
);

FILL FILL_5__15153_ (
);

FILL FILL_2_CLKBUF1_insert154 (
);

FILL FILL_0__7347_ (
);

INVX1 _9873_ (
    .A(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_1515_)
);

FILL FILL_2_CLKBUF1_insert155 (
);

FILL FILL_2_CLKBUF1_insert156 (
);

DFFSR _9453_ (
    .Q(\datapath_1.regfile_1.regOut[20] [23]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_1238_[23])
);

FILL FILL_2_CLKBUF1_insert157 (
);

OAI21X1 _9033_ (
    .A(_1096_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1097_),
    .Y(_1043_[27])
);

FILL FILL_2_CLKBUF1_insert158 (
);

FILL FILL_4__14986_ (
);

FILL FILL_2_CLKBUF1_insert159 (
);

FILL SFILL28840x35050 (
);

FILL FILL_4__14566_ (
);

FILL FILL_1__11701_ (
);

FILL FILL_4__14146_ (
);

FILL FILL_2__15180_ (
);

FILL SFILL103720x80050 (
);

FILL FILL_3__13979_ (
);

FILL FILL_2__8726_ (
);

FILL FILL_3__13559_ (
);

FILL FILL_1__14593_ (
);

FILL FILL_3__13139_ (
);

FILL FILL_1__14173_ (
);

FILL SFILL33800x18050 (
);

FILL FILL_6_BUFX2_insert1032 (
);

FILL FILL_0__13586_ (
);

OAI22X1 _13871_ (
    .A(_3884__bF$buf1),
    .B(_4373_),
    .C(_4374_),
    .D(_3967__bF$buf3),
    .Y(_4375_)
);

FILL FILL_0__13166_ (
);

NAND3X1 _13451_ (
    .A(_3946_),
    .B(_3951_),
    .C(_3962_),
    .Y(_3963_)
);

FILL FILL_6_BUFX2_insert1037 (
);

OAI21X1 _13031_ (
    .A(_3671_),
    .B(vdd),
    .C(_3672_),
    .Y(_3620_[26])
);

FILL FILL_3__14920_ (
);

FILL FILL_3__14500_ (
);

FILL FILL_6__12080_ (
);

FILL FILL_2__13913_ (
);

FILL FILL_5__16358_ (
);

FILL FILL_6__9519_ (
);

FILL FILL_5__11493_ (
);

FILL FILL_5__11073_ (
);

FILL FILL_1__12906_ (
);

FILL FILL_2__16385_ (
);

FILL FILL_4__10486_ (
);

FILL FILL_0__9913_ (
);

FILL FILL_4__10066_ (
);

FILL FILL_1__15798_ (
);

FILL FILL_1__15378_ (
);

FILL FILL_5__7936_ (
);

FILL SFILL13800x8050 (
);

AOI22X1 _14656_ (
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .B(_4129_),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_5143_)
);

INVX1 _14236_ (
    .A(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_4732_)
);

FILL FILL_3__15705_ (
);

FILL FILL_1__7928_ (
);

FILL FILL_1__7508_ (
);

FILL FILL_6__13285_ (
);

FILL FILL_3__10420_ (
);

FILL FILL_3__10000_ (
);

FILL FILL_0__15732_ (
);

FILL FILL_0__15312_ (
);

FILL FILL_5__12698_ (
);

FILL SFILL103640x42050 (
);

FILL FILL_5__12278_ (
);

DFFSR _6998_ (
    .Q(\datapath_1.regfile_1.regOut[1] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_3_[0])
);

FILL SFILL18840x33050 (
);

FILL FILL_1__11298_ (
);

FILL FILL_4__12632_ (
);

FILL FILL_4__12212_ (
);

NOR2X1 _10996_ (
    .A(\datapath_1.alu_1.ALUInA [30]),
    .B(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2115_)
);

INVX1 _10576_ (
    .A(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_1882_)
);

INVX1 _10156_ (
    .A(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_1663_)
);

FILL FILL_3_BUFX2_insert1090 (
);

FILL FILL_3_BUFX2_insert1091 (
);

FILL FILL_3_BUFX2_insert1092 (
);

FILL FILL_3__11625_ (
);

FILL FILL_3_BUFX2_insert1093 (
);

FILL FILL_3__11205_ (
);

FILL FILL_2__9684_ (
);

FILL FILL_2__10618_ (
);

FILL FILL_2__9264_ (
);

FILL FILL_0__11652_ (
);

FILL FILL_0__11232_ (
);

FILL FILL_3__14097_ (
);

FILL FILL_5__14844_ (
);

FILL FILL_5__14424_ (
);

FILL FILL_5__14004_ (
);

INVX1 _8724_ (
    .A(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_932_)
);

DFFSR _8304_ (
    .Q(\datapath_1.regfile_1.regOut[11] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_653_[26])
);

FILL FILL_1__7681_ (
);

FILL FILL_4__13837_ (
);

FILL FILL_2__14871_ (
);

FILL FILL_4__13417_ (
);

FILL FILL_2__14451_ (
);

FILL FILL_2__14031_ (
);

FILL FILL_3__7187_ (
);

FILL FILL_1__13864_ (
);

FILL FILL_1__13444_ (
);

FILL FILL_1__13024_ (
);

FILL FILL_4_CLKBUF1_insert190 (
);

FILL FILL_4_CLKBUF1_insert191 (
);

FILL FILL_4_CLKBUF1_insert192 (
);

FILL FILL_0__12857_ (
);

FILL FILL_4_CLKBUF1_insert193 (
);

FILL FILL_0__12437_ (
);

INVX1 _12722_ (
    .A(\datapath_1.PCJump [11]),
    .Y(_3507_)
);

FILL SFILL114520x81050 (
);

FILL FILL_4_CLKBUF1_insert194 (
);

FILL FILL_0__12017_ (
);

NAND3X1 _12302_ (
    .A(_3263_),
    .B(_3264_),
    .C(_3265_),
    .Y(\datapath_1.alu_1.ALUInB [21])
);

FILL SFILL53880x71050 (
);

FILL FILL_4_CLKBUF1_insert195 (
);

FILL FILL_5__8894_ (
);

FILL FILL_4_CLKBUF1_insert196 (
);

FILL FILL_5__8474_ (
);

FILL FILL_4_CLKBUF1_insert197 (
);

FILL FILL_4_CLKBUF1_insert198 (
);

FILL FILL_5__8054_ (
);

FILL FILL_4_CLKBUF1_insert199 (
);

OAI22X1 _15194_ (
    .A(_5489__bF$buf1),
    .B(_4095_),
    .C(_4121_),
    .D(_5504__bF$buf1),
    .Y(_5671_)
);

FILL FILL_5__15629_ (
);

FILL FILL_5__15209_ (
);

FILL FILL_3__16243_ (
);

OAI21X1 _9929_ (
    .A(_1551_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .C(_1552_),
    .Y(_1498_[27])
);

OAI21X1 _9509_ (
    .A(_1332_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .C(_1333_),
    .Y(_1303_[15])
);

FILL FILL_5__10764_ (
);

FILL FILL_1__8886_ (
);

FILL FILL_1__8466_ (
);

FILL FILL_2__15656_ (
);

FILL FILL_4__6891_ (
);

FILL FILL_2__15236_ (
);

FILL FILL_0__16270_ (
);

FILL FILL_2__10791_ (
);

FILL FILL_2__10371_ (
);

FILL FILL_1__14649_ (
);

FILL FILL_1__14229_ (
);

FILL FILL_3__9753_ (
);

AOI22X1 _13927_ (
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .B(_4005__bF$buf0),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_4430_)
);

OAI22X1 _13507_ (
    .A(_4017_),
    .B(_3971__bF$buf3),
    .C(_3924__bF$buf1),
    .D(_4016_),
    .Y(_4018_)
);

FILL FILL_5__9679_ (
);

FILL FILL_5__9259_ (
);

FILL FILL_6__12976_ (
);

FILL FILL_4__13590_ (
);

INVX1 _16399_ (
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .Y(_6820_)
);

FILL FILL_4__13170_ (
);

FILL FILL_5__11969_ (
);

FILL FILL_2__7750_ (
);

FILL FILL_5__11549_ (
);

FILL FILL_3__12583_ (
);

FILL FILL_2__7330_ (
);

FILL FILL_5__11129_ (
);

FILL FILL_3__12163_ (
);

FILL FILL_4__7676_ (
);

FILL FILL_2__11996_ (
);

FILL FILL_2__11576_ (
);

FILL FILL_2__11156_ (
);

FILL FILL_0__12190_ (
);

FILL FILL_5__12910_ (
);

FILL FILL_1__10989_ (
);

FILL FILL_1__10569_ (
);

FILL FILL_1__10149_ (
);

FILL FILL_4__11903_ (
);

FILL FILL_5__15382_ (
);

FILL FILL_0__7996_ (
);

FILL FILL_0__7576_ (
);

OAI21X1 _9682_ (
    .A(_1427_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .C(_1428_),
    .Y(_1368_[30])
);

FILL FILL_6__8123_ (
);

OAI21X1 _9262_ (
    .A(_1208_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1209_),
    .Y(_1173_[18])
);

FILL FILL_1_CLKBUF1_insert140 (
);

FILL FILL_1_CLKBUF1_insert141 (
);

FILL FILL_1_CLKBUF1_insert142 (
);

FILL FILL_4__14795_ (
);

FILL FILL_1__11930_ (
);

FILL FILL_1_CLKBUF1_insert143 (
);

FILL FILL_4__14375_ (
);

FILL FILL_1__11510_ (
);

FILL FILL_1_CLKBUF1_insert144 (
);

FILL FILL_1_CLKBUF1_insert145 (
);

FILL FILL_1_CLKBUF1_insert146 (
);

FILL FILL_1_CLKBUF1_insert147 (
);

FILL FILL_2__8955_ (
);

FILL FILL_1_CLKBUF1_insert148 (
);

FILL FILL_1_CLKBUF1_insert149 (
);

FILL FILL_0__10923_ (
);

FILL FILL_3__13788_ (
);

FILL SFILL7960x70050 (
);

FILL FILL_3__13368_ (
);

FILL FILL_2__8115_ (
);

FILL FILL_0__10503_ (
);

FILL SFILL59000x83050 (
);

FILL FILL_5__6960_ (
);

FILL FILL_6__14702_ (
);

FILL SFILL38120x42050 (
);

FILL SFILL3480x5050 (
);

FILL SFILL3560x69050 (
);

FILL SFILL59080x40050 (
);

OAI22X1 _13680_ (
    .A(_4186_),
    .B(_3893__bF$buf1),
    .C(_3967__bF$buf0),
    .D(_4187_),
    .Y(_4188_)
);

FILL FILL_0__13395_ (
);

NAND2X1 _13260_ (
    .A(_3750_),
    .B(_3775_),
    .Y(_3803_)
);

FILL SFILL38920x25050 (
);

FILL FILL_1__6952_ (
);

FILL FILL_4__9402_ (
);

FILL FILL_2__13722_ (
);

FILL FILL_2__13302_ (
);

FILL FILL_5__16167_ (
);

FILL FILL_3__6878_ (
);

FILL FILL_1__12715_ (
);

FILL FILL_2__16194_ (
);

FILL FILL_4__10295_ (
);

FILL FILL_0__9722_ (
);

FILL FILL_0__11708_ (
);

FILL FILL_1__15187_ (
);

FILL FILL_5__7745_ (
);

FILL SFILL113720x77050 (
);

FILL FILL_5__7325_ (
);

FILL FILL_4__16101_ (
);

INVX1 _14885_ (
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_5367_)
);

FILL SFILL49080x83050 (
);

INVX1 _14465_ (
    .A(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_4956_)
);

OAI22X1 _14045_ (
    .A(_3941_),
    .B(_4544_),
    .C(_3930__bF$buf0),
    .D(_4543_),
    .Y(_4545_)
);

FILL FILL_3__15934_ (
);

FILL FILL_3__15514_ (
);

FILL SFILL3560x24050 (
);

FILL FILL_1__7737_ (
);

FILL FILL_1__7317_ (
);

FILL FILL_2__14927_ (
);

FILL SFILL104440x41050 (
);

FILL FILL_2__14507_ (
);

FILL FILL_0__15961_ (
);

FILL FILL_0__15541_ (
);

FILL FILL_0__15121_ (
);

FILL FILL_5__12087_ (
);

FILL FILL112200x19050 (
);

FILL FILL_3__8604_ (
);

FILL FILL_4__12861_ (
);

FILL FILL_4__12441_ (
);

FILL FILL_4__12021_ (
);

INVX1 _10385_ (
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_1775_)
);

FILL SFILL49800x64050 (
);

FILL FILL_3__11854_ (
);

FILL FILL_3__11434_ (
);

FILL FILL_3__11014_ (
);

FILL SFILL28920x23050 (
);

FILL FILL_4__6947_ (
);

FILL FILL_0__16326_ (
);

FILL FILL_2__10427_ (
);

FILL FILL_0__11881_ (
);

FILL FILL_2__9493_ (
);

FILL FILL_2__10007_ (
);

FILL FILL_0__11461_ (
);

FILL FILL_0__11041_ (
);

FILL FILL_3__9809_ (
);

FILL FILL_5__14653_ (
);

FILL FILL_5__14233_ (
);

FILL FILL_0__6847_ (
);

INVX1 _8953_ (
    .A(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_1044_)
);

OAI21X1 _8533_ (
    .A(_844_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_845_),
    .Y(_783_[31])
);

OAI21X1 _8113_ (
    .A(_625_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_626_),
    .Y(_588_[19])
);

FILL FILL_1__7490_ (
);

FILL FILL_1__7070_ (
);

FILL FILL_4__13646_ (
);

FILL FILL_4__13226_ (
);

FILL FILL_2__14680_ (
);

FILL FILL_2__14260_ (
);

FILL FILL_2__7806_ (
);

FILL FILL_3__12639_ (
);

FILL FILL_1__13673_ (
);

FILL FILL_3__12219_ (
);

FILL FILL_1__13253_ (
);

FILL FILL_1_BUFX2_insert810 (
);

FILL FILL_1_BUFX2_insert811 (
);

FILL SFILL28440x16050 (
);

INVX1 _12951_ (
    .A(_2_[0]),
    .Y(_3683_)
);

FILL FILL_1_BUFX2_insert812 (
);

OAI21X1 _12531_ (
    .A(_3419_),
    .B(vdd),
    .C(_3420_),
    .Y(_3360_[30])
);

FILL FILL_0__12246_ (
);

FILL FILL_1_BUFX2_insert813 (
);

FILL FILL_1_BUFX2_insert814 (
);

NAND3X1 _12111_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[31]),
    .C(_3032__bF$buf1),
    .Y(_3129_)
);

FILL FILL_1_BUFX2_insert815 (
);

FILL FILL_1_BUFX2_insert816 (
);

FILL FILL_1_BUFX2_insert817 (
);

FILL FILL_1_BUFX2_insert818 (
);

FILL FILL_1_BUFX2_insert819 (
);

FILL FILL_5__15858_ (
);

FILL SFILL18520x52050 (
);

FILL SFILL73880x25050 (
);

FILL FILL_5__15438_ (
);

FILL FILL_5__15018_ (
);

OAI21X1 _9738_ (
    .A(_1444_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1445_),
    .Y(_1433_[6])
);

FILL FILL_3__16052_ (
);

DFFSR _9318_ (
    .Q(\datapath_1.regfile_1.regOut[19] [16]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_1173_[16])
);

FILL FILL_5__10993_ (
);

FILL FILL_5__10573_ (
);

FILL FILL_1__8695_ (
);

FILL FILL_5__10153_ (
);

FILL FILL_1__8275_ (
);

FILL FILL_2__15885_ (
);

FILL FILL_2__15465_ (
);

FILL FILL_2__15045_ (
);

FILL SFILL63960x61050 (
);

FILL SFILL94360x52050 (
);

FILL FILL_2__10180_ (
);

FILL FILL_1__14878_ (
);

FILL FILL_1__14458_ (
);

FILL FILL_1__14038_ (
);

FILL FILL_3__9982_ (
);

FILL FILL_3__9142_ (
);

AOI22X1 _13736_ (
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .B(_4102_),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_4243_)
);

NOR2X1 _13316_ (
    .A(_3790_),
    .B(_3847_),
    .Y(_3848_)
);

FILL FILL_5__9488_ (
);

FILL SFILL79160x32050 (
);

FILL FILL_0__14812_ (
);

FILL FILL_5__11778_ (
);

FILL FILL_5__11358_ (
);

FILL FILL_3__12392_ (
);

FILL FILL_4__7485_ (
);

FILL FILL_4__7065_ (
);

FILL SFILL18840x28050 (
);

FILL FILL_2__11385_ (
);

FILL FILL_1__10798_ (
);

FILL FILL_1__10378_ (
);

FILL FILL_4__11712_ (
);

FILL FILL_5__15191_ (
);

OAI21X1 _9491_ (
    .A(_1320_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1321_),
    .Y(_1303_[9])
);

DFFSR _9071_ (
    .Q(\datapath_1.regfile_1.regOut[17] [25]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_1043_[25])
);

FILL FILL_3__10705_ (
);

FILL FILL_4__14184_ (
);

FILL FILL_2__8764_ (
);

FILL FILL_3__13597_ (
);

FILL FILL_2__8344_ (
);

FILL FILL_0__10312_ (
);

FILL FILL_5__13924_ (
);

FILL FILL_5__13504_ (
);

FILL SFILL84360x50050 (
);

INVX1 _7804_ (
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_461_)
);

FILL FILL_4_BUFX2_insert320 (
);

FILL FILL_4_BUFX2_insert321 (
);

FILL FILL_4__9631_ (
);

FILL FILL_4_BUFX2_insert322 (
);

FILL FILL_4__12917_ (
);

FILL FILL_4__9211_ (
);

FILL FILL_4_BUFX2_insert323 (
);

FILL FILL_2__13951_ (
);

FILL FILL_4_BUFX2_insert324 (
);

FILL FILL_2__13531_ (
);

FILL FILL_5__16396_ (
);

FILL FILL_2__13111_ (
);

FILL FILL_4_BUFX2_insert325 (
);

FILL FILL_4_BUFX2_insert326 (
);

FILL FILL_4_BUFX2_insert327 (
);

FILL FILL_4_BUFX2_insert328 (
);

FILL FILL_4_BUFX2_insert329 (
);

FILL FILL_4__15389_ (
);

FILL FILL_1__12524_ (
);

FILL FILL_1__12104_ (
);

FILL FILL_2__9549_ (
);

FILL FILL_0__9531_ (
);

FILL FILL_0__11937_ (
);

FILL SFILL114520x76050 (
);

FILL FILL_0__9111_ (
);

FILL FILL_2__9129_ (
);

NAND3X1 _11802_ (
    .A(_2462__bF$buf0),
    .B(_2879_),
    .C(_2893_),
    .Y(_2894_)
);

FILL FILL_0__11517_ (
);

FILL SFILL53880x66050 (
);

FILL FILL_5__7974_ (
);

FILL FILL_5__7554_ (
);

FILL FILL_4__16330_ (
);

AOI22X1 _14694_ (
    .A(_3995__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[31] [26]),
    .C(\datapath_1.regfile_1.regOut[6] [26]),
    .D(_4001__bF$buf3),
    .Y(_5180_)
);

FILL FILL_6__10011_ (
);

AOI22X1 _14274_ (
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .B(_3942__bF$buf0),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_4769_)
);

FILL FILL_5__14709_ (
);

FILL FILL_3__15743_ (
);

FILL FILL_3__15323_ (
);

FILL FILL_1__7966_ (
);

FILL FILL_1__7546_ (
);

FILL SFILL69080x37050 (
);

FILL FILL_2__14736_ (
);

FILL FILL_2__14316_ (
);

FILL FILL_0__15770_ (
);

FILL FILL_0__15350_ (
);

FILL FILL_1__13729_ (
);

FILL FILL_1__13309_ (
);

FILL FILL_3__8833_ (
);

FILL FILL_5__8759_ (
);

FILL FILL_5__8339_ (
);

FILL SFILL114520x31050 (
);

OAI22X1 _15899_ (
    .A(_5530__bF$buf2),
    .B(_6357_),
    .C(_5532__bF$buf3),
    .D(_6356_),
    .Y(_6358_)
);

FILL FILL_6__11216_ (
);

OAI22X1 _15479_ (
    .A(_5948_),
    .B(_5545__bF$buf3),
    .C(_5485__bF$buf0),
    .D(_4445_),
    .Y(_5949_)
);

NAND3X1 _15059_ (
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5477_),
    .C(_5513_),
    .Y(_5539_)
);

FILL FILL_4__12250_ (
);

FILL SFILL3720x50050 (
);

FILL FILL_3__16108_ (
);

OAI21X1 _10194_ (
    .A(_1687_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .C(_1688_),
    .Y(_1628_[30])
);

FILL FILL_5__10629_ (
);

FILL FILL_3__11663_ (
);

FILL FILL_3__11243_ (
);

DFFSR _16420_ (
    .Q(\datapath_1.regfile_1.regOut[0] [3]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_6769_[3])
);

FILL FILL_0__16135_ (
);

OAI22X1 _16000_ (
    .A(_5495__bF$buf2),
    .B(_6456_),
    .C(_5080_),
    .D(_5534__bF$buf2),
    .Y(_6457_)
);

FILL FILL_2__10656_ (
);

FILL FILL_0__11690_ (
);

FILL FILL_2__10236_ (
);

FILL FILL_0__11270_ (
);

FILL FILL_3_BUFX2_insert340 (
);

FILL FILL_3__9618_ (
);

FILL FILL_3_BUFX2_insert341 (
);

FILL FILL_3_BUFX2_insert342 (
);

FILL FILL_5__14882_ (
);

FILL FILL_5__14462_ (
);

FILL FILL_3_BUFX2_insert343 (
);

FILL FILL_5__14042_ (
);

FILL FILL_3_BUFX2_insert344 (
);

OAI21X1 _8762_ (
    .A(_956_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_957_),
    .Y(_913_[22])
);

FILL FILL_3_BUFX2_insert345 (
);

FILL FILL_6__7203_ (
);

FILL FILL_3_BUFX2_insert346 (
);

OAI21X1 _8342_ (
    .A(_737_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_738_),
    .Y(_718_[10])
);

FILL FILL_3_BUFX2_insert347 (
);

FILL SFILL43880x64050 (
);

FILL FILL_3_BUFX2_insert348 (
);

FILL FILL_4__13875_ (
);

FILL FILL_3_BUFX2_insert349 (
);

FILL FILL_4__13455_ (
);

FILL FILL_4__13035_ (
);

INVX1 _11399_ (
    .A(_2214_),
    .Y(_2516_)
);

FILL SFILL7960x65050 (
);

FILL FILL_2__7615_ (
);

FILL FILL_3__12868_ (
);

FILL FILL_3__12448_ (
);

FILL SFILL59000x78050 (
);

FILL FILL_3__12028_ (
);

FILL FILL_1__13482_ (
);

FILL FILL_0__12895_ (
);

OAI21X1 _12760_ (
    .A(_3531_),
    .B(IRWrite_bF$buf1),
    .C(_3532_),
    .Y(_3490_[21])
);

FILL FILL_0__12475_ (
);

FILL FILL_0__12055_ (
);

NAND3X1 _12340_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf0),
    .Y(_3294_)
);

FILL FILL_5__8092_ (
);

FILL FILL_4__8902_ (
);

FILL FILL_5__15667_ (
);

FILL FILL_5__15247_ (
);

FILL FILL_3__16281_ (
);

DFFSR _9967_ (
    .Q(\datapath_1.regfile_1.regOut[24] [25]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_1498_[25])
);

NAND2X1 _9547_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1359_)
);

NAND2X1 _9127_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1140_)
);

FILL SFILL3640x12050 (
);

FILL FILL_5__10382_ (
);

FILL FILL_1__8084_ (
);

FILL SFILL64760x60050 (
);

FILL FILL_2__15694_ (
);

FILL FILL_2__15274_ (
);

FILL FILL_1__14687_ (
);

FILL FILL_1__14267_ (
);

FILL FILL_0_BUFX2_insert470 (
);

FILL FILL_0_BUFX2_insert471 (
);

FILL FILL_4__15601_ (
);

FILL FILL_0_BUFX2_insert472 (
);

FILL SFILL59000x33050 (
);

FILL FILL_3__9791_ (
);

FILL FILL_0_BUFX2_insert473 (
);

FILL SFILL49080x78050 (
);

FILL FILL_3__9371_ (
);

FILL FILL_0_BUFX2_insert474 (
);

INVX1 _13965_ (
    .A(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_4467_)
);

FILL FILL_0_BUFX2_insert475 (
);

INVX1 _13545_ (
    .A(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_4055_)
);

NAND2X1 _13125_ (
    .A(PCEn_bF$buf6),
    .B(\datapath_1.mux_pcsrc.dout [15]),
    .Y(_3715_)
);

FILL FILL_0_BUFX2_insert476 (
);

FILL FILL_0_BUFX2_insert477 (
);

FILL FILL_0_BUFX2_insert478 (
);

FILL SFILL3560x19050 (
);

FILL FILL_0_BUFX2_insert479 (
);

FILL FILL_5__9297_ (
);

FILL SFILL104440x36050 (
);

FILL FILL_0__14621_ (
);

FILL FILL_0__14201_ (
);

FILL FILL_5__11587_ (
);

FILL FILL_1__9289_ (
);

FILL FILL_5__11167_ (
);

FILL SFILL12920x64050 (
);

FILL FILL_2__16059_ (
);

FILL FILL_4__7294_ (
);

FILL SFILL33880x62050 (
);

FILL FILL_2__11194_ (
);

FILL FILL_1__10187_ (
);

FILL SFILL49000x76050 (
);

FILL FILL_4__11941_ (
);

FILL FILL_4__11521_ (
);

FILL FILL_4__11101_ (
);

FILL FILL_0__7194_ (
);

FILL SFILL49080x33050 (
);

FILL FILL_1__16413_ (
);

FILL FILL_3__10934_ (
);

FILL FILL_3__10514_ (
);

FILL SFILL28920x18050 (
);

FILL FILL_0__15826_ (
);

FILL FILL_0__15406_ (
);

FILL FILL_2__8993_ (
);

FILL FILL_0__10961_ (
);

FILL FILL_2__8573_ (
);

FILL FILL_0__10541_ (
);

FILL FILL_0__10121_ (
);

FILL SFILL115320x7050 (
);

FILL FILL_4__8499_ (
);

FILL SFILL49400x45050 (
);

FILL FILL_4__8079_ (
);

FILL FILL_2__12399_ (
);

FILL FILL_5__13733_ (
);

FILL FILL_5__13313_ (
);

OAI21X1 _7613_ (
    .A(_373_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_374_),
    .Y(_328_[23])
);

FILL FILL_1__6990_ (
);

FILL FILL_4__9860_ (
);

FILL FILL_4__9020_ (
);

FILL FILL_4__12726_ (
);

FILL FILL_2__13760_ (
);

FILL FILL_4__12306_ (
);

FILL FILL_2__13340_ (
);

FILL FILL_0__8399_ (
);

FILL SFILL49000x31050 (
);

FILL SFILL114600x9050 (
);

FILL SFILL39080x76050 (
);

FILL FILL_3__11719_ (
);

FILL FILL_1__12753_ (
);

FILL FILL_4__15198_ (
);

FILL FILL_1__12333_ (
);

FILL FILL_0__9760_ (
);

FILL FILL_2__9778_ (
);

FILL FILL_2__9358_ (
);

FILL FILL_0__11746_ (
);

FILL FILL_0__9340_ (
);

FILL FILL_0__11326_ (
);

OAI21X1 _11611_ (
    .A(_2716_),
    .B(_2458_),
    .C(_2714_),
    .Y(_2717_)
);

FILL FILL_6__15945_ (
);

FILL FILL_5__7363_ (
);

FILL FILL_5__14938_ (
);

OAI22X1 _14083_ (
    .A(_4581_),
    .B(_3890_),
    .C(_3944__bF$buf4),
    .D(_4580_),
    .Y(_4582_)
);

FILL FILL_3__15972_ (
);

FILL FILL_5__14518_ (
);

FILL FILL_3__15552_ (
);

DFFSR _8818_ (
    .Q(\datapath_1.regfile_1.regOut[15] [28]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_913_[28])
);

FILL FILL_3__15132_ (
);

FILL FILL_1__7355_ (
);

FILL FILL_2__14965_ (
);

FILL FILL111800x76050 (
);

FILL FILL_2__14545_ (
);

FILL FILL_2__14125_ (
);

FILL SFILL39000x74050 (
);

FILL SFILL94360x47050 (
);

FILL FILL_1__13958_ (
);

FILL FILL_1__13538_ (
);

FILL FILL_1__13118_ (
);

FILL SFILL39080x31050 (
);

FILL FILL_3__8642_ (
);

DFFSR _12816_ (
    .Q(\datapath_1.PCJump [27]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3490_[25])
);

FILL FILL_3__8222_ (
);

FILL FILL_5__8988_ (
);

FILL FILL_5__8568_ (
);

FILL FILL_5__8148_ (
);

FILL FILL_6__11865_ (
);

OAI22X1 _15288_ (
    .A(_5527__bF$buf3),
    .B(_4195_),
    .C(_5762_),
    .D(_5532__bF$buf1),
    .Y(_5763_)
);

FILL SFILL39400x43050 (
);

FILL FILL_3__16337_ (
);

FILL FILL_5__10438_ (
);

FILL FILL_3__11892_ (
);

FILL FILL_5__10018_ (
);

FILL FILL_3__11472_ (
);

FILL FILL_3__11052_ (
);

FILL FILL_4__6985_ (
);

FILL FILL_0__16364_ (
);

FILL FILL_2__10885_ (
);

FILL FILL_2__10045_ (
);

FILL FILL_1__9921_ (
);

FILL FILL_1__9501_ (
);

FILL FILL_3__9847_ (
);

FILL FILL_3__9427_ (
);

FILL FILL_3__9007_ (
);

FILL FILL_5__14691_ (
);

FILL FILL_0__6885_ (
);

FILL FILL_5__14271_ (
);

OAI21X1 _8991_ (
    .A(_1068_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1069_),
    .Y(_1043_[13])
);

OAI21X1 _8571_ (
    .A(_849_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .C(_850_),
    .Y(_848_[1])
);

FILL FILL111960x5050 (
);

DFFSR _8151_ (
    .Q(\datapath_1.regfile_1.regOut[10] [1]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_588_[1])
);

FILL FILL_4__13684_ (
);

FILL FILL_4__13264_ (
);

FILL SFILL8760x64050 (
);

FILL FILL111720x38050 (
);

FILL FILL_2__7844_ (
);

FILL FILL_2__7424_ (
);

FILL FILL_3__12257_ (
);

FILL FILL_1__13291_ (
);

FILL FILL_0__12284_ (
);

FILL SFILL114600x64050 (
);

FILL SFILL53960x54050 (
);

FILL SFILL84360x45050 (
);

FILL FILL_6__16063_ (
);

FILL FILL_4__8711_ (
);

FILL FILL_5__15896_ (
);

FILL FILL_2__12611_ (
);

FILL FILL_5__15476_ (
);

FILL FILL_5__15056_ (
);

FILL FILL_3__16090_ (
);

NAND2X1 _9776_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1471_)
);

NAND2X1 _9356_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1252_)
);

FILL FILL_5__10191_ (
);

FILL FILL_4__14889_ (
);

FILL FILL_4__14469_ (
);

FILL FILL_1__11604_ (
);

FILL FILL_4__14049_ (
);

FILL FILL_2__15083_ (
);

FILL FILL_2__8629_ (
);

FILL FILL_0__8611_ (
);

FILL FILL_2__8209_ (
);

FILL FILL_1__14496_ (
);

FILL FILL_1__14076_ (
);

FILL FILL_4__15830_ (
);

FILL FILL_4__15410_ (
);

INVX1 _13774_ (
    .A(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_4280_)
);

FILL FILL_0__13489_ (
);

OR2X2 _13354_ (
    .A(_3870_),
    .B(_3843_),
    .Y(_3871_)
);

FILL FILL_3__14823_ (
);

FILL FILL_3__14403_ (
);

FILL FILL_4__9916_ (
);

FILL FILL_2__13816_ (
);

FILL FILL_0__14850_ (
);

FILL FILL_0__14430_ (
);

FILL FILL_0__14010_ (
);

FILL FILL_5__11396_ (
);

FILL FILL_1__9098_ (
);

FILL FILL_2__16288_ (
);

FILL FILL_4__10389_ (
);

FILL FILL_5__7839_ (
);

FILL SFILL114520x26050 (
);

FILL FILL_5__7419_ (
);

INVX8 _14979_ (
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_5459_)
);

NAND3X1 _14559_ (
    .A(_5046_),
    .B(_5047_),
    .C(_5045_),
    .Y(_5048_)
);

FILL FILL_4__11750_ (
);

INVX1 _14139_ (
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_4637_)
);

FILL FILL_4__11330_ (
);

FILL FILL_3__15608_ (
);

FILL FILL_1__16222_ (
);

FILL FILL_3__10743_ (
);

FILL SFILL43960x52050 (
);

FILL FILL_3__10323_ (
);

FILL SFILL19000x70050 (
);

OAI22X1 _15920_ (
    .A(_6378_),
    .B(_5518__bF$buf2),
    .C(_5478__bF$buf1),
    .D(_4966_),
    .Y(_6379_)
);

FILL FILL_0__15635_ (
);

FILL FILL_0__15215_ (
);

NOR2X1 _15500_ (
    .A(_5967_),
    .B(_5968_),
    .Y(_5969_)
);

FILL FILL_2__8382_ (
);

FILL FILL_0__10770_ (
);

FILL FILL_5__13962_ (
);

FILL FILL_5__13542_ (
);

FILL FILL_5__13122_ (
);

OAI21X1 _7842_ (
    .A(_485_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .C(_486_),
    .Y(_458_[14])
);

FILL SFILL104520x69050 (
);

OAI21X1 _7422_ (
    .A(_266_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .C(_267_),
    .Y(_263_[2])
);

FILL SFILL43880x59050 (
);

DFFSR _7002_ (
    .Q(\datapath_1.regfile_1.regOut[1] [4]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_3_[4])
);

FILL FILL_4_BUFX2_insert700 (
);

FILL FILL_4_BUFX2_insert701 (
);

FILL FILL_4_BUFX2_insert702 (
);

FILL FILL_4__12955_ (
);

FILL FILL_4_BUFX2_insert703 (
);

FILL FILL_4__12115_ (
);

FILL FILL_4_BUFX2_insert704 (
);

FILL FILL_4_BUFX2_insert705 (
);

INVX1 _10899_ (
    .A(\control_1.reg_state.dout [1]),
    .Y(_2048_)
);

FILL FILL_4_BUFX2_insert706 (
);

FILL FILL_4_BUFX2_insert707 (
);

DFFSR _10479_ (
    .Q(\datapath_1.regfile_1.regOut[28] [25]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_1758_[25])
);

NAND2X1 _10059_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1619_)
);

FILL FILL_4_BUFX2_insert708 (
);

FILL FILL_3__11948_ (
);

FILL FILL_4_BUFX2_insert709 (
);

FILL FILL_1__12982_ (
);

FILL FILL_3__11528_ (
);

FILL FILL_3__11108_ (
);

FILL FILL_1__12142_ (
);

FILL FILL112280x63050 (
);

FILL FILL_0__11975_ (
);

FILL FILL_2__9167_ (
);

OAI21X1 _11840_ (
    .A(_2928_),
    .B(_2337_),
    .C(_2925_),
    .Y(_2929_)
);

FILL FILL_0__11555_ (
);

NAND3X1 _11420_ (
    .A(_2462__bF$buf2),
    .B(_2535_),
    .C(_2530_),
    .Y(_2536_)
);

FILL FILL_0__11135_ (
);

NOR2X1 _11000_ (
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2118_),
    .Y(_2119_)
);

FILL FILL_5__7592_ (
);

FILL FILL_5__7172_ (
);

FILL FILL_5__14747_ (
);

FILL FILL_3__15781_ (
);

FILL FILL_5__14327_ (
);

FILL FILL_3__15361_ (
);

NAND2X1 _8627_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_888_)
);

NAND2X1 _8207_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_669_)
);

FILL FILL_1__7584_ (
);

FILL FILL_1__7164_ (
);

FILL FILL_2__14774_ (
);

FILL SFILL104520x24050 (
);

FILL FILL_2__14354_ (
);

FILL SFILL43880x14050 (
);

FILL SFILL68280x80050 (
);

FILL FILL_1__13767_ (
);

FILL FILL_1__13347_ (
);

FILL FILL_3__8871_ (
);

FILL FILL_3__8451_ (
);

NAND2X1 _12625_ (
    .A(vdd),
    .B(memoryOutData[19]),
    .Y(_3463_)
);

INVX1 _12205_ (
    .A(\datapath_1.PCJump [30]),
    .Y(_3190_)
);

FILL SFILL84280x1050 (
);

FILL FILL_5__8377_ (
);

FILL FILL_6__16119_ (
);

INVX8 _15097_ (
    .A(_5463__bF$buf0),
    .Y(_5576_)
);

FILL FILL_0__13701_ (
);

FILL FILL_3__16146_ (
);

FILL FILL_5__10667_ (
);

FILL FILL_1__8789_ (
);

FILL FILL_1__8369_ (
);

FILL FILL_5__10247_ (
);

FILL FILL_3__11281_ (
);

FILL FILL_2__15979_ (
);

FILL FILL_2__15559_ (
);

FILL FILL_2__15139_ (
);

FILL FILL_0__16173_ (
);

FILL FILL_2__10694_ (
);

FILL FILL_2__10274_ (
);

FILL FILL_1__9730_ (
);

FILL FILL_3__9656_ (
);

FILL FILL_3_BUFX2_insert720 (
);

FILL FILL_3_BUFX2_insert721 (
);

FILL FILL_3__9236_ (
);

FILL FILL_3_BUFX2_insert722 (
);

FILL FILL_3_BUFX2_insert723 (
);

FILL FILL_3_BUFX2_insert724 (
);

FILL FILL_5__14080_ (
);

FILL FILL_1__15913_ (
);

FILL FILL_3_BUFX2_insert725 (
);

FILL FILL_3_BUFX2_insert726 (
);

NAND2X1 _8380_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_764_)
);

FILL FILL_3_BUFX2_insert727 (
);

FILL FILL_3_BUFX2_insert728 (
);

FILL FILL_6__12459_ (
);

FILL FILL_3_BUFX2_insert729 (
);

FILL FILL_6__12039_ (
);

FILL FILL_4__13493_ (
);

FILL FILL_0__14906_ (
);

FILL FILL_3__12486_ (
);

FILL FILL_2__7233_ (
);

FILL FILL_3__12066_ (
);

FILL FILL_4__7999_ (
);

FILL FILL_4__7579_ (
);

FILL FILL_4__7159_ (
);

FILL FILL_2__11899_ (
);

FILL FILL_2__11479_ (
);

FILL FILL_2__11059_ (
);

FILL FILL_0__12093_ (
);

FILL SFILL33880x12050 (
);

FILL FILL_4__8520_ (
);

FILL FILL_4__8100_ (
);

FILL FILL_4__11806_ (
);

FILL FILL_2__12840_ (
);

FILL FILL_2__12420_ (
);

FILL FILL_5__15285_ (
);

FILL SFILL49000x26050 (
);

FILL FILL_0__7479_ (
);

FILL FILL_2__12000_ (
);

DFFSR _9585_ (
    .Q(\datapath_1.regfile_1.regOut[21] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_1303_[27])
);

FILL FILL_0__7059_ (
);

INVX1 _9165_ (
    .A(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_1165_)
);

FILL FILL_4__14698_ (
);

FILL FILL_1__11833_ (
);

FILL FILL_4__14278_ (
);

FILL FILL_1__11413_ (
);

FILL SFILL94440x35050 (
);

FILL FILL_0__8840_ (
);

FILL FILL_2__8858_ (
);

FILL FILL_0__10826_ (
);

FILL FILL_2__8438_ (
);

FILL FILL_0__10406_ (
);

FILL FILL_0__8000_ (
);

FILL FILL_2__8018_ (
);

FILL FILL_6__14605_ (
);

FILL FILL_5__6863_ (
);

FILL FILL_0_BUFX2_insert850 (
);

FILL FILL_0_BUFX2_insert851 (
);

FILL FILL_0_BUFX2_insert852 (
);

FILL FILL_0_BUFX2_insert853 (
);

FILL FILL_0_BUFX2_insert854 (
);

FILL FILL_0__13298_ (
);

FILL FILL_0_BUFX2_insert855 (
);

NOR2X1 _13583_ (
    .A(_4081_),
    .B(_4092_),
    .Y(_4093_)
);

FILL FILL_0_BUFX2_insert856 (
);

INVX1 _13163_ (
    .A(\datapath_1.PCJump [28]),
    .Y(_3740_)
);

FILL SFILL23880x55050 (
);

FILL FILL_0_BUFX2_insert857 (
);

FILL FILL_3__14632_ (
);

FILL FILL_0_BUFX2_insert858 (
);

FILL FILL_3__14212_ (
);

FILL FILL_0_BUFX2_insert859 (
);

FILL FILL_1__6855_ (
);

FILL FILL_4__9725_ (
);

FILL FILL_2__13625_ (
);

FILL SFILL39000x69050 (
);

FILL FILL_1__12618_ (
);

FILL FILL_2__16097_ (
);

FILL FILL_0__9625_ (
);

FILL FILL_3__7722_ (
);

FILL FILL_3__7302_ (
);

FILL SFILL79640x8050 (
);

FILL FILL_5__7228_ (
);

FILL FILL_4__16004_ (
);

NOR2X1 _14788_ (
    .A(_5270_),
    .B(_5272_),
    .Y(_5273_)
);

INVX1 _14368_ (
    .A(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_4861_)
);

FILL SFILL23800x53050 (
);

FILL FILL_3__15837_ (
);

FILL FILL_3__15417_ (
);

FILL FILL_1__16451_ (
);

FILL FILL_1__16031_ (
);

FILL SFILL79320x2050 (
);

FILL FILL_3__10972_ (
);

FILL SFILL23880x10050 (
);

FILL FILL_3__10552_ (
);

FILL FILL_3__10132_ (
);

FILL FILL_0__15864_ (
);

FILL SFILL79240x7050 (
);

FILL FILL_0__15444_ (
);

FILL FILL_6_BUFX2_insert234 (
);

FILL FILL_0__15024_ (
);

FILL SFILL53960x3050 (
);

FILL FILL_2__8191_ (
);

FILL FILL_6_BUFX2_insert239 (
);

BUFX2 BUFX2_insert10 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf2 )
);

BUFX2 BUFX2_insert11 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf1 )
);

BUFX2 BUFX2_insert12 (
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf0 )
);

BUFX2 BUFX2_insert13 (
    .A(_5469_),
    .Y(_5469__bF$buf3)
);

BUFX2 BUFX2_insert14 (
    .A(_5469_),
    .Y(_5469__bF$buf2)
);

FILL FILL_3__8507_ (
);

BUFX2 BUFX2_insert15 (
    .A(_5469_),
    .Y(_5469__bF$buf1)
);

BUFX2 BUFX2_insert16 (
    .A(_5469_),
    .Y(_5469__bF$buf0)
);

FILL FILL_5__13771_ (
);

BUFX2 BUFX2_insert17 (
    .A(_3955_),
    .Y(_3955__bF$buf4)
);

FILL FILL_5__13351_ (
);

BUFX2 BUFX2_insert18 (
    .A(_3955_),
    .Y(_3955__bF$buf3)
);

BUFX2 BUFX2_insert19 (
    .A(_3955_),
    .Y(_3955__bF$buf2)
);

DFFSR _7651_ (
    .Q(\datapath_1.regfile_1.regOut[6] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_328_[13])
);

NAND2X1 _7231_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_181_)
);

FILL FILL_4__12764_ (
);

FILL SFILL8760x59050 (
);

FILL FILL_4__12344_ (
);

NAND2X1 _10288_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1731_)
);

FILL FILL_2__6924_ (
);

FILL FILL_3__11757_ (
);

FILL SFILL13880x53050 (
);

FILL FILL_3__11337_ (
);

FILL FILL_1__12371_ (
);

FILL FILL_0__16229_ (
);

FILL FILL_2__9396_ (
);

FILL FILL_0__11784_ (
);

FILL FILL_0__11364_ (
);

FILL SFILL53960x49050 (
);

FILL SFILL74120x50 (
);

FILL FILL_5__14976_ (
);

FILL SFILL103960x3050 (
);

FILL FILL_5__14556_ (
);

FILL FILL_5__14136_ (
);

FILL FILL_3__15590_ (
);

FILL FILL_3__15170_ (
);

NAND2X1 _8856_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1000_)
);

DFFSR _8436_ (
    .Q(\datapath_1.regfile_1.regOut[12] [30]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_718_[30])
);

INVX1 _8016_ (
    .A(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_582_)
);

FILL FILL_4__13969_ (
);

FILL FILL_4__13549_ (
);

FILL FILL_2__14583_ (
);

FILL FILL_4__13129_ (
);

FILL FILL_2__14163_ (
);

FILL SFILL48920x50 (
);

FILL FILL_2__7709_ (
);

FILL SFILL13800x51050 (
);

FILL FILL_1__13996_ (
);

FILL FILL_1__13576_ (
);

FILL FILL_1__13156_ (
);

FILL FILL_4__14910_ (
);

FILL FILL_0__12989_ (
);

FILL FILL_0__12569_ (
);

FILL FILL_3__8260_ (
);

NAND2X1 _12854_ (
    .A(vdd),
    .B(\datapath_1.rd1 [10]),
    .Y(_3575_)
);

NAND2X1 _12434_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [30]),
    .Y(_3355_)
);

FILL FILL_0__12149_ (
);

NAND3X1 _12014_ (
    .A(_3054_),
    .B(_3055_),
    .C(_3056_),
    .Y(\datapath_1.mux_pcsrc.dout [6])
);

FILL FILL_3__13903_ (
);

FILL FILL_5__8186_ (
);

FILL FILL_5_BUFX2_insert250 (
);

FILL FILL_5_BUFX2_insert251 (
);

FILL FILL_5_BUFX2_insert252 (
);

FILL FILL_0__13930_ (
);

FILL FILL_5_BUFX2_insert253 (
);

FILL FILL_3__16375_ (
);

FILL FILL_0__13510_ (
);

FILL FILL_5_BUFX2_insert254 (
);

FILL FILL_5_BUFX2_insert255 (
);

FILL FILL_5__10896_ (
);

FILL FILL_5_BUFX2_insert256 (
);

FILL FILL_1__8598_ (
);

FILL FILL_5_BUFX2_insert257 (
);

FILL FILL_5__10056_ (
);

FILL FILL_5_BUFX2_insert1040 (
);

FILL FILL_5_BUFX2_insert1041 (
);

FILL FILL_5_BUFX2_insert258 (
);

FILL FILL_3__11090_ (
);

FILL FILL_5_BUFX2_insert1042 (
);

FILL FILL_5_BUFX2_insert259 (
);

FILL FILL_2__15788_ (
);

FILL FILL_5_BUFX2_insert1043 (
);

FILL FILL_2__15368_ (
);

FILL FILL_5_BUFX2_insert1044 (
);

FILL FILL_5_BUFX2_insert1045 (
);

FILL FILL_5_BUFX2_insert1046 (
);

FILL FILL_5_BUFX2_insert1047 (
);

FILL FILL_5_BUFX2_insert1048 (
);

FILL FILL_5_BUFX2_insert1049 (
);

FILL FILL_5__6919_ (
);

FILL FILL_3__9885_ (
);

FILL FILL_3__9465_ (
);

FILL FILL_4__10830_ (
);

INVX1 _13639_ (
    .A(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_4147_)
);

FILL FILL_3__9045_ (
);

AOI21X1 _13219_ (
    .A(_3761_),
    .B(_3756_),
    .C(_3750_),
    .Y(_3762_)
);

FILL FILL_4__10410_ (
);

FILL FILL_6__7890_ (
);

FILL FILL_1__15722_ (
);

FILL FILL_1__15302_ (
);

FILL SFILL104600x57050 (
);

FILL FILL_0__14715_ (
);

FILL FILL_2__7882_ (
);

FILL FILL_2__7462_ (
);

FILL FILL_2__7042_ (
);

FILL FILL_3__12295_ (
);

FILL SFILL108920x65050 (
);

FILL FILL112360x51050 (
);

FILL FILL_2__11288_ (
);

FILL FILL_5__12622_ (
);

FILL FILL_5__12202_ (
);

OAI21X1 _6922_ (
    .A(_14_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_15_),
    .Y(_3_[6])
);

FILL FILL_2_BUFX2_insert380 (
);

FILL FILL_2_BUFX2_insert381 (
);

FILL FILL_2_BUFX2_insert382 (
);

FILL FILL_2_BUFX2_insert383 (
);

FILL FILL_2_BUFX2_insert384 (
);

FILL FILL_4__11615_ (
);

FILL FILL_2_BUFX2_insert385 (
);

FILL SFILL23880x7050 (
);

FILL FILL_2_BUFX2_insert386 (
);

FILL FILL_5__15094_ (
);

FILL FILL_0__7288_ (
);

FILL FILL_2_BUFX2_insert387 (
);

FILL FILL_2_BUFX2_insert388 (
);

INVX1 _9394_ (
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_1277_)
);

FILL FILL_2_BUFX2_insert389 (
);

FILL FILL_1__11642_ (
);

FILL FILL_1__11222_ (
);

FILL FILL_4__14087_ (
);

FILL FILL112280x58050 (
);

FILL FILL_0__10635_ (
);

FILL FILL_2__8247_ (
);

NOR2X1 _10920_ (
    .A(_2053_),
    .B(_2051_),
    .Y(MemToReg)
);

OAI21X1 _10500_ (
    .A(_1830_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .C(_1831_),
    .Y(_1823_[4])
);

NOR2X1 _13392_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3904_)
);

FILL FILL_5__13827_ (
);

FILL FILL_3__14861_ (
);

FILL FILL_5__13407_ (
);

FILL FILL_3__14441_ (
);

FILL FILL_3__14021_ (
);

NAND2X1 _7707_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_417_)
);

FILL FILL_4__9534_ (
);

FILL FILL_4__9114_ (
);

FILL FILL_2__13854_ (
);

FILL FILL_2__13434_ (
);

FILL FILL_5__16299_ (
);

FILL FILL_2__13014_ (
);

FILL SFILL24280x40050 (
);

FILL FILL_1__12847_ (
);

FILL FILL_1__12427_ (
);

FILL FILL_1__12007_ (
);

FILL FILL_3__7951_ (
);

FILL FILL_0__9854_ (
);

FILL FILL_0__9014_ (
);

FILL FILL_3__7111_ (
);

OAI21X1 _11705_ (
    .A(_2803_),
    .B(_2188_),
    .C(_2462__bF$buf3),
    .Y(_2804_)
);

FILL FILL112280x13050 (
);

FILL FILL_5__7877_ (
);

FILL FILL_5__7457_ (
);

FILL FILL_4__16233_ (
);

FILL FILL_5__7037_ (
);

AOI21X1 _14597_ (
    .A(_5085_),
    .B(_5059_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [23])
);

INVX1 _14177_ (
    .A(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_4674_)
);

FILL FILL_3__15646_ (
);

FILL FILL_3__15226_ (
);

FILL FILL_1__16260_ (
);

FILL FILL_1__7869_ (
);

FILL FILL_1__7449_ (
);

FILL FILL_3__10781_ (
);

FILL FILL_3__10361_ (
);

FILL SFILL94520x68050 (
);

FILL FILL_2__14639_ (
);

FILL FILL_0__15673_ (
);

FILL FILL_2__14219_ (
);

FILL FILL_0__15253_ (
);

FILL FILL_3__8736_ (
);

FILL SFILL98840x76050 (
);

FILL FILL_3__8316_ (
);

FILL FILL_5__13580_ (
);

FILL FILL_5__13160_ (
);

NAND2X1 _7880_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_512_)
);

NAND2X1 _7460_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_293_)
);

NAND2X1 _7040_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_74_)
);

FILL FILL_4__12993_ (
);

FILL FILL_4__12573_ (
);

FILL FILL_4__12153_ (
);

DFFSR _10097_ (
    .Q(\datapath_1.regfile_1.regOut[25] [27]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1563_[27])
);

FILL FILL_3__11986_ (
);

FILL FILL_5__9603_ (
);

FILL FILL_3__11566_ (
);

FILL FILL_3__11146_ (
);

FILL FILL_1__12180_ (
);

FILL FILL_0__16038_ (
);

OAI21X1 _16323_ (
    .A(_6832_),
    .B(gnd),
    .C(_6833_),
    .Y(_6769_[0])
);

FILL FILL_2__10979_ (
);

FILL FILL_2__10559_ (
);

FILL FILL_0__11593_ (
);

FILL FILL_2__10139_ (
);

FILL FILL_0__11173_ (
);

FILL FILL_6__15792_ (
);

FILL FILL_6__15372_ (
);

FILL FILL_4__7600_ (
);

FILL FILL_2__11920_ (
);

FILL FILL_5__14785_ (
);

FILL FILL_5__14365_ (
);

FILL FILL_2__11500_ (
);

FILL FILL_0__6979_ (
);

DFFSR _8665_ (
    .Q(\datapath_1.regfile_1.regOut[14] [3]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_848_[3])
);

INVX1 _8245_ (
    .A(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_694_)
);

FILL FILL_1__10913_ (
);

FILL FILL_4__13778_ (
);

FILL FILL_4__13358_ (
);

FILL FILL_2__14392_ (
);

FILL FILL_2__7938_ (
);

FILL FILL_0__7500_ (
);

FILL FILL_1__13385_ (
);

DFFSR _12663_ (
    .Q(\datapath_1.Data [0]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[0])
);

FILL FILL_0__12378_ (
);

NAND3X1 _12243_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3221_)
);

FILL FILL_3__13712_ (
);

FILL SFILL59080x2050 (
);

FILL FILL_6__11292_ (
);

FILL FILL_2__12705_ (
);

FILL FILL_3__16184_ (
);

FILL FILL_5__10285_ (
);

FILL FILL_2__15597_ (
);

FILL FILL_2__15177_ (
);

FILL FILL_0__8705_ (
);

FILL SFILL23000x65050 (
);

FILL FILL_4__15924_ (
);

FILL FILL_4__15504_ (
);

OAI22X1 _13868_ (
    .A(_4371_),
    .B(_3949_),
    .C(_3983__bF$buf0),
    .D(_4370_),
    .Y(_4372_)
);

FILL FILL_3__9274_ (
);

NAND3X1 _13448_ (
    .A(_3898_),
    .B(_3904_),
    .C(_3883_),
    .Y(_3960_)
);

OAI21X1 _13028_ (
    .A(_3669_),
    .B(vdd),
    .C(_3670_),
    .Y(_3620_[25])
);

FILL SFILL109480x3050 (
);

FILL FILL_3__14917_ (
);

FILL FILL_1__15951_ (
);

FILL FILL_1__15531_ (
);

FILL FILL_1__15111_ (
);

FILL FILL_0__14944_ (
);

FILL FILL_0__14524_ (
);

FILL FILL_0__14104_ (
);

FILL FILL_2__7691_ (
);

FILL SFILL39000x19050 (
);

FILL FILL_4__7197_ (
);

FILL FILL_2__11097_ (
);

FILL FILL_5__12851_ (
);

FILL FILL_5__12431_ (
);

FILL FILL_5__12011_ (
);

FILL FILL_4__11844_ (
);

FILL SFILL13080x65050 (
);

FILL FILL_4__11424_ (
);

FILL FILL_4__11004_ (
);

FILL FILL_0__7097_ (
);

FILL FILL_1__16316_ (
);

FILL SFILL13880x48050 (
);

FILL FILL_3__10837_ (
);

FILL FILL_1__11871_ (
);

FILL FILL_3__10417_ (
);

FILL SFILL88760x36050 (
);

FILL FILL_1__11451_ (
);

FILL FILL_1__11031_ (
);

FILL FILL_0__15729_ (
);

FILL FILL_0__15309_ (
);

FILL FILL_2__8896_ (
);

FILL FILL_2__8476_ (
);

FILL FILL_0__10444_ (
);

FILL FILL_2__8056_ (
);

FILL FILL_0__10024_ (
);

FILL SFILL74120x50050 (
);

FILL FILL_5__13636_ (
);

FILL FILL_5__13216_ (
);

FILL FILL_3__14670_ (
);

NAND2X1 _7936_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_529_)
);

FILL FILL_3__14250_ (
);

DFFSR _7516_ (
    .Q(\datapath_1.regfile_1.regOut[5] [6]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_263_[6])
);

FILL FILL_1__6893_ (
);

FILL FILL_4__9763_ (
);

FILL FILL_4__9343_ (
);

FILL FILL_4__12629_ (
);

FILL FILL_2__13663_ (
);

FILL FILL_4__12209_ (
);

FILL FILL_2__13243_ (
);

FILL SFILL13800x46050 (
);

FILL FILL_1__12656_ (
);

FILL FILL_1__12236_ (
);

FILL FILL_0__9663_ (
);

FILL FILL_3__7760_ (
);

OAI21X1 _11934_ (
    .A(_2996_),
    .B(IorD_bF$buf0),
    .C(_2997_),
    .Y(_1_[15])
);

FILL FILL_0__9243_ (
);

FILL FILL_3__7340_ (
);

FILL FILL_0__11649_ (
);

FILL FILL_0__11229_ (
);

OAI21X1 _11514_ (
    .A(_2625_),
    .B(_2624_),
    .C(_2623_),
    .Y(_2626_)
);

FILL FILL_6__15848_ (
);

FILL FILL_5__7686_ (
);

FILL FILL_4__16042_ (
);

FILL FILL_6__10563_ (
);

FILL FILL_3__15875_ (
);

FILL FILL_3__15455_ (
);

FILL FILL_3__15035_ (
);

FILL FILL_1__7678_ (
);

FILL FILL_3__10170_ (
);

FILL FILL_2__14868_ (
);

FILL FILL_6_BUFX2_insert613 (
);

FILL FILL_2__14448_ (
);

FILL FILL_2__14028_ (
);

FILL FILL_0__15482_ (
);

FILL FILL_0__15062_ (
);

FILL FILL_6_BUFX2_insert618 (
);

FILL FILL_3__8965_ (
);

FILL FILL_3__8125_ (
);

INVX1 _12719_ (
    .A(\datapath_1.PCJump [10]),
    .Y(_3505_)
);

FILL FILL_6__6970_ (
);

FILL FILL_1__14802_ (
);

FILL FILL_1_BUFX2_insert70 (
);

FILL FILL_1_BUFX2_insert71 (
);

FILL FILL_1_BUFX2_insert72 (
);

FILL FILL_6__11768_ (
);

FILL FILL_1_BUFX2_insert73 (
);

FILL FILL_1_BUFX2_insert74 (
);

FILL FILL_4__12382_ (
);

FILL FILL_1_BUFX2_insert75 (
);

FILL SFILL99240x61050 (
);

FILL FILL_1_BUFX2_insert76 (
);

FILL FILL_1_BUFX2_insert77 (
);

FILL FILL_1_BUFX2_insert78 (
);

FILL FILL_1_BUFX2_insert79 (
);

FILL FILL_2__6962_ (
);

FILL FILL_3__11795_ (
);

FILL FILL_5__9412_ (
);

FILL FILL_3__11375_ (
);

FILL FILL_4__6888_ (
);

FILL FILL_0__16267_ (
);

NAND2X1 _16132_ (
    .A(\datapath_1.regfile_1.regOut[7] [27]),
    .B(_5490_),
    .Y(_6585_)
);

FILL FILL112360x46050 (
);

FILL FILL_2__10788_ (
);

FILL FILL_2__10368_ (
);

FILL FILL_5__11702_ (
);

FILL FILL_1__9404_ (
);

FILL SFILL68760x77050 (
);

FILL SFILL64040x55050 (
);

FILL FILL_5__14594_ (
);

FILL FILL_5__14174_ (
);

INVX1 _8894_ (
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_1025_)
);

INVX1 _8474_ (
    .A(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_806_)
);

INVX1 _8054_ (
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_651_)
);

FILL FILL_4__13587_ (
);

FILL FILL_1__10302_ (
);

FILL FILL_4__13167_ (
);

FILL FILL_2__7747_ (
);

FILL FILL_2__7327_ (
);

FILL FILL_6__13914_ (
);

FILL SFILL114600x50 (
);

INVX1 _12892_ (
    .A(\datapath_1.a [23]),
    .Y(_3600_)
);

FILL FILL_0__12187_ (
);

INVX1 _12472_ (
    .A(ALUOut[11]),
    .Y(_3381_)
);

NAND3X1 _12052_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [16]),
    .C(_3034__bF$buf3),
    .Y(_3085_)
);

FILL FILL_5__12907_ (
);

FILL FILL_3__13941_ (
);

FILL FILL_3__13521_ (
);

FILL FILL_3__13101_ (
);

FILL FILL_4__8614_ (
);

FILL FILL_5_BUFX2_insert630 (
);

FILL FILL_5__15799_ (
);

FILL FILL_5_BUFX2_insert631 (
);

FILL FILL_5_BUFX2_insert632 (
);

FILL FILL_5__15379_ (
);

FILL FILL_2__12514_ (
);

FILL FILL_5_BUFX2_insert633 (
);

FILL FILL_5_BUFX2_insert634 (
);

OAI21X1 _9679_ (
    .A(_1425_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1426_),
    .Y(_1368_[29])
);

FILL FILL_5_BUFX2_insert635 (
);

OAI21X1 _9259_ (
    .A(_1206_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1207_),
    .Y(_1173_[17])
);

FILL FILL_5_BUFX2_insert636 (
);

FILL SFILL64040x10050 (
);

FILL FILL_5_BUFX2_insert637 (
);

FILL FILL_5_BUFX2_insert638 (
);

FILL FILL_1__11927_ (
);

FILL FILL_5_BUFX2_insert639 (
);

FILL FILL_1__11507_ (
);

FILL FILL_5__16320_ (
);

FILL FILL_6__9901_ (
);

FILL FILL_0__8514_ (
);

FILL FILL_1__14399_ (
);

FILL FILL_5__6957_ (
);

FILL FILL_4__15733_ (
);

FILL FILL_4__15313_ (
);

OAI22X1 _13677_ (
    .A(_4183_),
    .B(_3931__bF$buf2),
    .C(_3977__bF$buf3),
    .D(_4184_),
    .Y(_4185_)
);

FILL FILL_3__9083_ (
);

NAND2X1 _13257_ (
    .A(_3770_),
    .B(_3772_),
    .Y(_3800_)
);

FILL FILL_3__14726_ (
);

FILL FILL_1__15760_ (
);

FILL FILL_3__14306_ (
);

FILL FILL_1__15340_ (
);

FILL FILL_1__6949_ (
);

FILL FILL_2__13719_ (
);

FILL FILL_0__14753_ (
);

FILL FILL_0__14333_ (
);

FILL SFILL14280x78050 (
);

FILL FILL_5__11299_ (
);

FILL FILL_2__7080_ (
);

FILL FILL_3__7816_ (
);

FILL FILL_0__9719_ (
);

FILL FILL_5__12660_ (
);

FILL FILL_5__12240_ (
);

NAND2X1 _6960_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_41_)
);

FILL FILL_2_BUFX2_insert760 (
);

FILL SFILL58360x61050 (
);

FILL FILL_2_BUFX2_insert761 (
);

FILL FILL_2_BUFX2_insert762 (
);

FILL FILL_2_BUFX2_insert763 (
);

FILL FILL_2_BUFX2_insert764 (
);

FILL FILL_4__11653_ (
);

FILL FILL_2_BUFX2_insert765 (
);

FILL FILL_4__11233_ (
);

FILL FILL_2_BUFX2_insert766 (
);

FILL FILL_2_BUFX2_insert767 (
);

FILL FILL_2_BUFX2_insert768 (
);

FILL FILL_2_BUFX2_insert769 (
);

FILL FILL_1__16125_ (
);

FILL FILL_3__10646_ (
);

FILL FILL_1__11680_ (
);

FILL FILL_1__11260_ (
);

FILL FILL_0__15958_ (
);

FILL FILL_0__15538_ (
);

AOI22X1 _15823_ (
    .A(_5649_),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .C(\datapath_1.regfile_1.regOut[21] [19]),
    .D(_5685_),
    .Y(_6284_)
);

INVX1 _15403_ (
    .A(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_5875_)
);

FILL FILL_0__15118_ (
);

FILL SFILL94520x18050 (
);

FILL FILL_0__10673_ (
);

FILL FILL_0__10253_ (
);

FILL FILL_6__14452_ (
);

FILL FILL_6__14032_ (
);

FILL FILL_5__13865_ (
);

FILL FILL_5__13445_ (
);

FILL FILL_5__13025_ (
);

INVX1 _7745_ (
    .A(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_442_)
);

INVX1 _7325_ (
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_223_)
);

FILL FILL_4__9992_ (
);

FILL FILL_4__9152_ (
);

FILL FILL_4__12858_ (
);

FILL FILL_4__12438_ (
);

FILL FILL_2__13892_ (
);

FILL FILL_4__12018_ (
);

FILL FILL_2__13472_ (
);

FILL FILL_6__9498_ (
);

FILL FILL_1__12885_ (
);

FILL FILL_1__12465_ (
);

FILL FILL_1__12045_ (
);

FILL FILL_0__9892_ (
);

FILL FILL_6_CLKBUF1_insert214 (
);

FILL FILL_0__9472_ (
);

FILL FILL_0__11878_ (
);

FILL FILL_0__11458_ (
);

NAND2X1 _11743_ (
    .A(_2462__bF$buf3),
    .B(_2833_),
    .Y(_2839_)
);

FILL FILL_0__11038_ (
);

NOR2X1 _11323_ (
    .A(_2301_),
    .B(_2300_),
    .Y(_2442_)
);

FILL SFILL109400x83050 (
);

FILL FILL_6_CLKBUF1_insert219 (
);

FILL FILL_5__7495_ (
);

FILL FILL_5__7075_ (
);

FILL FILL_4__16271_ (
);

FILL SFILL44040x51050 (
);

FILL FILL_3__15684_ (
);

FILL FILL_3__15264_ (
);

FILL FILL_1__7487_ (
);

FILL FILL_1__7067_ (
);

FILL FILL_2__14677_ (
);

FILL FILL_2__14257_ (
);

FILL FILL_0__15291_ (
);

FILL SFILL104360x50 (
);

FILL FILL_1_BUFX2_insert780 (
);

FILL FILL_3__8774_ (
);

FILL FILL_1_BUFX2_insert781 (
);

FILL FILL_3__8354_ (
);

DFFSR _12948_ (
    .Q(\datapath_1.a [29]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3555_[29])
);

FILL FILL_1_BUFX2_insert782 (
);

OAI21X1 _12528_ (
    .A(_3417_),
    .B(vdd),
    .C(_3418_),
    .Y(_3360_[29])
);

FILL FILL_1_BUFX2_insert783 (
);

NAND3X1 _12108_ (
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump [30]),
    .C(_3034__bF$buf1),
    .Y(_3127_)
);

FILL FILL_1_BUFX2_insert784 (
);

FILL FILL_1_BUFX2_insert785 (
);

FILL FILL_1_BUFX2_insert786 (
);

FILL FILL_1__14611_ (
);

FILL FILL_1_BUFX2_insert787 (
);

FILL FILL_1_BUFX2_insert788 (
);

FILL FILL_1_BUFX2_insert789 (
);

FILL FILL_4__12191_ (
);

FILL FILL_0__13604_ (
);

FILL FILL_3__16049_ (
);

FILL FILL_5__9641_ (
);

FILL FILL_5__9221_ (
);

FILL FILL_3__11184_ (
);

NAND2X1 _16361_ (
    .A(gnd),
    .B(gnd),
    .Y(_6795_)
);

FILL FILL_0__16076_ (
);

FILL FILL_2__10177_ (
);

FILL SFILL8440x28050 (
);

FILL FILL_5__11931_ (
);

FILL FILL_1__9633_ (
);

FILL FILL_5__11511_ (
);

FILL FILL_1__9213_ (
);

FILL FILL_3__9979_ (
);

FILL FILL_2__16403_ (
);

FILL FILL_4__10924_ (
);

FILL FILL_3__9139_ (
);

FILL FILL_4__10504_ (
);

FILL FILL_1__15816_ (
);

DFFSR _8283_ (
    .Q(\datapath_1.regfile_1.regOut[11] [5]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_653_[5])
);

FILL FILL_1__10951_ (
);

FILL FILL_1__10531_ (
);

FILL FILL_4__13396_ (
);

FILL FILL_1__10111_ (
);

FILL SFILL69160x62050 (
);

FILL FILL_0__14809_ (
);

FILL FILL_2__7976_ (
);

FILL FILL_2__7556_ (
);

BUFX2 BUFX2_insert450 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf4 )
);

BUFX2 BUFX2_insert451 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf3 )
);

FILL FILL_3__12389_ (
);

BUFX2 BUFX2_insert452 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf2 )
);

BUFX2 BUFX2_insert453 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf1 )
);

BUFX2 BUFX2_insert454 (
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf0 )
);

BUFX2 BUFX2_insert455 (
    .A(_3954_),
    .Y(_3954__bF$buf4)
);

FILL SFILL74120x45050 (
);

BUFX2 BUFX2_insert456 (
    .A(_3954_),
    .Y(_3954__bF$buf3)
);

BUFX2 BUFX2_insert457 (
    .A(_3954_),
    .Y(_3954__bF$buf2)
);

BUFX2 BUFX2_insert458 (
    .A(_3954_),
    .Y(_3954__bF$buf1)
);

BUFX2 BUFX2_insert459 (
    .A(_3954_),
    .Y(_3954__bF$buf0)
);

AOI22X1 _12281_ (
    .A(_2_[16]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump [16]),
    .Y(_3250_)
);

FILL FILL_5__12716_ (
);

FILL FILL_3__13750_ (
);

FILL FILL_3__13330_ (
);

FILL FILL_4__8843_ (
);

FILL FILL_4__11709_ (
);

FILL FILL_4__8003_ (
);

FILL FILL_2__12743_ (
);

FILL FILL_5__15188_ (
);

FILL FILL_2__12323_ (
);

FILL FILL_6__8769_ (
);

OAI21X1 _9488_ (
    .A(_1318_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .C(_1319_),
    .Y(_1303_[8])
);

DFFSR _9068_ (
    .Q(\datapath_1.regfile_1.regOut[17] [22]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_1043_[22])
);

FILL FILL_1__11736_ (
);

FILL FILL_1__11316_ (
);

FILL FILL_0__8743_ (
);

FILL FILL_3__6840_ (
);

FILL FILL_0__8323_ (
);

FILL FILL_0__10309_ (
);

FILL FILL_6__14508_ (
);

FILL FILL_4__15962_ (
);

FILL FILL_4__15542_ (
);

FILL FILL_4__15122_ (
);

INVX8 _13486_ (
    .A(_3959_),
    .Y(_3997_)
);

DFFSR _13066_ (
    .Q(_2_[19]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_3620_[19])
);

FILL FILL_3__14955_ (
);

FILL FILL_3__14535_ (
);

FILL FILL_3__14115_ (
);

FILL FILL_4_BUFX2_insert290 (
);

FILL FILL_4__9628_ (
);

FILL FILL_4_BUFX2_insert291 (
);

FILL FILL_4_BUFX2_insert292 (
);

FILL FILL_4__9208_ (
);

FILL FILL_4_BUFX2_insert293 (
);

FILL FILL_2__13948_ (
);

FILL FILL_0__14982_ (
);

FILL FILL_4_BUFX2_insert294 (
);

FILL FILL_2__13528_ (
);

FILL FILL_4_BUFX2_insert295 (
);

FILL FILL_0__14562_ (
);

FILL FILL_2__13108_ (
);

FILL FILL_4_BUFX2_insert296 (
);

FILL FILL_0__14142_ (
);

FILL FILL_4_BUFX2_insert297 (
);

FILL FILL_4_BUFX2_insert298 (
);

FILL FILL_4_BUFX2_insert299 (
);

FILL FILL_0__9528_ (
);

FILL FILL_3__7625_ (
);

FILL FILL_3__7205_ (
);

FILL FILL_0__9108_ (
);

FILL SFILL59160x60050 (
);

FILL FILL_4__16327_ (
);

FILL FILL_4__11882_ (
);

FILL FILL_4__11462_ (
);

FILL FILL_4__11042_ (
);

FILL SFILL64120x43050 (
);

FILL FILL_1__16354_ (
);

FILL FILL_3__10875_ (
);

FILL FILL_5__8912_ (
);

FILL FILL_3__10035_ (
);

FILL FILL_0__15767_ (
);

FILL FILL_0__15347_ (
);

OAI21X1 _15632_ (
    .A(_5524__bF$buf1),
    .B(_4661_),
    .C(_6097_),
    .Y(_6098_)
);

NAND2X1 _15212_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5513_),
    .Y(_5688_)
);

FILL FILL_2__8094_ (
);

FILL FILL_0__10062_ (
);

FILL FILL_1__8904_ (
);

FILL SFILL99640x25050 (
);

FILL FILL_5__13674_ (
);

FILL FILL_5__13254_ (
);

INVX1 _7974_ (
    .A(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_554_)
);

INVX1 _7554_ (
    .A(\datapath_1.regfile_1.regOut[6] [4]),
    .Y(_335_)
);

DFFSR _7134_ (
    .Q(\datapath_1.regfile_1.regOut[2] [8]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_68_[8])
);

FILL FILL_4__9381_ (
);

FILL FILL_4__12247_ (
);

FILL FILL_2__13281_ (
);

FILL FILL_1__12274_ (
);

DFFSR _16417_ (
    .Q(\datapath_1.regfile_1.regOut[0] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_6769_[0])
);

NAND2X1 _11972_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[28]),
    .Y(_3023_)
);

FILL FILL_2__9299_ (
);

FILL FILL_0__11687_ (
);

FILL FILL_0__9281_ (
);

AND2X2 _11552_ (
    .A(_2660_),
    .B(_2231_),
    .Y(_2661_)
);

FILL FILL_0__11267_ (
);

FILL FILL_5_CLKBUF1_insert200 (
);

INVX1 _11132_ (
    .A(_2250_),
    .Y(_2251_)
);

FILL FILL_5_CLKBUF1_insert201 (
);

FILL FILL_3__12601_ (
);

FILL FILL_5_CLKBUF1_insert202 (
);

FILL FILL_5_CLKBUF1_insert203 (
);

FILL FILL_4__16080_ (
);

FILL FILL_5_CLKBUF1_insert204 (
);

FILL FILL_5_CLKBUF1_insert205 (
);

FILL FILL_5_CLKBUF1_insert206 (
);

FILL FILL_5_CLKBUF1_insert207 (
);

FILL FILL_6__10181_ (
);

FILL FILL_5_CLKBUF1_insert208 (
);

FILL FILL_5__14879_ (
);

FILL FILL_5__14459_ (
);

FILL FILL_5_CLKBUF1_insert209 (
);

FILL FILL_5__14039_ (
);

FILL FILL_3__15493_ (
);

OAI21X1 _8759_ (
    .A(_954_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_955_),
    .Y(_913_[21])
);

FILL FILL_3__15073_ (
);

OAI21X1 _8339_ (
    .A(_735_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_736_),
    .Y(_718_[9])
);

FILL FILL_1__7296_ (
);

FILL FILL_2__14486_ (
);

FILL FILL_2__14066_ (
);

FILL FILL_5__15820_ (
);

FILL FILL_5__15400_ (
);

FILL SFILL89240x54050 (
);

DFFSR _9700_ (
    .Q(\datapath_1.regfile_1.regOut[22] [14]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_1368_[14])
);

FILL FILL_1__13899_ (
);

FILL SFILL54120x41050 (
);

FILL FILL_1__13479_ (
);

FILL FILL_4__14813_ (
);

FILL FILL_3__8583_ (
);

OAI21X1 _12757_ (
    .A(_3529_),
    .B(IRWrite_bF$buf3),
    .C(_3530_),
    .Y(_3490_[20])
);

AOI22X1 _12337_ (
    .A(_2_[30]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3292_)
);

FILL FILL_3__13806_ (
);

FILL SFILL18680x74050 (
);

FILL FILL_1__14840_ (
);

FILL FILL_5__8089_ (
);

FILL FILL_1__14420_ (
);

FILL FILL_1__14000_ (
);

FILL FILL_0__13833_ (
);

FILL FILL_0__13413_ (
);

FILL FILL_3__16278_ (
);

FILL FILL_5__10799_ (
);

FILL FILL_5__10379_ (
);

FILL FILL_5__9870_ (
);

FILL FILL_5__9030_ (
);

OAI22X1 _16170_ (
    .A(_5530__bF$buf3),
    .B(_6621_),
    .C(_5472__bF$buf3),
    .D(_5297_),
    .Y(_6622_)
);

FILL FILL_5__11740_ (
);

FILL FILL_1__9862_ (
);

FILL FILL_5__11320_ (
);

FILL FILL_1__9022_ (
);

FILL FILL_3__9788_ (
);

FILL FILL_2__16212_ (
);

FILL FILL_3__9368_ (
);

FILL FILL_4__10313_ (
);

FILL FILL_6__7373_ (
);

FILL FILL_1__15625_ (
);

OAI21X1 _8092_ (
    .A(_611_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .C(_612_),
    .Y(_588_[12])
);

FILL FILL_1__15205_ (
);

FILL FILL_1__10760_ (
);

FILL FILL_0__14618_ (
);

INVX1 _14903_ (
    .A(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_5385_)
);

FILL FILL_2__7365_ (
);

FILL FILL_3__12198_ (
);

NAND3X1 _12090_ (
    .A(_3111_),
    .B(_3112_),
    .C(_3113_),
    .Y(\datapath_1.mux_pcsrc.dout [25])
);

FILL FILL_5__12525_ (
);

FILL FILL_5__12105_ (
);

FILL SFILL79240x52050 (
);

FILL FILL_4__8652_ (
);

FILL FILL_4__8232_ (
);

FILL FILL_4__11938_ (
);

FILL FILL_2__12972_ (
);

FILL FILL_4__11518_ (
);

FILL FILL_2__12132_ (
);

FILL FILL_6__8578_ (
);

NAND2X1 _9297_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1233_)
);

FILL FILL111880x65050 (
);

FILL FILL_1__11965_ (
);

FILL FILL_1__11545_ (
);

FILL FILL_1__11125_ (
);

FILL FILL_0__8972_ (
);

FILL FILL_0__10958_ (
);

FILL FILL_0__8132_ (
);

INVX1 _10823_ (
    .A(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_2006_)
);

FILL FILL_0__10538_ (
);

INVX1 _10403_ (
    .A(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_1787_)
);

FILL FILL_0__10118_ (
);

FILL SFILL109400x78050 (
);

FILL FILL_5__6995_ (
);

FILL FILL_4__15771_ (
);

FILL FILL_4__15351_ (
);

OAI21X1 _13295_ (
    .A(_3822_),
    .B(_3831_),
    .C(_3750_),
    .Y(_3832_)
);

FILL FILL_2__9931_ (
);

FILL FILL_2__9511_ (
);

FILL FILL_3__14764_ (
);

FILL FILL_3__14344_ (
);

FILL FILL_1__6987_ (
);

FILL FILL112200x6050 (
);

FILL FILL_4__9857_ (
);

FILL FILL_4__9017_ (
);

FILL FILL_2__13757_ (
);

FILL FILL_2__13337_ (
);

FILL FILL_0__14791_ (
);

FILL FILL_0__14371_ (
);

FILL FILL_3__7854_ (
);

FILL FILL_0__9757_ (
);

FILL FILL_3__7434_ (
);

FILL FILL_0__9337_ (
);

NOR2X1 _11608_ (
    .A(_2713_),
    .B(_2712_),
    .Y(_2714_)
);

FILL FILL_4__16136_ (
);

FILL FILL_6__10657_ (
);

FILL FILL_4__11691_ (
);

FILL FILL_4__11271_ (
);

FILL FILL_3__15969_ (
);

FILL FILL_3__15549_ (
);

FILL FILL_3__15129_ (
);

FILL FILL_1__16163_ (
);

FILL FILL_3__10684_ (
);

FILL FILL_5__8721_ (
);

FILL FILL_3__10264_ (
);

FILL FILL_0__15996_ (
);

OAI22X1 _15861_ (
    .A(_4898_),
    .B(_5539__bF$buf0),
    .C(_5469__bF$buf3),
    .D(_4924_),
    .Y(_6321_)
);

FILL FILL_0__15576_ (
);

FILL SFILL69240x50050 (
);

FILL FILL_0__15156_ (
);

NAND3X1 _15441_ (
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5912_)
);

NAND2X1 _15021_ (
    .A(_5500__bF$buf2),
    .B(_5471__bF$buf3),
    .Y(_5501_)
);

FILL FILL_0__10291_ (
);

FILL FILL_1__8713_ (
);

FILL FILL_2__15903_ (
);

FILL FILL_3__8639_ (
);

FILL FILL_3__8219_ (
);

FILL FILL_5__13483_ (
);

DFFSR _7783_ (
    .Q(\datapath_1.regfile_1.regOut[7] [17]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_393_[17])
);

OAI21X1 _7363_ (
    .A(_247_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .C(_248_),
    .Y(_198_[25])
);

FILL SFILL100040x5050 (
);

FILL SFILL99400x82050 (
);

FILL FILL_4__12896_ (
);

FILL FILL_4__12476_ (
);

FILL SFILL69160x57050 (
);

FILL FILL_4__12056_ (
);

FILL FILL_2__13090_ (
);

FILL FILL_5_BUFX2_insert20 (
);

FILL FILL_3__11889_ (
);

FILL FILL_5_BUFX2_insert21 (
);

FILL FILL_5__9926_ (
);

FILL FILL_5__9506_ (
);

FILL FILL_3__11469_ (
);

FILL FILL_5_BUFX2_insert22 (
);

FILL FILL_5_BUFX2_insert23 (
);

FILL FILL_3__11049_ (
);

FILL FILL_1__12083_ (
);

FILL FILL_5_BUFX2_insert24 (
);

FILL FILL_5_BUFX2_insert25 (
);

FILL FILL_5_BUFX2_insert26 (
);

NOR2X1 _16226_ (
    .A(_6676_),
    .B(_6674_),
    .Y(_6677_)
);

FILL FILL_5_BUFX2_insert27 (
);

FILL FILL_5_BUFX2_insert28 (
);

FILL FILL_5_BUFX2_insert29 (
);

FILL FILL_0__9090_ (
);

AND2X2 _11781_ (
    .A(_2863_),
    .B(_2558_),
    .Y(_2875_)
);

FILL FILL_0__11496_ (
);

INVX4 _11361_ (
    .A(_2344__bF$buf3),
    .Y(_2478_)
);

FILL FILL_0__11076_ (
);

FILL FILL_1__9918_ (
);

FILL FILL_6__15695_ (
);

FILL FILL_3__12830_ (
);

FILL FILL_3__12410_ (
);

FILL FILL_6__15275_ (
);

FILL FILL_4__7503_ (
);

FILL FILL_2__11823_ (
);

FILL FILL_5__14688_ (
);

FILL FILL_5__14268_ (
);

FILL FILL_2__11403_ (
);

OAI21X1 _8988_ (
    .A(_1066_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .C(_1067_),
    .Y(_1043_[12])
);

FILL FILL_6__7849_ (
);

OAI21X1 _8568_ (
    .A(_911_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_912_),
    .Y(_848_[0])
);

NAND2X1 _8148_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_650_)
);

FILL FILL_1__10816_ (
);

FILL FILL_2__14295_ (
);

FILL FILL_0__7823_ (
);

FILL SFILL69160x12050 (
);

FILL FILL_1__13288_ (
);

FILL FILL_4__14622_ (
);

FILL FILL_4__14202_ (
);

FILL SFILL78840x17050 (
);

OAI21X1 _12986_ (
    .A(_3641_),
    .B(vdd),
    .C(_3642_),
    .Y(_3620_[11])
);

FILL FILL_3__8392_ (
);

DFFSR _12566_ (
    .Q(ALUOut[31]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3360_[31])
);

NAND2X1 _12146_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.a [10]),
    .Y(_3151_)
);

FILL FILL_3__13615_ (
);

FILL FILL_4__8708_ (
);

FILL FILL_6__11195_ (
);

FILL FILL_2__12608_ (
);

FILL FILL_0__13642_ (
);

FILL FILL_0__13222_ (
);

FILL FILL_3__16087_ (
);

FILL FILL_5__10188_ (
);

FILL SFILL89400x80050 (
);

FILL FILL_5__16414_ (
);

FILL FILL_0__8608_ (
);

FILL SFILL59160x55050 (
);

FILL FILL_1__9671_ (
);

FILL FILL_1__9251_ (
);

FILL FILL_4__15827_ (
);

FILL FILL_4__15407_ (
);

BUFX2 BUFX2_insert1010 (
    .A(_4079_),
    .Y(_4079__bF$buf3)
);

BUFX2 BUFX2_insert1011 (
    .A(_4079_),
    .Y(_4079__bF$buf2)
);

FILL FILL_2__16021_ (
);

BUFX2 BUFX2_insert1012 (
    .A(_4079_),
    .Y(_4079__bF$buf1)
);

FILL FILL_3__9597_ (
);

FILL FILL_4__10962_ (
);

BUFX2 BUFX2_insert1013 (
    .A(_4079_),
    .Y(_4079__bF$buf0)
);

BUFX2 BUFX2_insert1014 (
    .A(_5534_),
    .Y(_5534__bF$buf4)
);

FILL FILL_4__10542_ (
);

FILL SFILL64120x38050 (
);

FILL FILL_4__10122_ (
);

BUFX2 BUFX2_insert1015 (
    .A(_5534_),
    .Y(_5534__bF$buf3)
);

BUFX2 BUFX2_insert1016 (
    .A(_5534_),
    .Y(_5534__bF$buf2)
);

FILL FILL_1__15854_ (
);

BUFX2 BUFX2_insert1017 (
    .A(_5534_),
    .Y(_5534__bF$buf1)
);

BUFX2 BUFX2_insert1018 (
    .A(_5534_),
    .Y(_5534__bF$buf0)
);

FILL FILL_1__15434_ (
);

FILL FILL_1__15014_ (
);

BUFX2 BUFX2_insert1019 (
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf7 )
);

FILL FILL_0__14847_ (
);

AOI21X1 _14712_ (
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .B(_4038__bF$buf0),
    .C(_5197_),
    .Y(_5198_)
);

FILL FILL_0__14427_ (
);

FILL FILL_0__14007_ (
);

BUFX2 BUFX2_insert830 (
    .A(_5526_),
    .Y(_5526__bF$buf4)
);

FILL FILL_2__7594_ (
);

BUFX2 BUFX2_insert831 (
    .A(_5526_),
    .Y(_5526__bF$buf3)
);

FILL FILL_2__7174_ (
);

BUFX2 BUFX2_insert832 (
    .A(_5526_),
    .Y(_5526__bF$buf2)
);

BUFX2 BUFX2_insert833 (
    .A(_5526_),
    .Y(_5526__bF$buf1)
);

FILL FILL_6__13761_ (
);

BUFX2 BUFX2_insert834 (
    .A(_5526_),
    .Y(_5526__bF$buf0)
);

FILL FILL_6__13341_ (
);

BUFX2 BUFX2_insert835 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf7 )
);

BUFX2 BUFX2_insert836 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf6 )
);

BUFX2 BUFX2_insert837 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf5 )
);

BUFX2 BUFX2_insert838 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf4 )
);

BUFX2 BUFX2_insert839 (
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf3 )
);

FILL FILL_5__12754_ (
);

FILL FILL_5__12334_ (
);

FILL SFILL59160x10050 (
);

FILL FILL_4__8881_ (
);

FILL FILL_4__8461_ (
);

FILL FILL_4__11747_ (
);

FILL FILL_2__12781_ (
);

FILL FILL_4__11327_ (
);

FILL FILL_2__12361_ (
);

FILL FILL_1__16219_ (
);

FILL FILL_1__11774_ (
);

FILL FILL_1__11354_ (
);

NAND3X1 _15917_ (
    .A(_6370_),
    .B(_6375_),
    .C(_6372_),
    .Y(_6376_)
);

FILL SFILL33960x82050 (
);

FILL FILL_0__8781_ (
);

FILL FILL_0__10767_ (
);

FILL FILL_2__8379_ (
);

FILL FILL_0__8361_ (
);

INVX1 _10632_ (
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_1899_)
);

FILL SFILL89320x42050 (
);

DFFSR _10212_ (
    .Q(\datapath_1.regfile_1.regOut[26] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_1628_[14])
);

FILL FILL_4__15580_ (
);

FILL FILL_4__15160_ (
);

FILL FILL_5__13959_ (
);

FILL SFILL113800x47050 (
);

FILL FILL_2__9740_ (
);

FILL FILL_3__14993_ (
);

FILL FILL_5__13539_ (
);

FILL FILL_3__14573_ (
);

FILL FILL_5__13119_ (
);

FILL FILL_3__14153_ (
);

OAI21X1 _7839_ (
    .A(_483_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_484_),
    .Y(_458_[13])
);

OAI21X1 _7419_ (
    .A(_264_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .C(_265_),
    .Y(_263_[1])
);

FILL SFILL49160x53050 (
);

FILL FILL_4_BUFX2_insert670 (
);

FILL FILL_4_BUFX2_insert671 (
);

FILL FILL_4__9666_ (
);

FILL FILL_4_BUFX2_insert672 (
);

FILL FILL_4__9246_ (
);

FILL FILL_2__13986_ (
);

FILL FILL_4_BUFX2_insert673 (
);

FILL FILL_4_BUFX2_insert674 (
);

FILL FILL_2__13566_ (
);

FILL FILL_2__13146_ (
);

FILL FILL_4_BUFX2_insert675 (
);

FILL FILL_0__14180_ (
);

FILL FILL_4_BUFX2_insert676 (
);

FILL FILL_4_BUFX2_insert677 (
);

FILL FILL_5__14900_ (
);

FILL FILL_4_BUFX2_insert678 (
);

FILL SFILL89240x49050 (
);

FILL FILL_4_BUFX2_insert679 (
);

FILL SFILL54120x36050 (
);

FILL FILL_1__12979_ (
);

FILL FILL_1__12139_ (
);

FILL FILL_0__9986_ (
);

FILL FILL_3__7243_ (
);

FILL FILL_0__9146_ (
);

NOR2X1 _11837_ (
    .A(\datapath_1.alu_1.ALUInA [0]),
    .B(_2490_),
    .Y(_2926_)
);

AOI21X1 _11417_ (
    .A(_2531_),
    .B(_2533_),
    .C(_2485_),
    .Y(_2534_)
);

FILL FILL_5__7589_ (
);

FILL FILL_1__13920_ (
);

FILL FILL_5__7169_ (
);

FILL FILL_4__16365_ (
);

FILL FILL_1__13500_ (
);

FILL FILL_6__10046_ (
);

FILL FILL_4__11080_ (
);

FILL FILL_3__15778_ (
);

FILL FILL_0__12913_ (
);

FILL FILL_3__15358_ (
);

FILL FILL_1__16392_ (
);

FILL FILL_5__8950_ (
);

FILL FILL_5__8530_ (
);

FILL FILL_3__10493_ (
);

FILL FILL_5__8110_ (
);

FILL FILL_0__15385_ (
);

INVX1 _15670_ (
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_6135_)
);

NOR2X1 _15250_ (
    .A(_5725_),
    .B(_5723_),
    .Y(_5726_)
);

FILL FILL_5__10820_ (
);

FILL FILL_5__10400_ (
);

FILL FILL_1__8522_ (
);

FILL FILL_1__8102_ (
);

FILL FILL_2__15712_ (
);

FILL FILL_3__8868_ (
);

FILL FILL_3__8448_ (
);

FILL FILL_5__13292_ (
);

FILL FILL_6__6873_ (
);

OAI21X1 _7592_ (
    .A(_359_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_360_),
    .Y(_328_[16])
);

FILL FILL_1__14705_ (
);

FILL FILL_4_BUFX2_insert1050 (
);

OAI21X1 _7172_ (
    .A(_140_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_141_),
    .Y(_133_[4])
);

FILL FILL_4_BUFX2_insert1051 (
);

FILL FILL_4_BUFX2_insert1052 (
);

FILL SFILL79320x40050 (
);

FILL FILL_4_BUFX2_insert1053 (
);

FILL SFILL18680x24050 (
);

FILL FILL_4_BUFX2_insert1054 (
);

FILL FILL_4_BUFX2_insert1055 (
);

FILL FILL_4__12285_ (
);

FILL FILL_4_BUFX2_insert1056 (
);

FILL FILL_4_BUFX2_insert1057 (
);

FILL FILL_4_BUFX2_insert1058 (
);

FILL FILL_4_BUFX2_insert1059 (
);

FILL FILL_2__6865_ (
);

FILL FILL_5__9735_ (
);

FILL FILL_3__11698_ (
);

FILL FILL_3__11278_ (
);

FILL FILL111960x53050 (
);

NAND3X1 _16035_ (
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .B(_5465_),
    .C(_5531__bF$buf4),
    .Y(_6491_)
);

OAI22X1 _11590_ (
    .A(_2247_),
    .B(_2480_),
    .C(_2248_),
    .D(_2344__bF$buf2),
    .Y(_2697_)
);

INVX4 _11170_ (
    .A(_2288_),
    .Y(_2289_)
);

FILL SFILL65000x75050 (
);

FILL FILL_1__9727_ (
);

FILL FILL_5__11605_ (
);

FILL SFILL79240x47050 (
);

FILL FILL_4__7732_ (
);

FILL FILL_3_BUFX2_insert690 (
);

FILL FILL_4__7312_ (
);

FILL FILL_3_BUFX2_insert691 (
);

FILL FILL_3_BUFX2_insert692 (
);

FILL FILL_5__14497_ (
);

FILL FILL_3_BUFX2_insert693 (
);

FILL FILL_2__11632_ (
);

FILL FILL_3_BUFX2_insert694 (
);

FILL FILL_2__11212_ (
);

FILL FILL_5__14077_ (
);

FILL FILL_3_BUFX2_insert695 (
);

DFFSR _8797_ (
    .Q(\datapath_1.regfile_1.regOut[15] [7]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_913_[7])
);

NAND2X1 _8377_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_762_)
);

FILL FILL_3_BUFX2_insert696 (
);

FILL FILL_3_BUFX2_insert697 (
);

FILL FILL_3_BUFX2_insert698 (
);

FILL FILL_3_BUFX2_insert699 (
);

FILL FILL_1__10625_ (
);

FILL FILL_0__7632_ (
);

FILL FILL_0__7212_ (
);

FILL FILL_1__13097_ (
);

FILL FILL_6__13817_ (
);

FILL SFILL54120x9050 (
);

FILL FILL_4__14851_ (
);

FILL FILL_4__14431_ (
);

FILL FILL_4__14011_ (
);

DFFSR _12795_ (
    .Q(\aluControl_1.inst [4]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3490_[4])
);

OAI21X1 _12375_ (
    .A(_3314_),
    .B(MemToReg_bF$buf4),
    .C(_3315_),
    .Y(\datapath_1.mux_wd3.dout [10])
);

FILL FILL_3__13844_ (
);

FILL FILL_3__13424_ (
);

FILL FILL_3__13004_ (
);

FILL FILL_4__8517_ (
);

FILL FILL_2__12837_ (
);

FILL FILL_0__13871_ (
);

FILL FILL_2__12417_ (
);

FILL FILL_0__13451_ (
);

FILL FILL_0__13031_ (
);

FILL FILL_5__16223_ (
);

FILL FILL_0__8837_ (
);

FILL FILL_3__6934_ (
);

FILL FILL_1__9480_ (
);

FILL FILL_4__15636_ (
);

FILL FILL_4__15216_ (
);

FILL FILL_2__16250_ (
);

FILL FILL_4__10771_ (
);

FILL FILL_3__14629_ (
);

FILL FILL_1__15663_ (
);

FILL FILL_3__14209_ (
);

FILL FILL_1__15243_ (
);

FILL FILL_5__7801_ (
);

FILL SFILL69240x45050 (
);

NOR2X1 _14941_ (
    .A(_5421_),
    .B(_3955__bF$buf1),
    .Y(_5422_)
);

FILL FILL_0__14656_ (
);

FILL FILL_0__14236_ (
);

NOR2X1 _14521_ (
    .A(_5010_),
    .B(_3935__bF$buf1),
    .Y(_5011_)
);

OAI22X1 _14101_ (
    .A(_4598_),
    .B(_3930__bF$buf2),
    .C(_3931__bF$buf3),
    .D(_4599_),
    .Y(_4600_)
);

FILL FILL_3__7719_ (
);

FILL FILL_5__12983_ (
);

FILL FILL_5__12143_ (
);

BUFX2 _6863_ (
    .A(_1_[25]),
    .Y(memoryAddress[25])
);

FILL FILL_4__8270_ (
);

FILL FILL_4__11976_ (
);

FILL FILL_4__11556_ (
);

FILL SFILL34040x39050 (
);

FILL FILL_2__12590_ (
);

FILL FILL_4__11136_ (
);

FILL FILL_2__12170_ (
);

FILL FILL_6__8196_ (
);

FILL FILL_1__16028_ (
);

FILL FILL_3__10969_ (
);

FILL FILL_3__10549_ (
);

FILL FILL_3__10129_ (
);

FILL FILL_1__11583_ (
);

FILL FILL_1__11163_ (
);

OAI22X1 _15726_ (
    .A(_5523_),
    .B(_4744_),
    .C(_4754_),
    .D(_5524__bF$buf3),
    .Y(_6190_)
);

OAI22X1 _15306_ (
    .A(_5526__bF$buf3),
    .B(_4280_),
    .C(_4283_),
    .D(_5527__bF$buf4),
    .Y(_5780_)
);

FILL FILL_0__8590_ (
);

FILL FILL_0__10996_ (
);

DFFSR _10861_ (
    .Q(\datapath_1.regfile_1.regOut[31] [23]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_1953_[23])
);

FILL FILL_0__10576_ (
);

FILL FILL_2__8188_ (
);

FILL SFILL104360x70050 (
);

FILL FILL_0__10156_ (
);

OAI21X1 _10441_ (
    .A(_1811_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .C(_1812_),
    .Y(_1758_[27])
);

OAI21X1 _10021_ (
    .A(_1592_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .C(_1593_),
    .Y(_1563_[15])
);

FILL FILL_3__11910_ (
);

FILL FILL_2__10903_ (
);

FILL FILL_5__13768_ (
);

FILL FILL_5__13348_ (
);

FILL FILL_3__14382_ (
);

FILL FILL_6__6929_ (
);

DFFSR _7648_ (
    .Q(\datapath_1.regfile_1.regOut[6] [10]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_328_[10])
);

NAND2X1 _7228_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_179_)
);

FILL FILL_4__9895_ (
);

FILL FILL_4__9475_ (
);

FILL FILL_2__13795_ (
);

FILL FILL_2__13375_ (
);

FILL SFILL99400x32050 (
);

FILL FILL_0__6903_ (
);

FILL FILL_1__12788_ (
);

FILL FILL_1__12368_ (
);

FILL FILL_4__13702_ (
);

FILL FILL_3__7892_ (
);

FILL FILL_0__9795_ (
);

FILL FILL_3__7472_ (
);

FILL FILL_0__9375_ (
);

FILL FILL_3__7052_ (
);

OAI21X1 _11646_ (
    .A(_2404_),
    .B(_2480_),
    .C(_2748_),
    .Y(_2749_)
);

OAI21X1 _11226_ (
    .A(_2111_),
    .B(_2344__bF$buf0),
    .C(_2342_),
    .Y(_2345_)
);

FILL FILL_4__16174_ (
);

FILL SFILL99320x39050 (
);

FILL FILL_0__12722_ (
);

FILL FILL_3__15587_ (
);

FILL FILL_0__12302_ (
);

FILL FILL_3__15167_ (
);

FILL FILL_0__15194_ (
);

FILL FILL_5__15914_ (
);

FILL SFILL28760x59050 (
);

FILL FILL_1__8751_ (
);

FILL FILL_1__8331_ (
);

FILL SFILL3720x7050 (
);

FILL FILL_4__14907_ (
);

FILL FILL_2__15941_ (
);

FILL FILL_2__15521_ (
);

FILL FILL_2__15101_ (
);

FILL FILL_3__8257_ (
);

FILL FILL_1__14934_ (
);

FILL FILL_1__14514_ (
);

FILL FILL_4__12094_ (
);

FILL FILL_0__13927_ (
);

FILL FILL_0__13507_ (
);

FILL FILL_5__9544_ (
);

FILL FILL_5__9124_ (
);

FILL FILL_3__11087_ (
);

FILL FILL_6__12841_ (
);

FILL FILL_0__16399_ (
);

NOR2X1 _16264_ (
    .A(_5378_),
    .B(_5549__bF$buf0),
    .Y(_6714_)
);

FILL SFILL114440x1050 (
);

FILL FILL_5__11834_ (
);

FILL FILL_1__9536_ (
);

FILL FILL_5__11414_ (
);

FILL SFILL28760x14050 (
);

FILL FILL_1__9116_ (
);

FILL SFILL94280x81050 (
);

FILL FILL_4__7961_ (
);

FILL FILL_2__16306_ (
);

FILL FILL_4__10827_ (
);

FILL FILL_4__7121_ (
);

FILL FILL_4__10407_ (
);

FILL FILL_2__11861_ (
);

FILL FILL_2__11441_ (
);

FILL FILL_2__11021_ (
);

FILL FILL_1__15719_ (
);

FILL FILL_6__7467_ (
);

NAND2X1 _8186_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_655_)
);

FILL FILL_4__13299_ (
);

FILL FILL_1__10434_ (
);

FILL FILL_1__10014_ (
);

FILL SFILL113640x8050 (
);

FILL SFILL33960x77050 (
);

FILL FILL_0__7861_ (
);

FILL FILL_2__7879_ (
);

FILL FILL_2__7459_ (
);

FILL FILL_0__7441_ (
);

FILL SFILL89320x37050 (
);

FILL FILL_2__7039_ (
);

FILL FILL_4__14660_ (
);

FILL FILL_4__14240_ (
);

INVX1 _12184_ (
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3176_)
);

FILL FILL_5__12619_ (
);

FILL FILL_3__13653_ (
);

FILL FILL_2__8400_ (
);

FILL SFILL18760x57050 (
);

FILL FILL_3__13233_ (
);

OAI21X1 _6919_ (
    .A(_12_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .C(_13_),
    .Y(_3_[5])
);

FILL SFILL33560x63050 (
);

FILL FILL_4__8746_ (
);

FILL FILL_4__8326_ (
);

FILL FILL_2__12646_ (
);

FILL FILL_0__13680_ (
);

FILL FILL_2__12226_ (
);

FILL FILL_0__13260_ (
);

FILL FILL_1__11639_ (
);

FILL FILL_1__11219_ (
);

FILL FILL_6_BUFX2_insert70 (
);

FILL FILL_5__16032_ (
);

FILL FILL_0__8646_ (
);

NOR2X1 _10917_ (
    .A(_2051_),
    .B(_2059_),
    .Y(PCWrite)
);

FILL FILL_0__8226_ (
);

FILL FILL_6_BUFX2_insert75 (
);

FILL SFILL33960x32050 (
);

FILL FILL_4__15865_ (
);

FILL FILL_4__15445_ (
);

FILL FILL_4__15025_ (
);

NOR2X1 _13389_ (
    .A(_3899_),
    .B(_3900_),
    .Y(_3901_)
);

FILL FILL_4__10580_ (
);

FILL FILL_4__10160_ (
);

FILL FILL_3__14858_ (
);

FILL FILL_2__9605_ (
);

FILL FILL_1__15892_ (
);

FILL FILL_3__14438_ (
);

FILL FILL_3__14018_ (
);

FILL FILL_1__15472_ (
);

FILL FILL_1__15052_ (
);

FILL FILL_5__7610_ (
);

FILL SFILL18760x12050 (
);

FILL FILL_0__14885_ (
);

FILL FILL_0__14465_ (
);

INVX1 _14750_ (
    .A(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_5235_)
);

FILL FILL_0__14045_ (
);

OAI22X1 _14330_ (
    .A(_4822_),
    .B(_3884__bF$buf3),
    .C(_3920_),
    .D(_4823_),
    .Y(_4824_)
);

FILL SFILL79720x49050 (
);

FILL FILL_1__7602_ (
);

FILL FILL_3__7948_ (
);

FILL FILL_3__7108_ (
);

FILL FILL_5__12372_ (
);

FILL SFILL18680x19050 (
);

FILL FILL_4__11785_ (
);

FILL FILL_4__11365_ (
);

FILL FILL_1__16257_ (
);

FILL FILL_3__10778_ (
);

FILL FILL111960x48050 (
);

FILL FILL_3__10358_ (
);

FILL FILL_1__11392_ (
);

NAND2X1 _15955_ (
    .A(_6407_),
    .B(_6412_),
    .Y(_6413_)
);

NOR3X1 _15535_ (
    .A(_5992_),
    .B(_5981_),
    .C(_6003_),
    .Y(_6004_)
);

OAI21X1 _15115_ (
    .A(_5524__bF$buf2),
    .B(_4002_),
    .C(_5593_),
    .Y(_5594_)
);

OAI21X1 _10670_ (
    .A(_1923_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .C(_1924_),
    .Y(_1888_[18])
);

FILL FILL_0__10385_ (
);

OAI21X1 _10250_ (
    .A(_1704_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1705_),
    .Y(_1693_[6])
);

FILL FILL_5__13997_ (
);

FILL FILL_5__13577_ (
);

FILL FILL_5__13157_ (
);

FILL FILL_3__14191_ (
);

NAND2X1 _7877_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_510_)
);

NAND2X1 _7457_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_291_)
);

NAND2X1 _7037_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_72_)
);

FILL FILL_4__9284_ (
);

FILL SFILL114440x60050 (
);

FILL FILL_1__12597_ (
);

FILL FILL_1__12177_ (
);

FILL FILL_4__13931_ (
);

FILL FILL_4__13511_ (
);

INVX1 _11875_ (
    .A(\datapath_1.PCJump [19]),
    .Y(_2960_)
);

NAND3X1 _11455_ (
    .A(_2324_),
    .B(_2449_),
    .C(_2570_),
    .Y(_2571_)
);

XNOR2X1 _11035_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2154_)
);

FILL FILL_3__12504_ (
);

FILL SFILL114360x67050 (
);

FILL FILL_2__11917_ (
);

FILL FILL_0__12951_ (
);

FILL FILL_3__15396_ (
);

FILL FILL_0__12531_ (
);

FILL FILL_0__12111_ (
);

FILL FILL_1__7199_ (
);

FILL FILL_2__14389_ (
);

FILL FILL_5__15723_ (
);

FILL FILL_5__15303_ (
);

NAND2X1 _9603_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1376_)
);

FILL FILL_1__8980_ (
);

FILL FILL_1__8140_ (
);

FILL FILL_4__14716_ (
);

FILL FILL_2__15750_ (
);

FILL FILL_2__15330_ (
);

FILL FILL_3__8486_ (
);

FILL FILL_3__8066_ (
);

FILL FILL_3__13709_ (
);

FILL FILL_1__14743_ (
);

FILL FILL_1__14323_ (
);

FILL FILL_0__13736_ (
);

FILL FILL_0__13316_ (
);

OAI22X1 _13601_ (
    .A(_4108_),
    .B(_3905__bF$buf1),
    .C(_3977__bF$buf1),
    .D(_4109_),
    .Y(_4110_)
);

FILL FILL_5__9773_ (
);

FILL FILL_5__9353_ (
);

OAI22X1 _16073_ (
    .A(_6526_),
    .B(_5545__bF$buf3),
    .C(_5485__bF$buf0),
    .D(_6527_),
    .Y(_6528_)
);

FILL FILL_1__9765_ (
);

FILL FILL_5__11643_ (
);

FILL FILL_1__9345_ (
);

FILL FILL_5__11223_ (
);

FILL FILL_2__16115_ (
);

FILL FILL_4__7350_ (
);

FILL FILL_4__10636_ (
);

FILL FILL_2__11670_ (
);

FILL FILL_2__11250_ (
);

FILL FILL_1__15948_ (
);

FILL SFILL114280x29050 (
);

FILL FILL_1__15528_ (
);

FILL FILL_1__15108_ (
);

FILL FILL_1__10663_ (
);

FILL FILL_1__10243_ (
);

OAI22X1 _14806_ (
    .A(_5289_),
    .B(_3949_),
    .C(_3983__bF$buf0),
    .D(_5288_),
    .Y(_5290_)
);

FILL FILL_2__7688_ (
);

FILL FILL_0__7670_ (
);

FILL SFILL104360x65050 (
);

FILL FILL_0__7250_ (
);

FILL SFILL69160x8050 (
);

FILL SFILL43880x4050 (
);

FILL FILL_5__12848_ (
);

FILL FILL_5__12428_ (
);

FILL FILL_3__13882_ (
);

FILL FILL_3__13462_ (
);

FILL FILL_5__12008_ (
);

FILL FILL_3__13042_ (
);

FILL FILL_4__8975_ (
);

FILL SFILL8600x4050 (
);

FILL FILL_4__8135_ (
);

FILL FILL_2__12875_ (
);

FILL FILL_2__12455_ (
);

FILL SFILL99400x27050 (
);

FILL FILL_2__12035_ (
);

FILL FILL_1__11868_ (
);

FILL FILL_1__11448_ (
);

FILL FILL_1__11028_ (
);

FILL FILL_3__6972_ (
);

FILL FILL_0__8875_ (
);

FILL FILL_5__16261_ (
);

FILL FILL_0__8455_ (
);

FILL FILL112440x71050 (
);

DFFSR _10726_ (
    .Q(\datapath_1.regfile_1.regOut[30] [16]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_1888_[16])
);

FILL FILL_6__9002_ (
);

NAND2X1 _10306_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1743_)
);

FILL FILL_5__6898_ (
);

FILL FILL_4__15674_ (
);

FILL SFILL104360x20050 (
);

FILL FILL_4__15254_ (
);

FILL SFILL83720x49050 (
);

DFFSR _13198_ (
    .Q(\datapath_1.mux_iord.din0 [23]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3685_[23])
);

FILL FILL_2__9414_ (
);

FILL FILL_0__11802_ (
);

FILL FILL_3__14667_ (
);

FILL FILL_3__14247_ (
);

FILL FILL_1__15281_ (
);

FILL FILL_0__14694_ (
);

FILL FILL_0__14274_ (
);

FILL FILL_1__7831_ (
);

FILL SFILL104280x27050 (
);

FILL FILL_2__14601_ (
);

FILL FILL_3__7757_ (
);

FILL FILL_3__7337_ (
);

FILL FILL_5__12181_ (
);

FILL FILL_4__16039_ (
);

FILL FILL_4__11594_ (
);

FILL FILL_4__11174_ (
);

FILL FILL_1__16066_ (
);

FILL FILL_5__8624_ (
);

FILL FILL_3__10167_ (
);

FILL FILL_5__8204_ (
);

FILL FILL_6_BUFX2_insert582 (
);

FILL FILL_0__15899_ (
);

NAND3X1 _15764_ (
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .B(_5471__bF$buf4),
    .C(_5531__bF$buf3),
    .Y(_6227_)
);

FILL FILL_0__15479_ (
);

INVX1 _15344_ (
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_5817_)
);

FILL FILL_0__15059_ (
);

FILL FILL_6_BUFX2_insert587 (
);

FILL FILL_0__10194_ (
);

FILL SFILL89400x25050 (
);

FILL FILL_5__10914_ (
);

FILL FILL_1__8616_ (
);

FILL SFILL94280x76050 (
);

FILL FILL_2__15806_ (
);

FILL FILL_0__16000_ (
);

FILL FILL_2__10941_ (
);

FILL FILL_5__13386_ (
);

FILL FILL_2__10521_ (
);

NAND2X1 _7686_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_403_)
);

DFFSR _7266_ (
    .Q(\datapath_1.regfile_1.regOut[3] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_133_[12])
);

FILL FILL_4__9093_ (
);

FILL FILL_4__12379_ (
);

FILL FILL_3__9903_ (
);

FILL FILL_2__6959_ (
);

FILL FILL_0__6941_ (
);

FILL FILL_5__9409_ (
);

FILL FILL_4__13740_ (
);

FILL FILL_4__13320_ (
);

AOI22X1 _16129_ (
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [27]),
    .C(\datapath_1.regfile_1.regOut[22] [27]),
    .D(_5650_),
    .Y(_6582_)
);

FILL FILL_3__7090_ (
);

NOR2X1 _11684_ (
    .A(_2165_),
    .B(_2764_),
    .Y(_2785_)
);

FILL FILL_0__11399_ (
);

NAND2X1 _11264_ (
    .A(_2379_),
    .B(_2382_),
    .Y(_2383_)
);

FILL SFILL63800x83050 (
);

FILL SFILL79400x68050 (
);

FILL SFILL94200x74050 (
);

FILL FILL_3__12733_ (
);

FILL FILL_6__15598_ (
);

FILL FILL_6__15178_ (
);

FILL FILL_3__12313_ (
);

FILL FILL_4__7826_ (
);

FILL FILL_2__11726_ (
);

FILL FILL_0__12760_ (
);

FILL FILL_2__11306_ (
);

FILL FILL_0__12340_ (
);

FILL FILL_2__14198_ (
);

FILL FILL_5__15952_ (
);

FILL FILL_5__15532_ (
);

FILL FILL_0__7726_ (
);

FILL FILL_5__15112_ (
);

FILL FILL_0__7306_ (
);

DFFSR _9832_ (
    .Q(\datapath_1.regfile_1.regOut[23] [18]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_1433_[18])
);

INVX1 _9412_ (
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_1289_)
);

FILL SFILL33960x27050 (
);

FILL FILL_4__14945_ (
);

FILL FILL_4__14525_ (
);

FILL FILL_4__14105_ (
);

INVX1 _12889_ (
    .A(\datapath_1.a [22]),
    .Y(_3598_)
);

INVX1 _12469_ (
    .A(ALUOut[10]),
    .Y(_3379_)
);

AOI22X1 _12049_ (
    .A(\datapath_1.ALUResult [15]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3083_)
);

FILL FILL_3__13938_ (
);

FILL FILL_1__14972_ (
);

FILL FILL_3__13518_ (
);

FILL FILL_1__14552_ (
);

FILL FILL_1__14132_ (
);

FILL SFILL79400x23050 (
);

FILL FILL_6__11098_ (
);

FILL SFILL115160x21050 (
);

FILL FILL_0__13965_ (
);

AOI21X1 _13830_ (
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .B(_4040_),
    .C(_4334_),
    .Y(_4335_)
);

FILL FILL_0__13545_ (
);

FILL FILL_0__13125_ (
);

INVX1 _13410_ (
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_3922_)
);

FILL FILL_5__9162_ (
);

FILL FILL_5__16317_ (
);

FILL FILL_5__11872_ (
);

FILL FILL_1__9994_ (
);

FILL FILL_5__11452_ (
);

FILL FILL_5__11032_ (
);

FILL FILL_1__9154_ (
);

FILL FILL_2__16344_ (
);

FILL FILL_4__10445_ (
);

FILL FILL_4__10025_ (
);

FILL FILL_1__15757_ (
);

FILL FILL_1__15337_ (
);

FILL FILL_1__10892_ (
);

FILL SFILL23560x56050 (
);

FILL FILL_1__10052_ (
);

OAI22X1 _14615_ (
    .A(_5102_),
    .B(_3902__bF$buf1),
    .C(_3954__bF$buf1),
    .D(_5101_),
    .Y(_5103_)
);

FILL FILL_2__7497_ (
);

FILL FILL_2__7077_ (
);

FILL SFILL114840x69050 (
);

FILL FILL_6__13664_ (
);

FILL FILL_6__13244_ (
);

FILL FILL_5__12657_ (
);

FILL FILL_5__12237_ (
);

FILL FILL_3__13691_ (
);

FILL FILL_3__13271_ (
);

NAND2X1 _6957_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_39_)
);

FILL FILL_4__8784_ (
);

FILL FILL_4__8364_ (
);

FILL FILL_2__12264_ (
);

FILL FILL_1__11677_ (
);

FILL FILL_1__11257_ (
);

FILL SFILL69400x21050 (
);

FILL FILL_5__16070_ (
);

FILL SFILL74280x72050 (
);

NAND3X1 _10955_ (
    .A(_2084_),
    .B(_2072_),
    .C(_2087_),
    .Y(_2088_)
);

FILL FILL_0__8264_ (
);

NAND2X1 _10535_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1855_)
);

NAND2X1 _10115_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1636_)
);

FILL FILL_4__15483_ (
);

FILL FILL_4__15063_ (
);

FILL FILL_2__9643_ (
);

FILL FILL_3__14896_ (
);

FILL FILL_3__14476_ (
);

FILL FILL_2__9223_ (
);

FILL FILL_0__11611_ (
);

FILL FILL_3__14056_ (
);

FILL FILL_1__15090_ (
);

FILL FILL_4__9989_ (
);

FILL FILL_4__9149_ (
);

FILL FILL_2__13889_ (
);

FILL FILL_2__13469_ (
);

FILL FILL_0__14083_ (
);

FILL FILL_5__14803_ (
);

FILL SFILL114440x10050 (
);

FILL FILL_1__7220_ (
);

FILL FILL_2__14830_ (
);

FILL FILL_6_CLKBUF1_insert183 (
);

FILL FILL_0__9889_ (
);

FILL FILL_2__14410_ (
);

FILL FILL_3__7986_ (
);

FILL SFILL74200x70050 (
);

FILL FILL_3__7566_ (
);

FILL FILL_0__9469_ (
);

FILL FILL_6_CLKBUF1_insert188 (
);

FILL FILL_1__13823_ (
);

FILL FILL_1__13403_ (
);

FILL FILL_4__16268_ (
);

FILL FILL_1__16295_ (
);

FILL SFILL17880x62050 (
);

FILL FILL_5__8853_ (
);

FILL FILL_3__10396_ (
);

FILL FILL_5__8013_ (
);

NOR2X1 _15993_ (
    .A(_6448_),
    .B(_6449_),
    .Y(_6450_)
);

AOI21X1 _15573_ (
    .A(_6017_),
    .B(_6040_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [12])
);

FILL FILL_0__15288_ (
);

INVX1 _15153_ (
    .A(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_5631_)
);

FILL FILL_3__16202_ (
);

FILL FILL_1__8845_ (
);

FILL FILL_5__10303_ (
);

FILL FILL_1__8005_ (
);

FILL FILL_4_CLKBUF1_insert1080 (
);

FILL FILL_4_CLKBUF1_insert1081 (
);

FILL FILL_2__15615_ (
);

FILL FILL_4_CLKBUF1_insert1082 (
);

FILL FILL_4_CLKBUF1_insert1083 (
);

FILL FILL_4__6850_ (
);

FILL FILL_2__10750_ (
);

FILL FILL_1__14608_ (
);

INVX1 _7495_ (
    .A(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_316_)
);

INVX1 _7075_ (
    .A(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_97_)
);

FILL FILL_4__12188_ (
);

FILL FILL_5__9638_ (
);

FILL FILL_5__9218_ (
);

FILL FILL_6__12515_ (
);

NAND2X1 _16358_ (
    .A(gnd),
    .B(gnd),
    .Y(_6793_)
);

OAI21X1 _11493_ (
    .A(_2604_),
    .B(_2297_),
    .C(_2470__bF$buf2),
    .Y(_2606_)
);

FILL FILL_5__11928_ (
);

NOR2X1 _11073_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2192_)
);

FILL FILL_3__12962_ (
);

FILL FILL_5__11508_ (
);

FILL SFILL95080x30050 (
);

FILL FILL_3__12122_ (
);

FILL FILL_4__7635_ (
);

FILL FILL_4__7215_ (
);

FILL FILL_2__11955_ (
);

FILL FILL_2__11535_ (
);

FILL FILL_2__11115_ (
);

FILL FILL_3_CLKBUF1_insert130 (
);

FILL FILL_3_CLKBUF1_insert131 (
);

FILL FILL_3_CLKBUF1_insert132 (
);

FILL FILL_3_CLKBUF1_insert133 (
);

FILL FILL_3_CLKBUF1_insert134 (
);

FILL FILL_1__10948_ (
);

FILL FILL_3_CLKBUF1_insert135 (
);

FILL FILL_1__10528_ (
);

FILL FILL_3_CLKBUF1_insert136 (
);

FILL FILL_3_CLKBUF1_insert137 (
);

FILL FILL_1__10108_ (
);

FILL FILL_3_CLKBUF1_insert138 (
);

FILL FILL_3_CLKBUF1_insert139 (
);

FILL FILL_5__15761_ (
);

FILL FILL_5__15341_ (
);

FILL FILL_0__7955_ (
);

FILL FILL112440x66050 (
);

FILL FILL_0__7115_ (
);

INVX1 _9641_ (
    .A(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_1401_)
);

INVX1 _9221_ (
    .A(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_1182_)
);

FILL SFILL104360x15050 (
);

FILL FILL_4__14754_ (
);

FILL FILL_4__14334_ (
);

INVX1 _12698_ (
    .A(\aluControl_1.inst [1]),
    .Y(_3491_)
);

NAND3X1 _12278_ (
    .A(_3245_),
    .B(_3246_),
    .C(_3247_),
    .Y(\datapath_1.alu_1.ALUInB [15])
);

FILL FILL_2__8914_ (
);

FILL FILL_3__13747_ (
);

FILL SFILL108600x66050 (
);

FILL FILL_3__13327_ (
);

FILL FILL_1__14781_ (
);

FILL FILL_1__14361_ (
);

FILL FILL112040x52050 (
);

FILL FILL_0__13774_ (
);

FILL FILL_0__13354_ (
);

FILL FILL_5__9391_ (
);

FILL FILL_1__6911_ (
);

FILL FILL_3__6837_ (
);

FILL FILL_5__16126_ (
);

FILL FILL_5__11681_ (
);

FILL FILL_1__9383_ (
);

FILL FILL_5__11261_ (
);

FILL FILL_4__15959_ (
);

FILL FILL112440x21050 (
);

FILL FILL_4__15539_ (
);

FILL FILL_4__15119_ (
);

FILL FILL_2__16153_ (
);

FILL FILL_4__10674_ (
);

FILL FILL_4__10254_ (
);

FILL FILL_1__15986_ (
);

FILL FILL_1__15566_ (
);

FILL FILL_1__15146_ (
);

FILL FILL_5__7704_ (
);

FILL FILL_1__10281_ (
);

FILL FILL_0__14979_ (
);

FILL FILL_0__14559_ (
);

OAI22X1 _14844_ (
    .A(_5325_),
    .B(_3893__bF$buf2),
    .C(_3959_),
    .D(_5326_),
    .Y(_5327_)
);

FILL FILL_0__14139_ (
);

INVX1 _14424_ (
    .A(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_4916_)
);

AOI21X1 _14004_ (
    .A(\datapath_1.regfile_1.regOut[24] [11]),
    .B(_4079__bF$buf3),
    .C(_4504_),
    .Y(_4505_)
);

FILL FILL_0__15920_ (
);

FILL FILL_0__15500_ (
);

FILL FILL_5__12886_ (
);

FILL FILL_5__12466_ (
);

FILL FILL_5__12046_ (
);

FILL FILL_3__13080_ (
);

FILL FILL_4__8593_ (
);

FILL FILL_4__11879_ (
);

FILL FILL_4__11459_ (
);

FILL FILL_2__12493_ (
);

FILL FILL_4__11039_ (
);

FILL FILL_2__12073_ (
);

FILL FILL_5__8909_ (
);

FILL FILL_1__11486_ (
);

FILL FILL_1__11066_ (
);

NOR2X1 _15629_ (
    .A(_6084_),
    .B(_6094_),
    .Y(_6095_)
);

FILL FILL_4__12400_ (
);

INVX4 _15209_ (
    .A(_5472__bF$buf2),
    .Y(_5685_)
);

FILL FILL_0__10899_ (
);

FILL FILL_0__8493_ (
);

NAND2X1 _10764_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1967_)
);

FILL FILL_0__8073_ (
);

FILL FILL_0__10059_ (
);

DFFSR _10344_ (
    .Q(\datapath_1.regfile_1.regOut[27] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_1693_[18])
);

FILL FILL_3__11813_ (
);

FILL FILL_4__15292_ (
);

FILL FILL_4__6906_ (
);

FILL SFILL94280x26050 (
);

FILL FILL_2__9872_ (
);

FILL FILL_2__10806_ (
);

FILL FILL_0__11840_ (
);

FILL FILL_3__14285_ (
);

FILL FILL_0__11420_ (
);

FILL FILL_2__9032_ (
);

FILL FILL_0__11000_ (
);

FILL FILL_4__9798_ (
);

FILL FILL_4__9378_ (
);

FILL FILL_2__13698_ (
);

FILL FILL_2__13278_ (
);

FILL FILL_5__14612_ (
);

INVX1 _8912_ (
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_1037_)
);

FILL FILL_4__13605_ (
);

FILL FILL_0__9278_ (
);

FILL FILL_3__7375_ (
);

NAND2X1 _11969_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[27]),
    .Y(_3021_)
);

NAND3X1 _11549_ (
    .A(_2653_),
    .B(_2656_),
    .C(_2658_),
    .Y(\datapath_1.ALUResult [22])
);

FILL FILL_5_CLKBUF1_insert170 (
);

NAND2X1 _11129_ (
    .A(_2247_),
    .B(_2245_),
    .Y(_2248_)
);

FILL FILL_5_CLKBUF1_insert171 (
);

FILL FILL_5_CLKBUF1_insert172 (
);

FILL FILL_1__13632_ (
);

FILL FILL_5_CLKBUF1_insert173 (
);

FILL FILL_1__13212_ (
);

FILL FILL_5_CLKBUF1_insert174 (
);

FILL FILL_4__16077_ (
);

FILL FILL_5_CLKBUF1_insert175 (
);

FILL FILL_5_CLKBUF1_insert176 (
);

FILL SFILL84280x69050 (
);

FILL FILL_5_CLKBUF1_insert177 (
);

FILL FILL_5_CLKBUF1_insert178 (
);

FILL FILL_1_BUFX2_insert400 (
);

FILL FILL_1_BUFX2_insert401 (
);

FILL FILL_5_CLKBUF1_insert179 (
);

FILL FILL_1_BUFX2_insert402 (
);

FILL FILL_0__12625_ (
);

INVX1 _12910_ (
    .A(\datapath_1.a [29]),
    .Y(_3612_)
);

FILL FILL_1_BUFX2_insert403 (
);

FILL FILL_0__12205_ (
);

FILL FILL_1_BUFX2_insert404 (
);

FILL FILL_1_BUFX2_insert405 (
);

FILL FILL_1_BUFX2_insert406 (
);

FILL FILL_6_BUFX2_insert960 (
);

FILL FILL_1_BUFX2_insert407 (
);

FILL FILL_5__8242_ (
);

FILL FILL_1_BUFX2_insert408 (
);

FILL FILL_1_BUFX2_insert409 (
);

AOI22X1 _15382_ (
    .A(\datapath_1.regfile_1.regOut[1] [8]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_5854_)
);

FILL FILL_0__15097_ (
);

FILL FILL_6_BUFX2_insert966 (
);

FILL FILL_5__15817_ (
);

FILL FILL_3__16011_ (
);

FILL FILL_5__10952_ (
);

FILL FILL_1__8654_ (
);

FILL FILL_5__10532_ (
);

FILL FILL_5__10112_ (
);

FILL FILL_1__8234_ (
);

FILL SFILL8680x43050 (
);

FILL FILL_2__15844_ (
);

FILL FILL_2__15424_ (
);

FILL FILL_2__15004_ (
);

FILL SFILL109560x60050 (
);

FILL FILL_1__14837_ (
);

FILL FILL_1__14417_ (
);

FILL SFILL84200x67050 (
);

FILL FILL_3__9941_ (
);

FILL FILL_3__9521_ (
);

FILL FILL_3__9101_ (
);

FILL SFILL84280x24050 (
);

FILL FILL_2__6997_ (
);

FILL FILL_5__9867_ (
);

FILL FILL_5__9027_ (
);

INVX1 _16167_ (
    .A(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_6619_)
);

FILL FILL_1__9859_ (
);

FILL FILL_5__11737_ (
);

FILL FILL_3__12771_ (
);

FILL FILL_5__11317_ (
);

FILL FILL_1__9019_ (
);

FILL FILL_3__12351_ (
);

FILL SFILL8600x41050 (
);

FILL SFILL84600x36050 (
);

FILL FILL_2__16209_ (
);

FILL FILL_4__7864_ (
);

FILL FILL_4__7444_ (
);

FILL FILL_2__11764_ (
);

FILL FILL_2__11344_ (
);

OAI21X1 _8089_ (
    .A(_609_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .C(_610_),
    .Y(_588_[11])
);

FILL FILL_1__10757_ (
);

FILL FILL_2_CLKBUF1_insert120 (
);

FILL FILL_2_CLKBUF1_insert121 (
);

FILL FILL_5__15990_ (
);

FILL FILL_2_CLKBUF1_insert122 (
);

FILL FILL_2_CLKBUF1_insert123 (
);

FILL FILL_5__15570_ (
);

FILL FILL_0__7764_ (
);

FILL FILL_2_CLKBUF1_insert124 (
);

FILL FILL_5__15150_ (
);

INVX1 _9870_ (
    .A(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_1513_)
);

FILL FILL_0__7344_ (
);

FILL FILL_2_CLKBUF1_insert125 (
);

FILL FILL_2_CLKBUF1_insert126 (
);

DFFSR _9450_ (
    .Q(\datapath_1.regfile_1.regOut[20] [20]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_1238_[20])
);

OAI21X1 _9030_ (
    .A(_1094_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .C(_1095_),
    .Y(_1043_[26])
);

FILL FILL_2_CLKBUF1_insert127 (
);

FILL FILL_2_CLKBUF1_insert128 (
);

FILL FILL_4__14983_ (
);

FILL FILL_2_CLKBUF1_insert129 (
);

FILL FILL_4__14563_ (
);

FILL FILL_4__14143_ (
);

FILL SFILL13640x42050 (
);

NAND3X1 _12087_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[25]),
    .C(_3032__bF$buf2),
    .Y(_3111_)
);

FILL FILL_3__13976_ (
);

FILL FILL_2__8723_ (
);

FILL FILL_3__13556_ (
);

FILL FILL_1__14590_ (
);

FILL FILL_3__13136_ (
);

FILL FILL_1__14170_ (
);

FILL FILL_6_BUFX2_insert1001 (
);

FILL FILL_4__8649_ (
);

FILL FILL_4__8229_ (
);

FILL FILL_5_BUFX2_insert980 (
);

FILL FILL_2__12969_ (
);

FILL FILL_5_BUFX2_insert981 (
);

FILL SFILL53720x38050 (
);

FILL FILL_5_BUFX2_insert982 (
);

FILL FILL_5_BUFX2_insert983 (
);

FILL FILL_2__12129_ (
);

FILL FILL_0__13583_ (
);

FILL FILL_0__13163_ (
);

FILL FILL_5_BUFX2_insert984 (
);

FILL FILL_6_BUFX2_insert1007 (
);

FILL FILL_5_BUFX2_insert985 (
);

FILL FILL_5_BUFX2_insert986 (
);

FILL FILL_5_BUFX2_insert987 (
);

FILL FILL_5_BUFX2_insert988 (
);

FILL FILL_5_BUFX2_insert989 (
);

FILL FILL_2__13910_ (
);

FILL SFILL74200x65050 (
);

FILL FILL_0__8969_ (
);

FILL FILL_5__16355_ (
);

FILL FILL_0__8129_ (
);

FILL FILL_5__11490_ (
);

FILL FILL_5__11070_ (
);

FILL SFILL74280x22050 (
);

FILL FILL_1__12903_ (
);

FILL FILL_4__15768_ (
);

FILL FILL_4__15348_ (
);

FILL FILL_2__16382_ (
);

FILL FILL_0__9910_ (
);

FILL FILL_4__10063_ (
);

FILL FILL_2__9928_ (
);

FILL FILL_2__9508_ (
);

FILL FILL_1__15795_ (
);

FILL FILL_1__15375_ (
);

FILL FILL_5__7933_ (
);

FILL FILL_0__14788_ (
);

FILL FILL_0__14368_ (
);

OAI22X1 _14653_ (
    .A(_5138_),
    .B(_3893__bF$buf3),
    .C(_3944__bF$buf1),
    .D(_5139_),
    .Y(_5140_)
);

OAI22X1 _14233_ (
    .A(_3959_),
    .B(_4728_),
    .C(_3954__bF$buf1),
    .D(_4727_),
    .Y(_4729_)
);

FILL FILL_3__15702_ (
);

FILL FILL_1__7505_ (
);

FILL FILL_5__12695_ (
);

FILL FILL_5__12275_ (
);

FILL SFILL74200x20050 (
);

INVX1 _6995_ (
    .A(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_64_)
);

FILL FILL_4__11688_ (
);

FILL FILL_4__11268_ (
);

FILL FILL_5__8718_ (
);

FILL FILL_1__11295_ (
);

NAND2X1 _15858_ (
    .A(\datapath_1.regfile_1.regOut[8] [20]),
    .B(_5579_),
    .Y(_6318_)
);

OAI22X1 _15438_ (
    .A(_4425_),
    .B(_5545__bF$buf3),
    .C(_5485__bF$buf0),
    .D(_4422_),
    .Y(_5909_)
);

INVX1 _15018_ (
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_5498_)
);

INVX1 _10993_ (
    .A(\datapath_1.alu_1.ALUInA [30]),
    .Y(_2112_)
);

INVX1 _10573_ (
    .A(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_1880_)
);

FILL FILL_0__10288_ (
);

FILL FILL_3_BUFX2_insert1060 (
);

INVX1 _10153_ (
    .A(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_1661_)
);

FILL FILL_3_BUFX2_insert1061 (
);

FILL FILL_6__14487_ (
);

FILL FILL_3_BUFX2_insert1062 (
);

FILL FILL_3__11622_ (
);

FILL FILL_3__11202_ (
);

FILL FILL_3_BUFX2_insert1063 (
);

FILL FILL_3_BUFX2_insert1064 (
);

FILL FILL_3_BUFX2_insert1065 (
);

FILL FILL_3_BUFX2_insert1066 (
);

FILL FILL_3_BUFX2_insert1067 (
);

FILL FILL_3_BUFX2_insert1068 (
);

FILL FILL_2__10615_ (
);

FILL FILL_2__9681_ (
);

FILL FILL_3_BUFX2_insert1069 (
);

FILL SFILL33800x72050 (
);

FILL FILL_2__9261_ (
);

FILL SFILL64200x63050 (
);

FILL FILL_3__14094_ (
);

FILL FILL_2__13087_ (
);

FILL FILL_5__14841_ (
);

FILL FILL_5__14421_ (
);

FILL FILL_5__14001_ (
);

INVX1 _8721_ (
    .A(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_930_)
);

DFFSR _8301_ (
    .Q(\datapath_1.regfile_1.regOut[11] [23]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_653_[23])
);

FILL FILL_4__13834_ (
);

FILL FILL_4__13414_ (
);

FILL FILL_3__7184_ (
);

FILL FILL_0__9087_ (
);

OAI21X1 _11778_ (
    .A(_2558_),
    .B(_2344__bF$buf3),
    .C(_2871_),
    .Y(_2872_)
);

AOI21X1 _11358_ (
    .A(_2474_),
    .B(_2450_),
    .C(_2321_),
    .Y(_2475_)
);

FILL FILL_3__12827_ (
);

FILL FILL_3__12407_ (
);

FILL FILL_1__13861_ (
);

FILL SFILL113960x74050 (
);

FILL FILL_1__13441_ (
);

FILL FILL_1__13021_ (
);

FILL FILL_4_CLKBUF1_insert160 (
);

FILL FILL_4_CLKBUF1_insert161 (
);

FILL FILL_4_CLKBUF1_insert162 (
);

FILL FILL_0__12854_ (
);

FILL FILL_0__12434_ (
);

FILL FILL_3__15299_ (
);

FILL FILL_4_CLKBUF1_insert163 (
);

FILL FILL_0__12014_ (
);

FILL FILL_4_CLKBUF1_insert164 (
);

FILL FILL_4_CLKBUF1_insert165 (
);

FILL FILL_4_CLKBUF1_insert166 (
);

FILL FILL_5__8891_ (
);

FILL FILL_5__8471_ (
);

FILL FILL_4_CLKBUF1_insert167 (
);

FILL FILL_4_CLKBUF1_insert168 (
);

FILL FILL_4_CLKBUF1_insert169 (
);

OAI22X1 _15191_ (
    .A(_5478__bF$buf0),
    .B(_5667_),
    .C(_5666_),
    .D(_5480__bF$buf0),
    .Y(_5668_)
);

FILL FILL_5__15626_ (
);

FILL FILL_5__15206_ (
);

FILL FILL_3__16240_ (
);

OAI21X1 _9926_ (
    .A(_1549_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1550_),
    .Y(_1498_[26])
);

FILL SFILL9480x42050 (
);

OAI21X1 _9506_ (
    .A(_1330_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1331_),
    .Y(_1303_[14])
);

FILL FILL_5__10761_ (
);

FILL FILL_1__8883_ (
);

FILL FILL_1__8463_ (
);

FILL FILL112440x16050 (
);

FILL FILL_4__14619_ (
);

FILL FILL_2__15653_ (
);

FILL FILL_2__15233_ (
);

FILL FILL_3__8389_ (
);

FILL FILL_1__14646_ (
);

FILL FILL_1__14226_ (
);

FILL SFILL49320x19050 (
);

FILL FILL_3__9750_ (
);

FILL FILL_0__13639_ (
);

OAI22X1 _13924_ (
    .A(_4425_),
    .B(_3925_),
    .C(_3971__bF$buf2),
    .D(_4426_),
    .Y(_4427_)
);

FILL FILL_0__13219_ (
);

NOR2X1 _13504_ (
    .A(_4014_),
    .B(_4000_),
    .Y(_4015_)
);

FILL FILL_5__9676_ (
);

FILL FILL_5__9256_ (
);

INVX1 _16396_ (
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .Y(_6818_)
);

FILL FILL_5__11966_ (
);

FILL FILL_1__9668_ (
);

FILL FILL_5__11546_ (
);

FILL FILL_3__12580_ (
);

FILL FILL_1__9248_ (
);

FILL FILL_5__11126_ (
);

FILL FILL_3__12160_ (
);

FILL FILL_2__16018_ (
);

FILL FILL_4__7673_ (
);

FILL FILL_4__10959_ (
);

FILL FILL_4__7253_ (
);

FILL FILL_4__10539_ (
);

FILL FILL_2__11993_ (
);

FILL FILL_2__11573_ (
);

FILL FILL_4__10119_ (
);

FILL FILL_2__11153_ (
);

FILL SFILL23720x77050 (
);

FILL FILL_1__10566_ (
);

FILL FILL_1__10146_ (
);

FILL FILL_4__11900_ (
);

NOR2X1 _14709_ (
    .A(_5194_),
    .B(_5191_),
    .Y(_5195_)
);

FILL FILL_0__7993_ (
);

FILL FILL_0__7573_ (
);

FILL FILL_1_CLKBUF1_insert111 (
);

FILL FILL_1_CLKBUF1_insert112 (
);

FILL FILL_4__14792_ (
);

FILL FILL_4__14372_ (
);

FILL FILL_1_CLKBUF1_insert113 (
);

FILL FILL_1_CLKBUF1_insert114 (
);

FILL FILL_1_CLKBUF1_insert115 (
);

FILL FILL_1_CLKBUF1_insert116 (
);

FILL FILL_1_CLKBUF1_insert117 (
);

FILL FILL_1_CLKBUF1_insert118 (
);

FILL FILL_2__8952_ (
);

FILL FILL_1_CLKBUF1_insert119 (
);

FILL FILL_0__10920_ (
);

FILL FILL_3__13785_ (
);

FILL FILL_2__8532_ (
);

FILL FILL_3__13365_ (
);

FILL FILL_0__10500_ (
);

FILL FILL_2__8112_ (
);

FILL FILL_4__8878_ (
);

FILL FILL_4__8458_ (
);

FILL FILL_2__12778_ (
);

FILL FILL_2__12358_ (
);

FILL FILL_0__13392_ (
);

FILL FILL_0__8778_ (
);

FILL FILL_3__6875_ (
);

FILL FILL_5__16164_ (
);

FILL FILL_0__8358_ (
);

INVX1 _10629_ (
    .A(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_1897_)
);

DFFSR _10209_ (
    .Q(\datapath_1.regfile_1.regOut[26] [11]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_1628_[11])
);

FILL FILL_4__15997_ (
);

FILL FILL_1__12712_ (
);

FILL FILL_4__15577_ (
);

FILL FILL_4__15157_ (
);

FILL SFILL48920x81050 (
);

FILL FILL_2__16191_ (
);

FILL FILL_4__10292_ (
);

FILL FILL_2__9737_ (
);

FILL FILL_0__11705_ (
);

FILL FILL_1__15184_ (
);

FILL FILL_5__7742_ (
);

FILL FILL_5__7322_ (
);

FILL SFILL23640x39050 (
);

FILL FILL_0__14597_ (
);

INVX1 _14882_ (
    .A(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_5364_)
);

FILL SFILL59720x5050 (
);

INVX1 _14462_ (
    .A(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_4953_)
);

FILL FILL_0__14177_ (
);

NOR2X1 _14042_ (
    .A(_4541_),
    .B(_3890_),
    .Y(_4542_)
);

FILL FILL_3__15931_ (
);

FILL FILL_3__15511_ (
);

FILL FILL_1__7734_ (
);

FILL FILL_1__7314_ (
);

FILL SFILL13720x75050 (
);

FILL FILL_2__14924_ (
);

FILL FILL_2__14504_ (
);

FILL SFILL109560x55050 (
);

FILL FILL_5__12084_ (
);

FILL FILL_1__13917_ (
);

FILL SFILL99560x2050 (
);

FILL FILL_4__11497_ (
);

FILL FILL_4__11077_ (
);

FILL FILL_3__8601_ (
);

FILL SFILL84280x19050 (
);

FILL FILL_1__16389_ (
);

FILL FILL_5__8527_ (
);

FILL FILL_5__8107_ (
);

FILL FILL_6__11824_ (
);

NAND3X1 _15667_ (
    .A(_6126_),
    .B(_6127_),
    .C(_6131_),
    .Y(_6132_)
);

OAI22X1 _15247_ (
    .A(_4176_),
    .B(_5518__bF$buf2),
    .C(_5478__bF$buf1),
    .D(_4175_),
    .Y(_5723_)
);

FILL SFILL99160x1050 (
);

FILL SFILL109960x24050 (
);

INVX1 _10382_ (
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_1773_)
);

FILL FILL_5__10817_ (
);

FILL FILL_1__8519_ (
);

FILL FILL_3__11851_ (
);

FILL SFILL8600x36050 (
);

FILL FILL_3__11431_ (
);

FILL FILL_3__11011_ (
);

FILL FILL_2__15709_ (
);

FILL FILL_4__6944_ (
);

FILL FILL_0__16323_ (
);

FILL SFILL13240x68050 (
);

FILL SFILL13720x30050 (
);

FILL FILL_5__13289_ (
);

FILL FILL_2__10424_ (
);

FILL FILL_2__9490_ (
);

FILL FILL_2__10004_ (
);

OAI21X1 _7589_ (
    .A(_357_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .C(_358_),
    .Y(_328_[15])
);

OAI21X1 _7169_ (
    .A(_138_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .C(_139_),
    .Y(_133_[3])
);

FILL SFILL109560x10050 (
);

FILL FILL_3__9806_ (
);

FILL FILL_5__14650_ (
);

FILL FILL_5__14230_ (
);

FILL FILL_0__6844_ (
);

INVX1 _8950_ (
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_1106_)
);

OAI21X1 _8530_ (
    .A(_842_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .C(_843_),
    .Y(_783_[30])
);

OAI21X1 _8110_ (
    .A(_623_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .C(_624_),
    .Y(_588_[18])
);

FILL FILL_6__12609_ (
);

FILL FILL_4__13643_ (
);

FILL FILL_4__13223_ (
);

FILL SFILL13640x37050 (
);

OAI21X1 _11587_ (
    .A(_2693_),
    .B(_2269_),
    .C(_2692_),
    .Y(_2694_)
);

NAND2X1 _11167_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2286_)
);

FILL FILL_2__7803_ (
);

FILL FILL_3__12636_ (
);

FILL SFILL109480x17050 (
);

FILL FILL_1__13670_ (
);

FILL FILL_3__12216_ (
);

FILL FILL_1__13250_ (
);

FILL FILL_4__7729_ (
);

FILL FILL_4__7309_ (
);

FILL FILL_2__11629_ (
);

FILL FILL_2__11209_ (
);

FILL FILL_0__12243_ (
);

FILL FILL_6__16022_ (
);

FILL FILL_5__15855_ (
);

FILL FILL_5__15435_ (
);

FILL FILL_0__7629_ (
);

FILL FILL_5__15015_ (
);

FILL FILL_0__7209_ (
);

OAI21X1 _9735_ (
    .A(_1442_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1443_),
    .Y(_1433_[5])
);

FILL FILL_5__10990_ (
);

DFFSR _9315_ (
    .Q(\datapath_1.regfile_1.regOut[19] [13]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_1173_[13])
);

FILL FILL_5__10570_ (
);

FILL SFILL74280x17050 (
);

FILL FILL_5__10150_ (
);

FILL FILL_1__8272_ (
);

FILL FILL_4__14848_ (
);

FILL FILL_2__15882_ (
);

FILL FILL_4__14428_ (
);

FILL FILL_4__14008_ (
);

FILL FILL_2__15462_ (
);

FILL FILL_2__15042_ (
);

FILL FILL_3__8198_ (
);

FILL FILL112200x73050 (
);

FILL FILL_1__14875_ (
);

FILL SFILL99480x66050 (
);

FILL FILL_1__14455_ (
);

FILL FILL_1__14035_ (
);

FILL FILL_0__13868_ (
);

FILL FILL_0__13448_ (
);

OAI22X1 _13733_ (
    .A(_4239_),
    .B(_3936__bF$buf4),
    .C(_3972__bF$buf3),
    .D(_4238_),
    .Y(_4240_)
);

NAND3X1 _13313_ (
    .A(_3841_),
    .B(_3845_),
    .C(_3788_),
    .Y(_3846_)
);

FILL FILL_0__13028_ (
);

FILL SFILL38840x41050 (
);

FILL FILL_5__9485_ (
);

FILL FILL_6__12362_ (
);

FILL FILL_5__11775_ (
);

FILL FILL_1__9897_ (
);

FILL SFILL74200x15050 (
);

FILL FILL_5__11355_ (
);

FILL FILL_1__9477_ (
);

FILL FILL_2__16247_ (
);

FILL FILL_4__7482_ (
);

FILL FILL_4__10768_ (
);

FILL FILL_4__7062_ (
);

FILL FILL_2__11382_ (
);

FILL FILL_1__10795_ (
);

FILL FILL_1__10375_ (
);

FILL SFILL99480x21050 (
);

NOR2X1 _14938_ (
    .A(_5415_),
    .B(_5418_),
    .Y(_5419_)
);

OAI22X1 _14518_ (
    .A(_5006_),
    .B(_3905__bF$buf2),
    .C(_3977__bF$buf3),
    .D(_5007_),
    .Y(_5008_)
);

FILL FILL_3__10702_ (
);

FILL FILL_6__13567_ (
);

FILL FILL_4__14181_ (
);

FILL SFILL33800x67050 (
);

FILL FILL_2__8761_ (
);

FILL SFILL64200x58050 (
);

FILL FILL_3__13594_ (
);

FILL FILL_2__8341_ (
);

FILL FILL_3__13174_ (
);

FILL FILL_4__8267_ (
);

FILL FILL_2__12587_ (
);

FILL FILL_2__12167_ (
);

FILL FILL_5__13921_ (
);

FILL FILL_5__13501_ (
);

INVX1 _7801_ (
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_459_)
);

FILL FILL_4__12914_ (
);

FILL FILL_5__16393_ (
);

FILL FILL_0__8587_ (
);

FILL FILL_6__9974_ (
);

DFFSR _10858_ (
    .Q(\datapath_1.regfile_1.regOut[31] [20]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_1953_[20])
);

FILL FILL_6__9554_ (
);

OAI21X1 _10438_ (
    .A(_1809_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .C(_1810_),
    .Y(_1758_[26])
);

OAI21X1 _10018_ (
    .A(_1590_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1591_),
    .Y(_1563_[14])
);

FILL FILL_3__11907_ (
);

FILL FILL_4__15386_ (
);

FILL FILL_1__12521_ (
);

FILL FILL_1__12101_ (
);

FILL FILL_2__9546_ (
);

FILL FILL_0__11934_ (
);

FILL FILL_3__14799_ (
);

FILL FILL_2__9126_ (
);

FILL FILL_3__14379_ (
);

FILL FILL_0__11514_ (
);

FILL FILL_5__7971_ (
);

FILL FILL_5__7551_ (
);

FILL SFILL64200x13050 (
);

NOR2X1 _14691_ (
    .A(_5177_),
    .B(_5167_),
    .Y(_5178_)
);

OAI22X1 _14271_ (
    .A(_4765_),
    .B(_3902__bF$buf2),
    .C(_3966__bF$buf2),
    .D(_4764_),
    .Y(_4766_)
);

FILL FILL_5__14706_ (
);

FILL FILL_3__15740_ (
);

FILL FILL_3__15320_ (
);

FILL FILL_1__7963_ (
);

FILL FILL_1__7543_ (
);

FILL FILL_1__7123_ (
);

FILL FILL_2__14733_ (
);

FILL FILL_2__14313_ (
);

FILL FILL_3__7889_ (
);

FILL FILL_3__7469_ (
);

FILL FILL_3__7049_ (
);

FILL FILL_1__13726_ (
);

FILL FILL_1__13306_ (
);

FILL SFILL18840x82050 (
);

FILL FILL_3__8830_ (
);

FILL FILL_0__12719_ (
);

FILL FILL_1__16198_ (
);

FILL FILL_5__8756_ (
);

FILL FILL_5__8336_ (
);

FILL FILL_3__10299_ (
);

NOR3X1 _15896_ (
    .A(_6352_),
    .B(_6354_),
    .C(_6353_),
    .Y(_6355_)
);

OAI22X1 _15476_ (
    .A(_5466__bF$buf1),
    .B(_5945_),
    .C(_4434_),
    .D(_5483__bF$buf0),
    .Y(_5946_)
);

OAI22X1 _15056_ (
    .A(_3896_),
    .B(_5535__bF$buf2),
    .C(_5534__bF$buf4),
    .D(_3980_),
    .Y(_5536_)
);

FILL FILL_3__16105_ (
);

OAI21X1 _10191_ (
    .A(_1685_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .C(_1686_),
    .Y(_1628_[29])
);

FILL FILL_5__10626_ (
);

FILL FILL_1__8748_ (
);

FILL FILL_1__8328_ (
);

FILL FILL_3__11660_ (
);

FILL FILL_3__11240_ (
);

FILL FILL_2__15938_ (
);

FILL FILL_2__15518_ (
);

FILL FILL_0__16132_ (
);

FILL FILL_2__10653_ (
);

FILL FILL_5__13098_ (
);

FILL FILL_2__10233_ (
);

DFFSR _7398_ (
    .Q(\datapath_1.regfile_1.regOut[4] [16]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_198_[16])
);

FILL FILL_3__9615_ (
);

FILL FILL_3_BUFX2_insert310 (
);

FILL FILL_3_BUFX2_insert311 (
);

FILL FILL_3_BUFX2_insert312 (
);

FILL FILL_3_BUFX2_insert313 (
);

FILL FILL_3_BUFX2_insert314 (
);

FILL FILL_3_BUFX2_insert315 (
);

FILL FILL_3_BUFX2_insert316 (
);

FILL FILL_3_BUFX2_insert317 (
);

FILL FILL_3_BUFX2_insert318 (
);

FILL FILL_4__13872_ (
);

FILL FILL_6__12418_ (
);

FILL FILL_3_BUFX2_insert319 (
);

FILL FILL_4__13452_ (
);

FILL FILL_4__13032_ (
);

AOI21X1 _11396_ (
    .A(_2173_),
    .B(_2509_),
    .C(_2512_),
    .Y(_2513_)
);

FILL FILL_2__7612_ (
);

FILL FILL_3__12865_ (
);

FILL FILL_3__12445_ (
);

FILL FILL_3__12025_ (
);

FILL FILL_4__7958_ (
);

FILL FILL_4__7118_ (
);

FILL FILL_2__11858_ (
);

FILL FILL_0__12892_ (
);

FILL FILL_2__11438_ (
);

FILL FILL_0__12472_ (
);

FILL FILL_2__11018_ (
);

FILL FILL_0__12052_ (
);

FILL SFILL74120x6050 (
);

FILL SFILL23720x27050 (
);

FILL FILL_5__15664_ (
);

FILL FILL_5__15244_ (
);

FILL FILL_0__7858_ (
);

FILL SFILL38840x2050 (
);

FILL FILL_0__7438_ (
);

DFFSR _9964_ (
    .Q(\datapath_1.regfile_1.regOut[24] [22]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1498_[22])
);

NAND2X1 _9544_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1357_)
);

NAND2X1 _9124_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1138_)
);

FILL FILL_1__8081_ (
);

FILL FILL_4__14657_ (
);

FILL FILL_2__15691_ (
);

FILL FILL_4__14237_ (
);

FILL FILL_2__15271_ (
);

FILL FILL_1__14684_ (
);

FILL FILL_1__14264_ (
);

FILL FILL_0_BUFX2_insert440 (
);

FILL FILL_0_BUFX2_insert441 (
);

FILL FILL_0_BUFX2_insert442 (
);

FILL FILL_0_BUFX2_insert443 (
);

FILL FILL_0_BUFX2_insert444 (
);

FILL FILL_0__13677_ (
);

AOI22X1 _13962_ (
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .B(_4005__bF$buf0),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_4464_)
);

FILL FILL_0__13257_ (
);

FILL FILL_0_BUFX2_insert445 (
);

AOI22X1 _13542_ (
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .B(_3891__bF$buf2),
    .C(_4051__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_4052_)
);

FILL FILL_0_BUFX2_insert446 (
);

NAND2X1 _13122_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [14]),
    .Y(_3713_)
);

FILL FILL_0_BUFX2_insert447 (
);

FILL FILL_0_BUFX2_insert448 (
);

FILL FILL_5__9294_ (
);

FILL FILL_0_BUFX2_insert449 (
);

FILL FILL_5__16449_ (
);

FILL FILL_5__16029_ (
);

FILL FILL_5__11584_ (
);

FILL FILL_1__9286_ (
);

FILL FILL_5__11164_ (
);

FILL FILL_2__16056_ (
);

FILL FILL_4__10997_ (
);

FILL FILL_4__7291_ (
);

FILL FILL_4__10577_ (
);

FILL FILL_4__10157_ (
);

FILL SFILL48920x31050 (
);

FILL FILL_2__11191_ (
);

FILL FILL_1__15889_ (
);

FILL FILL_1__15469_ (
);

FILL FILL_1__15049_ (
);

FILL SFILL109160x36050 (
);

FILL FILL_5__7607_ (
);

FILL FILL_1__10184_ (
);

INVX1 _14747_ (
    .A(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_5232_)
);

OAI22X1 _14327_ (
    .A(_3916_),
    .B(_4819_),
    .C(_3977__bF$buf4),
    .D(_4820_),
    .Y(_4821_)
);

FILL FILL_0__7191_ (
);

FILL FILL_1__16410_ (
);

FILL FILL_3__10931_ (
);

FILL FILL_3__10511_ (
);

FILL FILL_0__15823_ (
);

FILL FILL_0__15403_ (
);

FILL SFILL13720x25050 (
);

FILL FILL_5__12789_ (
);

FILL FILL_2__8990_ (
);

FILL FILL_5__12369_ (
);

FILL FILL_2__8570_ (
);

FILL FILL_4__8496_ (
);

FILL FILL_4__8076_ (
);

FILL FILL_2__12396_ (
);

FILL SFILL38920x74050 (
);

FILL FILL_5__13730_ (
);

FILL FILL_5__13310_ (
);

OAI21X1 _7610_ (
    .A(_371_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_372_),
    .Y(_328_[22])
);

FILL FILL_1__11389_ (
);

FILL FILL_4__12723_ (
);

FILL FILL_4__12303_ (
);

FILL FILL_0__8396_ (
);

OAI21X1 _10667_ (
    .A(_1921_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .C(_1922_),
    .Y(_1888_[17])
);

OAI21X1 _10247_ (
    .A(_1702_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .C(_1703_),
    .Y(_1693_[5])
);

FILL FILL_3__11716_ (
);

FILL FILL_1__12750_ (
);

FILL FILL_4__15195_ (
);

FILL FILL_1__12330_ (
);

FILL FILL_2__10709_ (
);

FILL FILL_2__9775_ (
);

FILL FILL_2__9355_ (
);

FILL FILL_0__11743_ (
);

FILL FILL_3__14188_ (
);

FILL FILL_0__11323_ (
);

FILL FILL_5__7360_ (
);

FILL SFILL3560x73050 (
);

FILL FILL_5__14935_ (
);

OAI22X1 _14080_ (
    .A(_4577_),
    .B(_3893__bF$buf3),
    .C(_3977__bF$buf2),
    .D(_4578_),
    .Y(_4579_)
);

FILL FILL_5__14515_ (
);

DFFSR _8815_ (
    .Q(\datapath_1.regfile_1.regOut[15] [25]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_913_[25])
);

FILL FILL_1__7352_ (
);

FILL FILL_4__13928_ (
);

FILL FILL_2__14962_ (
);

FILL FILL_4__13508_ (
);

FILL FILL_2__14542_ (
);

FILL FILL_3__7698_ (
);

FILL FILL_2__14122_ (
);

FILL SFILL34520x28050 (
);

FILL FILL112200x68050 (
);

FILL FILL_1__13955_ (
);

FILL FILL_1__13535_ (
);

FILL FILL_1__13115_ (
);

DFFSR _12813_ (
    .Q(\datapath_1.PCJump [24]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3490_[22])
);

FILL FILL_0__12528_ (
);

FILL FILL_0__12108_ (
);

FILL SFILL38840x36050 (
);

FILL FILL_5__8985_ (
);

FILL FILL_5__8145_ (
);

NAND2X1 _15285_ (
    .A(_5755_),
    .B(_5759_),
    .Y(_5760_)
);

FILL FILL_3__16334_ (
);

FILL SFILL28920x72050 (
);

FILL FILL_1__8977_ (
);

FILL FILL_5__10435_ (
);

FILL FILL_1__8137_ (
);

FILL FILL_5__10015_ (
);

FILL FILL_2__15747_ (
);

FILL FILL_2__15327_ (
);

FILL FILL_4__6982_ (
);

FILL FILL_0__16361_ (
);

FILL FILL_2__10882_ (
);

FILL FILL_2__10042_ (
);

FILL SFILL99480x16050 (
);

FILL FILL_3__9424_ (
);

FILL FILL_3__9004_ (
);

FILL FILL_0__6882_ (
);

FILL SFILL28840x79050 (
);

FILL FILL_4__13681_ (
);

FILL FILL_4__13261_ (
);

FILL FILL_2__7841_ (
);

FILL FILL_2__7421_ (
);

FILL FILL_3__12254_ (
);

FILL FILL_4__7347_ (
);

FILL FILL_2__11667_ (
);

FILL FILL_2__11247_ (
);

FILL FILL_0__12281_ (
);

FILL FILL_5__15893_ (
);

FILL FILL_5__15473_ (
);

FILL FILL_5__15053_ (
);

FILL FILL_0__7247_ (
);

NAND2X1 _9773_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1469_)
);

NAND2X1 _9353_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1250_)
);

FILL FILL_4__14886_ (
);

FILL SFILL28840x34050 (
);

FILL FILL_4__14466_ (
);

FILL FILL_1__11601_ (
);

FILL FILL_4__14046_ (
);

FILL FILL_2__15080_ (
);

FILL FILL_3__13879_ (
);

FILL FILL_2__8626_ (
);

FILL FILL_2__8206_ (
);

FILL FILL_3__13459_ (
);

FILL FILL_1__14493_ (
);

FILL FILL_3__13039_ (
);

FILL FILL_1__14073_ (
);

FILL SFILL33800x17050 (
);

FILL SFILL18920x70050 (
);

AOI22X1 _13771_ (
    .A(_3882__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [6]),
    .C(\datapath_1.regfile_1.regOut[13] [6]),
    .D(_4051__bF$buf3),
    .Y(_4277_)
);

FILL FILL_0__13486_ (
);

FILL SFILL28440x20050 (
);

NOR2X1 _13351_ (
    .A(_3869_),
    .B(_3867_),
    .Y(\datapath_1.regfile_1.regEn [25])
);

FILL FILL_3__14820_ (
);

FILL FILL_3__14400_ (
);

FILL SFILL79960x64050 (
);

FILL FILL_4__9913_ (
);

FILL FILL_2__13813_ (
);

FILL FILL_3__6969_ (
);

FILL FILL_5__16258_ (
);

FILL FILL_5__11393_ (
);

FILL FILL_1__9095_ (
);

FILL SFILL18840x77050 (
);

FILL FILL_2__16285_ (
);

FILL FILL_4__10386_ (
);

FILL FILL_0__9813_ (
);

FILL FILL_1__15698_ (
);

FILL FILL_1__15278_ (
);

FILL FILL_5__7836_ (
);

FILL FILL_5__7416_ (
);

NAND3X1 _14976_ (
    .A(_5446_),
    .B(_5449_),
    .C(_5456_),
    .Y(_5457_)
);

FILL SFILL13800x7050 (
);

NOR2X1 _14556_ (
    .A(_5044_),
    .B(_5041_),
    .Y(_5045_)
);

INVX1 _14136_ (
    .A(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_4634_)
);

FILL FILL_3__15605_ (
);

FILL FILL_1__7828_ (
);

FILL FILL_3__10320_ (
);

FILL FILL_0__15632_ (
);

FILL FILL_0__15212_ (
);

FILL FILL_5__12598_ (
);

FILL FILL_5__12178_ (
);

BUFX2 _6898_ (
    .A(_2_[28]),
    .Y(memoryWriteData[28])
);

FILL SFILL18840x32050 (
);

FILL FILL_1__11198_ (
);

FILL FILL_4__12952_ (
);

FILL FILL_4__12532_ (
);

FILL FILL_4__12112_ (
);

OAI21X1 _10896_ (
    .A(_2041_),
    .B(_2036_),
    .C(_2025_),
    .Y(ALUControl[2])
);

DFFSR _10476_ (
    .Q(\datapath_1.regfile_1.regOut[28] [22]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1758_[22])
);

FILL FILL_6__9172_ (
);

NAND2X1 _10056_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1617_)
);

FILL FILL_3__11945_ (
);

FILL FILL_3__11525_ (
);

FILL FILL_3__11105_ (
);

FILL FILL_2__10938_ (
);

FILL FILL_0__11972_ (
);

FILL FILL_2__10518_ (
);

FILL FILL_2__9164_ (
);

FILL FILL_0__11552_ (
);

FILL FILL_0__11132_ (
);

FILL FILL_6__15751_ (
);

FILL FILL_5__14744_ (
);

FILL FILL_0__6938_ (
);

FILL FILL_5__14324_ (
);

NAND2X1 _8624_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_886_)
);

NAND2X1 _8204_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_667_)
);

FILL FILL_1__7581_ (
);

FILL FILL_1__7161_ (
);

FILL FILL_4__13737_ (
);

FILL FILL_4__13317_ (
);

FILL FILL_2__14771_ (
);

FILL FILL_2__14351_ (
);

FILL FILL_3__7087_ (
);

FILL FILL_1__13764_ (
);

FILL FILL_1__13344_ (
);

FILL FILL_0__12757_ (
);

NAND2X1 _12622_ (
    .A(vdd),
    .B(memoryOutData[18]),
    .Y(_3461_)
);

FILL FILL_0__12337_ (
);

FILL SFILL114520x80050 (
);

INVX1 _12202_ (
    .A(\datapath_1.PCJump [29]),
    .Y(_3188_)
);

FILL SFILL53880x70050 (
);

FILL FILL_5__8374_ (
);

FILL FILL_6__11671_ (
);

FILL FILL_6__11251_ (
);

FILL FILL_5__15949_ (
);

NAND3X1 _15094_ (
    .A(_5566_),
    .B(_5568_),
    .C(_5572_),
    .Y(_5573_)
);

FILL FILL_5__15529_ (
);

FILL FILL_5__15109_ (
);

DFFSR _9829_ (
    .Q(\datapath_1.regfile_1.regOut[23] [15]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_1433_[15])
);

FILL FILL_3__16143_ (
);

INVX1 _9409_ (
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_1287_)
);

FILL FILL_5__10664_ (
);

FILL FILL_1__8786_ (
);

FILL FILL_5__10244_ (
);

FILL FILL_1__8366_ (
);

FILL FILL_2__15976_ (
);

FILL SFILL69080x41050 (
);

FILL FILL_2__15556_ (
);

FILL FILL_2__15136_ (
);

FILL FILL_0__16170_ (
);

FILL SFILL48920x26050 (
);

FILL FILL_2__10691_ (
);

FILL FILL_2__10271_ (
);

FILL FILL_1__14969_ (
);

FILL FILL_1__14549_ (
);

FILL FILL_1__14129_ (
);

FILL FILL_3__9653_ (
);

AOI22X1 _13827_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [7]),
    .C(\datapath_1.regfile_1.regOut[31] [7]),
    .D(_3995__bF$buf1),
    .Y(_4332_)
);

FILL FILL_3__9233_ (
);

NOR2X1 _13407_ (
    .A(\datapath_1.PCJump [20]),
    .B(_3918_),
    .Y(_3919_)
);

FILL FILL_5__9999_ (
);

FILL FILL_1__15910_ (
);

FILL FILL_5__9159_ (
);

FILL FILL_4__13490_ (
);

OAI21X1 _16299_ (
    .A(_5524__bF$buf0),
    .B(_5442_),
    .C(_6747_),
    .Y(_6748_)
);

FILL FILL_0__14903_ (
);

FILL FILL_5__11869_ (
);

FILL FILL_5__11449_ (
);

FILL FILL_2__7230_ (
);

FILL FILL_3__12483_ (
);

FILL FILL_5__11029_ (
);

FILL FILL_3__12063_ (
);

FILL FILL_4__7996_ (
);

FILL FILL_4__7576_ (
);

FILL FILL_2__11896_ (
);

FILL SFILL38920x69050 (
);

FILL FILL_2__11476_ (
);

FILL FILL_2__11056_ (
);

FILL FILL_0__12090_ (
);

FILL FILL_1__10889_ (
);

FILL FILL_1__10049_ (
);

FILL FILL_4__11803_ (
);

FILL SFILL3640x61050 (
);

FILL FILL_5__15282_ (
);

FILL FILL_0__7476_ (
);

FILL FILL_0__7056_ (
);

DFFSR _9582_ (
    .Q(\datapath_1.regfile_1.regOut[21] [24]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_1303_[24])
);

INVX1 _9162_ (
    .A(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_1163_)
);

FILL FILL_1__11830_ (
);

FILL FILL_4__14695_ (
);

FILL FILL_4__14275_ (
);

FILL FILL_1__11410_ (
);

FILL FILL_2__8855_ (
);

FILL FILL_0__10823_ (
);

FILL FILL_3__13688_ (
);

FILL FILL_2__8015_ (
);

FILL FILL_3__13268_ (
);

FILL FILL_0__10403_ (
);

FILL SFILL59000x82050 (
);

FILL FILL_5__6860_ (
);

FILL FILL_0_BUFX2_insert820 (
);

FILL FILL_0_BUFX2_insert821 (
);

FILL FILL_0_BUFX2_insert822 (
);

FILL FILL_0_BUFX2_insert823 (
);

FILL FILL_0_BUFX2_insert824 (
);

FILL SFILL3560x68050 (
);

FILL FILL_0__13295_ (
);

FILL FILL_0_BUFX2_insert825 (
);

INVX8 _13580_ (
    .A(_3931__bF$buf3),
    .Y(_4090_)
);

INVX1 _13160_ (
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3738_)
);

FILL FILL_0_BUFX2_insert826 (
);

FILL FILL_0_BUFX2_insert827 (
);

FILL FILL_0_BUFX2_insert828 (
);

FILL FILL_0_BUFX2_insert829 (
);

FILL FILL_1__6852_ (
);

FILL FILL_4__9722_ (
);

FILL FILL_2__13622_ (
);

FILL FILL_5__16067_ (
);

FILL FILL_6__9648_ (
);

FILL FILL_1__12615_ (
);

FILL FILL_2__16094_ (
);

FILL FILL_4__10195_ (
);

FILL FILL_0__9622_ (
);

FILL FILL_0__11608_ (
);

FILL FILL_1__15087_ (
);

FILL FILL_6__15807_ (
);

FILL FILL_5__7225_ (
);

FILL FILL_4__16001_ (
);

FILL FILL_6__10522_ (
);

NOR2X1 _14785_ (
    .A(_5269_),
    .B(_3971__bF$buf2),
    .Y(_5270_)
);

FILL SFILL49080x82050 (
);

OAI22X1 _14365_ (
    .A(_4856_),
    .B(_3931__bF$buf2),
    .C(_3960_),
    .D(_4857_),
    .Y(_4858_)
);

FILL FILL_3__15834_ (
);

FILL FILL_3__15414_ (
);

FILL SFILL28920x67050 (
);

FILL SFILL3560x23050 (
);

FILL FILL_1__7637_ (
);

FILL FILL_1__7217_ (
);

FILL FILL_2__14827_ (
);

FILL SFILL104440x40050 (
);

FILL FILL_2__14407_ (
);

FILL FILL_0__15861_ (
);

FILL FILL_0__15441_ (
);

FILL FILL_0__15021_ (
);

FILL FILL112200x18050 (
);

FILL FILL_3__8504_ (
);

FILL SFILL89560x47050 (
);

FILL FILL_6__11727_ (
);

FILL FILL_4__12761_ (
);

FILL FILL_4__12341_ (
);

NAND2X1 _10285_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1729_)
);

FILL FILL_2__6921_ (
);

FILL FILL_3__11754_ (
);

FILL FILL_3__11334_ (
);

FILL SFILL28920x22050 (
);

FILL FILL_4__6847_ (
);

FILL FILL_0__16226_ (
);

FILL FILL_2__10747_ (
);

FILL FILL_2__9393_ (
);

FILL FILL_0__11781_ (
);

FILL FILL_0__11361_ (
);

FILL FILL_5__14973_ (
);

FILL FILL_5__14553_ (
);

FILL FILL_5__14133_ (
);

NAND2X1 _8853_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_998_)
);

DFFSR _8433_ (
    .Q(\datapath_1.regfile_1.regOut[12] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_718_[27])
);

INVX1 _8013_ (
    .A(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_580_)
);

FILL FILL_4__13966_ (
);

FILL FILL_4__13546_ (
);

FILL FILL_2__14580_ (
);

FILL FILL_4__13126_ (
);

FILL SFILL103720x74050 (
);

FILL FILL_2__14160_ (
);

FILL FILL_2__7706_ (
);

FILL FILL_3__12959_ (
);

FILL FILL_1__13993_ (
);

FILL FILL_3__12119_ (
);

FILL FILL_1__13573_ (
);

FILL FILL_1__13153_ (
);

FILL FILL_0__12986_ (
);

NAND2X1 _12851_ (
    .A(vdd),
    .B(\datapath_1.rd1 [9]),
    .Y(_3573_)
);

NAND2X1 _12431_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [29]),
    .Y(_3353_)
);

FILL FILL_0__12146_ (
);

NAND3X1 _12011_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[6]),
    .C(_3032__bF$buf4),
    .Y(_3054_)
);

FILL FILL_3__13900_ (
);

FILL FILL_6__16345_ (
);

FILL FILL_5__8183_ (
);

FILL FILL_5__15758_ (
);

FILL FILL_5__15338_ (
);

FILL FILL_3__16372_ (
);

INVX1 _9638_ (
    .A(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_1399_)
);

FILL FILL_5_BUFX2_insert225 (
);

INVX1 _9218_ (
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_1180_)
);

FILL FILL_5__10893_ (
);

FILL FILL_5_BUFX2_insert226 (
);

FILL FILL_1__8595_ (
);

FILL FILL_5_BUFX2_insert227 (
);

FILL FILL_5_BUFX2_insert1010 (
);

FILL FILL_5__10053_ (
);

FILL FILL_5_BUFX2_insert228 (
);

FILL FILL_5_BUFX2_insert1011 (
);

FILL FILL_5_BUFX2_insert229 (
);

FILL FILL_5_BUFX2_insert1012 (
);

FILL FILL_2__15785_ (
);

FILL FILL_2__15365_ (
);

FILL FILL_5_BUFX2_insert1013 (
);

FILL FILL_5_BUFX2_insert1014 (
);

FILL FILL_5_BUFX2_insert1015 (
);

FILL FILL_5_BUFX2_insert1016 (
);

FILL SFILL94360x51050 (
);

FILL FILL_5_BUFX2_insert1017 (
);

FILL FILL_5_BUFX2_insert1018 (
);

FILL FILL_1__14778_ (
);

FILL FILL_5_BUFX2_insert1019 (
);

FILL FILL_1__14358_ (
);

FILL FILL_5__6916_ (
);

FILL FILL_3__9882_ (
);

FILL FILL_3__9462_ (
);

NOR2X1 _13636_ (
    .A(_4131_),
    .B(_4144_),
    .Y(_4145_)
);

FILL FILL_3__9042_ (
);

NAND2X1 _13216_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_3759_)
);

FILL FILL_5__9388_ (
);

FILL SFILL79160x31050 (
);

FILL FILL_1__6908_ (
);

FILL FILL_0__14712_ (
);

FILL FILL_5__11678_ (
);

FILL FILL_5__11258_ (
);

FILL FILL_3__12292_ (
);

FILL FILL_2__11285_ (
);

FILL FILL_1__10698_ (
);

FILL FILL_2_BUFX2_insert350 (
);

FILL FILL_1__10278_ (
);

FILL FILL_2_BUFX2_insert351 (
);

FILL FILL_2_BUFX2_insert352 (
);

FILL FILL_2_BUFX2_insert353 (
);

FILL FILL_2_BUFX2_insert354 (
);

FILL FILL_4__11612_ (
);

FILL FILL_2_BUFX2_insert355 (
);

FILL FILL_2_BUFX2_insert356 (
);

FILL FILL_5__15091_ (
);

FILL FILL_2_BUFX2_insert357 (
);

FILL FILL_6__8252_ (
);

FILL FILL_2_BUFX2_insert358 (
);

INVX1 _9391_ (
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_1275_)
);

FILL FILL_2_BUFX2_insert359 (
);

FILL FILL_4__14084_ (
);

FILL FILL_0__15917_ (
);

FILL FILL_0__10632_ (
);

FILL FILL_2__8244_ (
);

FILL FILL_3__13497_ (
);

FILL FILL_6__14411_ (
);

FILL FILL_5__13824_ (
);

FILL FILL_5__13404_ (
);

FILL FILL_2_BUFX2_insert1070 (
);

FILL FILL_2_BUFX2_insert1071 (
);

FILL FILL_2_BUFX2_insert1072 (
);

NAND2X1 _7704_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_415_)
);

FILL FILL_2_BUFX2_insert1073 (
);

FILL FILL_4__9531_ (
);

FILL FILL_4__9111_ (
);

FILL FILL_2__13851_ (
);

FILL SFILL110200x67050 (
);

FILL FILL_2__13431_ (
);

FILL FILL_5__16296_ (
);

FILL FILL_2__13011_ (
);

FILL FILL_1__12844_ (
);

FILL FILL_1__12424_ (
);

FILL FILL_4__15289_ (
);

FILL FILL_1__12004_ (
);

FILL FILL_2__9869_ (
);

FILL FILL_0__9851_ (
);

FILL FILL_0__11837_ (
);

FILL SFILL114520x75050 (
);

FILL FILL_2__9029_ (
);

FILL FILL_0__11417_ (
);

FILL FILL_0__9011_ (
);

AOI21X1 _11702_ (
    .A(_2502_),
    .B(_2496_),
    .C(_2504_),
    .Y(_2801_)
);

FILL FILL_5__7874_ (
);

FILL FILL_5__7454_ (
);

FILL FILL_4__16230_ (
);

FILL FILL_5__7034_ (
);

NOR2X1 _14594_ (
    .A(_5082_),
    .B(_5079_),
    .Y(_5083_)
);

OAI22X1 _14174_ (
    .A(_3893__bF$buf2),
    .B(_4670_),
    .C(_3930__bF$buf3),
    .D(_4669_),
    .Y(_4671_)
);

FILL SFILL95000x1050 (
);

FILL FILL_5__14609_ (
);

FILL FILL_3__15643_ (
);

INVX1 _8909_ (
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_1035_)
);

FILL FILL_3__15223_ (
);

FILL FILL_1__7866_ (
);

FILL FILL_1__7446_ (
);

FILL SFILL69080x36050 (
);

FILL FILL_2__14636_ (
);

FILL FILL_0__15670_ (
);

FILL FILL_2__14216_ (
);

FILL FILL_0__15250_ (
);

FILL FILL_1__13629_ (
);

FILL FILL_1__13209_ (
);

FILL FILL_1_BUFX2_insert370 (
);

FILL FILL_1_BUFX2_insert371 (
);

FILL FILL_3__8733_ (
);

FILL FILL_1_BUFX2_insert372 (
);

INVX1 _12907_ (
    .A(\datapath_1.a [28]),
    .Y(_3610_)
);

FILL FILL_3__8313_ (
);

FILL FILL_1_BUFX2_insert373 (
);

FILL FILL_1_BUFX2_insert374 (
);

FILL FILL_1_BUFX2_insert375 (
);

FILL FILL_1_BUFX2_insert376 (
);

FILL FILL_5__8659_ (
);

FILL FILL_1_BUFX2_insert377 (
);

FILL FILL_5__8239_ (
);

FILL SFILL114520x30050 (
);

FILL FILL_1_BUFX2_insert378 (
);

FILL FILL_1_BUFX2_insert379 (
);

NOR2X1 _15799_ (
    .A(_6257_),
    .B(_6260_),
    .Y(_6261_)
);

FILL FILL_4__12990_ (
);

FILL FILL_4__12570_ (
);

NOR3X1 _15379_ (
    .A(_5847_),
    .B(_5850_),
    .C(_5848_),
    .Y(_5851_)
);

FILL FILL_4__12150_ (
);

FILL FILL_3__16008_ (
);

FILL FILL_5__10949_ (
);

DFFSR _10094_ (
    .Q(\datapath_1.regfile_1.regOut[25] [24]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1563_[24])
);

FILL FILL_3__11983_ (
);

FILL FILL_5__10529_ (
);

FILL FILL_5__9600_ (
);

FILL FILL_3__11563_ (
);

FILL FILL_5__10109_ (
);

FILL FILL_3__11143_ (
);

FILL FILL_0__16035_ (
);

AOI21X1 _16320_ (
    .A(_6745_),
    .B(_6768_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [31])
);

FILL FILL_2__10976_ (
);

FILL FILL_2__10556_ (
);

FILL FILL_2__10136_ (
);

FILL FILL_0__11590_ (
);

FILL FILL_0__11170_ (
);

FILL FILL_3__9938_ (
);

FILL FILL_3__9518_ (
);

FILL SFILL43080x80050 (
);

FILL SFILL3640x56050 (
);

FILL FILL_5__14782_ (
);

FILL FILL_0__6976_ (
);

FILL FILL_5__14362_ (
);

DFFSR _8662_ (
    .Q(\datapath_1.regfile_1.regOut[14] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_848_[0])
);

FILL SFILL22920x65050 (
);

INVX1 _8242_ (
    .A(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_692_)
);

FILL SFILL104520x73050 (
);

FILL SFILL43880x63050 (
);

FILL FILL_1__10910_ (
);

FILL FILL_4__13775_ (
);

FILL FILL_4__13355_ (
);

INVX1 _11299_ (
    .A(_2252_),
    .Y(_2418_)
);

FILL FILL_2__7935_ (
);

FILL FILL_3__12768_ (
);

FILL FILL_3__12348_ (
);

FILL SFILL59000x77050 (
);

FILL FILL_1__13382_ (
);

INVX1 _12660_ (
    .A(\datapath_1.Data [31]),
    .Y(_3486_)
);

FILL FILL_0__12375_ (
);

NAND3X1 _12240_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [8]),
    .C(_3198__bF$buf2),
    .Y(_3219_)
);

FILL SFILL38920x19050 (
);

FILL FILL_5__15987_ (
);

FILL FILL_2__12702_ (
);

FILL FILL_5__15567_ (
);

FILL FILL_5__15147_ (
);

INVX1 _9867_ (
    .A(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_1511_)
);

FILL FILL_3__16181_ (
);

FILL FILL_6__8728_ (
);

DFFSR _9447_ (
    .Q(\datapath_1.regfile_1.regOut[20] [17]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_1238_[17])
);

OAI21X1 _9027_ (
    .A(_1092_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1093_),
    .Y(_1043_[25])
);

FILL SFILL3640x11050 (
);

FILL FILL_5__10282_ (
);

FILL FILL_2__15594_ (
);

FILL FILL_2__15174_ (
);

FILL FILL_0__8702_ (
);

FILL FILL_1__14587_ (
);

FILL FILL_1__14167_ (
);

FILL FILL_4__15921_ (
);

FILL FILL_4__15501_ (
);

FILL SFILL59000x32050 (
);

AOI22X1 _13865_ (
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .B(_4090_),
    .C(_3948_),
    .D(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_4369_)
);

FILL FILL_3__9271_ (
);

INVX1 _13445_ (
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_3957_)
);

OAI21X1 _13025_ (
    .A(_3667_),
    .B(vdd),
    .C(_3668_),
    .Y(_3620_[24])
);

FILL FILL_3__14914_ (
);

FILL SFILL3560x18050 (
);

FILL SFILL104440x35050 (
);

FILL FILL_2__13907_ (
);

FILL FILL_0__14941_ (
);

FILL FILL_0__14521_ (
);

FILL FILL_0__14101_ (
);

FILL FILL_5__11487_ (
);

FILL FILL_5__11067_ (
);

FILL FILL_2__16379_ (
);

FILL FILL_4__7194_ (
);

FILL SFILL33880x61050 (
);

FILL FILL_0__9907_ (
);

FILL FILL_2__11094_ (
);

FILL SFILL64600x8050 (
);

FILL SFILL49000x75050 (
);

FILL FILL_4__11841_ (
);

FILL FILL_4__11421_ (
);

FILL FILL_4__11001_ (
);

FILL FILL_0__7094_ (
);

FILL FILL_1__16313_ (
);

FILL FILL_6__8061_ (
);

FILL FILL_3__10834_ (
);

FILL FILL_3__10414_ (
);

FILL FILL_0__15726_ (
);

FILL FILL_0__15306_ (
);

FILL FILL_2__8893_ (
);

FILL FILL_2__8473_ (
);

FILL FILL_0__10441_ (
);

FILL FILL_0__10021_ (
);

FILL FILL_4__8399_ (
);

FILL FILL_2__12299_ (
);

FILL FILL_5__13633_ (
);

FILL FILL_5__13213_ (
);

NAND2X1 _7933_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_527_)
);

DFFSR _7513_ (
    .Q(\datapath_1.regfile_1.regOut[5] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_263_[3])
);

FILL FILL_1__6890_ (
);

FILL FILL_4__9760_ (
);

FILL SFILL94840x53050 (
);

FILL FILL_4__9340_ (
);

FILL FILL_4__12626_ (
);

FILL FILL_2__13660_ (
);

FILL FILL_4__12206_ (
);

FILL FILL_2__13240_ (
);

FILL SFILL49000x30050 (
);

FILL SFILL39080x75050 (
);

FILL FILL_3__11619_ (
);

FILL FILL_1__12653_ (
);

FILL FILL_4__15098_ (
);

FILL FILL_1__12233_ (
);

FILL FILL_0__9660_ (
);

FILL FILL_2__9678_ (
);

FILL FILL_0__9240_ (
);

OAI21X1 _11931_ (
    .A(_2994_),
    .B(IorD_bF$buf4),
    .C(_2995_),
    .Y(_1_[14])
);

FILL FILL_2__9258_ (
);

FILL FILL_0__11646_ (
);

FILL FILL_0__11226_ (
);

AOI21X1 _11511_ (
    .A(_2602_),
    .B(_2620_),
    .C(_2622_),
    .Y(_2623_)
);

FILL FILL_5__7683_ (
);

FILL FILL_6__10140_ (
);

FILL FILL_5__14838_ (
);

FILL FILL_5__14418_ (
);

FILL FILL_3__15872_ (
);

FILL FILL_3__15452_ (
);

INVX1 _8718_ (
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_928_)
);

FILL FILL_3__15032_ (
);

FILL FILL_1__7675_ (
);

FILL FILL_2__14865_ (
);

FILL FILL111800x75050 (
);

FILL FILL_2__14445_ (
);

FILL FILL_2__14025_ (
);

FILL SFILL63960x55050 (
);

FILL SFILL39000x73050 (
);

FILL SFILL94360x46050 (
);

FILL FILL_1__13858_ (
);

FILL FILL_1__13438_ (
);

FILL FILL_1__13018_ (
);

FILL FILL_3__8962_ (
);

INVX1 _12716_ (
    .A(\datapath_1.PCJump [9]),
    .Y(_3503_)
);

FILL FILL_3__8122_ (
);

FILL FILL_5__8888_ (
);

FILL SFILL79160x26050 (
);

FILL FILL_5__8468_ (
);

FILL FILL_1_BUFX2_insert40 (
);

FILL FILL_1_BUFX2_insert41 (
);

FILL FILL_1_BUFX2_insert42 (
);

FILL FILL_1_BUFX2_insert43 (
);

OAI22X1 _15188_ (
    .A(_4137_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf4),
    .D(_4138_),
    .Y(_5665_)
);

FILL FILL_1_BUFX2_insert44 (
);

FILL FILL_1_BUFX2_insert45 (
);

FILL FILL_1_BUFX2_insert46 (
);

FILL FILL_3__16237_ (
);

FILL FILL_1_BUFX2_insert47 (
);

FILL FILL_1_BUFX2_insert48 (
);

FILL FILL_1_BUFX2_insert49 (
);

FILL FILL_5__10758_ (
);

FILL FILL_3__11792_ (
);

FILL FILL_3__11372_ (
);

FILL FILL_4__6885_ (
);

FILL FILL_0__16264_ (
);

FILL FILL_2__10785_ (
);

FILL FILL_2__10365_ (
);

FILL FILL_1__9401_ (
);

FILL FILL_3__9747_ (
);

FILL FILL_5__14591_ (
);

FILL FILL_5__14171_ (
);

INVX1 _8891_ (
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_1023_)
);

FILL FILL112280x1050 (
);

FILL FILL_6__7332_ (
);

INVX1 _8471_ (
    .A(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_804_)
);

DFFSR _8051_ (
    .Q(\datapath_1.regfile_1.regOut[9] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_523_[29])
);

FILL FILL_4__13584_ (
);

FILL FILL_4__13164_ (
);

FILL SFILL8760x63050 (
);

FILL FILL_2__7744_ (
);

FILL FILL_3__12997_ (
);

FILL FILL_3__12577_ (
);

FILL FILL_2__7324_ (
);

FILL FILL_3__12157_ (
);

FILL FILL_0__12184_ (
);

FILL SFILL114600x63050 (
);

FILL FILL_5__12904_ (
);

FILL SFILL84360x44050 (
);

FILL FILL_4__8611_ (
);

FILL FILL_5_BUFX2_insert600 (
);

FILL FILL_5__15796_ (
);

FILL FILL_5_BUFX2_insert601 (
);

FILL FILL_5__15376_ (
);

FILL FILL_2__12511_ (
);

FILL FILL_5_BUFX2_insert602 (
);

FILL FILL_5_BUFX2_insert603 (
);

FILL FILL_5_BUFX2_insert604 (
);

OAI21X1 _9676_ (
    .A(_1423_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1424_),
    .Y(_1368_[28])
);

FILL FILL_5_BUFX2_insert605 (
);

OAI21X1 _9256_ (
    .A(_1204_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1205_),
    .Y(_1173_[16])
);

FILL FILL_5_BUFX2_insert606 (
);

FILL FILL_5_BUFX2_insert607 (
);

FILL FILL_5_BUFX2_insert608 (
);

FILL FILL_1__11924_ (
);

FILL FILL_4__14789_ (
);

FILL FILL_4__14369_ (
);

FILL FILL_5_BUFX2_insert609 (
);

FILL FILL_1__11504_ (
);

FILL FILL_0__10917_ (
);

FILL FILL_0__8511_ (
);

FILL FILL_2__8529_ (
);

FILL FILL_2__8109_ (
);

FILL FILL_1__14396_ (
);

FILL FILL_5__6954_ (
);

FILL FILL_4__15730_ (
);

FILL FILL_4__15310_ (
);

NAND3X1 _13674_ (
    .A(_4173_),
    .B(_4174_),
    .C(_4181_),
    .Y(_4182_)
);

FILL FILL_0__13389_ (
);

FILL FILL_3__9080_ (
);

INVX4 _13254_ (
    .A(RegWrite_bF$buf0),
    .Y(_3797_)
);

FILL FILL_3__14723_ (
);

FILL FILL_3__14303_ (
);

FILL FILL_1__6946_ (
);

FILL FILL_2__13716_ (
);

FILL FILL_0__14750_ (
);

FILL FILL_0__14330_ (
);

FILL FILL_5__11296_ (
);

FILL FILL_1__12709_ (
);

FILL FILL_2__16188_ (
);

FILL FILL_4__10289_ (
);

FILL FILL_3__7813_ (
);

FILL FILL_5__7739_ (
);

FILL SFILL114520x25050 (
);

FILL FILL_5__7319_ (
);

FILL FILL_2_BUFX2_insert730 (
);

FILL FILL_2_BUFX2_insert731 (
);

FILL FILL_2_BUFX2_insert732 (
);

NAND3X1 _14879_ (
    .A(_5360_),
    .B(_5361_),
    .C(_5359_),
    .Y(_5362_)
);

FILL FILL_6__10616_ (
);

FILL FILL_2_BUFX2_insert733 (
);

AOI22X1 _14459_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [21]),
    .C(\datapath_1.regfile_1.regOut[7] [21]),
    .D(_3948_),
    .Y(_4950_)
);

FILL FILL_2_BUFX2_insert734 (
);

FILL FILL_4__11650_ (
);

INVX1 _14039_ (
    .A(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_4539_)
);

FILL FILL_2_BUFX2_insert735 (
);

FILL FILL_4__11230_ (
);

FILL FILL_3__15928_ (
);

FILL FILL_2_BUFX2_insert736 (
);

FILL FILL_3__15508_ (
);

FILL FILL_2_BUFX2_insert737 (
);

FILL FILL_2_BUFX2_insert738 (
);

FILL FILL_1__16122_ (
);

FILL FILL_2_BUFX2_insert739 (
);

FILL FILL_3__10643_ (
);

FILL SFILL43960x51050 (
);

FILL FILL_0__15955_ (
);

FILL FILL_0__15535_ (
);

OAI22X1 _15820_ (
    .A(_4877_),
    .B(_5539__bF$buf1),
    .C(_5552__bF$buf0),
    .D(_4853_),
    .Y(_6281_)
);

INVX1 _15400_ (
    .A(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_5872_)
);

FILL FILL_0__15115_ (
);

FILL FILL_0__10670_ (
);

FILL FILL_0__10250_ (
);

FILL FILL_5__13862_ (
);

FILL FILL_5__13442_ (
);

FILL FILL_5__13022_ (
);

INVX1 _7742_ (
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_440_)
);

INVX1 _7322_ (
    .A(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_221_)
);

FILL SFILL43880x58050 (
);

FILL FILL_4__12855_ (
);

FILL FILL_4__12435_ (
);

FILL FILL_4__12015_ (
);

INVX1 _10799_ (
    .A(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_1990_)
);

INVX1 _10379_ (
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .Y(_1771_)
);

FILL FILL_3__11848_ (
);

FILL FILL_1__12882_ (
);

FILL FILL_3__11428_ (
);

FILL FILL_1__12462_ (
);

FILL FILL_3__11008_ (
);

FILL FILL_1__12042_ (
);

FILL SFILL59080x29050 (
);

FILL FILL112280x62050 (
);

FILL FILL_2__9487_ (
);

FILL FILL_0__11875_ (
);

AOI21X1 _11740_ (
    .A(_2836_),
    .B(_2834_),
    .C(_2832_),
    .Y(_2837_)
);

FILL FILL_0__11455_ (
);

FILL FILL_0__11035_ (
);

INVX2 _11320_ (
    .A(_2438_),
    .Y(_2439_)
);

FILL FILL_6__15654_ (
);

FILL FILL_6__15234_ (
);

FILL FILL_5__7492_ (
);

FILL FILL_5__7072_ (
);

FILL FILL_5__14647_ (
);

FILL FILL_3__15681_ (
);

FILL FILL_5__14227_ (
);

DFFSR _8947_ (
    .Q(\datapath_1.regfile_1.regOut[16] [29]),
    .CLK(clk_bF$buf21),
    .R(rst_bF$buf106),
    .S(vdd),
    .D(_978_[29])
);

FILL FILL_6__7808_ (
);

FILL FILL_3__15261_ (
);

OAI21X1 _8527_ (
    .A(_840_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_841_),
    .Y(_783_[29])
);

OAI21X1 _8107_ (
    .A(_621_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_622_),
    .Y(_588_[17])
);

FILL FILL_1__7484_ (
);

FILL FILL_1__7064_ (
);

FILL FILL_2__14674_ (
);

FILL FILL_2__14254_ (
);

FILL SFILL43880x13050 (
);

FILL FILL_1__13667_ (
);

FILL FILL_1__13247_ (
);

FILL SFILL59000x27050 (
);

FILL FILL_1_BUFX2_insert750 (
);

FILL FILL_1_BUFX2_insert751 (
);

FILL FILL_3__8771_ (
);

FILL FILL_1_BUFX2_insert752 (
);

DFFSR _12945_ (
    .Q(\datapath_1.a [26]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3555_[26])
);

FILL FILL_3__8351_ (
);

OAI21X1 _12525_ (
    .A(_3415_),
    .B(vdd),
    .C(_3416_),
    .Y(_3360_[28])
);

FILL FILL_1_BUFX2_insert753 (
);

AOI22X1 _12105_ (
    .A(\datapath_1.ALUResult [29]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3125_)
);

FILL FILL_1_BUFX2_insert754 (
);

FILL FILL_1_BUFX2_insert755 (
);

FILL FILL_1_BUFX2_insert756 (
);

FILL FILL_5__8697_ (
);

FILL FILL_1_BUFX2_insert757 (
);

FILL FILL_5__8277_ (
);

FILL FILL_1_BUFX2_insert758 (
);

FILL FILL_1_BUFX2_insert759 (
);

FILL FILL_6__11574_ (
);

FILL FILL_6__11154_ (
);

FILL FILL_0__13601_ (
);

FILL FILL_3__16046_ (
);

FILL FILL_5__10567_ (
);

FILL FILL_1__8269_ (
);

FILL FILL_5__10147_ (
);

FILL FILL_3__11181_ (
);

FILL FILL_2__15879_ (
);

FILL FILL_2__15459_ (
);

FILL FILL_2__15039_ (
);

FILL SFILL33880x56050 (
);

FILL FILL_0__16073_ (
);

FILL FILL_2__10174_ (
);

FILL FILL_1__9630_ (
);

FILL FILL_1__9210_ (
);

FILL SFILL18600x79050 (
);

FILL FILL_3__9976_ (
);

FILL FILL_2__16400_ (
);

FILL FILL_3__9556_ (
);

FILL FILL_4__10921_ (
);

FILL FILL_3__9136_ (
);

FILL FILL_4__10501_ (
);

FILL FILL_1__15813_ (
);

DFFSR _8280_ (
    .Q(\datapath_1.regfile_1.regOut[11] [2]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_653_[2])
);

FILL FILL_6__12779_ (
);

FILL SFILL94440x79050 (
);

FILL FILL_4__13393_ (
);

FILL FILL_0__14806_ (
);

FILL FILL_2__7973_ (
);

FILL FILL_2__7553_ (
);

BUFX2 BUFX2_insert420 (
    .A(_5471_),
    .Y(_5471__bF$buf4)
);

FILL FILL_3__12386_ (
);

BUFX2 BUFX2_insert421 (
    .A(_5471_),
    .Y(_5471__bF$buf3)
);

BUFX2 BUFX2_insert422 (
    .A(_5471_),
    .Y(_5471__bF$buf2)
);

BUFX2 BUFX2_insert423 (
    .A(_5471_),
    .Y(_5471__bF$buf1)
);

BUFX2 BUFX2_insert424 (
    .A(_5471_),
    .Y(_5471__bF$buf0)
);

FILL FILL_6__13720_ (
);

FILL FILL_4__7479_ (
);

BUFX2 BUFX2_insert425 (
    .A(_5527_),
    .Y(_5527__bF$buf4)
);

BUFX2 BUFX2_insert426 (
    .A(_5527_),
    .Y(_5527__bF$buf3)
);

FILL FILL_4__7059_ (
);

BUFX2 BUFX2_insert427 (
    .A(_5527_),
    .Y(_5527__bF$buf2)
);

FILL FILL_2__11799_ (
);

BUFX2 BUFX2_insert428 (
    .A(_5527_),
    .Y(_5527__bF$buf1)
);

FILL FILL_2__11379_ (
);

BUFX2 BUFX2_insert429 (
    .A(_5527_),
    .Y(_5527__bF$buf0)
);

FILL SFILL33880x11050 (
);

FILL FILL_5__12713_ (
);

FILL FILL_4__8840_ (
);

FILL FILL_4__8000_ (
);

FILL FILL_4__11706_ (
);

FILL FILL_2__12740_ (
);

FILL FILL_5__15185_ (
);

FILL FILL_0__7799_ (
);

FILL FILL_2__12320_ (
);

FILL SFILL49000x25050 (
);

FILL FILL_0__7379_ (
);

OAI21X1 _9485_ (
    .A(_1316_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .C(_1317_),
    .Y(_1303_[7])
);

DFFSR _9065_ (
    .Q(\datapath_1.regfile_1.regOut[17] [19]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_1043_[19])
);

FILL FILL_4__14598_ (
);

FILL FILL_1__11733_ (
);

FILL FILL_4__14178_ (
);

FILL FILL_1__11313_ (
);

FILL FILL_0__8740_ (
);

FILL FILL_2__8758_ (
);

FILL FILL_0__8320_ (
);

FILL FILL_2__8338_ (
);

FILL FILL_0__10306_ (
);

NOR2X1 _13483_ (
    .A(_3993_),
    .B(_3990_),
    .Y(_3994_)
);

DFFSR _13063_ (
    .Q(_2_[16]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3620_[16])
);

FILL FILL_5__13918_ (
);

FILL FILL_3__14952_ (
);

FILL FILL_3__14532_ (
);

FILL FILL_3__14112_ (
);

FILL FILL_4_BUFX2_insert260 (
);

FILL FILL_4__9625_ (
);

FILL FILL_4_BUFX2_insert261 (
);

FILL FILL_4_BUFX2_insert262 (
);

FILL FILL_4_BUFX2_insert263 (
);

FILL FILL_2__13945_ (
);

FILL FILL_4_BUFX2_insert264 (
);

FILL FILL_2__13525_ (
);

FILL FILL_2__13105_ (
);

FILL FILL_4_BUFX2_insert265 (
);

FILL SFILL39000x68050 (
);

FILL FILL_4_BUFX2_insert266 (
);

FILL FILL_4_BUFX2_insert267 (
);

FILL FILL_4_BUFX2_insert268 (
);

FILL FILL_4_BUFX2_insert269 (
);

FILL FILL_1__12518_ (
);

FILL FILL_0__9525_ (
);

FILL FILL_3__7622_ (
);

FILL FILL_3__7202_ (
);

FILL FILL_0__9105_ (
);

FILL FILL_5__7968_ (
);

FILL FILL_5__7548_ (
);

FILL FILL_4__16324_ (
);

AOI22X1 _14688_ (
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .B(_3995__bF$buf2),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_5175_)
);

OAI22X1 _14268_ (
    .A(_4761_),
    .B(_3910_),
    .C(_3935__bF$buf2),
    .D(_4762_),
    .Y(_4763_)
);

FILL FILL_6__10005_ (
);

FILL SFILL23800x52050 (
);

FILL FILL_3__15737_ (
);

FILL FILL_3__15317_ (
);

FILL FILL_1__16351_ (
);

FILL SFILL79320x1050 (
);

FILL FILL_3__10872_ (
);

FILL FILL_3__10452_ (
);

FILL FILL_3__10032_ (
);

FILL FILL_0__15764_ (
);

FILL FILL_0__15344_ (
);

FILL SFILL53960x2050 (
);

FILL FILL_2__8091_ (
);

FILL FILL_1__8901_ (
);

FILL FILL_3__8827_ (
);

FILL FILL_5__13671_ (
);

FILL FILL_5__13251_ (
);

INVX1 _7971_ (
    .A(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_552_)
);

FILL SFILL84440x32050 (
);

INVX1 _7551_ (
    .A(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_333_)
);

DFFSR _7131_ (
    .Q(\datapath_1.regfile_1.regOut[2] [5]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_68_[5])
);

FILL SFILL8760x58050 (
);

FILL FILL_4__12244_ (
);

OAI21X1 _10188_ (
    .A(_1683_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .C(_1684_),
    .Y(_1628_[28])
);

FILL FILL_3__11657_ (
);

FILL FILL_3__11237_ (
);

FILL FILL_1__12271_ (
);

INVX1 _16414_ (
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_6830_)
);

FILL FILL_0__16129_ (
);

FILL FILL_0__11684_ (
);

FILL FILL_2__9296_ (
);

FILL FILL_0__11264_ (
);

FILL SFILL53960x48050 (
);

FILL SFILL84360x39050 (
);

FILL FILL_3_BUFX2_insert280 (
);

FILL FILL_3_BUFX2_insert281 (
);

FILL FILL_5__14876_ (
);

FILL FILL_3_BUFX2_insert282 (
);

FILL FILL_5__14456_ (
);

FILL FILL_3_BUFX2_insert283 (
);

FILL FILL_5__14036_ (
);

FILL FILL_3_BUFX2_insert284 (
);

FILL FILL_3__15490_ (
);

FILL FILL_3__15070_ (
);

FILL FILL_3_BUFX2_insert285 (
);

OAI21X1 _8756_ (
    .A(_952_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .C(_953_),
    .Y(_913_[20])
);

OAI21X1 _8336_ (
    .A(_733_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .C(_734_),
    .Y(_718_[8])
);

FILL FILL_3_BUFX2_insert286 (
);

FILL FILL_3_BUFX2_insert287 (
);

FILL FILL_3_BUFX2_insert288 (
);

FILL FILL_1__7293_ (
);

FILL FILL_4__13869_ (
);

FILL FILL_3_BUFX2_insert289 (
);

FILL FILL_4__13449_ (
);

FILL FILL_2__14483_ (
);

FILL FILL_4__13029_ (
);

FILL FILL_2__14063_ (
);

FILL SFILL8760x13050 (
);

FILL FILL_2__7609_ (
);

FILL SFILL13800x50050 (
);

FILL FILL_1__13896_ (
);

FILL FILL_1__13476_ (
);

FILL FILL_4__14810_ (
);

FILL FILL_3__8580_ (
);

FILL FILL_0__12889_ (
);

OAI21X1 _12754_ (
    .A(_3527_),
    .B(IRWrite_bF$buf0),
    .C(_3528_),
    .Y(_3490_[19])
);

FILL FILL_0__12469_ (
);

FILL FILL_0__12049_ (
);

NAND3X1 _12334_ (
    .A(_3287_),
    .B(_3288_),
    .C(_3289_),
    .Y(\datapath_1.alu_1.ALUInB [29])
);

FILL FILL_3__13803_ (
);

FILL FILL_5__8086_ (
);

FILL SFILL114600x13050 (
);

FILL FILL_0__13830_ (
);

FILL FILL_0__13410_ (
);

FILL FILL_3__16275_ (
);

FILL FILL_5__10796_ (
);

FILL FILL_5__10376_ (
);

FILL FILL_1__8498_ (
);

FILL FILL_1__8078_ (
);

FILL FILL_2__15688_ (
);

FILL FILL_2__15268_ (
);

FILL FILL_3__9785_ (
);

OAI22X1 _13959_ (
    .A(_4459_),
    .B(_3936__bF$buf1),
    .C(_3935__bF$buf0),
    .D(_4460_),
    .Y(_4461_)
);

FILL FILL_3__9365_ (
);

OAI22X1 _13539_ (
    .A(_3967__bF$buf1),
    .B(_4047_),
    .C(_4048_),
    .D(_3902__bF$buf2),
    .Y(_4049_)
);

FILL SFILL3720x39050 (
);

FILL FILL_4__10310_ (
);

NAND2X1 _13119_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [13]),
    .Y(_3711_)
);

FILL FILL_1__15622_ (
);

FILL FILL_1__15202_ (
);

FILL FILL_6__12588_ (
);

FILL FILL_0__14615_ (
);

NAND2X1 _14900_ (
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .B(_4102_),
    .Y(_5382_)
);

FILL FILL_2__7362_ (
);

FILL FILL_3__12195_ (
);

FILL FILL_4__7288_ (
);

FILL FILL112360x50050 (
);

FILL FILL_2__11188_ (
);

FILL FILL_5__12522_ (
);

FILL FILL_5__12102_ (
);

FILL FILL_4__11935_ (
);

FILL FILL_4__11515_ (
);

FILL SFILL23880x6050 (
);

FILL FILL_2_BUFX2_insert90 (
);

FILL FILL_0__7188_ (
);

NAND2X1 _9294_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1231_)
);

FILL FILL_2_BUFX2_insert91 (
);

FILL FILL_1__16407_ (
);

FILL FILL_2_BUFX2_insert92 (
);

FILL FILL_3__10928_ (
);

FILL FILL_2_BUFX2_insert93 (
);

FILL FILL_3__10508_ (
);

FILL FILL_1__11962_ (
);

FILL FILL_2_BUFX2_insert94 (
);

FILL FILL_2_BUFX2_insert95 (
);

FILL FILL_1__11542_ (
);

FILL FILL_2_BUFX2_insert96 (
);

FILL FILL_1__11122_ (
);

FILL FILL_2_BUFX2_insert97 (
);

FILL FILL_2_BUFX2_insert98 (
);

FILL FILL112280x57050 (
);

FILL FILL_2_BUFX2_insert99 (
);

FILL FILL_2__8987_ (
);

FILL FILL_2__8567_ (
);

FILL FILL_0__10955_ (
);

FILL FILL_0__10535_ (
);

FILL FILL_2__8147_ (
);

INVX1 _10820_ (
    .A(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_2004_)
);

FILL FILL_0__10115_ (
);

INVX1 _10400_ (
    .A(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_1785_)
);

FILL FILL_5__6992_ (
);

FILL FILL_6__14314_ (
);

OR2X2 _13292_ (
    .A(_3796_),
    .B(_3829_),
    .Y(_3830_)
);

FILL FILL_5__13727_ (
);

FILL FILL_5__13307_ (
);

FILL FILL_3__14761_ (
);

FILL FILL_3__14341_ (
);

OAI21X1 _7607_ (
    .A(_369_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_370_),
    .Y(_328_[21])
);

FILL FILL_1__6984_ (
);

FILL FILL_4__9854_ (
);

FILL FILL_4__9014_ (
);

FILL SFILL104520x18050 (
);

FILL FILL_2__13754_ (
);

FILL FILL_2__13334_ (
);

FILL FILL_5__16199_ (
);

FILL FILL_1__12747_ (
);

FILL FILL_1__12327_ (
);

FILL FILL_0__9754_ (
);

FILL FILL_3__7851_ (
);

FILL SFILL108840x26050 (
);

FILL FILL_0__9334_ (
);

FILL FILL_3__7431_ (
);

NAND2X1 _11605_ (
    .A(_2239_),
    .B(_2341__bF$buf1),
    .Y(_2711_)
);

FILL FILL112280x12050 (
);

FILL FILL_5__7357_ (
);

FILL FILL_4__16133_ (
);

NOR2X1 _14497_ (
    .A(_4987_),
    .B(_4984_),
    .Y(_4988_)
);

AOI22X1 _14077_ (
    .A(_3998__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[2] [13]),
    .C(\datapath_1.regfile_1.regOut[27] [13]),
    .D(_4129_),
    .Y(_4576_)
);

FILL FILL_3__15966_ (
);

FILL FILL_3__15546_ (
);

FILL FILL_3__15126_ (
);

FILL FILL_1__16160_ (
);

FILL FILL_1__7349_ (
);

FILL FILL_3__10681_ (
);

FILL FILL_3__10261_ (
);

FILL FILL_2__14959_ (
);

FILL SFILL94520x67050 (
);

FILL FILL_0__15993_ (
);

FILL FILL_2__14539_ (
);

FILL FILL_0__15573_ (
);

FILL FILL_2__14119_ (
);

FILL FILL_0__15153_ (
);

FILL FILL_1__8710_ (
);

FILL FILL_2__15900_ (
);

FILL FILL_3__8636_ (
);

FILL FILL_3__8216_ (
);

FILL FILL_5__13480_ (
);

DFFSR _7780_ (
    .Q(\datapath_1.regfile_1.regOut[7] [14]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_393_[14])
);

OAI21X1 _7360_ (
    .A(_245_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .C(_246_),
    .Y(_198_[24])
);

FILL FILL_4__12893_ (
);

FILL FILL_4__12473_ (
);

FILL FILL_4__12053_ (
);

FILL SFILL33000x66050 (
);

FILL FILL_3__11886_ (
);

FILL FILL_5__9923_ (
);

FILL FILL_3__11466_ (
);

FILL FILL_5__9503_ (
);

FILL FILL_3__11046_ (
);

FILL FILL_1__12080_ (
);

FILL FILL_4__6979_ (
);

FILL FILL_0__16358_ (
);

OAI22X1 _16223_ (
    .A(_5534__bF$buf2),
    .B(_5343_),
    .C(_6673_),
    .D(_5549__bF$buf4),
    .Y(_6674_)
);

FILL FILL_2__10879_ (
);

FILL FILL_2__10039_ (
);

FILL FILL_0__11493_ (
);

FILL FILL_0__11073_ (
);

FILL FILL_1__9915_ (
);

FILL FILL_4__7500_ (
);

FILL FILL_2__11820_ (
);

FILL FILL_5__14685_ (
);

FILL FILL_5__14265_ (
);

FILL FILL_2__11400_ (
);

FILL FILL_0__6879_ (
);

OAI21X1 _8985_ (
    .A(_1064_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .C(_1065_),
    .Y(_1043_[11])
);

FILL FILL_6__7426_ (
);

DFFSR _8565_ (
    .Q(\datapath_1.regfile_1.regOut[13] [31]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_783_[31])
);

NAND2X1 _8145_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_648_)
);

FILL FILL_1__10813_ (
);

FILL FILL_4__13678_ (
);

FILL SFILL4200x62050 (
);

FILL FILL_4__13258_ (
);

FILL FILL_2__14292_ (
);

FILL SFILL94440x29050 (
);

FILL FILL_0__7820_ (
);

FILL FILL_2__7838_ (
);

FILL FILL_2__7418_ (
);

FILL FILL_1__13285_ (
);

FILL FILL_0__12698_ (
);

OAI21X1 _12983_ (
    .A(_3639_),
    .B(vdd),
    .C(_3640_),
    .Y(_3620_[10])
);

DFFSR _12563_ (
    .Q(ALUOut[28]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3360_[28])
);

FILL FILL_0__12278_ (
);

FILL SFILL23880x49050 (
);

NAND2X1 _12143_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.a [9]),
    .Y(_3149_)
);

FILL FILL_3__13612_ (
);

FILL FILL_4__8705_ (
);

FILL FILL_2__12605_ (
);

FILL FILL_3__16084_ (
);

FILL FILL_5__10185_ (
);

FILL FILL_2__15497_ (
);

FILL FILL_2__15077_ (
);

FILL FILL_5__16411_ (
);

FILL FILL_0__8605_ (
);

FILL FILL_4__15824_ (
);

FILL FILL_4__15404_ (
);

FILL FILL_3__9594_ (
);

OAI22X1 _13768_ (
    .A(_3941_),
    .B(_4273_),
    .C(_3930__bF$buf3),
    .D(_4272_),
    .Y(_4274_)
);

FILL SFILL23800x47050 (
);

OR2X2 _13348_ (
    .A(_3866_),
    .B(_3762_),
    .Y(_3867_)
);

FILL SFILL109480x2050 (
);

FILL FILL_3__14817_ (
);

FILL FILL_1__15851_ (
);

FILL FILL_1__15431_ (
);

FILL FILL_1__15011_ (
);

FILL FILL_6__12397_ (
);

FILL FILL_0__14844_ (
);

FILL FILL_0__14424_ (
);

FILL FILL_0__14004_ (
);

FILL FILL_2__7591_ (
);

BUFX2 BUFX2_insert800 (
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf0 )
);

FILL FILL_2__7171_ (
);

BUFX2 BUFX2_insert801 (
    .A(_5570_),
    .Y(_5570__bF$buf3)
);

FILL SFILL23400x33050 (
);

FILL SFILL39000x18050 (
);

BUFX2 BUFX2_insert802 (
    .A(_5570_),
    .Y(_5570__bF$buf2)
);

BUFX2 BUFX2_insert803 (
    .A(_5570_),
    .Y(_5570__bF$buf1)
);

BUFX2 BUFX2_insert804 (
    .A(_5570_),
    .Y(_5570__bF$buf0)
);

BUFX2 BUFX2_insert805 (
    .A(_4001_),
    .Y(_4001__bF$buf3)
);

FILL FILL_4__7097_ (
);

BUFX2 BUFX2_insert806 (
    .A(_4001_),
    .Y(_4001__bF$buf2)
);

BUFX2 BUFX2_insert807 (
    .A(_4001_),
    .Y(_4001__bF$buf1)
);

BUFX2 BUFX2_insert808 (
    .A(_4001_),
    .Y(_4001__bF$buf0)
);

BUFX2 BUFX2_insert809 (
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf7 )
);

FILL FILL_5__12751_ (
);

FILL FILL_5__12331_ (
);

FILL FILL_4__11744_ (
);

FILL FILL_4__11324_ (
);

FILL FILL_1__16216_ (
);

FILL FILL_3__10317_ (
);

FILL FILL_1__11771_ (
);

FILL FILL_1__11351_ (
);

INVX1 _15914_ (
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_6373_)
);

FILL FILL_0__15629_ (
);

FILL FILL_0__15209_ (
);

FILL FILL_0__10764_ (
);

FILL FILL_2__8376_ (
);

FILL FILL_6__14963_ (
);

FILL FILL_5__13956_ (
);

FILL FILL_3__14990_ (
);

FILL FILL_5__13536_ (
);

FILL FILL_3__14570_ (
);

FILL FILL_5__13116_ (
);

FILL FILL_3__14150_ (
);

OAI21X1 _7836_ (
    .A(_481_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .C(_482_),
    .Y(_458_[12])
);

OAI21X1 _7416_ (
    .A(_326_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_327_),
    .Y(_263_[0])
);

FILL FILL_4_BUFX2_insert640 (
);

FILL FILL_4__9663_ (
);

FILL FILL_4_BUFX2_insert641 (
);

FILL FILL_4__9243_ (
);

FILL FILL_4_BUFX2_insert642 (
);

FILL FILL_2__13983_ (
);

FILL FILL_4_BUFX2_insert643 (
);

FILL FILL_4__12529_ (
);

FILL FILL_4_BUFX2_insert644 (
);

FILL FILL_4__12109_ (
);

FILL FILL_2__13563_ (
);

FILL FILL_2__13143_ (
);

FILL FILL_4_BUFX2_insert645 (
);

FILL FILL_4_BUFX2_insert646 (
);

FILL FILL_4_BUFX2_insert647 (
);

FILL FILL_4_BUFX2_insert648 (
);

FILL SFILL13800x45050 (
);

FILL FILL_4_BUFX2_insert649 (
);

FILL FILL_1__12976_ (
);

FILL FILL_1__12136_ (
);

FILL FILL_0__9983_ (
);

FILL FILL_0__11969_ (
);

FILL FILL_0__9143_ (
);

NAND2X1 _11834_ (
    .A(_2922_),
    .B(_2921_),
    .Y(_2923_)
);

FILL FILL_3__7240_ (
);

FILL FILL_0__11549_ (
);

NAND3X1 _11414_ (
    .A(_2451_),
    .B(_2486_),
    .C(_2530_),
    .Y(_2531_)
);

FILL FILL_0__11129_ (
);

FILL FILL_5__7586_ (
);

FILL FILL_5__7166_ (
);

FILL FILL_4__16362_ (
);

FILL FILL_0__12910_ (
);

FILL FILL_3__15775_ (
);

FILL FILL_3__15355_ (
);

FILL SFILL64920x75050 (
);

FILL FILL_1__7998_ (
);

FILL FILL_1__7578_ (
);

FILL FILL_1__7158_ (
);

FILL FILL_3__10490_ (
);

FILL FILL_2__14768_ (
);

FILL FILL_2__14348_ (
);

FILL FILL_0__15382_ (
);

FILL SFILL28760x3050 (
);

FILL FILL_3__8865_ (
);

FILL FILL_3__8445_ (
);

NAND2X1 _12619_ (
    .A(vdd),
    .B(memoryOutData[17]),
    .Y(_3459_)
);

FILL FILL_4_BUFX2_insert1020 (
);

FILL FILL_1__14702_ (
);

FILL FILL_4_BUFX2_insert1021 (
);

FILL FILL_4_BUFX2_insert1022 (
);

FILL FILL_4_BUFX2_insert1023 (
);

FILL FILL_4_BUFX2_insert1024 (
);

FILL FILL_4_BUFX2_insert1025 (
);

FILL FILL_4__12282_ (
);

FILL FILL_4_BUFX2_insert1026 (
);

FILL FILL_4_BUFX2_insert1027 (
);

FILL FILL_4_BUFX2_insert1028 (
);

FILL FILL_4_BUFX2_insert1029 (
);

FILL FILL_2__6862_ (
);

FILL FILL_5__9732_ (
);

FILL FILL_3__11695_ (
);

FILL FILL_3__11275_ (
);

FILL FILL_0__16167_ (
);

NOR2X1 _16032_ (
    .A(_6486_),
    .B(_6487_),
    .Y(_6488_)
);

FILL FILL_2__10688_ (
);

FILL FILL_2__10268_ (
);

FILL FILL_1__9724_ (
);

FILL FILL_5__11602_ (
);

FILL FILL_6__15081_ (
);

FILL FILL_3_BUFX2_insert660 (
);

FILL FILL_3_BUFX2_insert661 (
);

FILL FILL_3_BUFX2_insert662 (
);

FILL SFILL64040x54050 (
);

FILL FILL_5__14494_ (
);

FILL FILL_3_BUFX2_insert663 (
);

FILL FILL_5__14074_ (
);

FILL FILL_3_BUFX2_insert664 (
);

FILL FILL_1__15907_ (
);

DFFSR _8794_ (
    .Q(\datapath_1.regfile_1.regOut[15] [4]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_913_[4])
);

FILL FILL_3_BUFX2_insert665 (
);

NAND2X1 _8374_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_760_)
);

FILL FILL_3_BUFX2_insert666 (
);

FILL FILL_3_BUFX2_insert667 (
);

FILL FILL_3_BUFX2_insert668 (
);

FILL FILL_3_BUFX2_insert669 (
);

FILL FILL_4__13487_ (
);

FILL FILL_1__10622_ (
);

FILL FILL_2__7227_ (
);

FILL FILL_1__13094_ (
);

DFFSR _12792_ (
    .Q(\aluControl_1.inst [1]),
    .CLK(clk_bF$buf105),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[1])
);

OAI21X1 _12372_ (
    .A(_3312_),
    .B(MemToReg_bF$buf0),
    .C(_3313_),
    .Y(\datapath_1.mux_wd3.dout [9])
);

FILL FILL_0__12087_ (
);

FILL FILL_3__13841_ (
);

FILL FILL_3__13421_ (
);

FILL FILL_3__13001_ (
);

FILL FILL_4__8514_ (
);

FILL FILL_5__15699_ (
);

FILL FILL_2__12834_ (
);

FILL FILL_2__12414_ (
);

FILL FILL_5__15279_ (
);

NAND2X1 _9999_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1579_)
);

DFFSR _9579_ (
    .Q(\datapath_1.regfile_1.regOut[21] [21]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1303_[21])
);

INVX1 _9159_ (
    .A(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_1161_)
);

FILL FILL_1__11827_ (
);

FILL FILL_1__11407_ (
);

FILL FILL_5__16220_ (
);

FILL FILL_0__8834_ (
);

FILL FILL_3__6931_ (
);

FILL FILL_1__14299_ (
);

FILL FILL_5__6857_ (
);

FILL FILL_0_BUFX2_insert790 (
);

FILL FILL_4__15633_ (
);

FILL FILL_0_BUFX2_insert791 (
);

FILL FILL_4__15213_ (
);

FILL FILL_0_BUFX2_insert792 (
);

FILL FILL_0_BUFX2_insert793 (
);

FILL FILL_0_BUFX2_insert794 (
);

NAND3X1 _13997_ (
    .A(_4489_),
    .B(_4490_),
    .C(_4497_),
    .Y(_4498_)
);

FILL FILL_0_BUFX2_insert795 (
);

OAI22X1 _13577_ (
    .A(_3983__bF$buf2),
    .B(_4085_),
    .C(_3977__bF$buf2),
    .D(_4086_),
    .Y(_4087_)
);

INVX1 _13157_ (
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3736_)
);

FILL FILL_0_BUFX2_insert796 (
);

FILL FILL_0_BUFX2_insert797 (
);

FILL FILL_3__14626_ (
);

FILL FILL_0_BUFX2_insert798 (
);

FILL FILL_0_BUFX2_insert799 (
);

FILL FILL_1__15660_ (
);

FILL FILL_3__14206_ (
);

FILL FILL_1__15240_ (
);

FILL FILL_1__6849_ (
);

FILL FILL_4__9719_ (
);

FILL FILL_2__13619_ (
);

FILL FILL_0__14653_ (
);

FILL FILL_0__14233_ (
);

FILL FILL_5__11199_ (
);

FILL SFILL54040x52050 (
);

FILL FILL_3__7716_ (
);

FILL FILL_0__9619_ (
);

FILL FILL_5__12980_ (
);

FILL FILL_5__12140_ (
);

BUFX2 _6860_ (
    .A(_1_[22]),
    .Y(memoryAddress[22])
);

FILL FILL_4__11973_ (
);

FILL FILL_4__11553_ (
);

FILL FILL_4__11133_ (
);

FILL FILL_1__16025_ (
);

FILL FILL_3__10966_ (
);

FILL FILL_3__10546_ (
);

FILL FILL_3__10126_ (
);

FILL FILL_1__11580_ (
);

FILL FILL_1__11160_ (
);

FILL FILL_0__15858_ (
);

INVX1 _15723_ (
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_6187_)
);

FILL FILL_0__15438_ (
);

NAND3X1 _15303_ (
    .A(_5771_),
    .B(_5772_),
    .C(_5776_),
    .Y(_5777_)
);

FILL FILL_0__15018_ (
);

FILL FILL_0__10993_ (
);

FILL FILL_0__10573_ (
);

FILL FILL_2__8185_ (
);

FILL FILL_0__10153_ (
);

FILL FILL_2__10900_ (
);

FILL FILL_5__13765_ (
);

FILL FILL_5__13345_ (
);

FILL SFILL54360x28050 (
);

DFFSR _7645_ (
    .Q(\datapath_1.regfile_1.regOut[6] [7]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_328_[7])
);

NAND2X1 _7225_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_177_)
);

FILL FILL_4__9892_ (
);

FILL FILL_4__9472_ (
);

FILL FILL_4__12758_ (
);

FILL FILL_2__13792_ (
);

FILL FILL_4__12338_ (
);

FILL FILL_2__13372_ (
);

FILL FILL_0__6900_ (
);

FILL FILL_2__6918_ (
);

FILL FILL_1__12785_ (
);

FILL FILL_1__12365_ (
);

FILL FILL_0__9792_ (
);

FILL FILL_0__9372_ (
);

FILL FILL_0__11778_ (
);

FILL FILL_0__11358_ (
);

AOI21X1 _11643_ (
    .A(_2161_),
    .B(_2745_),
    .C(_2337_),
    .Y(_2746_)
);

NAND2X1 _11223_ (
    .A(_2107_),
    .B(_2341__bF$buf2),
    .Y(_2342_)
);

FILL FILL_6__15557_ (
);

FILL FILL_6__15137_ (
);

FILL FILL_4__16171_ (
);

FILL SFILL44040x50050 (
);

FILL FILL_6__10692_ (
);

FILL FILL_3__15584_ (
);

FILL FILL_3__15164_ (
);

FILL FILL_2__14997_ (
);

FILL FILL_2__14577_ (
);

FILL FILL_2__14157_ (
);

FILL FILL_0__15191_ (
);

FILL FILL_5__15911_ (
);

FILL SFILL23000x59050 (
);

FILL FILL_4__14904_ (
);

FILL FILL_3__8254_ (
);

NAND2X1 _12848_ (
    .A(vdd),
    .B(\datapath_1.rd1 [8]),
    .Y(_3571_)
);

NAND2X1 _12428_ (
    .A(MemToReg_bF$buf2),
    .B(\datapath_1.Data [28]),
    .Y(_3351_)
);

NAND3X1 _12008_ (
    .A(PCSource_1_bF$buf4),
    .B(\aluControl_1.inst [3]),
    .C(_3034__bF$buf1),
    .Y(_3052_)
);

FILL FILL_1__14931_ (
);

FILL FILL_1__14511_ (
);

FILL FILL_6__11477_ (
);

FILL FILL_6__11057_ (
);

FILL FILL_4__12091_ (
);

FILL FILL_0__13924_ (
);

FILL FILL_3__16369_ (
);

FILL FILL_0__13504_ (
);

FILL FILL_5__9541_ (
);

FILL FILL_5__9121_ (
);

FILL FILL_3__11084_ (
);

FILL FILL_0__16396_ (
);

OAI22X1 _16261_ (
    .A(_5472__bF$buf0),
    .B(_5393_),
    .C(_5392_),
    .D(_5552__bF$buf1),
    .Y(_6711_)
);

FILL FILL_2__10497_ (
);

FILL FILL_5__11831_ (
);

FILL FILL_1__9533_ (
);

FILL FILL_5__11411_ (
);

FILL FILL_1__9113_ (
);

FILL FILL_3__9879_ (
);

FILL FILL_2__16303_ (
);

FILL FILL_3__9039_ (
);

FILL FILL_4__10824_ (
);

FILL FILL_4__10404_ (
);

FILL FILL_1__15716_ (
);

NAND2X1 _8183_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .Y(_717_)
);

FILL FILL_4__13296_ (
);

FILL FILL_1__10431_ (
);

FILL FILL_1__10011_ (
);

FILL SFILL69160x61050 (
);

FILL FILL_0__14709_ (
);

FILL FILL_2__7876_ (
);

FILL FILL_2__7456_ (
);

FILL FILL_3__12289_ (
);

FILL FILL_2__7036_ (
);

FILL FILL_6__13623_ (
);

FILL SFILL74120x44050 (
);

INVX1 _12181_ (
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3174_)
);

FILL FILL_5__12616_ (
);

FILL FILL_3__13650_ (
);

FILL FILL_3__13230_ (
);

OAI21X1 _6916_ (
    .A(_10_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .C(_11_),
    .Y(_3_[4])
);

FILL FILL_4__8743_ (
);

FILL FILL_4__8323_ (
);

FILL FILL_4__11609_ (
);

FILL FILL_2__12643_ (
);

FILL FILL_5__15088_ (
);

FILL FILL_2__12223_ (
);

INVX1 _9388_ (
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_1273_)
);

FILL FILL_1__11636_ (
);

FILL FILL_1__11216_ (
);

FILL FILL_6_BUFX2_insert40 (
);

FILL FILL_0__8643_ (
);

NAND2X1 _10914_ (
    .A(\control_1.reg_state.dout [2]),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2058_)
);

FILL FILL_0__10629_ (
);

FILL FILL_0__8223_ (
);

FILL FILL_6_BUFX2_insert45 (
);

FILL FILL_4__15862_ (
);

FILL FILL_4__15442_ (
);

FILL FILL_4__15022_ (
);

INVX4 _13386_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_3898_)
);

FILL FILL_3__14855_ (
);

FILL FILL_2__9602_ (
);

FILL FILL_3__14435_ (
);

FILL FILL_3__14015_ (
);

FILL FILL_4__9528_ (
);

FILL FILL_4__9108_ (
);

FILL FILL_2__13848_ (
);

FILL SFILL24440x60050 (
);

FILL FILL_2__13428_ (
);

FILL FILL_0__14882_ (
);

FILL FILL_0__14462_ (
);

FILL FILL_2__13008_ (
);

FILL FILL_0__14042_ (
);

FILL FILL_3__7945_ (
);

FILL FILL_0__9848_ (
);

FILL FILL_0__9428_ (
);

FILL FILL_0__9008_ (
);

FILL FILL_3__7105_ (
);

FILL FILL_4__16227_ (
);

FILL FILL_4__11782_ (
);

FILL FILL_4__11362_ (
);

FILL SFILL64120x42050 (
);

FILL FILL_1__16254_ (
);

FILL FILL_3__10775_ (
);

FILL FILL_0__15667_ (
);

INVX1 _15952_ (
    .A(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_6410_)
);

FILL FILL_0__15247_ (
);

OAI22X1 _15532_ (
    .A(_4494_),
    .B(_5544__bF$buf1),
    .C(_5523_),
    .D(_6000_),
    .Y(_6001_)
);

NOR2X1 _15112_ (
    .A(_5590_),
    .B(_5589_),
    .Y(_5591_)
);

FILL FILL_0__10382_ (
);

FILL SFILL64040x49050 (
);

FILL FILL_5__13994_ (
);

FILL FILL_5__13574_ (
);

FILL FILL_5__13154_ (
);

NAND2X1 _7874_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_508_)
);

NAND2X1 _7454_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_289_)
);

NAND2X1 _7034_ (
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_70_)
);

FILL FILL_4__12987_ (
);

FILL FILL_4__9281_ (
);

FILL FILL_4__12567_ (
);

FILL FILL_4__12147_ (
);

FILL FILL_1__12594_ (
);

FILL FILL_1__12174_ (
);

NOR2X1 _16317_ (
    .A(_6763_),
    .B(_6765_),
    .Y(_6766_)
);

INVX1 _11872_ (
    .A(\datapath_1.PCJump [18]),
    .Y(_2958_)
);

FILL FILL_0__11587_ (
);

FILL FILL_0__11167_ (
);

NAND2X1 _11452_ (
    .A(_2551_),
    .B(_2567_),
    .Y(_2568_)
);

INVX1 _11032_ (
    .A(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2151_)
);

FILL FILL_3__12501_ (
);

FILL FILL_2__11914_ (
);

FILL FILL_5__14779_ (
);

FILL FILL_5__14359_ (
);

FILL FILL_3__15393_ (
);

INVX1 _8659_ (
    .A(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_909_)
);

INVX1 _8239_ (
    .A(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_690_)
);

FILL FILL_1__7196_ (
);

FILL FILL_1__10907_ (
);

FILL FILL_2__14386_ (
);

FILL FILL_5__15720_ (
);

FILL FILL_5__15300_ (
);

FILL FILL_1__13799_ (
);

NAND2X1 _9600_ (
    .A(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1374_)
);

FILL SFILL54120x40050 (
);

FILL FILL_1__13379_ (
);

FILL SFILL39000x50 (
);

FILL FILL_4__14713_ (
);

FILL FILL_3__8483_ (
);

INVX1 _12657_ (
    .A(\datapath_1.Data [30]),
    .Y(_3484_)
);

FILL FILL_3__8063_ (
);

AOI22X1 _12237_ (
    .A(_2_[5]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf3),
    .D(\aluControl_1.inst [3]),
    .Y(_3217_)
);

FILL FILL_3__13706_ (
);

FILL SFILL18680x73050 (
);

FILL FILL_1__14740_ (
);

FILL FILL_1__14320_ (
);

FILL FILL_0__13733_ (
);

FILL FILL_0__13313_ (
);

FILL FILL_3__16178_ (
);

FILL FILL_5__10699_ (
);

FILL FILL_5__9770_ (
);

FILL FILL_5__10279_ (
);

FILL FILL_5__9350_ (
);

AOI21X1 _16070_ (
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .B(_5567_),
    .C(_6524_),
    .Y(_6525_)
);

FILL FILL_1__9762_ (
);

FILL FILL_5__11640_ (
);

FILL FILL_5__11220_ (
);

FILL FILL_1__9342_ (
);

FILL FILL_4__15918_ (
);

FILL FILL_2__16112_ (
);

FILL FILL_3__9268_ (
);

FILL FILL_4__10633_ (
);

FILL FILL_1__15945_ (
);

FILL FILL_1__15525_ (
);

FILL FILL_1__15105_ (
);

FILL FILL_1__10660_ (
);

FILL FILL_1__10240_ (
);

FILL FILL_0__14938_ (
);

AOI22X1 _14803_ (
    .A(_4129_),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .C(\datapath_1.regfile_1.regOut[18] [28]),
    .D(_4135_),
    .Y(_5287_)
);

FILL FILL_0__14518_ (
);

FILL FILL_2__7685_ (
);

FILL FILL_3__12098_ (
);

FILL FILL_5__12845_ (
);

FILL FILL_5__12425_ (
);

FILL FILL_5__12005_ (
);

FILL SFILL79240x51050 (
);

FILL FILL_4__8972_ (
);

FILL FILL_4__8132_ (
);

FILL FILL_4__11838_ (
);

FILL FILL_2__12872_ (
);

FILL FILL_4__11418_ (
);

FILL FILL_2__12452_ (
);

FILL FILL_2__12032_ (
);

FILL FILL_6__8898_ (
);

DFFSR _9197_ (
    .Q(\datapath_1.regfile_1.regOut[18] [23]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1108_[23])
);

FILL FILL111880x64050 (
);

FILL FILL_1__11865_ (
);

FILL FILL_1__11445_ (
);

FILL FILL_1__11025_ (
);

FILL FILL_0__8872_ (
);

FILL FILL_0__8452_ (
);

FILL FILL_0__10438_ (
);

DFFSR _10723_ (
    .Q(\datapath_1.regfile_1.regOut[30] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_1888_[13])
);

NAND2X1 _10303_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1741_)
);

FILL FILL_0__10018_ (
);

FILL FILL_5__6895_ (
);

FILL FILL_4__15671_ (
);

FILL SFILL44040x45050 (
);

FILL FILL_4__15251_ (
);

DFFSR _13195_ (
    .Q(\datapath_1.mux_iord.din0 [20]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3685_[20])
);

FILL FILL_2__9411_ (
);

FILL FILL_3__14664_ (
);

FILL FILL_3__14244_ (
);

FILL FILL_1__6887_ (
);

FILL FILL112200x5050 (
);

FILL FILL_4__9757_ (
);

FILL FILL_4__9337_ (
);

FILL FILL_2__13657_ (
);

FILL FILL_2__13237_ (
);

FILL FILL_0__14691_ (
);

FILL FILL_0__14271_ (
);

FILL FILL_3__7754_ (
);

FILL FILL_0__9657_ (
);

FILL FILL_3__7334_ (
);

OAI21X1 _11928_ (
    .A(_2992_),
    .B(IorD_bF$buf3),
    .C(_2993_),
    .Y(_1_[13])
);

FILL FILL_0__9237_ (
);

INVX8 _11508_ (
    .A(_2347__bF$buf1),
    .Y(_2620_)
);

FILL FILL_4__16036_ (
);

FILL SFILL109400x32050 (
);

FILL FILL_4__11591_ (
);

FILL FILL_4__11171_ (
);

FILL FILL_3__15869_ (
);

FILL FILL_3__15449_ (
);

FILL FILL_3__15029_ (
);

FILL FILL_1__16063_ (
);

FILL FILL_5__8621_ (
);

FILL FILL_5__8201_ (
);

FILL FILL_3__10164_ (
);

FILL FILL_6_BUFX2_insert551 (
);

FILL FILL_0__15896_ (
);

OAI22X1 _15761_ (
    .A(_5480__bF$buf1),
    .B(_4789_),
    .C(_4775_),
    .D(_5499__bF$buf0),
    .Y(_6224_)
);

FILL FILL_0__15476_ (
);

NOR2X1 _15341_ (
    .A(_4339_),
    .B(_5534__bF$buf0),
    .Y(_5814_)
);

FILL FILL_0__15056_ (
);

FILL FILL_6_BUFX2_insert556 (
);

FILL FILL_0__10191_ (
);

FILL FILL_5__10911_ (
);

FILL FILL_1__8613_ (
);

FILL FILL_6__14390_ (
);

FILL FILL_2__15803_ (
);

FILL FILL_3__8959_ (
);

FILL FILL_3__8119_ (
);

FILL FILL_5__13383_ (
);

NAND2X1 _7683_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_401_)
);

DFFSR _7263_ (
    .Q(\datapath_1.regfile_1.regOut[3] [9]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_133_[9])
);

FILL SFILL99400x81050 (
);

FILL FILL_4__9090_ (
);

FILL FILL_4__12376_ (
);

FILL FILL_3__9900_ (
);

FILL FILL_2__6956_ (
);

FILL FILL_3__11789_ (
);

FILL FILL_5__9406_ (
);

FILL FILL_3__11369_ (
);

OAI22X1 _16126_ (
    .A(_5252_),
    .B(_5469__bF$buf2),
    .C(_5463__bF$buf0),
    .D(_6578_),
    .Y(_6579_)
);

NAND2X1 _11681_ (
    .A(_2397_),
    .B(_2481__bF$buf3),
    .Y(_2782_)
);

FILL FILL_0__11396_ (
);

NAND2X1 _11261_ (
    .A(_2168_),
    .B(_2169_),
    .Y(_2380_)
);

FILL FILL_3__12730_ (
);

FILL FILL_3__12310_ (
);

FILL FILL_4__7823_ (
);

FILL FILL_5__14588_ (
);

FILL FILL_2__11723_ (
);

FILL FILL_5__14168_ (
);

FILL FILL_2__11303_ (
);

INVX1 _8888_ (
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_1021_)
);

INVX1 _8468_ (
    .A(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_802_)
);

DFFSR _8048_ (
    .Q(\datapath_1.regfile_1.regOut[9] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_523_[26])
);

FILL FILL_2__14195_ (
);

FILL SFILL38760x20050 (
);

FILL FILL_0__7723_ (
);

FILL SFILL69160x11050 (
);

FILL FILL_0__7303_ (
);

FILL FILL_4__14942_ (
);

FILL FILL_4__14522_ (
);

FILL FILL_4__14102_ (
);

INVX1 _12886_ (
    .A(\datapath_1.a [21]),
    .Y(_3596_)
);

INVX1 _12466_ (
    .A(ALUOut[9]),
    .Y(_3377_)
);

NAND3X1 _12046_ (
    .A(_3078_),
    .B(_3079_),
    .C(_3080_),
    .Y(\datapath_1.mux_pcsrc.dout [14])
);

FILL FILL_3__13935_ (
);

FILL FILL_3__13515_ (
);

FILL FILL_4__8608_ (
);

FILL FILL_5_BUFX2_insert570 (
);

FILL FILL_5_BUFX2_insert571 (
);

FILL FILL_5_BUFX2_insert572 (
);

FILL FILL_2__12508_ (
);

FILL FILL_0__13962_ (
);

FILL SFILL99320x43050 (
);

FILL FILL_5_BUFX2_insert573 (
);

FILL FILL_0__13542_ (
);

FILL SFILL38680x27050 (
);

FILL FILL_0__13122_ (
);

FILL FILL_5_BUFX2_insert574 (
);

FILL FILL_5_BUFX2_insert575 (
);

FILL FILL_5_BUFX2_insert576 (
);

FILL FILL_5_BUFX2_insert577 (
);

FILL FILL_5_BUFX2_insert578 (
);

FILL FILL_5_BUFX2_insert579 (
);

FILL FILL_5__16314_ (
);

FILL SFILL28760x63050 (
);

FILL FILL_0__8508_ (
);

FILL FILL_1__9991_ (
);

FILL FILL_1__9151_ (
);

FILL FILL_4__15727_ (
);

FILL FILL_4__15307_ (
);

FILL FILL_2__16341_ (
);

FILL FILL_3__9497_ (
);

FILL FILL_4__10442_ (
);

FILL SFILL64120x37050 (
);

FILL FILL_4__10022_ (
);

FILL FILL_1__15754_ (
);

FILL FILL_1__15334_ (
);

FILL FILL_0__14747_ (
);

OAI22X1 _14612_ (
    .A(_3893__bF$buf2),
    .B(_5099_),
    .C(_3930__bF$buf3),
    .D(_5098_),
    .Y(_5100_)
);

FILL FILL_0__14327_ (
);

FILL FILL_2__7494_ (
);

FILL FILL_2__7074_ (
);

FILL FILL_5__12654_ (
);

FILL FILL_5__12234_ (
);

NAND2X1 _6954_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_37_)
);

FILL SFILL84200x4050 (
);

FILL FILL_4__8781_ (
);

FILL FILL_4__8361_ (
);

FILL FILL_4__11647_ (
);

FILL FILL_4__11227_ (
);

FILL FILL_2__12261_ (
);

FILL FILL_1__16119_ (
);

FILL FILL_1__11674_ (
);

FILL FILL_1__11254_ (
);

AOI22X1 _15817_ (
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .B(_5494_),
    .C(_5479_),
    .D(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_6278_)
);

FILL SFILL33960x81050 (
);

FILL FILL_2__8699_ (
);

NOR2X1 _10952_ (
    .A(\control_1.op [2]),
    .B(\control_1.op [3]),
    .Y(_2085_)
);

FILL FILL_0__8261_ (
);

FILL FILL_0__10667_ (
);

NAND2X1 _10532_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1853_)
);

FILL FILL_0__10247_ (
);

NAND2X1 _10112_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1634_)
);

FILL FILL_6__14866_ (
);

FILL FILL_4__15480_ (
);

FILL FILL_4__15060_ (
);

FILL FILL_5__13859_ (
);

FILL FILL_2__9640_ (
);

FILL FILL_5__13439_ (
);

FILL FILL_3__14893_ (
);

FILL FILL_3__14473_ (
);

FILL FILL_2__9220_ (
);

FILL FILL_5__13019_ (
);

INVX1 _7739_ (
    .A(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_438_)
);

FILL FILL_3__14053_ (
);

FILL SFILL18760x61050 (
);

INVX1 _7319_ (
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_219_)
);

FILL FILL_4__9986_ (
);

FILL FILL_4__9146_ (
);

FILL FILL_2__13886_ (
);

FILL FILL_2__13466_ (
);

FILL FILL_2__13046_ (
);

FILL FILL_0__14080_ (
);

FILL FILL_5__14800_ (
);

FILL SFILL54120x35050 (
);

FILL FILL_1__12879_ (
);

FILL FILL_1__12459_ (
);

FILL FILL_1__12039_ (
);

FILL FILL_6_CLKBUF1_insert152 (
);

FILL FILL_3__7983_ (
);

FILL FILL_0__9886_ (
);

FILL FILL_3__7563_ (
);

FILL FILL_0__9466_ (
);

NAND3X1 _11737_ (
    .A(_2168_),
    .B(_2198_),
    .C(_2833_),
    .Y(_2834_)
);

FILL FILL_6_CLKBUF1_insert157 (
);

OAI21X1 _11317_ (
    .A(_2415_),
    .B(_2428_),
    .C(_2435_),
    .Y(_2436_)
);

FILL FILL_1__13820_ (
);

FILL FILL_5__7489_ (
);

FILL FILL_1__13400_ (
);

FILL FILL_4__16265_ (
);

FILL FILL_5__7069_ (
);

FILL FILL_6__10786_ (
);

FILL FILL_3__15678_ (
);

FILL FILL_3__15258_ (
);

FILL FILL_1__16292_ (
);

FILL FILL_5__8850_ (
);

FILL FILL_3__10393_ (
);

FILL FILL_5__8010_ (
);

NAND3X1 _15990_ (
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf2),
    .Y(_6447_)
);

NOR3X1 _15570_ (
    .A(_6037_),
    .B(_6033_),
    .C(_6036_),
    .Y(_6038_)
);

FILL FILL_0__15285_ (
);

NOR2X1 _15150_ (
    .A(_5625_),
    .B(_5627_),
    .Y(_5628_)
);

FILL FILL_1__8842_ (
);

FILL FILL_5__10300_ (
);

FILL FILL_1__8002_ (
);

FILL FILL_2__15612_ (
);

FILL FILL_3__8768_ (
);

FILL FILL_3__8348_ (
);

FILL FILL_1__14605_ (
);

INVX1 _7492_ (
    .A(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_314_)
);

INVX1 _7072_ (
    .A(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_95_)
);

FILL SFILL18680x23050 (
);

FILL FILL_4__12185_ (
);

FILL FILL_5__9635_ (
);

FILL FILL_3__11598_ (
);

FILL FILL_5__9215_ (
);

FILL FILL_3__11178_ (
);

FILL FILL111960x52050 (
);

NAND2X1 _16355_ (
    .A(gnd),
    .B(gnd),
    .Y(_6791_)
);

NAND2X1 _11490_ (
    .A(_2554_),
    .B(_2549_),
    .Y(_2603_)
);

FILL FILL_5__11925_ (
);

INVX1 _11070_ (
    .A(\datapath_1.alu_1.ALUInB [10]),
    .Y(_2189_)
);

FILL FILL_1__9627_ (
);

FILL FILL_5__11505_ (
);

FILL FILL_1__9207_ (
);

FILL SFILL79240x46050 (
);

FILL FILL_4__7632_ (
);

FILL FILL_4__10918_ (
);

FILL FILL_4__7212_ (
);

FILL FILL_2__11952_ (
);

FILL FILL_5__14397_ (
);

FILL FILL_2__11532_ (
);

FILL FILL_6__7978_ (
);

FILL FILL_2__11112_ (
);

INVX1 _8697_ (
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_914_)
);

OAI21X1 _8277_ (
    .A(_714_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_715_),
    .Y(_653_[31])
);

FILL FILL_1__10945_ (
);

FILL FILL_1__10525_ (
);

FILL FILL_1__10105_ (
);

FILL FILL_0__7952_ (
);

BUFX2 BUFX2_insert390 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf3 )
);

BUFX2 BUFX2_insert391 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf2 )
);

FILL FILL_0__7112_ (
);

BUFX2 BUFX2_insert392 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf1 )
);

BUFX2 BUFX2_insert393 (
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf0 )
);

BUFX2 BUFX2_insert394 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf7 )
);

FILL SFILL54120x8050 (
);

FILL FILL_4__14751_ (
);

BUFX2 BUFX2_insert395 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf6 )
);

BUFX2 BUFX2_insert396 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf5 )
);

FILL FILL_4__14331_ (
);

FILL SFILL94360x6050 (
);

BUFX2 BUFX2_insert397 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf4 )
);

BUFX2 BUFX2_insert398 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf3 )
);

INVX1 _12695_ (
    .A(\aluControl_1.inst [0]),
    .Y(_3553_)
);

BUFX2 BUFX2_insert399 (
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf2 )
);

NAND3X1 _12275_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3245_)
);

FILL FILL_2__8911_ (
);

FILL FILL_3__13744_ (
);

FILL FILL_3__13324_ (
);

FILL FILL_4__8837_ (
);

FILL FILL_2__12737_ (
);

FILL SFILL114360x71050 (
);

FILL FILL_0__13771_ (
);

FILL FILL_2__12317_ (
);

FILL FILL_0__13351_ (
);

FILL FILL111880x14050 (
);

FILL FILL_0__8737_ (
);

FILL FILL_5__16123_ (
);

FILL FILL_0__8317_ (
);

FILL SFILL104520x9050 (
);

FILL FILL_1__9380_ (
);

FILL FILL_4__15956_ (
);

FILL FILL_4__15536_ (
);

FILL FILL_4__15116_ (
);

FILL SFILL109400x27050 (
);

FILL FILL_2__16150_ (
);

FILL FILL_4__10671_ (
);

FILL FILL_4__10251_ (
);

FILL FILL_3__14949_ (
);

FILL FILL_1__15983_ (
);

FILL FILL_3__14529_ (
);

FILL FILL_1__15563_ (
);

FILL FILL_3__14109_ (
);

FILL FILL_1__15143_ (
);

FILL FILL_5__7701_ (
);

FILL FILL_0__14976_ (
);

FILL FILL_0__14556_ (
);

OAI22X1 _14841_ (
    .A(_5322_),
    .B(_3944__bF$buf2),
    .C(_3954__bF$buf3),
    .D(_5323_),
    .Y(_5324_)
);

FILL FILL_0__14136_ (
);

NOR2X1 _14421_ (
    .A(_4909_),
    .B(_4912_),
    .Y(_4913_)
);

AOI21X1 _14001_ (
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .B(_4225_),
    .C(_4501_),
    .Y(_4502_)
);

FILL FILL_3__7619_ (
);

FILL FILL_5__12883_ (
);

FILL FILL_5__12463_ (
);

FILL FILL_5__12043_ (
);

FILL FILL_4__8590_ (
);

FILL FILL_4__11876_ (
);

FILL SFILL104760x83050 (
);

FILL FILL_4__11456_ (
);

FILL FILL_2__12490_ (
);

FILL FILL_4__11036_ (
);

FILL FILL_2__12070_ (
);

FILL FILL_1__16348_ (
);

FILL FILL_5__8906_ (
);

FILL FILL_3__10449_ (
);

FILL FILL_3__10029_ (
);

FILL FILL_1__11483_ (
);

FILL FILL_1__11063_ (
);

NOR2X1 _15626_ (
    .A(_6091_),
    .B(_5530__bF$buf2),
    .Y(_6092_)
);

NAND2X1 _15206_ (
    .A(_5678_),
    .B(_5682_),
    .Y(_5683_)
);

FILL FILL_0__10896_ (
);

FILL FILL_0__8490_ (
);

NAND2X1 _10761_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1965_)
);

FILL FILL_2__8088_ (
);

FILL FILL_0__8070_ (
);

DFFSR _10341_ (
    .Q(\datapath_1.regfile_1.regOut[27] [15]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_1693_[15])
);

FILL FILL_0__10056_ (
);

FILL FILL_3__11810_ (
);

FILL FILL_4__6903_ (
);

FILL FILL_5__13668_ (
);

FILL FILL_2__10803_ (
);

FILL FILL_5__13248_ (
);

INVX1 _7968_ (
    .A(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_550_)
);

FILL FILL_3__14282_ (
);

INVX1 _7548_ (
    .A(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_331_)
);

DFFSR _7128_ (
    .Q(\datapath_1.regfile_1.regOut[2] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_68_[2])
);

FILL FILL_4__9795_ (
);

FILL FILL_4__9375_ (
);

FILL FILL_2__13695_ (
);

FILL FILL_2__13275_ (
);

FILL SFILL99400x31050 (
);

FILL FILL_1__12268_ (
);

FILL FILL_4__13602_ (
);

FILL FILL_3__7372_ (
);

FILL FILL_0__9275_ (
);

NAND2X1 _11966_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[26]),
    .Y(_3019_)
);

AOI21X1 _11546_ (
    .A(_2409_),
    .B(_2620_),
    .C(_2655_),
    .Y(_2656_)
);

FILL FILL_5_CLKBUF1_insert140 (
);

INVX2 _11126_ (
    .A(_2244_),
    .Y(_2245_)
);

FILL FILL_5_CLKBUF1_insert141 (
);

FILL FILL_5_CLKBUF1_insert142 (
);

FILL FILL_5__7298_ (
);

FILL FILL_5_CLKBUF1_insert143 (
);

FILL FILL_5_CLKBUF1_insert144 (
);

FILL FILL_4__16074_ (
);

FILL FILL_5_CLKBUF1_insert145 (
);

FILL FILL_5_CLKBUF1_insert146 (
);

FILL FILL_5_CLKBUF1_insert147 (
);

FILL FILL_5_CLKBUF1_insert148 (
);

FILL SFILL99320x38050 (
);

FILL FILL_5_CLKBUF1_insert149 (
);

FILL FILL_0__12622_ (
);

FILL FILL_3__15487_ (
);

FILL FILL_0__12202_ (
);

FILL FILL_3__15067_ (
);

FILL FILL_6__16401_ (
);

FILL FILL_6_BUFX2_insert930 (
);

FILL FILL_6_BUFX2_insert935 (
);

FILL FILL_0__15094_ (
);

FILL FILL_5__15814_ (
);

FILL FILL_1__8651_ (
);

FILL FILL_1__8231_ (
);

FILL SFILL3720x6050 (
);

FILL FILL_4__14807_ (
);

FILL FILL_2__15841_ (
);

FILL FILL_3__8997_ (
);

FILL FILL_2__15421_ (
);

FILL FILL_3__8577_ (
);

FILL FILL_2__15001_ (
);

FILL FILL_1__14834_ (
);

FILL FILL_1__14414_ (
);

FILL SFILL28360x44050 (
);

FILL FILL_0__13827_ (
);

FILL FILL_0__13407_ (
);

FILL FILL_2__6994_ (
);

FILL FILL_5__9864_ (
);

FILL FILL_5__9024_ (
);

FILL FILL_0__16299_ (
);

FILL FILL_6__12321_ (
);

AOI21X1 _16164_ (
    .A(_6593_),
    .B(_6616_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [27])
);

FILL FILL_1__9856_ (
);

FILL FILL_5__11734_ (
);

FILL FILL_5__11314_ (
);

FILL SFILL28760x13050 (
);

FILL FILL_1__9016_ (
);

FILL SFILL94280x80050 (
);

FILL FILL_4__7861_ (
);

FILL FILL_2__16206_ (
);

FILL FILL_4__7441_ (
);

FILL FILL_2__11761_ (
);

FILL FILL_4__10307_ (
);

FILL FILL_2__11341_ (
);

FILL FILL_1__15619_ (
);

OAI21X1 _8086_ (
    .A(_607_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_608_),
    .Y(_588_[10])
);

FILL SFILL113720x2050 (
);

FILL FILL_1__10754_ (
);

FILL FILL_0__7761_ (
);

FILL FILL_2__7359_ (
);

FILL FILL_0__7341_ (
);

FILL FILL_4__14980_ (
);

FILL FILL_6__13526_ (
);

FILL FILL_4__14560_ (
);

FILL FILL_4__14140_ (
);

NAND3X1 _12084_ (
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [24]),
    .C(_3034__bF$buf0),
    .Y(_3109_)
);

FILL FILL_2__8720_ (
);

FILL FILL_5__12519_ (
);

FILL FILL_3__13973_ (
);

FILL FILL_3__13553_ (
);

FILL SFILL18760x56050 (
);

FILL FILL_3__13133_ (
);

FILL FILL_4__8646_ (
);

FILL FILL_4__8226_ (
);

FILL FILL_5_BUFX2_insert950 (
);

FILL FILL_5_BUFX2_insert951 (
);

FILL FILL_2__12966_ (
);

FILL FILL_5_BUFX2_insert952 (
);

FILL FILL_2__12126_ (
);

FILL FILL_0__13580_ (
);

FILL FILL_5_BUFX2_insert953 (
);

FILL FILL_5_BUFX2_insert954 (
);

FILL FILL_0__13160_ (
);

FILL FILL_5_BUFX2_insert955 (
);

FILL SFILL73640x58050 (
);

FILL FILL_5_BUFX2_insert956 (
);

FILL FILL_5_BUFX2_insert957 (
);

FILL FILL_1__11959_ (
);

FILL FILL_5_BUFX2_insert958 (
);

FILL FILL_5_BUFX2_insert959 (
);

FILL FILL_1__11539_ (
);

FILL FILL_1__11119_ (
);

FILL FILL_0__8966_ (
);

FILL FILL_5__16352_ (
);

FILL FILL_0__8126_ (
);

FILL FILL_6__9513_ (
);

INVX1 _10817_ (
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_2002_)
);

FILL SFILL33960x31050 (
);

FILL FILL_5__6989_ (
);

FILL FILL_4__15765_ (
);

FILL FILL_1__12900_ (
);

FILL FILL_4__15345_ (
);

OR2X2 _13289_ (
    .A(_3826_),
    .B(\datapath_1.a3 [4]),
    .Y(_3827_)
);

FILL FILL_4__10060_ (
);

FILL FILL_2__9925_ (
);

FILL FILL_2__9505_ (
);

FILL FILL_3__14758_ (
);

FILL FILL_3__14338_ (
);

FILL FILL_1__15792_ (
);

FILL FILL_1__15372_ (
);

FILL FILL_5__7930_ (
);

FILL SFILL18760x11050 (
);

FILL FILL_0__14785_ (
);

FILL FILL_0__14365_ (
);

OAI22X1 _14650_ (
    .A(_5135_),
    .B(_3890_),
    .C(_3960_),
    .D(_5136_),
    .Y(_5137_)
);

OAI22X1 _14230_ (
    .A(_3982__bF$buf3),
    .B(_4724_),
    .C(_3971__bF$buf4),
    .D(_4725_),
    .Y(_4726_)
);

FILL FILL_1__7502_ (
);

FILL FILL_3__7848_ (
);

FILL FILL_3__7428_ (
);

FILL FILL_5__12272_ (
);

INVX1 _6992_ (
    .A(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_62_)
);

FILL SFILL79320x34050 (
);

FILL SFILL18680x18050 (
);

FILL FILL_4__11685_ (
);

FILL FILL_4__11265_ (
);

FILL FILL_1__16157_ (
);

FILL FILL_3__10678_ (
);

FILL FILL_5__8715_ (
);

FILL FILL_3__10258_ (
);

FILL FILL_1__11292_ (
);

AOI22X1 _15855_ (
    .A(_5490_),
    .B(\datapath_1.regfile_1.regOut[7] [20]),
    .C(\datapath_1.regfile_1.regOut[10] [20]),
    .D(_6314_),
    .Y(_6315_)
);

NAND2X1 _15435_ (
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .B(_5570__bF$buf1),
    .Y(_5906_)
);

NAND3X1 _15015_ (
    .A(_5459__bF$buf2),
    .B(_5468_),
    .C(_5465_),
    .Y(_5495_)
);

INVX1 _10990_ (
    .A(_2108_),
    .Y(_2109_)
);

INVX1 _10570_ (
    .A(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_1878_)
);

FILL FILL_0__10285_ (
);

INVX1 _10150_ (
    .A(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_1659_)
);

FILL FILL_3_BUFX2_insert1030 (
);

FILL FILL_1__8707_ (
);

FILL FILL_3_BUFX2_insert1031 (
);

FILL FILL_3_BUFX2_insert1032 (
);

FILL FILL_3_BUFX2_insert1033 (
);

FILL FILL_3_BUFX2_insert1034 (
);

FILL FILL_3_BUFX2_insert1035 (
);

FILL FILL_3_BUFX2_insert1036 (
);

FILL FILL_3_BUFX2_insert1037 (
);

FILL FILL_3_BUFX2_insert1038 (
);

FILL FILL_5__13897_ (
);

FILL FILL_3_BUFX2_insert1039 (
);

FILL FILL_5__13477_ (
);

DFFSR _7777_ (
    .Q(\datapath_1.regfile_1.regOut[7] [11]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_393_[11])
);

FILL FILL_3__14091_ (
);

OAI21X1 _7357_ (
    .A(_243_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_244_),
    .Y(_198_[23])
);

FILL FILL_2__13084_ (
);

FILL FILL_1__12497_ (
);

FILL FILL_1__12077_ (
);

FILL SFILL110040x58050 (
);

FILL FILL_4__13831_ (
);

FILL FILL_4__13411_ (
);

FILL FILL_3__7181_ (
);

NOR2X1 _11775_ (
    .A(_2337_),
    .B(_2852_),
    .Y(_2869_)
);

FILL FILL_0__9084_ (
);

NOR2X1 _11355_ (
    .A(_2472_),
    .B(_2464_),
    .Y(_2473_)
);

FILL FILL_3__12824_ (
);

FILL FILL_3__12404_ (
);

FILL FILL_4_CLKBUF1_insert130 (
);

FILL FILL_4_CLKBUF1_insert131 (
);

FILL FILL_2__11817_ (
);

FILL FILL_4_CLKBUF1_insert132 (
);

FILL FILL_0__12851_ (
);

FILL FILL_0__12431_ (
);

FILL FILL_4_CLKBUF1_insert133 (
);

FILL FILL_3__15296_ (
);

FILL FILL_0__12011_ (
);

FILL FILL_4_CLKBUF1_insert134 (
);

FILL FILL_4_CLKBUF1_insert135 (
);

FILL FILL_4_CLKBUF1_insert136 (
);

FILL FILL_1__7099_ (
);

FILL FILL_4_CLKBUF1_insert137 (
);

FILL FILL_4_CLKBUF1_insert138 (
);

FILL FILL_4_CLKBUF1_insert139 (
);

FILL FILL_2__14289_ (
);

FILL FILL_5__15623_ (
);

FILL FILL_5__15203_ (
);

FILL FILL_0__7817_ (
);

OAI21X1 _9923_ (
    .A(_1547_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .C(_1548_),
    .Y(_1498_[25])
);

OAI21X1 _9503_ (
    .A(_1328_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .C(_1329_),
    .Y(_1303_[13])
);

FILL FILL_1__8880_ (
);

FILL FILL_1__8460_ (
);

FILL FILL_4__14616_ (
);

FILL FILL_2__15650_ (
);

FILL FILL_2__15230_ (
);

FILL FILL_3__8386_ (
);

FILL FILL_3__13609_ (
);

FILL FILL_1__14643_ (
);

FILL FILL_1__14223_ (
);

FILL FILL_0__13636_ (
);

OAI22X1 _13921_ (
    .A(_4423_),
    .B(_3967__bF$buf1),
    .C(_3881_),
    .D(_4422_),
    .Y(_4424_)
);

FILL FILL_0__13216_ (
);

OAI22X1 _13501_ (
    .A(_4011_),
    .B(_3902__bF$buf2),
    .C(_3954__bF$buf2),
    .D(_4010_),
    .Y(_4012_)
);

FILL FILL_5__9673_ (
);

FILL FILL_5__9253_ (
);

INVX1 _16393_ (
    .A(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_6816_)
);

FILL FILL_5__16408_ (
);

FILL FILL_5__11963_ (
);

FILL FILL_5__11543_ (
);

FILL FILL_1__9665_ (
);

FILL FILL_1__9245_ (
);

FILL FILL_5__11123_ (
);

FILL FILL_2__16015_ (
);

FILL FILL_4__7670_ (
);

FILL FILL_4__10956_ (
);

FILL FILL_4__7250_ (
);

FILL FILL_4__10536_ (
);

FILL FILL_2__11990_ (
);

FILL FILL_4__10116_ (
);

FILL FILL_2__11570_ (
);

FILL FILL_2__11150_ (
);

FILL FILL_1__15848_ (
);

FILL FILL_6__7596_ (
);

FILL FILL_1__15428_ (
);

FILL FILL_1__15008_ (
);

FILL FILL_1__10983_ (
);

FILL FILL_1__10563_ (
);

FILL FILL_1__10143_ (
);

INVX1 _14706_ (
    .A(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_5192_)
);

FILL FILL_0__7990_ (
);

FILL FILL_2__7588_ (
);

BUFX2 BUFX2_insert770 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf6 )
);

FILL FILL_0__7570_ (
);

FILL FILL_2__7168_ (
);

BUFX2 BUFX2_insert771 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf5 )
);

FILL SFILL29000x4050 (
);

BUFX2 BUFX2_insert772 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf4 )
);

BUFX2 BUFX2_insert773 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf3 )
);

BUFX2 BUFX2_insert774 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf2 )
);

BUFX2 BUFX2_insert775 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf1 )
);

BUFX2 BUFX2_insert776 (
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf0 )
);

BUFX2 BUFX2_insert777 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf7)
);

BUFX2 BUFX2_insert778 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf6)
);

FILL SFILL69160x7050 (
);

BUFX2 BUFX2_insert779 (
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf5)
);

FILL FILL_5__12748_ (
);

FILL FILL_3__13782_ (
);

FILL FILL_5__12328_ (
);

FILL FILL_3__13362_ (
);

FILL FILL_4__8875_ (
);

FILL FILL_4__8455_ (
);

FILL FILL_2__12775_ (
);

FILL FILL_2__12355_ (
);

FILL SFILL99400x26050 (
);

FILL SFILL68520x4050 (
);

FILL FILL_1__11768_ (
);

FILL FILL_1__11348_ (
);

FILL FILL_3__6872_ (
);

FILL FILL_0__8775_ (
);

FILL FILL_5__16161_ (
);

FILL FILL_0__8355_ (
);

FILL FILL112440x70050 (
);

INVX1 _10626_ (
    .A(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_1895_)
);

DFFSR _10206_ (
    .Q(\datapath_1.regfile_1.regOut[26] [8]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_1628_[8])
);

FILL FILL_4__15994_ (
);

FILL FILL_4__15574_ (
);

FILL FILL_4__15154_ (
);

NAND2X1 _13098_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [6]),
    .Y(_3697_)
);

FILL FILL_3__14987_ (
);

FILL FILL_2__9734_ (
);

FILL FILL_3__14567_ (
);

FILL FILL_0__11702_ (
);

FILL FILL_3__14147_ (
);

FILL FILL_1__15181_ (
);

FILL FILL_0__14594_ (
);

FILL SFILL89400x69050 (
);

FILL FILL_0__14174_ (
);

FILL FILL_1__7731_ (
);

FILL FILL_1__7311_ (
);

FILL FILL_2__14921_ (
);

FILL FILL_2__14501_ (
);

FILL FILL_3__7237_ (
);

FILL FILL_5__12081_ (
);

FILL FILL_1__13914_ (
);

FILL FILL_4__16359_ (
);

FILL FILL_4__11494_ (
);

FILL FILL_4__11074_ (
);

FILL FILL_0__12907_ (
);

FILL FILL_1__16386_ (
);

FILL FILL_3__10487_ (
);

FILL FILL_5__8524_ (
);

FILL FILL_5__8104_ (
);

FILL FILL_3__10067_ (
);

FILL FILL_0__15799_ (
);

INVX1 _15664_ (
    .A(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_6129_)
);

FILL FILL_0__15379_ (
);

OAI21X1 _15244_ (
    .A(_5719_),
    .B(_5511_),
    .C(_5459__bF$buf3),
    .Y(_5720_)
);

FILL FILL_5__10814_ (
);

FILL FILL_1__8516_ (
);

FILL SFILL94280x75050 (
);

FILL FILL_6__14293_ (
);

FILL FILL_2__15706_ (
);

FILL FILL_4__6941_ (
);

FILL FILL_0__16320_ (
);

FILL FILL_2__10421_ (
);

FILL FILL_5__13286_ (
);

FILL FILL_2__10001_ (
);

OAI21X1 _7586_ (
    .A(_355_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_356_),
    .Y(_328_[14])
);

OAI21X1 _7166_ (
    .A(_136_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_137_),
    .Y(_133_[2])
);

FILL FILL_4__12699_ (
);

FILL FILL_4__12279_ (
);

FILL FILL_3__9803_ (
);

FILL FILL_0__6841_ (
);

FILL FILL_2__6859_ (
);

FILL FILL_5__9729_ (
);

INVX1 _16449_ (
    .A(BranchNe),
    .Y(_6834_)
);

FILL FILL_4__13640_ (
);

FILL FILL_4__13220_ (
);

NAND3X1 _16029_ (
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf4),
    .Y(_6485_)
);

FILL FILL_0__11299_ (
);

INVX1 _11584_ (
    .A(_2272_),
    .Y(_2691_)
);

AOI21X1 _11164_ (
    .A(_2226_),
    .B(_2278_),
    .C(_2282_),
    .Y(_2283_)
);

FILL FILL_2__7800_ (
);

FILL FILL_3__12633_ (
);

FILL FILL_3__12213_ (
);

FILL FILL_4__7726_ (
);

FILL FILL_4__7306_ (
);

FILL FILL_2__11626_ (
);

FILL FILL_0__12660_ (
);

FILL FILL_2__11206_ (
);

FILL FILL_0__12240_ (
);

FILL SFILL39240x78050 (
);

FILL FILL_1__10619_ (
);

FILL FILL_2__14098_ (
);

FILL FILL_5__15852_ (
);

FILL FILL_5__15432_ (
);

FILL FILL_0__7626_ (
);

FILL FILL_5__15012_ (
);

OAI21X1 _9732_ (
    .A(_1440_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1441_),
    .Y(_1433_[4])
);

FILL FILL_0__7206_ (
);

DFFSR _9312_ (
    .Q(\datapath_1.regfile_1.regOut[19] [10]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_1173_[10])
);

FILL SFILL33960x26050 (
);

FILL FILL_4__14845_ (
);

FILL FILL_4__14425_ (
);

FILL FILL_4__14005_ (
);

NAND2X1 _12789_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[31]),
    .Y(_3552_)
);

FILL FILL_3__8195_ (
);

OAI21X1 _12369_ (
    .A(_3310_),
    .B(MemToReg_bF$buf2),
    .C(_3311_),
    .Y(\datapath_1.mux_wd3.dout [8])
);

FILL FILL_3__13838_ (
);

FILL FILL_1__14872_ (
);

FILL FILL_3__13418_ (
);

FILL FILL_1__14452_ (
);

FILL FILL_1__14032_ (
);

FILL SFILL84280x73050 (
);

FILL FILL_0__13865_ (
);

FILL FILL_0__13445_ (
);

OAI22X1 _13730_ (
    .A(_4235_),
    .B(_3905__bF$buf3),
    .C(_3977__bF$buf2),
    .D(_4236_),
    .Y(_4237_)
);

NOR2X1 _13310_ (
    .A(_3789_),
    .B(_3812_),
    .Y(_3843_)
);

FILL FILL_0__13025_ (
);

FILL FILL_5__9482_ (
);

FILL FILL_3__6928_ (
);

FILL FILL_5__16217_ (
);

FILL FILL_1__9894_ (
);

FILL FILL_5__11772_ (
);

FILL FILL_1__9474_ (
);

FILL FILL_5__11352_ (
);

FILL SFILL79320x29050 (
);

FILL FILL_2__16244_ (
);

FILL FILL_4__10765_ (
);

FILL FILL_1__15657_ (
);

FILL FILL_1__15237_ (
);

FILL FILL_1__10792_ (
);

FILL FILL_1__10372_ (
);

INVX1 _14935_ (
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_5416_)
);

OAI22X1 _14515_ (
    .A(_5004_),
    .B(_3936__bF$buf0),
    .C(_3930__bF$buf1),
    .D(_5003_),
    .Y(_5005_)
);

FILL SFILL109480x71050 (
);

FILL FILL_5__12977_ (
);

FILL FILL_3__13591_ (
);

FILL FILL_5__12137_ (
);

BUFX2 _6857_ (
    .A(_1_[19]),
    .Y(memoryAddress[19])
);

FILL FILL_3__13171_ (
);

FILL FILL_4__8264_ (
);

FILL FILL_2__12584_ (
);

FILL SFILL114440x54050 (
);

FILL FILL_2__12164_ (
);

FILL FILL_1__11997_ (
);

FILL FILL_1__11577_ (
);

FILL FILL_1__11157_ (
);

FILL FILL_4__12911_ (
);

FILL FILL_5__16390_ (
);

FILL FILL_0__8584_ (
);

DFFSR _10855_ (
    .Q(\datapath_1.regfile_1.regOut[31] [17]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_1953_[17])
);

FILL FILL_6__9131_ (
);

OAI21X1 _10435_ (
    .A(_1807_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1808_),
    .Y(_1758_[25])
);

OAI21X1 _10015_ (
    .A(_1588_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .C(_1589_),
    .Y(_1563_[13])
);

FILL FILL_3__11904_ (
);

FILL FILL_6__14769_ (
);

FILL FILL_6__14349_ (
);

FILL FILL_4__15383_ (
);

FILL FILL_3__14796_ (
);

FILL FILL_0__11931_ (
);

FILL FILL_2__9543_ (
);

FILL FILL_2__9123_ (
);

FILL FILL_3__14376_ (
);

FILL FILL_0__11511_ (
);

FILL FILL_6__15710_ (
);

FILL FILL_4__9889_ (
);

FILL FILL_4__9469_ (
);

FILL FILL_2__13789_ (
);

FILL FILL_2__13369_ (
);

FILL FILL_5__14703_ (
);

FILL FILL_1__7960_ (
);

FILL FILL_1__7120_ (
);

FILL FILL_2__14730_ (
);

FILL FILL_0__9789_ (
);

FILL FILL_3__7886_ (
);

FILL FILL_2__14310_ (
);

FILL FILL_0__9369_ (
);

FILL FILL_3__7466_ (
);

FILL SFILL29160x38050 (
);

FILL FILL_3__7046_ (
);

FILL FILL_1__13723_ (
);

FILL FILL_1__13303_ (
);

FILL FILL_4__16168_ (
);

FILL FILL_6__10269_ (
);

FILL FILL_0__12716_ (
);

FILL FILL_1__16195_ (
);

FILL FILL_5__8753_ (
);

FILL FILL_5__8333_ (
);

FILL FILL_3__10296_ (
);

NOR2X1 _15893_ (
    .A(_4986_),
    .B(_5549__bF$buf4),
    .Y(_6352_)
);

FILL FILL_6__11630_ (
);

FILL FILL_0__15188_ (
);

NOR2X1 _15473_ (
    .A(_5942_),
    .B(_5936_),
    .Y(_5943_)
);

FILL FILL_5__15908_ (
);

OAI22X1 _15053_ (
    .A(_5530__bF$buf3),
    .B(_3915_),
    .C(_5532__bF$buf0),
    .D(_3914_),
    .Y(_5533_)
);

FILL FILL_3__16102_ (
);

FILL FILL_5__10623_ (
);

FILL FILL_1__8745_ (
);

FILL FILL_1__8325_ (
);

FILL FILL_2__15935_ (
);

FILL FILL_2__15515_ (
);

FILL FILL_2__10650_ (
);

FILL FILL_2__10230_ (
);

FILL FILL_5__13095_ (
);

FILL FILL_1__14928_ (
);

FILL FILL_1__14508_ (
);

DFFSR _7395_ (
    .Q(\datapath_1.regfile_1.regOut[4] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf55),
    .S(vdd),
    .D(_198_[13])
);

FILL FILL_4__12088_ (
);

FILL FILL_3__9612_ (
);

FILL SFILL104360x59050 (
);

FILL FILL_5__9538_ (
);

FILL FILL_5__9118_ (
);

NAND3X1 _16258_ (
    .A(_6702_),
    .B(_6703_),
    .C(_6707_),
    .Y(_6708_)
);

INVX1 _11393_ (
    .A(_2201_),
    .Y(_2510_)
);

FILL FILL_5__11828_ (
);

FILL FILL_3__12862_ (
);

FILL FILL_5__11408_ (
);

FILL FILL_3__12442_ (
);

FILL FILL_3__12022_ (
);

FILL FILL_4__7955_ (
);

FILL FILL_4__7115_ (
);

FILL FILL_2__11855_ (
);

FILL FILL_2__11435_ (
);

FILL FILL_2__11015_ (
);

FILL FILL_1__10428_ (
);

FILL FILL_1__10008_ (
);

FILL FILL_5__15661_ (
);

FILL FILL_5__15241_ (
);

FILL FILL_0__7855_ (
);

FILL FILL112440x65050 (
);

FILL FILL_0__7435_ (
);

DFFSR _9961_ (
    .Q(\datapath_1.regfile_1.regOut[24] [19]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_1498_[19])
);

NAND2X1 _9541_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1355_)
);

FILL FILL_6__8402_ (
);

NAND2X1 _9121_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1136_)
);

FILL SFILL104360x14050 (
);

FILL FILL_4__14654_ (
);

FILL FILL_4__14234_ (
);

NAND2X1 _12598_ (
    .A(vdd),
    .B(memoryOutData[10]),
    .Y(_3445_)
);

INVX1 _12178_ (
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3172_)
);

FILL FILL_3__13647_ (
);

FILL FILL_3__13227_ (
);

FILL FILL_1__14681_ (
);

FILL FILL_1__14261_ (
);

FILL FILL112040x51050 (
);

FILL FILL_0_BUFX2_insert410 (
);

FILL FILL_0_BUFX2_insert411 (
);

FILL FILL_0_BUFX2_insert412 (
);

FILL FILL_0_BUFX2_insert413 (
);

FILL FILL_0__13674_ (
);

FILL FILL_0_BUFX2_insert414 (
);

FILL FILL_0__13254_ (
);

FILL FILL_0_BUFX2_insert415 (
);

FILL FILL_0_BUFX2_insert416 (
);

FILL FILL_0_BUFX2_insert417 (
);

FILL FILL_0_BUFX2_insert418 (
);

FILL FILL_5__9291_ (
);

FILL FILL_0_BUFX2_insert419 (
);

FILL FILL_5__16026_ (
);

FILL FILL_6__9607_ (
);

FILL FILL_5__11581_ (
);

FILL FILL_5__11161_ (
);

FILL FILL_1__9283_ (
);

FILL FILL_4__15859_ (
);

FILL FILL112440x20050 (
);

FILL FILL_4__15439_ (
);

FILL FILL_4__15019_ (
);

FILL FILL_2__16053_ (
);

FILL FILL_4__10994_ (
);

FILL FILL_4__10574_ (
);

FILL FILL_4__10154_ (
);

FILL FILL_1__15886_ (
);

FILL FILL_1__15466_ (
);

FILL FILL_1__15046_ (
);

FILL FILL_5__7604_ (
);

FILL FILL_1__10181_ (
);

FILL FILL_0__14879_ (
);

FILL FILL_0__14459_ (
);

NOR2X1 _14744_ (
    .A(_5228_),
    .B(_3977__bF$buf2),
    .Y(_5229_)
);

FILL FILL_0__14039_ (
);

AOI22X1 _14324_ (
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .B(_4005__bF$buf1),
    .C(_3995__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_4818_)
);

FILL FILL_0__15820_ (
);

FILL FILL_0__15400_ (
);

FILL FILL_5__12786_ (
);

FILL FILL_5__12366_ (
);

FILL FILL_4__8493_ (
);

FILL FILL_4__8073_ (
);

FILL FILL_4__11779_ (
);

FILL FILL_4__11359_ (
);

FILL FILL_2__12393_ (
);

FILL SFILL23720x81050 (
);

FILL FILL_1__11386_ (
);

NOR2X1 _15949_ (
    .A(_6404_),
    .B(_6406_),
    .Y(_6407_)
);

FILL FILL_4__12720_ (
);

INVX1 _15529_ (
    .A(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_5998_)
);

FILL FILL_4__12300_ (
);

NOR2X1 _15109_ (
    .A(_5587_),
    .B(_5585_),
    .Y(_5588_)
);

FILL FILL_0__10799_ (
);

FILL FILL_0__8393_ (
);

FILL FILL_0__10379_ (
);

OAI21X1 _10664_ (
    .A(_1919_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1920_),
    .Y(_1888_[16])
);

OAI21X1 _10244_ (
    .A(_1700_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .C(_1701_),
    .Y(_1693_[4])
);

FILL FILL_3__11713_ (
);

FILL FILL_4__15192_ (
);

FILL SFILL58440x80050 (
);

FILL SFILL94280x25050 (
);

FILL FILL_2__9772_ (
);

FILL FILL_2__10706_ (
);

FILL FILL_2__9352_ (
);

FILL FILL_0__11740_ (
);

FILL FILL_3__14185_ (
);

FILL FILL_0__11320_ (
);

FILL FILL_4_BUFX2_insert990 (
);

FILL FILL_4_BUFX2_insert991 (
);

FILL FILL_4__9278_ (
);

FILL FILL_4_BUFX2_insert992 (
);

FILL FILL_4_BUFX2_insert993 (
);

FILL FILL_4_BUFX2_insert994 (
);

FILL FILL_2__13598_ (
);

FILL FILL_4_BUFX2_insert995 (
);

FILL FILL_4_BUFX2_insert996 (
);

FILL FILL_4_BUFX2_insert997 (
);

FILL FILL_5__14932_ (
);

FILL FILL_4_BUFX2_insert998 (
);

FILL FILL_5__14512_ (
);

FILL FILL_4_BUFX2_insert999 (
);

DFFSR _8812_ (
    .Q(\datapath_1.regfile_1.regOut[15] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_913_[22])
);

FILL FILL_4__13925_ (
);

FILL FILL_4__13505_ (
);

FILL FILL_3__7695_ (
);

FILL FILL_0__9598_ (
);

NOR2X1 _11869_ (
    .A(\datapath_1.ALUResult [27]),
    .B(\datapath_1.ALUResult [23]),
    .Y(_2956_)
);

OAI21X1 _11449_ (
    .A(_2563_),
    .B(_2375_),
    .C(_2564_),
    .Y(_2565_)
);

XNOR2X1 _11029_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2148_)
);

FILL FILL_3__12918_ (
);

FILL FILL_1__13952_ (
);

FILL FILL_1__13532_ (
);

FILL FILL_4__16397_ (
);

FILL SFILL98920x45050 (
);

FILL FILL_1__13112_ (
);

FILL SFILL94200x23050 (
);

DFFSR _12810_ (
    .Q(\datapath_1.PCJump [21]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3490_[19])
);

FILL FILL_0__12525_ (
);

FILL FILL_0__12105_ (
);

FILL FILL_5__8982_ (
);

FILL FILL_6__16304_ (
);

FILL FILL_5__8142_ (
);

OAI21X1 _15282_ (
    .A(_4235_),
    .B(_5535__bF$buf1),
    .C(_5756_),
    .Y(_5757_)
);

FILL FILL_5__15717_ (
);

FILL FILL_3__16331_ (
);

FILL FILL_1__8974_ (
);

FILL FILL_5__10432_ (
);

FILL FILL_5__10012_ (
);

FILL FILL_1__8134_ (
);

FILL FILL_2__15744_ (
);

FILL FILL_2__15324_ (
);

FILL FILL_1__14737_ (
);

FILL FILL_1__14317_ (
);

FILL SFILL84200x66050 (
);

FILL FILL_3__9421_ (
);

FILL FILL_3__9001_ (
);

FILL FILL_2__6897_ (
);

FILL FILL_5__9767_ (
);

FILL FILL_5__9347_ (
);

FILL FILL_6__12644_ (
);

FILL FILL_6__12224_ (
);

NOR2X1 _16067_ (
    .A(_6521_),
    .B(_6514_),
    .Y(_6522_)
);

FILL FILL_1__9759_ (
);

FILL FILL_5__11637_ (
);

FILL FILL_5__11217_ (
);

FILL FILL_1__9339_ (
);

FILL FILL_3__12251_ (
);

FILL SFILL8600x40050 (
);

FILL FILL_4__7764_ (
);

FILL FILL_2__16109_ (
);

FILL FILL_4__7344_ (
);

FILL FILL_2__11664_ (
);

FILL FILL_2__11244_ (
);

FILL FILL_1__10657_ (
);

FILL FILL_1__10237_ (
);

FILL FILL_5__15890_ (
);

FILL SFILL84200x21050 (
);

FILL FILL_5__15470_ (
);

FILL FILL_5__15050_ (
);

NAND2X1 _9770_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1467_)
);

FILL FILL_0__7244_ (
);

NAND2X1 _9350_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1248_)
);

FILL FILL_6__8211_ (
);

FILL FILL_4__14883_ (
);

FILL FILL_4__14463_ (
);

FILL FILL_4__14043_ (
);

FILL SFILL13160x79050 (
);

FILL FILL_3__13876_ (
);

FILL FILL_2__8623_ (
);

FILL FILL_2__8203_ (
);

FILL FILL_3__13456_ (
);

FILL FILL_1__14490_ (
);

FILL FILL_3__13036_ (
);

FILL FILL_1__14070_ (
);

FILL FILL_4__8969_ (
);

FILL FILL_4__8129_ (
);

FILL FILL_2__12869_ (
);

FILL FILL_2__12449_ (
);

FILL FILL_2__12029_ (
);

FILL FILL_0__13483_ (
);

FILL FILL_4__9910_ (
);

FILL FILL_2__13810_ (
);

FILL SFILL74200x64050 (
);

FILL FILL_0__8869_ (
);

FILL FILL_3__6966_ (
);

FILL FILL_5__16255_ (
);

FILL FILL_0__8449_ (
);

FILL FILL_5__11390_ (
);

FILL FILL_1__9092_ (
);

FILL SFILL74280x21050 (
);

FILL FILL_4__15668_ (
);

FILL FILL_4__15248_ (
);

FILL FILL_2__16282_ (
);

FILL FILL_4__10383_ (
);

FILL FILL_0__9810_ (
);

FILL FILL_2__9408_ (
);

FILL FILL_1__15695_ (
);

FILL FILL_1__15275_ (
);

FILL SFILL99480x70050 (
);

FILL FILL_5__7833_ (
);

INVX1 _14973_ (
    .A(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_5454_)
);

FILL FILL_0__14688_ (
);

INVX1 _14553_ (
    .A(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_5042_)
);

FILL FILL_0__14268_ (
);

NAND3X1 _14133_ (
    .A(_4628_),
    .B(_4630_),
    .C(_4627_),
    .Y(_4631_)
);

FILL FILL_3__15602_ (
);

FILL FILL_1__7825_ (
);

FILL FILL_5__12595_ (
);

FILL FILL_5__12175_ (
);

BUFX2 _6895_ (
    .A(_2_[25]),
    .Y(memoryWriteData[25])
);

FILL FILL_4__11588_ (
);

FILL FILL_4__11168_ (
);

FILL FILL_5__8618_ (
);

FILL FILL_1__11195_ (
);

NAND2X1 _15758_ (
    .A(_6216_),
    .B(_6220_),
    .Y(_6221_)
);

AOI21X1 _15338_ (
    .A(_5784_),
    .B(_5811_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [6])
);

INVX1 _10893_ (
    .A(\aluControl_1.inst [2]),
    .Y(_2039_)
);

FILL FILL_0__10188_ (
);

DFFSR _10473_ (
    .Q(\datapath_1.regfile_1.regOut[28] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_1758_[19])
);

FILL FILL_5__10908_ (
);

NAND2X1 _10053_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1615_)
);

FILL FILL_3__11942_ (
);

FILL FILL_3__11522_ (
);

FILL FILL_3__11102_ (
);

FILL FILL_0__16414_ (
);

FILL FILL_2__10935_ (
);

FILL FILL_2__10515_ (
);

FILL SFILL33800x71050 (
);

FILL FILL_2__9161_ (
);

FILL FILL_4__9087_ (
);

FILL FILL_5__14741_ (
);

FILL FILL_0__6935_ (
);

FILL FILL_5__14321_ (
);

NAND2X1 _8621_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_884_)
);

NAND2X1 _8201_ (
    .A(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_665_)
);

FILL FILL_4__13734_ (
);

FILL FILL_4__13314_ (
);

FILL FILL_3__7084_ (
);

OR2X2 _11678_ (
    .A(_2778_),
    .B(_2164_),
    .Y(_2779_)
);

NAND2X1 _11258_ (
    .A(_2161_),
    .B(_2162_),
    .Y(_2377_)
);

FILL FILL_3__12727_ (
);

FILL SFILL89720x5050 (
);

FILL FILL_1__13761_ (
);

FILL FILL_3__12307_ (
);

FILL FILL_1__13341_ (
);

FILL FILL112040x46050 (
);

FILL FILL_0__12754_ (
);

FILL FILL_3__15199_ (
);

FILL FILL_0__12334_ (
);

FILL FILL_5__8371_ (
);

FILL FILL_5__15946_ (
);

INVX8 _15091_ (
    .A(_5569_),
    .Y(_5570_)
);

FILL FILL_5__15526_ (
);

FILL FILL_5__15106_ (
);

DFFSR _9826_ (
    .Q(\datapath_1.regfile_1.regOut[23] [12]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_1433_[12])
);

FILL FILL_3__16140_ (
);

INVX1 _9406_ (
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_1285_)
);

FILL FILL_5__10661_ (
);

FILL FILL_1__8783_ (
);

FILL FILL_5__10241_ (
);

FILL FILL_1__8363_ (
);

FILL FILL112440x15050 (
);

FILL FILL_4__14939_ (
);

FILL FILL_2__15973_ (
);

FILL FILL_4__14519_ (
);

FILL FILL_2__15553_ (
);

FILL FILL_2__15133_ (
);

FILL FILL_1__14966_ (
);

FILL FILL_1__14546_ (
);

FILL FILL_1__14126_ (
);

FILL SFILL85080x22050 (
);

FILL FILL_3__9650_ (
);

FILL FILL_0__13959_ (
);

FILL FILL_3__9230_ (
);

OAI22X1 _13824_ (
    .A(_4327_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf3),
    .D(_4328_),
    .Y(_4329_)
);

FILL FILL_0__13539_ (
);

NAND3X1 _13404_ (
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3903_),
    .C(_3888_),
    .Y(_3916_)
);

FILL FILL_0__13119_ (
);

FILL FILL_5__9996_ (
);

FILL FILL_5__9156_ (
);

FILL SFILL54200x60050 (
);

NOR3X1 _16296_ (
    .A(_6739_),
    .B(_6735_),
    .C(_6744_),
    .Y(_6745_)
);

FILL FILL_0__14900_ (
);

FILL FILL_1__9988_ (
);

FILL FILL_5__11866_ (
);

FILL FILL_5__11446_ (
);

FILL FILL_1__9148_ (
);

FILL FILL_3__12480_ (
);

FILL FILL_5__11026_ (
);

FILL FILL_3__12060_ (
);

FILL FILL_4__7993_ (
);

FILL FILL_2__16338_ (
);

FILL FILL_4__7573_ (
);

FILL FILL_2__11893_ (
);

FILL FILL_4__10439_ (
);

FILL FILL_4__10019_ (
);

FILL FILL_2__11473_ (
);

FILL FILL_2__11053_ (
);

FILL FILL_6__7079_ (
);

FILL SFILL23720x76050 (
);

FILL FILL_1__10886_ (
);

FILL FILL_1__10046_ (
);

AOI22X1 _14609_ (
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .B(_3942__bF$buf1),
    .C(_3995__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_5097_)
);

FILL FILL_4__11800_ (
);

FILL FILL_0__7893_ (
);

FILL FILL_0__7473_ (
);

FILL FILL_0__7053_ (
);

FILL FILL_4__14692_ (
);

FILL FILL_4__14272_ (
);

FILL SFILL23320x62050 (
);

FILL FILL_2__8852_ (
);

FILL FILL_3__13685_ (
);

FILL FILL_0__10820_ (
);

FILL FILL_3__13265_ (
);

FILL FILL_2__8012_ (
);

FILL FILL_0__10400_ (
);

FILL FILL_4__8778_ (
);

FILL FILL_4__8358_ (
);

FILL FILL_2__12258_ (
);

FILL FILL_0__13292_ (
);

FILL FILL_5__16064_ (
);

OAI21X1 _10949_ (
    .A(_2074_),
    .B(_2075_),
    .C(_2081_),
    .Y(_2082_)
);

FILL FILL_0__8258_ (
);

NAND2X1 _10529_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1851_)
);

NAND2X1 _10109_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1632_)
);

FILL FILL_4__15897_ (
);

FILL FILL_1__12612_ (
);

FILL FILL_4__15477_ (
);

FILL FILL_4__15057_ (
);

FILL FILL_2__16091_ (
);

FILL FILL_4__10192_ (
);

FILL FILL_2__9637_ (
);

FILL FILL_2__9217_ (
);

FILL FILL_0__11605_ (
);

FILL FILL_1__15084_ (
);

FILL FILL_5__7222_ (
);

FILL SFILL23640x38050 (
);

FILL FILL_0__14497_ (
);

NOR2X1 _14782_ (
    .A(_5266_),
    .B(_5263_),
    .Y(_5267_)
);

OAI22X1 _14362_ (
    .A(_4854_),
    .B(_3890_),
    .C(_3955__bF$buf4),
    .D(_4853_),
    .Y(_4855_)
);

FILL FILL_0__14077_ (
);

FILL FILL_3__15831_ (
);

FILL FILL_3__15411_ (
);

FILL FILL_1__7634_ (
);

FILL SFILL99880x7050 (
);

FILL FILL_1__7214_ (
);

FILL SFILL8680x37050 (
);

FILL SFILL13720x74050 (
);

FILL FILL_2__14824_ (
);

FILL SFILL44120x65050 (
);

FILL FILL_2__14404_ (
);

FILL FILL_1__13817_ (
);

FILL FILL_4__11397_ (
);

FILL SFILL99480x6050 (
);

FILL FILL_3__8501_ (
);

FILL SFILL84280x18050 (
);

FILL FILL_1__16289_ (
);

FILL FILL_5__8847_ (
);

FILL FILL_5__8007_ (
);

OAI22X1 _15987_ (
    .A(_5499__bF$buf2),
    .B(_5043_),
    .C(_5532__bF$buf3),
    .D(_5039_),
    .Y(_6444_)
);

NAND3X1 _15567_ (
    .A(\datapath_1.PCJump [24]),
    .B(_5460_),
    .C(_5462_),
    .Y(_6035_)
);

OAI21X1 _15147_ (
    .A(_5524__bF$buf2),
    .B(_4086_),
    .C(_5624_),
    .Y(_5625_)
);

NAND2X1 _10282_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1727_)
);

FILL FILL_1__8839_ (
);

FILL FILL_3__11751_ (
);

FILL SFILL8600x35050 (
);

FILL FILL_6__14196_ (
);

FILL FILL_3__11331_ (
);

FILL FILL_2__15609_ (
);

FILL FILL_4__6844_ (
);

FILL FILL_0__16223_ (
);

FILL FILL_2__10744_ (
);

FILL FILL_2__9390_ (
);

FILL FILL_2__10324_ (
);

INVX1 _7489_ (
    .A(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_312_)
);

INVX1 _7069_ (
    .A(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_93_)
);

FILL SFILL84200x16050 (
);

FILL FILL_5__14970_ (
);

FILL FILL_5__14550_ (
);

FILL FILL_5__14130_ (
);

NAND2X1 _8850_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_996_)
);

DFFSR _8430_ (
    .Q(\datapath_1.regfile_1.regOut[12] [24]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_718_[24])
);

INVX1 _8010_ (
    .A(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_578_)
);

FILL FILL_4__13963_ (
);

FILL FILL_4__13543_ (
);

FILL FILL_4__13123_ (
);

FILL SFILL13640x36050 (
);

NAND3X1 _11487_ (
    .A(_2470__bF$buf3),
    .B(_2587_),
    .C(_2600_),
    .Y(_2601_)
);

OAI21X1 _11067_ (
    .A(_2184_),
    .B(_2185_),
    .C(_2181_),
    .Y(_2186_)
);

FILL FILL_2__7703_ (
);

FILL FILL_3__12956_ (
);

FILL FILL_1__13990_ (
);

FILL SFILL109480x16050 (
);

FILL FILL_3__12116_ (
);

FILL FILL_1__13570_ (
);

FILL FILL_1__13150_ (
);

FILL FILL_4__7629_ (
);

FILL FILL_4__7209_ (
);

FILL FILL_2__11949_ (
);

FILL FILL_0__12983_ (
);

FILL FILL_2__11529_ (
);

FILL FILL_2__11109_ (
);

FILL FILL_0__12143_ (
);

FILL SFILL78600x60050 (
);

FILL SFILL74200x59050 (
);

FILL FILL_5__15755_ (
);

FILL FILL_0__7949_ (
);

FILL FILL_5__15335_ (
);

INVX1 _9635_ (
    .A(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_1397_)
);

FILL FILL_0__7109_ (
);

INVX1 _9215_ (
    .A(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_1178_)
);

FILL FILL_5__10890_ (
);

FILL FILL_1__8592_ (
);

FILL SFILL74280x16050 (
);

FILL FILL_5__10050_ (
);

FILL FILL_4__14748_ (
);

FILL FILL_2__15782_ (
);

FILL FILL_4__14328_ (
);

FILL FILL_2__15362_ (
);

FILL FILL_3__8098_ (
);

FILL FILL_2__8908_ (
);

FILL FILL_1__14775_ (
);

FILL SFILL99480x65050 (
);

FILL FILL_1__14355_ (
);

FILL FILL_5__6913_ (
);

FILL FILL_0__13768_ (
);

FILL FILL_0__13348_ (
);

OAI22X1 _13633_ (
    .A(_4141_),
    .B(_3971__bF$buf4),
    .C(_3924__bF$buf3),
    .D(_4140_),
    .Y(_4142_)
);

INVX2 _13213_ (
    .A(_3755_),
    .Y(_3756_)
);

FILL FILL_5__9385_ (
);

FILL FILL_1__6905_ (
);

FILL FILL_1__9797_ (
);

FILL FILL_5__11675_ (
);

FILL SFILL74200x14050 (
);

FILL FILL_1__9377_ (
);

FILL FILL_5__11255_ (
);

FILL FILL_2__16147_ (
);

FILL FILL_4__10668_ (
);

FILL FILL_4__10248_ (
);

FILL FILL_2__11282_ (
);

FILL FILL_2_BUFX2_insert320 (
);

FILL FILL_1__10695_ (
);

FILL FILL_1__10275_ (
);

FILL FILL_2_BUFX2_insert321 (
);

FILL SFILL99480x20050 (
);

FILL FILL_2_BUFX2_insert322 (
);

AOI21X1 _14838_ (
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .B(_4115_),
    .C(_5320_),
    .Y(_5321_)
);

FILL FILL_2_BUFX2_insert323 (
);

FILL FILL_2_BUFX2_insert324 (
);

INVX1 _14418_ (
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_4910_)
);

FILL FILL_2_BUFX2_insert325 (
);

FILL FILL_2_BUFX2_insert326 (
);

FILL FILL_2_BUFX2_insert327 (
);

FILL SFILL28840x83050 (
);

FILL FILL_2_BUFX2_insert328 (
);

FILL FILL_2_BUFX2_insert329 (
);

FILL FILL_4__14081_ (
);

FILL FILL_0__15914_ (
);

FILL SFILL68920x79050 (
);

FILL FILL_2__8661_ (
);

FILL SFILL64200x57050 (
);

FILL FILL_3__13494_ (
);

FILL FILL_2__8241_ (
);

FILL FILL112120x34050 (
);

FILL FILL_4__8587_ (
);

FILL FILL_2__12487_ (
);

FILL FILL_2__12067_ (
);

FILL FILL_5__13821_ (
);

FILL FILL_5__13401_ (
);

FILL FILL_2_BUFX2_insert1040 (
);

FILL FILL_2_BUFX2_insert1041 (
);

FILL FILL_2_BUFX2_insert1042 (
);

NAND2X1 _7701_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_413_)
);

FILL FILL_2_BUFX2_insert1043 (
);

FILL FILL_2_BUFX2_insert1044 (
);

FILL FILL_2_BUFX2_insert1045 (
);

FILL FILL_2_BUFX2_insert1046 (
);

FILL FILL_2_BUFX2_insert1047 (
);

FILL FILL_2_BUFX2_insert1048 (
);

FILL FILL_5__16293_ (
);

FILL FILL_0__8487_ (
);

FILL FILL_2_BUFX2_insert1049 (
);

FILL FILL_0__8067_ (
);

NAND2X1 _10758_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1963_)
);

DFFSR _10338_ (
    .Q(\datapath_1.regfile_1.regOut[27] [12]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_1693_[12])
);

FILL FILL_3__11807_ (
);

FILL FILL_1__12841_ (
);

FILL FILL_1__12421_ (
);

FILL FILL_4__15286_ (
);

FILL FILL_1__12001_ (
);

FILL FILL_2__9866_ (
);

FILL FILL_3__14699_ (
);

FILL FILL_0__11834_ (
);

FILL FILL_3__14279_ (
);

FILL FILL_0__11414_ (
);

FILL FILL_2__9026_ (
);

FILL FILL_5__7871_ (
);

FILL FILL_6__15613_ (
);

FILL SFILL33800x21050 (
);

FILL FILL_5__7451_ (
);

FILL FILL_5__7031_ (
);

INVX1 _14591_ (
    .A(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_5080_)
);

AOI21X1 _14171_ (
    .A(_4668_),
    .B(_4642_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [14])
);

FILL FILL_5__14606_ (
);

FILL FILL_3__15640_ (
);

INVX1 _8906_ (
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_1033_)
);

FILL FILL_3__15220_ (
);

FILL FILL_1__7863_ (
);

FILL FILL_1__7443_ (
);

FILL FILL_2__14633_ (
);

FILL FILL_2__14213_ (
);

FILL FILL_3__7369_ (
);

FILL FILL_1__13626_ (
);

FILL SFILL18840x81050 (
);

FILL FILL_1_BUFX2_insert340 (
);

FILL FILL_1_BUFX2_insert341 (
);

FILL FILL_3__8730_ (
);

FILL FILL_0__12619_ (
);

FILL FILL_3__8310_ (
);

INVX1 _12904_ (
    .A(\datapath_1.a [27]),
    .Y(_3608_)
);

FILL FILL_1_BUFX2_insert342 (
);

FILL FILL_1_BUFX2_insert343 (
);

FILL FILL_1__16098_ (
);

FILL FILL_1_BUFX2_insert344 (
);

FILL FILL_1_BUFX2_insert345 (
);

FILL SFILL58920x77050 (
);

FILL FILL_1_BUFX2_insert346 (
);

FILL FILL_5__8656_ (
);

FILL FILL_5__8236_ (
);

FILL FILL_1_BUFX2_insert347 (
);

FILL FILL_1_BUFX2_insert348 (
);

FILL FILL_1_BUFX2_insert349 (
);

INVX1 _15796_ (
    .A(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_6258_)
);

FILL FILL_6__11533_ (
);

NOR2X1 _15376_ (
    .A(_4370_),
    .B(_5534__bF$buf4),
    .Y(_5848_)
);

FILL FILL_6__11113_ (
);

FILL FILL_3__16005_ (
);

DFFSR _10091_ (
    .Q(\datapath_1.regfile_1.regOut[25] [21]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_1563_[21])
);

FILL FILL_5__10946_ (
);

FILL FILL_3__11980_ (
);

FILL FILL_1__8648_ (
);

FILL FILL_5__10526_ (
);

FILL FILL_1__8228_ (
);

FILL FILL_3__11560_ (
);

FILL FILL_5__10106_ (
);

FILL FILL_3__11140_ (
);

FILL FILL_2__15838_ (
);

FILL FILL_2__15418_ (
);

FILL FILL_0__16032_ (
);

FILL FILL_2__10973_ (
);

FILL FILL_2__10553_ (
);

FILL FILL_2__10133_ (
);

INVX1 _7298_ (
    .A(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_205_)
);

FILL SFILL105320x79050 (
);

FILL FILL_3__9935_ (
);

FILL FILL_3__9515_ (
);

FILL FILL_0__6973_ (
);

FILL FILL_6__12738_ (
);

FILL FILL_4__13772_ (
);

FILL FILL_4__13352_ (
);

NAND2X1 _11296_ (
    .A(_2412_),
    .B(_2414_),
    .Y(_2415_)
);

FILL FILL_2__7932_ (
);

FILL FILL_3__12765_ (
);

FILL FILL_3__12345_ (
);

FILL FILL_4__7858_ (
);

FILL FILL_4__7438_ (
);

FILL FILL_2__11758_ (
);

FILL FILL_2__11338_ (
);

FILL FILL_0__12372_ (
);

FILL SFILL74120x5050 (
);

FILL FILL_5__15984_ (
);

FILL FILL_5__15564_ (
);

FILL FILL_0__7758_ (
);

FILL FILL_5__15144_ (
);

FILL SFILL38840x1050 (
);

INVX1 _9864_ (
    .A(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_1509_)
);

FILL FILL_0__7338_ (
);

DFFSR _9444_ (
    .Q(\datapath_1.regfile_1.regOut[20] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_1238_[14])
);

OAI21X1 _9024_ (
    .A(_1090_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .C(_1091_),
    .Y(_1043_[24])
);

FILL FILL_4__14977_ (
);

FILL FILL_4__14557_ (
);

FILL SFILL48920x75050 (
);

FILL FILL_4__14137_ (
);

FILL FILL_2__15591_ (
);

FILL FILL_2__15171_ (
);

FILL SFILL109640x42050 (
);

FILL FILL_2__8717_ (
);

FILL FILL_1__14584_ (
);

FILL FILL_1__14164_ (
);

FILL FILL_0__13997_ (
);

NAND3X1 _13862_ (
    .A(_4357_),
    .B(_4358_),
    .C(_4365_),
    .Y(_4366_)
);

FILL FILL_0__13577_ (
);

NAND3X1 _13442_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3888_),
    .C(_3879_),
    .Y(_3954_)
);

FILL FILL_0__13157_ (
);

OAI21X1 _13022_ (
    .A(_3665_),
    .B(vdd),
    .C(_3666_),
    .Y(_3620_[23])
);

FILL FILL_3__14911_ (
);

FILL SFILL13720x69050 (
);

FILL FILL_2__13904_ (
);

FILL FILL_5__16349_ (
);

FILL SFILL109560x49050 (
);

FILL FILL_5__11484_ (
);

FILL FILL_5__11064_ (
);

FILL FILL_2__16376_ (
);

FILL FILL_4__10897_ (
);

FILL FILL_4__7191_ (
);

FILL FILL_0__9904_ (
);

FILL FILL_4__10057_ (
);

FILL SFILL48920x30050 (
);

FILL FILL_2__11091_ (
);

FILL FILL_1__15789_ (
);

FILL FILL_1__15369_ (
);

FILL FILL_5__7927_ (
);

FILL FILL_5__7507_ (
);

AOI21X1 _14647_ (
    .A(_5106_),
    .B(_5134_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [24])
);

NAND3X1 _14227_ (
    .A(_4721_),
    .B(_4722_),
    .C(_4720_),
    .Y(_4723_)
);

FILL FILL_0__7091_ (
);

FILL FILL_1__16310_ (
);

FILL FILL_3__10831_ (
);

FILL FILL_3__10411_ (
);

FILL FILL_0__15723_ (
);

FILL FILL_0__15303_ (
);

FILL SFILL13720x24050 (
);

FILL FILL_2__8890_ (
);

FILL FILL_5__12269_ (
);

FILL FILL_2__8470_ (
);

INVX1 _6989_ (
    .A(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_60_)
);

FILL FILL_4__8396_ (
);

FILL FILL_2__12296_ (
);

FILL SFILL38920x73050 (
);

FILL FILL_5__13630_ (
);

FILL FILL_5__13210_ (
);

NAND2X1 _7930_ (
    .A(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_525_)
);

DFFSR _7510_ (
    .Q(\datapath_1.regfile_1.regOut[5] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_263_[0])
);

FILL FILL_1__11289_ (
);

FILL FILL_4__12623_ (
);

FILL FILL_4__12203_ (
);

DFFSR _10987_ (
    .Q(\control_1.reg_state.dout [3]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_2098_[3])
);

INVX1 _10567_ (
    .A(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_1876_)
);

INVX1 _10147_ (
    .A(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_1657_)
);

FILL FILL_3__11616_ (
);

FILL FILL_1__12650_ (
);

FILL FILL_1__12230_ (
);

FILL FILL_4__15095_ (
);

FILL FILL_2__9675_ (
);

FILL FILL_2__9255_ (
);

FILL FILL_0__11643_ (
);

FILL FILL_0__11223_ (
);

FILL FILL_3__14088_ (
);

FILL FILL_5__7680_ (
);

FILL SFILL3560x72050 (
);

FILL FILL_5__14835_ (
);

FILL FILL_5__14415_ (
);

INVX1 _8715_ (
    .A(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_926_)
);

FILL FILL_1__7672_ (
);

FILL FILL_1__7252_ (
);

FILL FILL_4__13828_ (
);

FILL FILL_2__14862_ (
);

FILL FILL_4__13408_ (
);

FILL FILL_2__14442_ (
);

FILL FILL_2__14022_ (
);

FILL FILL_3__7598_ (
);

FILL FILL_3__7178_ (
);

FILL FILL112200x67050 (
);

FILL FILL_1__13855_ (
);

FILL FILL_1__13435_ (
);

FILL FILL_1__13015_ (
);

FILL SFILL44040x9050 (
);

FILL FILL_0__12848_ (
);

FILL FILL_0__12428_ (
);

INVX1 _12713_ (
    .A(\datapath_1.PCJump [8]),
    .Y(_3501_)
);

FILL FILL_0__12008_ (
);

FILL SFILL38840x35050 (
);

FILL FILL_5__8885_ (
);

FILL FILL_5__8465_ (
);

FILL SFILL34120x13050 (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1_BUFX2_insert12 (
);

FILL FILL_1_BUFX2_insert13 (
);

NOR2X1 _15185_ (
    .A(_5661_),
    .B(_5653_),
    .Y(_5662_)
);

FILL FILL_1_BUFX2_insert14 (
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_1_BUFX2_insert16 (
);

FILL FILL_3__16234_ (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_1_BUFX2_insert18 (
);

FILL SFILL28920x71050 (
);

FILL FILL_5__10755_ (
);

FILL FILL_1__8877_ (
);

FILL FILL_1_BUFX2_insert19 (
);

FILL FILL_1__8457_ (
);

FILL FILL_2__15647_ (
);

FILL FILL_2__15227_ (
);

FILL FILL_4__6882_ (
);

FILL FILL_0__16261_ (
);

FILL FILL_2__10782_ (
);

FILL FILL_2__10362_ (
);

FILL FILL112200x22050 (
);

FILL SFILL99480x15050 (
);

FILL FILL_3__9744_ (
);

NAND3X1 _13918_ (
    .A(_4412_),
    .B(_4413_),
    .C(_4420_),
    .Y(_4421_)
);

FILL SFILL28840x78050 (
);

FILL FILL_4__13581_ (
);

FILL FILL_4__13161_ (
);

FILL FILL_2__7741_ (
);

FILL FILL_3__12994_ (
);

FILL FILL_3__12574_ (
);

FILL FILL_2__7321_ (
);

FILL FILL_3__12154_ (
);

FILL FILL112120x29050 (
);

FILL FILL_4__7247_ (
);

FILL FILL_2__11987_ (
);

FILL FILL_2__11567_ (
);

FILL FILL_2__11147_ (
);

FILL FILL_0__12181_ (
);

FILL FILL_5__12901_ (
);

FILL FILL_6__16380_ (
);

FILL FILL_5__15793_ (
);

FILL FILL_5__15373_ (
);

FILL FILL_0__7987_ (
);

FILL FILL_0__7567_ (
);

OAI21X1 _9673_ (
    .A(_1421_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1422_),
    .Y(_1368_[27])
);

OAI21X1 _9253_ (
    .A(_1202_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1203_),
    .Y(_1173_[15])
);

FILL FILL_1__11921_ (
);

FILL FILL_4__14786_ (
);

FILL SFILL28840x33050 (
);

FILL FILL_4__14366_ (
);

FILL FILL_1__11501_ (
);

FILL FILL_0__10914_ (
);

FILL FILL_2__8526_ (
);

FILL FILL_3__13779_ (
);

FILL FILL_3__13359_ (
);

FILL FILL_2__8106_ (
);

FILL FILL_1__14393_ (
);

FILL SFILL33800x16050 (
);

FILL FILL_5__6951_ (
);

INVX1 _13671_ (
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_4179_)
);

FILL FILL_0__13386_ (
);

AOI21X1 _13251_ (
    .A(_3793_),
    .B(_3761_),
    .C(\datapath_1.a3 [4]),
    .Y(_3794_)
);

FILL FILL_3__14720_ (
);

FILL FILL_3__14300_ (
);

FILL FILL_1__6943_ (
);

FILL FILL_4__9813_ (
);

FILL FILL_2__13713_ (
);

FILL FILL_3__6869_ (
);

FILL FILL_5__16158_ (
);

FILL FILL_5__11293_ (
);

FILL FILL_1__12706_ (
);

FILL SFILL18840x76050 (
);

FILL FILL_2__16185_ (
);

FILL SFILL113960x18050 (
);

FILL FILL_4__10286_ (
);

FILL FILL_3__7810_ (
);

FILL FILL_1__15598_ (
);

FILL FILL_1__15178_ (
);

FILL FILL_5__7736_ (
);

FILL FILL_5__7316_ (
);

FILL FILL_2_BUFX2_insert700 (
);

FILL FILL_2_BUFX2_insert701 (
);

FILL FILL_2_BUFX2_insert702 (
);

NOR2X1 _14876_ (
    .A(_5358_),
    .B(_5355_),
    .Y(_5359_)
);

FILL FILL_2_BUFX2_insert703 (
);

FILL SFILL13800x6050 (
);

OAI22X1 _14456_ (
    .A(_4946_),
    .B(_3909_),
    .C(_3881_),
    .D(_4945_),
    .Y(_4947_)
);

FILL FILL_2_BUFX2_insert704 (
);

NAND3X1 _14036_ (
    .A(_4532_),
    .B(_4535_),
    .C(_4531_),
    .Y(_4536_)
);

FILL FILL_2_BUFX2_insert705 (
);

FILL FILL_3__15925_ (
);

FILL FILL_2_BUFX2_insert706 (
);

FILL FILL_3__15505_ (
);

FILL FILL_2_BUFX2_insert707 (
);

FILL FILL_2_BUFX2_insert708 (
);

FILL FILL_2_BUFX2_insert709 (
);

FILL FILL_1__7728_ (
);

FILL FILL_3__10640_ (
);

FILL FILL_1__7308_ (
);

FILL FILL_2__14918_ (
);

FILL FILL_0__15952_ (
);

FILL FILL_0__15532_ (
);

FILL FILL_0__15112_ (
);

FILL FILL_5__12498_ (
);

FILL FILL_5__12078_ (
);

FILL SFILL18840x31050 (
);

FILL FILL_1__11098_ (
);

FILL FILL_4__12852_ (
);

FILL FILL_4__12432_ (
);

FILL FILL_4__12012_ (
);

INVX1 _10796_ (
    .A(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_1988_)
);

INVX1 _10376_ (
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_1769_)
);

FILL FILL_3__11845_ (
);

FILL FILL_3__11425_ (
);

FILL FILL_3__11005_ (
);

FILL FILL_4__6938_ (
);

FILL FILL_0__16317_ (
);

FILL FILL_2__9484_ (
);

FILL FILL_0__11872_ (
);

FILL FILL_2__10418_ (
);

FILL FILL_0__11452_ (
);

FILL FILL_0__11032_ (
);

FILL FILL_5__14644_ (
);

FILL FILL_5__14224_ (
);

FILL FILL_0__6838_ (
);

DFFSR _8944_ (
    .Q(\datapath_1.regfile_1.regOut[16] [26]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_978_[26])
);

OAI21X1 _8524_ (
    .A(_838_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_839_),
    .Y(_783_[28])
);

OAI21X1 _8104_ (
    .A(_619_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .C(_620_),
    .Y(_588_[16])
);

FILL FILL_1__7481_ (
);

FILL FILL_1__7061_ (
);

FILL FILL_4__13637_ (
);

FILL FILL_4__13217_ (
);

FILL FILL_2__14671_ (
);

FILL FILL_2__14251_ (
);

FILL FILL_1__13664_ (
);

FILL FILL_1__13244_ (
);

FILL FILL_1_BUFX2_insert720 (
);

FILL FILL_1_BUFX2_insert721 (
);

FILL FILL_0__12657_ (
);

DFFSR _12942_ (
    .Q(\datapath_1.a [23]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3555_[23])
);

FILL FILL_1_BUFX2_insert722 (
);

FILL FILL_1_BUFX2_insert723 (
);

OAI21X1 _12522_ (
    .A(_3413_),
    .B(vdd),
    .C(_3414_),
    .Y(_3360_[27])
);

FILL FILL_0__12237_ (
);

FILL FILL_1_BUFX2_insert724 (
);

NAND3X1 _12102_ (
    .A(_3120_),
    .B(_3121_),
    .C(_3122_),
    .Y(\datapath_1.mux_pcsrc.dout [28])
);

FILL FILL_1_BUFX2_insert725 (
);

FILL FILL_1_BUFX2_insert726 (
);

FILL FILL_5__8694_ (
);

FILL FILL_1_BUFX2_insert727 (
);

FILL FILL_5__8274_ (
);

FILL FILL_1_BUFX2_insert728 (
);

FILL FILL_1_BUFX2_insert729 (
);

FILL FILL_5__15849_ (
);

FILL FILL_5__15429_ (
);

FILL FILL_5__15009_ (
);

OAI21X1 _9729_ (
    .A(_1438_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .C(_1439_),
    .Y(_1433_[3])
);

FILL FILL_3__16043_ (
);

DFFSR _9309_ (
    .Q(\datapath_1.regfile_1.regOut[19] [7]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_1173_[7])
);

FILL FILL_5__10564_ (
);

FILL FILL_1__8266_ (
);

FILL FILL_5__10144_ (
);

FILL FILL_2__15876_ (
);

FILL SFILL69080x40050 (
);

FILL FILL_2__15456_ (
);

FILL FILL_2__15036_ (
);

FILL FILL_0__16070_ (
);

FILL SFILL48920x25050 (
);

FILL FILL_2__10171_ (
);

FILL FILL_1__14869_ (
);

FILL FILL_1__14449_ (
);

FILL FILL_1__14029_ (
);

FILL FILL_3__9553_ (
);

FILL FILL_3__9133_ (
);

NAND3X1 _13727_ (
    .A(_4224_),
    .B(_4226_),
    .C(_4233_),
    .Y(_4234_)
);

AOI21X1 _13307_ (
    .A(_3763_),
    .B(_3790_),
    .C(_3835_),
    .Y(_3841_)
);

FILL FILL_5__9899_ (
);

FILL FILL_1__15810_ (
);

FILL FILL_5__9479_ (
);

OAI22X1 _16199_ (
    .A(_5549__bF$buf2),
    .B(_6650_),
    .C(_5466__bF$buf2),
    .D(_6649_),
    .Y(_6651_)
);

FILL FILL_4__13390_ (
);

FILL FILL_0__14803_ (
);

FILL FILL_2__7970_ (
);

FILL FILL_5__11769_ (
);

FILL FILL_5__11349_ (
);

FILL FILL_2__7550_ (
);

FILL FILL_3__12383_ (
);

FILL SFILL59080x83050 (
);

FILL FILL_4__7476_ (
);

FILL FILL_4__7056_ (
);

FILL FILL_2__11796_ (
);

FILL SFILL38920x68050 (
);

FILL FILL_2__11376_ (
);

FILL FILL_5__12710_ (
);

FILL FILL_1__10789_ (
);

FILL FILL_1__10369_ (
);

FILL FILL_4__11703_ (
);

FILL SFILL3640x60050 (
);

FILL FILL_5__15182_ (
);

FILL FILL_0__7376_ (
);

OAI21X1 _9482_ (
    .A(_1314_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1315_),
    .Y(_1303_[6])
);

DFFSR _9062_ (
    .Q(\datapath_1.regfile_1.regOut[17] [16]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1043_[16])
);

FILL FILL_4__14595_ (
);

FILL FILL_1__11730_ (
);

FILL FILL_4__14175_ (
);

FILL FILL_1__11310_ (
);

FILL FILL_2__8755_ (
);

FILL FILL_3__13588_ (
);

FILL FILL_2__8335_ (
);

FILL FILL_0__10303_ (
);

FILL FILL_3__13168_ (
);

FILL SFILL59000x81050 (
);

FILL FILL_6__14922_ (
);

FILL SFILL3480x3050 (
);

FILL SFILL3560x67050 (
);

INVX1 _13480_ (
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_3991_)
);

FILL FILL_5__13915_ (
);

DFFSR _13060_ (
    .Q(_2_[13]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_3620_[13])
);

FILL FILL_4_BUFX2_insert230 (
);

FILL FILL_4_BUFX2_insert231 (
);

FILL FILL_4__9622_ (
);

FILL FILL_4__12908_ (
);

FILL FILL_4_BUFX2_insert232 (
);

FILL FILL_4_BUFX2_insert233 (
);

FILL FILL_2__13942_ (
);

FILL FILL_5__16387_ (
);

FILL FILL_2__13522_ (
);

FILL FILL_4_BUFX2_insert234 (
);

FILL FILL_2__13102_ (
);

FILL FILL_4_BUFX2_insert235 (
);

FILL FILL_4_BUFX2_insert236 (
);

FILL FILL_4_BUFX2_insert237 (
);

FILL FILL_4_BUFX2_insert238 (
);

FILL FILL_4_BUFX2_insert239 (
);

FILL FILL_1__12515_ (
);

FILL FILL_0__11928_ (
);

FILL FILL_0__9522_ (
);

FILL FILL_0__9102_ (
);

FILL FILL_0__11508_ (
);

FILL FILL_5__7965_ (
);

FILL FILL_5__7545_ (
);

FILL FILL_4__16321_ (
);

FILL FILL_5__7125_ (
);

INVX1 _14685_ (
    .A(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_5172_)
);

AOI21X1 _14265_ (
    .A(_4739_),
    .B(_4760_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [16])
);

FILL FILL_3__15734_ (
);

FILL FILL_3__15314_ (
);

FILL SFILL28920x66050 (
);

FILL SFILL3560x22050 (
);

FILL FILL_1__7957_ (
);

FILL FILL_1__7117_ (
);

FILL FILL_2__14727_ (
);

FILL FILL_2__14307_ (
);

FILL FILL_0__15761_ (
);

FILL FILL_0__15341_ (
);

FILL FILL_3__8824_ (
);

FILL FILL_3__8404_ (
);

FILL FILL_4__12661_ (
);

FILL FILL_4__12241_ (
);

OAI21X1 _10185_ (
    .A(_1681_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1682_),
    .Y(_1628_[27])
);

FILL FILL_3__11654_ (
);

FILL FILL_3__11234_ (
);

FILL FILL_6__14099_ (
);

FILL SFILL28920x21050 (
);

FILL FILL_0__16126_ (
);

INVX1 _16411_ (
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_6828_)
);

FILL FILL_2__10647_ (
);

FILL FILL_2__9293_ (
);

FILL FILL_0__11681_ (
);

FILL FILL_0__11261_ (
);

FILL FILL_6__15040_ (
);

FILL FILL_3__9609_ (
);

FILL FILL_3_BUFX2_insert250 (
);

FILL FILL_3_BUFX2_insert251 (
);

FILL FILL_5__14873_ (
);

FILL FILL_3_BUFX2_insert252 (
);

FILL SFILL28040x45050 (
);

FILL FILL_5__14453_ (
);

FILL FILL_3_BUFX2_insert253 (
);

FILL FILL_3_BUFX2_insert254 (
);

FILL FILL_5__14033_ (
);

FILL FILL_3_BUFX2_insert255 (
);

OAI21X1 _8753_ (
    .A(_950_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_951_),
    .Y(_913_[19])
);

OAI21X1 _8333_ (
    .A(_731_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_732_),
    .Y(_718_[7])
);

FILL FILL_3_BUFX2_insert256 (
);

FILL FILL_3_BUFX2_insert257 (
);

FILL FILL_3_BUFX2_insert258 (
);

FILL FILL_1__7290_ (
);

FILL SFILL28840x28050 (
);

FILL FILL_4__13866_ (
);

FILL FILL_3_BUFX2_insert259 (
);

FILL FILL_4__13446_ (
);

FILL FILL_2__14480_ (
);

FILL FILL_4__13026_ (
);

FILL FILL_2__14060_ (
);

FILL SFILL89080x39050 (
);

FILL FILL_2__7606_ (
);

FILL FILL_3__12859_ (
);

FILL FILL_3__12439_ (
);

FILL FILL_1__13893_ (
);

FILL FILL_3__12019_ (
);

FILL FILL_1__13473_ (
);

FILL FILL_0__12886_ (
);

OAI21X1 _12751_ (
    .A(_3525_),
    .B(IRWrite_bF$buf7),
    .C(_3526_),
    .Y(_3490_[18])
);

FILL FILL_0__12466_ (
);

FILL FILL_0__12046_ (
);

NAND3X1 _12331_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3287_)
);

FILL FILL_3__13800_ (
);

FILL FILL_5__8083_ (
);

FILL FILL_5__15658_ (
);

FILL FILL_5__15238_ (
);

DFFSR _9958_ (
    .Q(\datapath_1.regfile_1.regOut[24] [16]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_1498_[16])
);

FILL FILL_3__16272_ (
);

NAND2X1 _9538_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1353_)
);

FILL FILL_5__10793_ (
);

NAND2X1 _9118_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1134_)
);

FILL FILL_1__8495_ (
);

FILL FILL_5__10373_ (
);

FILL FILL_1__8075_ (
);

FILL FILL_2__15685_ (
);

FILL FILL_2__15265_ (
);

FILL SFILL94360x50050 (
);

FILL FILL_1__14678_ (
);

FILL FILL_1__14258_ (
);

FILL FILL_0_BUFX2_insert380 (
);

FILL FILL_0_BUFX2_insert381 (
);

FILL FILL_0_BUFX2_insert382 (
);

FILL FILL_3__9782_ (
);

FILL FILL_0_BUFX2_insert383 (
);

FILL FILL_0_BUFX2_insert384 (
);

OAI22X1 _13956_ (
    .A(_4456_),
    .B(_3902__bF$buf3),
    .C(_3971__bF$buf2),
    .D(_4457_),
    .Y(_4458_)
);

FILL FILL_3__9362_ (
);

FILL FILL_0_BUFX2_insert385 (
);

OAI22X1 _13536_ (
    .A(_4044_),
    .B(_3910_),
    .C(_3935__bF$buf2),
    .D(_4045_),
    .Y(_4046_)
);

FILL FILL_0_BUFX2_insert386 (
);

NAND2X1 _13116_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_pcsrc.dout [12]),
    .Y(_3709_)
);

FILL FILL_0_BUFX2_insert387 (
);

FILL FILL_0_BUFX2_insert388 (
);

FILL FILL_0_BUFX2_insert389 (
);

FILL FILL_5__9288_ (
);

FILL SFILL79160x30050 (
);

FILL FILL_0__14612_ (
);

FILL FILL_5__11998_ (
);

FILL FILL_5__11578_ (
);

FILL FILL_5__11158_ (
);

FILL FILL_3__12192_ (
);

FILL SFILL18840x26050 (
);

FILL FILL_2__11185_ (
);

FILL FILL_1__10178_ (
);

FILL FILL_4__11932_ (
);

FILL FILL_4__11512_ (
);

FILL FILL_2_BUFX2_insert60 (
);

FILL FILL_0__7185_ (
);

FILL FILL_2_BUFX2_insert61 (
);

NAND2X1 _9291_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1229_)
);

FILL FILL_1__16404_ (
);

FILL FILL_2_BUFX2_insert62 (
);

FILL FILL_3__10925_ (
);

FILL FILL_2_BUFX2_insert63 (
);

FILL FILL_3__10505_ (
);

FILL FILL_2_BUFX2_insert64 (
);

FILL FILL_2_BUFX2_insert65 (
);

FILL FILL_2_BUFX2_insert66 (
);

FILL FILL_0__15817_ (
);

FILL FILL_2_BUFX2_insert67 (
);

FILL FILL_2_BUFX2_insert68 (
);

FILL FILL_2_BUFX2_insert69 (
);

FILL FILL_2__8984_ (
);

FILL FILL_0__10952_ (
);

FILL FILL_0__10532_ (
);

FILL FILL_3__13397_ (
);

FILL FILL_2__8144_ (
);

FILL FILL_0__10112_ (
);

FILL FILL_5__13724_ (
);

FILL FILL_5__13304_ (
);

OAI21X1 _7604_ (
    .A(_367_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_368_),
    .Y(_328_[20])
);

FILL FILL_1__6981_ (
);

FILL FILL_4__9851_ (
);

FILL FILL_4__12717_ (
);

FILL FILL_4__9011_ (
);

FILL FILL_2__13751_ (
);

FILL FILL_2__13331_ (
);

FILL FILL_5__16196_ (
);

FILL FILL_6__9777_ (
);

FILL FILL_1__12744_ (
);

FILL FILL_4__15189_ (
);

FILL FILL_1__12324_ (
);

FILL FILL_0__9751_ (
);

FILL FILL_2__9769_ (
);

FILL FILL_2__9349_ (
);

FILL FILL_0__11737_ (
);

INVX1 _11602_ (
    .A(_2707_),
    .Y(_2708_)
);

FILL FILL_0__11317_ (
);

FILL FILL_6__15516_ (
);

FILL FILL_5__7354_ (
);

FILL FILL_4__16130_ (
);

FILL FILL_6__10651_ (
);

INVX1 _14494_ (
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_4985_)
);

NOR2X1 _14074_ (
    .A(_4563_),
    .B(_4573_),
    .Y(_4574_)
);

FILL FILL_5__14929_ (
);

FILL FILL_5__14509_ (
);

FILL FILL_3__15963_ (
);

FILL SFILL69000x78050 (
);

FILL FILL_3__15543_ (
);

DFFSR _8809_ (
    .Q(\datapath_1.regfile_1.regOut[15] [19]),
    .CLK(clk_bF$buf61),
    .R(rst_bF$buf87),
    .S(vdd),
    .D(_913_[19])
);

FILL FILL_3__15123_ (
);

FILL FILL_1__7346_ (
);

FILL SFILL69080x35050 (
);

FILL FILL_2__14956_ (
);

FILL FILL_0__15990_ (
);

FILL FILL_2__14536_ (
);

FILL FILL_0__15570_ (
);

FILL FILL_2__14116_ (
);

FILL FILL_0__15150_ (
);

FILL FILL_1__13949_ (
);

FILL FILL_1__13529_ (
);

FILL FILL_1__13109_ (
);

FILL FILL_3__8633_ (
);

DFFSR _12807_ (
    .Q(\datapath_1.PCJump [18]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3490_[16])
);

FILL FILL_3__8213_ (
);

FILL FILL_5__8979_ (
);

FILL FILL_5__8139_ (
);

NOR2X1 _15699_ (
    .A(_6162_),
    .B(_5544__bF$buf3),
    .Y(_6163_)
);

FILL FILL_4__12890_ (
);

FILL FILL_6__11436_ (
);

FILL FILL_4__12470_ (
);

FILL FILL_6__11016_ (
);

OAI22X1 _15279_ (
    .A(_5480__bF$buf1),
    .B(_4209_),
    .C(_4199_),
    .D(_5499__bF$buf0),
    .Y(_5754_)
);

FILL FILL_4__12050_ (
);

FILL FILL_3__16328_ (
);

FILL FILL_5__10429_ (
);

FILL FILL_3__11883_ (
);

FILL FILL_5__9920_ (
);

FILL FILL_5__10009_ (
);

FILL FILL_5__9500_ (
);

FILL FILL_3__11463_ (
);

FILL FILL_3__11043_ (
);

FILL SFILL59080x78050 (
);

FILL FILL_4__6976_ (
);

FILL FILL_0__16355_ (
);

NOR2X1 _16220_ (
    .A(_6670_),
    .B(_6661_),
    .Y(_6671_)
);

FILL FILL_2__10876_ (
);

FILL FILL_0__11490_ (
);

FILL FILL_2__10036_ (
);

FILL FILL_0__11070_ (
);

FILL FILL_1__9912_ (
);

FILL FILL_3__9418_ (
);

FILL SFILL3640x55050 (
);

FILL FILL_5__14682_ (
);

FILL FILL_5__14262_ (
);

FILL FILL_0__6876_ (
);

OAI21X1 _8982_ (
    .A(_1062_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1063_),
    .Y(_1043_[10])
);

DFFSR _8562_ (
    .Q(\datapath_1.regfile_1.regOut[13] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_783_[28])
);

NAND2X1 _8142_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_646_)
);

FILL SFILL43880x62050 (
);

FILL FILL_4__13675_ (
);

FILL FILL_1__10810_ (
);

FILL FILL_4__13255_ (
);

INVX1 _11199_ (
    .A(\datapath_1.alu_1.ALUInB [29]),
    .Y(_2318_)
);

FILL FILL_2__7835_ (
);

FILL FILL_2__7415_ (
);

FILL FILL_3__12248_ (
);

FILL SFILL59000x76050 (
);

FILL FILL_1__13282_ (
);

FILL SFILL59080x33050 (
);

FILL FILL_0__12695_ (
);

OAI21X1 _12980_ (
    .A(_3637_),
    .B(vdd),
    .C(_3638_),
    .Y(_3620_[9])
);

DFFSR _12560_ (
    .Q(ALUOut[25]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3360_[25])
);

FILL FILL_0__12275_ (
);

NAND2X1 _12140_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [8]),
    .Y(_3147_)
);

FILL SFILL38920x18050 (
);

FILL FILL_4__8702_ (
);

FILL FILL_5__15887_ (
);

FILL FILL_2__12602_ (
);

FILL FILL_5__15467_ (
);

FILL FILL_5__15047_ (
);

NAND2X1 _9767_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1465_)
);

FILL FILL_3__16081_ (
);

NAND2X1 _9347_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1246_)
);

FILL SFILL3640x10050 (
);

FILL FILL_5__10182_ (
);

FILL FILL_2__15494_ (
);

FILL FILL_2__15074_ (
);

FILL FILL_0__8602_ (
);

FILL FILL_1__14487_ (
);

FILL FILL_1__14067_ (
);

FILL FILL_4__15821_ (
);

FILL FILL_4__15401_ (
);

FILL FILL_3__9591_ (
);

FILL SFILL49080x76050 (
);

NOR2X1 _13765_ (
    .A(_4270_),
    .B(_3931__bF$buf0),
    .Y(_4271_)
);

FILL FILL_3__9171_ (
);

NOR2X1 _13345_ (
    .A(_3798_),
    .B(_3774_),
    .Y(\datapath_1.regfile_1.regEn [24])
);

FILL FILL_3__14814_ (
);

FILL SFILL3560x17050 (
);

FILL FILL_5__9097_ (
);

FILL FILL_4__9907_ (
);

FILL SFILL104440x34050 (
);

FILL FILL_2__13807_ (
);

FILL FILL_0__14841_ (
);

FILL FILL_0__14421_ (
);

FILL FILL_0__14001_ (
);

FILL FILL_5__11387_ (
);

FILL FILL_1__9089_ (
);

FILL SFILL28840x50 (
);

FILL FILL_2__16279_ (
);

FILL FILL_4__7094_ (
);

FILL FILL_0__9807_ (
);

FILL FILL_4__11741_ (
);

FILL FILL_4__11321_ (
);

FILL FILL_6__8381_ (
);

FILL SFILL49080x31050 (
);

FILL FILL_1__16213_ (
);

FILL FILL_3__10314_ (
);

FILL SFILL94440x83050 (
);

NAND2X1 _15911_ (
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .B(_5570__bF$buf3),
    .Y(_6370_)
);

FILL FILL_0__15626_ (
);

FILL FILL_0__15206_ (
);

FILL FILL_2__8373_ (
);

FILL FILL_0__10761_ (
);

FILL FILL_2__12199_ (
);

FILL FILL_5__13953_ (
);

FILL FILL_5__13533_ (
);

FILL FILL_5__13113_ (
);

OAI21X1 _7833_ (
    .A(_479_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .C(_480_),
    .Y(_458_[11])
);

DFFSR _7413_ (
    .Q(\datapath_1.regfile_1.regOut[4] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_198_[31])
);

FILL FILL_4_BUFX2_insert610 (
);

FILL FILL_4__9660_ (
);

FILL FILL_4_BUFX2_insert611 (
);

FILL FILL_4__9240_ (
);

FILL FILL_4_BUFX2_insert612 (
);

FILL FILL_4__12526_ (
);

FILL FILL_2__13980_ (
);

FILL FILL_4_BUFX2_insert613 (
);

FILL SFILL90120x30050 (
);

FILL FILL_4_BUFX2_insert614 (
);

FILL FILL_4__12106_ (
);

FILL FILL_2__13560_ (
);

FILL FILL_4_BUFX2_insert615 (
);

FILL FILL_2__13140_ (
);

FILL FILL_4_BUFX2_insert616 (
);

FILL FILL_0__8199_ (
);

FILL FILL_4_BUFX2_insert617 (
);

FILL FILL_4_BUFX2_insert618 (
);

FILL FILL_3__11939_ (
);

FILL FILL_4_BUFX2_insert619 (
);

FILL FILL_1__12973_ (
);

FILL FILL_3__11519_ (
);

FILL FILL_1__12133_ (
);

FILL FILL_2__9998_ (
);

FILL FILL_0__9980_ (
);

FILL FILL_0__11966_ (
);

FILL FILL_2__9158_ (
);

FILL FILL_0__9140_ (
);

NOR2X1 _11831_ (
    .A(_2357_),
    .B(_2491_),
    .Y(_2920_)
);

FILL FILL_0__11546_ (
);

AOI21X1 _11411_ (
    .A(_2526_),
    .B(_2522_),
    .C(_2527_),
    .Y(_2528_)
);

FILL FILL_0__11126_ (
);

FILL FILL_5__7583_ (
);

FILL FILL_5__7163_ (
);

FILL FILL_5__14738_ (
);

FILL FILL_5__14318_ (
);

FILL FILL_3__15772_ (
);

FILL SFILL39480x43050 (
);

FILL FILL_3__15352_ (
);

NAND2X1 _8618_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_882_)
);

FILL FILL_1__7995_ (
);

FILL FILL_1__7575_ (
);

FILL FILL_2__14765_ (
);

FILL FILL_2__14345_ (
);

FILL SFILL39000x72050 (
);

FILL FILL_1__13758_ (
);

FILL FILL_1__13338_ (
);

FILL FILL_3__8862_ (
);

FILL FILL_3__8442_ (
);

NAND2X1 _12616_ (
    .A(vdd),
    .B(memoryOutData[16]),
    .Y(_3457_)
);

FILL FILL_5__8788_ (
);

FILL SFILL79160x25050 (
);

FILL FILL_5__8368_ (
);

INVX8 _15088_ (
    .A(_5544__bF$buf3),
    .Y(_5567_)
);

FILL FILL_3__16137_ (
);

FILL FILL_5__10658_ (
);

FILL FILL_5__10238_ (
);

FILL FILL_3__11692_ (
);

FILL FILL_3__11272_ (
);

FILL FILL_0__16164_ (
);

FILL FILL_2__10685_ (
);

FILL FILL_2__10265_ (
);

FILL FILL_1__9721_ (
);

FILL FILL_1__9301_ (
);

FILL FILL_3_BUFX2_insert630 (
);

FILL FILL_3__9647_ (
);

FILL FILL_3__9227_ (
);

FILL FILL_3_BUFX2_insert631 (
);

FILL FILL_3_BUFX2_insert632 (
);

FILL FILL_3_BUFX2_insert633 (
);

FILL FILL_5__14491_ (
);

FILL FILL_3_BUFX2_insert634 (
);

FILL FILL_5__14071_ (
);

FILL FILL_3_BUFX2_insert635 (
);

FILL FILL_1__15904_ (
);

DFFSR _8791_ (
    .Q(\datapath_1.regfile_1.regOut[15] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_913_[1])
);

FILL FILL_3_BUFX2_insert636 (
);

NAND2X1 _8371_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_758_)
);

FILL FILL111960x3050 (
);

FILL FILL_3_BUFX2_insert637 (
);

FILL FILL_3_BUFX2_insert638 (
);

FILL FILL_3_BUFX2_insert639 (
);

FILL FILL_4__13484_ (
);

FILL SFILL8760x62050 (
);

FILL FILL_3__12897_ (
);

FILL SFILL63880x16050 (
);

FILL FILL_2__7224_ (
);

FILL FILL_3__12477_ (
);

FILL FILL_3__12057_ (
);

FILL FILL_1__13091_ (
);

FILL FILL_0__12084_ (
);

FILL SFILL114600x62050 (
);

FILL SFILL53960x52050 (
);

FILL SFILL84360x43050 (
);

FILL FILL_6__16283_ (
);

FILL FILL_4__8511_ (
);

FILL FILL_5__15696_ (
);

FILL FILL_2__12831_ (
);

FILL FILL_2__12411_ (
);

FILL FILL_5__15276_ (
);

NAND2X1 _9996_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1577_)
);

FILL FILL_6__8857_ (
);

DFFSR _9576_ (
    .Q(\datapath_1.regfile_1.regOut[21] [18]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_1303_[18])
);

INVX1 _9156_ (
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_1159_)
);

FILL FILL_1__11824_ (
);

FILL FILL_4__14689_ (
);

FILL FILL_4__14269_ (
);

FILL FILL_1__11404_ (
);

FILL FILL_0__8831_ (
);

FILL FILL_2__8849_ (
);

FILL FILL_0__10817_ (
);

FILL FILL_2__8009_ (
);

FILL FILL_1__14296_ (
);

FILL FILL_0_BUFX2_insert760 (
);

FILL FILL_5__6854_ (
);

FILL FILL_4__15630_ (
);

FILL FILL_0_BUFX2_insert761 (
);

FILL FILL_4__15210_ (
);

FILL FILL_0_BUFX2_insert762 (
);

FILL FILL_0_BUFX2_insert763 (
);

FILL FILL_0_BUFX2_insert764 (
);

INVX1 _13994_ (
    .A(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_4495_)
);

FILL FILL_0__13289_ (
);

FILL FILL_0_BUFX2_insert765 (
);

OAI22X1 _13574_ (
    .A(_4083_),
    .B(_3936__bF$buf4),
    .C(_3944__bF$buf4),
    .D(_4082_),
    .Y(_4084_)
);

FILL FILL_0_BUFX2_insert766 (
);

INVX1 _13154_ (
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3734_)
);

FILL FILL_0_BUFX2_insert767 (
);

FILL FILL_0_BUFX2_insert768 (
);

FILL FILL_3__14623_ (
);

FILL FILL_0_BUFX2_insert769 (
);

FILL FILL_3__14203_ (
);

FILL FILL_1__6846_ (
);

FILL SFILL114120x55050 (
);

FILL FILL_2__13616_ (
);

FILL FILL_0__14650_ (
);

FILL FILL_0__14230_ (
);

FILL FILL_5__11196_ (
);

FILL FILL_1__12609_ (
);

FILL FILL_2__16088_ (
);

FILL FILL_4__10189_ (
);

FILL FILL_0__9616_ (
);

FILL FILL_3__7713_ (
);

FILL SFILL114520x24050 (
);

FILL FILL_4__16415_ (
);

FILL FILL_5__7219_ (
);

FILL FILL_4__11970_ (
);

INVX1 _14779_ (
    .A(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_5264_)
);

AOI22X1 _14359_ (
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .B(_4102_),
    .C(_4129_),
    .D(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_4852_)
);

FILL FILL_4__11550_ (
);

FILL FILL_4__11130_ (
);

FILL SFILL3720x43050 (
);

FILL FILL_3__15828_ (
);

FILL FILL_3__15408_ (
);

FILL FILL_1__16022_ (
);

FILL FILL_3__10963_ (
);

FILL FILL_3__10543_ (
);

FILL SFILL43960x50050 (
);

FILL FILL_3__10123_ (
);

FILL FILL_0__15855_ (
);

NAND2X1 _15720_ (
    .A(_6183_),
    .B(_6178_),
    .Y(_6184_)
);

FILL FILL_0__15435_ (
);

INVX1 _15300_ (
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_5774_)
);

FILL FILL_0__15015_ (
);

FILL FILL_0__10990_ (
);

FILL FILL_0__10570_ (
);

FILL FILL_2__8182_ (
);

FILL FILL_0__10150_ (
);

FILL FILL_5__13762_ (
);

FILL FILL_5__13342_ (
);

DFFSR _7642_ (
    .Q(\datapath_1.regfile_1.regOut[6] [4]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_328_[4])
);

FILL SFILL104520x67050 (
);

NAND2X1 _7222_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_175_)
);

FILL SFILL43880x57050 (
);

FILL FILL_4__12755_ (
);

FILL FILL_4__12335_ (
);

NAND2X1 _10699_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1944_)
);

NAND2X1 _10279_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1725_)
);

FILL FILL_2__6915_ (
);

FILL FILL_3__11748_ (
);

FILL FILL_1__12782_ (
);

FILL FILL_3__11328_ (
);

FILL FILL_1__12362_ (
);

FILL SFILL59080x28050 (
);

FILL FILL112280x61050 (
);

FILL FILL_2__9387_ (
);

FILL FILL_0__11775_ (
);

FILL FILL_0__11355_ (
);

OAI21X1 _11640_ (
    .A(_2742_),
    .B(_2205_),
    .C(_2166_),
    .Y(_2743_)
);

OAI21X1 _11220_ (
    .A(_2111_),
    .B(_2332_),
    .C(_2338_),
    .Y(_2339_)
);

FILL FILL_5__14967_ (
);

FILL FILL_5__14547_ (
);

FILL FILL_5__14127_ (
);

FILL FILL_3__15581_ (
);

NAND2X1 _8847_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_994_)
);

FILL FILL_3__15161_ (
);

DFFSR _8427_ (
    .Q(\datapath_1.regfile_1.regOut[12] [21]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_718_[21])
);

INVX1 _8007_ (
    .A(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_576_)
);

FILL FILL_2__14994_ (
);

FILL FILL_2__14574_ (
);

FILL FILL_2__14154_ (
);

FILL SFILL43880x12050 (
);

FILL FILL_1__13987_ (
);

FILL FILL_1__13567_ (
);

FILL FILL_1__13147_ (
);

FILL FILL_4__14901_ (
);

FILL SFILL59000x26050 (
);

FILL FILL_3__8251_ (
);

NAND2X1 _12845_ (
    .A(vdd),
    .B(\datapath_1.rd1 [7]),
    .Y(_3569_)
);

FILL SFILL108840x30050 (
);

NAND2X1 _12425_ (
    .A(MemToReg_bF$buf6),
    .B(\datapath_1.Data [27]),
    .Y(_3349_)
);

AOI22X1 _12005_ (
    .A(\datapath_1.ALUResult [4]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3050_)
);

FILL FILL_6__16339_ (
);

FILL FILL_5__8597_ (
);

FILL FILL_0__13921_ (
);

FILL FILL_3__16366_ (
);

FILL FILL_0__13501_ (
);

FILL FILL_5__10887_ (
);

FILL FILL_1__8589_ (
);

FILL FILL_5__10047_ (
);

FILL FILL_3__11081_ (
);

FILL FILL_2__15779_ (
);

FILL FILL_2__15359_ (
);

FILL FILL_0__16393_ (
);

FILL FILL_2__10494_ (
);

FILL FILL_1__9530_ (
);

FILL FILL_1__9110_ (
);

FILL SFILL49000x69050 (
);

FILL FILL_2__16300_ (
);

FILL FILL_3__9876_ (
);

FILL FILL_3__9036_ (
);

FILL FILL_4__10821_ (
);

FILL FILL_4__10401_ (
);

FILL SFILL49080x26050 (
);

FILL FILL_1__15713_ (
);

FILL FILL_6__7461_ (
);

DFFSR _8180_ (
    .Q(\datapath_1.regfile_1.regOut[10] [30]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_588_[30])
);

FILL FILL_6__12259_ (
);

FILL FILL_4__13293_ (
);

FILL FILL_0__14706_ (
);

FILL FILL_2__7873_ (
);

FILL FILL_2__7453_ (
);

FILL FILL_3__12286_ (
);

FILL FILL_2__7033_ (
);

FILL FILL_4__7799_ (
);

FILL FILL_4__7379_ (
);

FILL FILL_2__11699_ (
);

FILL FILL_2__11279_ (
);

FILL SFILL33880x10050 (
);

FILL FILL_5__12613_ (
);

OAI21X1 _6913_ (
    .A(_8_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .C(_9_),
    .Y(_3_[3])
);

FILL FILL_2_BUFX2_insert290 (
);

FILL FILL_2_BUFX2_insert291 (
);

FILL FILL_4__8740_ (
);

FILL FILL_2_BUFX2_insert292 (
);

FILL FILL_4__8320_ (
);

FILL FILL_2_BUFX2_insert293 (
);

FILL FILL_2_BUFX2_insert294 (
);

FILL FILL_4__11606_ (
);

FILL FILL_2__12640_ (
);

FILL FILL_2_BUFX2_insert295 (
);

FILL FILL_2_BUFX2_insert296 (
);

FILL FILL_2__12220_ (
);

FILL FILL_5__15085_ (
);

FILL FILL_0__7699_ (
);

FILL FILL_2_BUFX2_insert297 (
);

FILL SFILL39080x69050 (
);

INVX1 _9385_ (
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_1271_)
);

FILL FILL_2_BUFX2_insert298 (
);

FILL FILL_2_BUFX2_insert299 (
);

FILL FILL_4__14498_ (
);

FILL FILL_1__11633_ (
);

FILL FILL_1__11213_ (
);

FILL FILL_4__14078_ (
);

FILL SFILL94440x33050 (
);

FILL FILL_0__8640_ (
);

FILL FILL_2__8658_ (
);

OAI21X1 _10911_ (
    .A(\control_1.reg_state.dout [1]),
    .B(_2047_),
    .C(_2056_),
    .Y(ALUSrcA)
);

FILL FILL_0__10626_ (
);

FILL FILL_0__8220_ (
);

FILL FILL_2__8238_ (
);

FILL FILL_6_BUFX2_insert14 (
);

FILL FILL_6__14825_ (
);

FILL FILL_6_BUFX2_insert19 (
);

AOI22X1 _13383_ (
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .B(_3894_),
    .C(_3891__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_3895_)
);

FILL FILL_0__13098_ (
);

FILL FILL_5__13818_ (
);

FILL SFILL23880x53050 (
);

FILL FILL_3__14852_ (
);

FILL FILL_3__14432_ (
);

FILL FILL_3__14012_ (
);

FILL FILL_4__9525_ (
);

FILL FILL_4__9105_ (
);

FILL FILL111800x69050 (
);

FILL FILL_2__13845_ (
);

FILL FILL_2__13425_ (
);

FILL SFILL63960x49050 (
);

FILL FILL_2__13005_ (
);

FILL SFILL39000x67050 (
);

FILL FILL_1__12838_ (
);

FILL FILL_1__12418_ (
);

FILL FILL_3__7942_ (
);

FILL FILL_0__9425_ (
);

FILL FILL_3__7102_ (
);

FILL FILL_0__9005_ (
);

FILL FILL_5__7868_ (
);

FILL FILL_5__7448_ (
);

FILL FILL_4__16224_ (
);

FILL FILL_6__10745_ (
);

INVX1 _14588_ (
    .A(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_5077_)
);

FILL FILL_6__10325_ (
);

NOR2X1 _14168_ (
    .A(_4665_),
    .B(_4662_),
    .Y(_4666_)
);

FILL SFILL23800x51050 (
);

FILL FILL_3__15637_ (
);

FILL FILL_3__15217_ (
);

FILL FILL_1__16251_ (
);

FILL FILL_3__10772_ (
);

FILL FILL_0__15664_ (
);

FILL SFILL79240x5050 (
);

FILL FILL_0__15244_ (
);

FILL SFILL53960x1050 (
);

FILL SFILL39000x22050 (
);

FILL FILL_3__8727_ (
);

FILL FILL_5__13991_ (
);

FILL FILL_5__13571_ (
);

FILL FILL_5__13151_ (
);

NAND2X1 _7871_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_506_)
);

NAND2X1 _7451_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_287_)
);

NAND2X1 _7031_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .Y(_132_)
);

FILL FILL_4__12984_ (
);

FILL FILL_4__12144_ (
);

DFFSR _10088_ (
    .Q(\datapath_1.regfile_1.regOut[25] [18]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf10),
    .S(vdd),
    .D(_1563_[18])
);

FILL FILL_3__11977_ (
);

FILL FILL_3__11557_ (
);

FILL FILL_1__12591_ (
);

FILL FILL_3__11137_ (
);

FILL FILL_1__12171_ (
);

FILL FILL_0__16449_ (
);

FILL FILL_0__16029_ (
);

OAI22X1 _16314_ (
    .A(_5534__bF$buf3),
    .B(_5434_),
    .C(_6762_),
    .D(_5549__bF$buf1),
    .Y(_6763_)
);

FILL FILL_0__11584_ (
);

FILL SFILL114600x57050 (
);

FILL FILL_0__11164_ (
);

FILL SFILL53960x47050 (
);

FILL SFILL84360x38050 (
);

FILL FILL_2__11911_ (
);

FILL FILL_5__14776_ (
);

FILL FILL_5__14356_ (
);

FILL FILL_6__7937_ (
);

FILL FILL_3__15390_ (
);

INVX1 _8656_ (
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_907_)
);

INVX1 _8236_ (
    .A(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_688_)
);

FILL FILL_1__7193_ (
);

FILL FILL_1__10904_ (
);

FILL FILL_4__13769_ (
);

FILL FILL_4__13349_ (
);

FILL FILL_2__14383_ (
);

FILL FILL_2__7929_ (
);

FILL SFILL8760x12050 (
);

FILL FILL_2__7509_ (
);

FILL FILL_1__13796_ (
);

FILL FILL_1__13376_ (
);

FILL FILL_4__14710_ (
);

FILL SFILL74040x60050 (
);

FILL FILL_0__12789_ (
);

FILL FILL_3__8480_ (
);

INVX1 _12654_ (
    .A(\datapath_1.Data [29]),
    .Y(_3482_)
);

FILL FILL_0__12369_ (
);

FILL FILL_3__8060_ (
);

NAND3X1 _12234_ (
    .A(_3212_),
    .B(_3213_),
    .C(_3214_),
    .Y(\datapath_1.alu_1.ALUInB [4])
);

FILL FILL_3__13703_ (
);

FILL FILL_0__13730_ (
);

FILL FILL_0__13310_ (
);

FILL FILL_3__16175_ (
);

FILL FILL_5__10696_ (
);

FILL FILL_1__8398_ (
);

FILL FILL_5__10276_ (
);

FILL FILL_2__15588_ (
);

FILL FILL_2__15168_ (
);

FILL FILL_4__15915_ (
);

FILL FILL_3__9685_ (
);

INVX1 _13859_ (
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_4363_)
);

FILL FILL_3__9265_ (
);

AOI22X1 _13439_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [0]),
    .C(\datapath_1.regfile_1.regOut[11] [0]),
    .D(_3950__bF$buf3),
    .Y(_3951_)
);

FILL FILL_4__10630_ (
);

OAI21X1 _13019_ (
    .A(_3663_),
    .B(vdd),
    .C(_3664_),
    .Y(_3620_[22])
);

FILL FILL_3__14908_ (
);

FILL FILL_1__15942_ (
);

FILL FILL_1__15522_ (
);

FILL FILL_1__15102_ (
);

FILL SFILL43960x45050 (
);

FILL FILL_0__14935_ (
);

NOR2X1 _14800_ (
    .A(_5280_),
    .B(_5283_),
    .Y(_5284_)
);

FILL FILL_0__14515_ (
);

FILL SFILL49640x5050 (
);

FILL FILL_2__7682_ (
);

FILL FILL_3__12095_ (
);

FILL FILL_4__7188_ (
);

FILL FILL_2__11088_ (
);

FILL FILL_5__12842_ (
);

FILL FILL_5__12422_ (
);

FILL FILL_5__12002_ (
);

FILL SFILL48920x7050 (
);

FILL FILL_4__11835_ (
);

FILL FILL_4__11415_ (
);

FILL FILL_6__8475_ (
);

FILL FILL_0__7088_ (
);

FILL FILL_1__16307_ (
);

DFFSR _9194_ (
    .Q(\datapath_1.regfile_1.regOut[18] [20]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_1108_[20])
);

FILL FILL_3__10828_ (
);

FILL FILL_3__10408_ (
);

FILL FILL_1__11862_ (
);

FILL FILL_1__11442_ (
);

FILL FILL_1__11022_ (
);

FILL FILL112280x56050 (
);

FILL FILL_2__8887_ (
);

FILL SFILL88760x4050 (
);

FILL FILL_2__8467_ (
);

DFFSR _10720_ (
    .Q(\datapath_1.regfile_1.regOut[30] [10]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1888_[10])
);

FILL FILL_0__10435_ (
);

NAND2X1 _10300_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1739_)
);

FILL FILL_0__10015_ (
);

FILL FILL_5__6892_ (
);

DFFSR _13192_ (
    .Q(\datapath_1.mux_iord.din0 [17]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[17])
);

FILL FILL_5__13627_ (
);

FILL FILL_5__13207_ (
);

FILL FILL_3__14661_ (
);

FILL FILL_3__14241_ (
);

NAND2X1 _7927_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .Y(_587_)
);

INVX1 _7507_ (
    .A(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_324_)
);

FILL FILL_1__6884_ (
);

FILL FILL_4__9754_ (
);

FILL FILL_4__9334_ (
);

FILL SFILL104520x17050 (
);

FILL FILL_2__13654_ (
);

FILL FILL_2__13234_ (
);

FILL FILL_5__16099_ (
);

FILL FILL_1__12647_ (
);

FILL FILL_1__12227_ (
);

FILL FILL_0__9654_ (
);

FILL FILL_3__7751_ (
);

FILL SFILL108840x25050 (
);

FILL FILL_3__7331_ (
);

OAI21X1 _11925_ (
    .A(_2990_),
    .B(IorD_bF$buf4),
    .C(_2991_),
    .Y(_1_[12])
);

FILL FILL_0__9234_ (
);

NOR2X1 _11505_ (
    .A(_2284_),
    .B(_2261_),
    .Y(_2617_)
);

FILL FILL112280x11050 (
);

FILL FILL_6__15419_ (
);

FILL FILL_5__7677_ (
);

FILL FILL_4__16033_ (
);

NOR2X1 _14397_ (
    .A(_4886_),
    .B(_4889_),
    .Y(_4890_)
);

FILL FILL_3__15866_ (
);

FILL FILL_3__15446_ (
);

FILL FILL_3__15026_ (
);

FILL FILL_1__16060_ (
);

FILL FILL_3__10581_ (
);

FILL FILL_1__7249_ (
);

FILL FILL_6_BUFX2_insert521 (
);

FILL FILL_3__10161_ (
);

FILL FILL_2__14859_ (
);

FILL FILL_0__15893_ (
);

FILL FILL_2__14439_ (
);

FILL FILL_2__14019_ (
);

FILL FILL_0__15473_ (
);

FILL FILL_0__15053_ (
);

FILL FILL_6_BUFX2_insert526 (
);

FILL FILL_1__8610_ (
);

FILL FILL_2__15800_ (
);

FILL FILL_3__8956_ (
);

FILL FILL_3__8116_ (
);

FILL FILL_5__13380_ (
);

NAND2X1 _7680_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_399_)
);

DFFSR _7260_ (
    .Q(\datapath_1.regfile_1.regOut[3] [6]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_133_[6])
);

FILL FILL_4__12373_ (
);

FILL FILL_2__6953_ (
);

FILL FILL_3__11786_ (
);

FILL FILL_5__9403_ (
);

FILL FILL_3__11366_ (
);

FILL FILL_4__6879_ (
);

FILL FILL_0__16258_ (
);

NOR2X1 _16123_ (
    .A(_6565_),
    .B(_6576_),
    .Y(_6577_)
);

FILL FILL_2__10779_ (
);

FILL FILL_2__10359_ (
);

FILL FILL_0__11393_ (
);

FILL FILL_6__15592_ (
);

FILL FILL_4__7820_ (
);

FILL FILL_5__14585_ (
);

FILL FILL_2__11720_ (
);

FILL FILL_5__14165_ (
);

FILL FILL_2__11300_ (
);

INVX1 _8885_ (
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_1019_)
);

INVX1 _8465_ (
    .A(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_800_)
);

DFFSR _8045_ (
    .Q(\datapath_1.regfile_1.regOut[9] [23]),
    .CLK(clk_bF$buf23),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_523_[23])
);

FILL FILL_4__13998_ (
);

FILL FILL_4__13578_ (
);

FILL FILL_4__13158_ (
);

FILL FILL_2__14192_ (
);

FILL SFILL94440x28050 (
);

FILL FILL_0__7720_ (
);

FILL FILL_2__7738_ (
);

FILL FILL_0__7300_ (
);

FILL FILL_2__7318_ (
);

FILL FILL_0__12598_ (
);

INVX1 _12883_ (
    .A(\datapath_1.a [20]),
    .Y(_3594_)
);

FILL FILL_0__12178_ (
);

INVX1 _12463_ (
    .A(ALUOut[8]),
    .Y(_3375_)
);

FILL SFILL23880x48050 (
);

NAND3X1 _12043_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[14]),
    .C(_3032__bF$buf3),
    .Y(_3078_)
);

FILL FILL_3__13932_ (
);

FILL FILL_3__13512_ (
);

FILL FILL_4__8605_ (
);

FILL FILL_5_BUFX2_insert540 (
);

FILL FILL_5_BUFX2_insert541 (
);

FILL FILL_2__12505_ (
);

FILL FILL_5_BUFX2_insert542 (
);

FILL FILL_5_BUFX2_insert543 (
);

FILL FILL_5_BUFX2_insert544 (
);

FILL FILL_5_BUFX2_insert545 (
);

FILL FILL_5_BUFX2_insert546 (
);

FILL FILL_5_BUFX2_insert547 (
);

FILL FILL_5_BUFX2_insert548 (
);

FILL FILL_1__11918_ (
);

FILL FILL_5_BUFX2_insert549 (
);

FILL FILL_2__15397_ (
);

FILL FILL_5__16311_ (
);

FILL FILL_0__8505_ (
);

FILL FILL_5__6948_ (
);

FILL FILL_4__15724_ (
);

FILL FILL_1_BUFX2_insert1070 (
);

FILL FILL_1_BUFX2_insert1071 (
);

FILL FILL_4__15304_ (
);

FILL FILL_1_BUFX2_insert1072 (
);

FILL FILL_1_BUFX2_insert1073 (
);

FILL FILL_3__9494_ (
);

INVX1 _13668_ (
    .A(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_4176_)
);

INVX1 _13248_ (
    .A(_3790_),
    .Y(_3791_)
);

FILL SFILL109480x1050 (
);

FILL FILL_3__14717_ (
);

FILL FILL_1__15751_ (
);

FILL FILL_1__15331_ (
);

FILL FILL_0__14744_ (
);

FILL FILL_0__14324_ (
);

FILL FILL_2__7491_ (
);

FILL FILL_2__7071_ (
);

FILL FILL_3__7807_ (
);

FILL SFILL108680x8050 (
);

FILL FILL_5__12651_ (
);

FILL FILL_5__12231_ (
);

NAND2X1 _6951_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_35_)
);

FILL FILL_2_BUFX2_insert670 (
);

FILL FILL_2_BUFX2_insert671 (
);

FILL FILL_2_BUFX2_insert672 (
);

FILL FILL_2_BUFX2_insert673 (
);

FILL FILL_2_BUFX2_insert674 (
);

FILL FILL_4__11644_ (
);

FILL FILL_2_BUFX2_insert675 (
);

FILL FILL_4__11224_ (
);

FILL FILL_2_BUFX2_insert676 (
);

FILL FILL_2_BUFX2_insert677 (
);

FILL FILL_2_BUFX2_insert678 (
);

FILL FILL_1__16116_ (
);

FILL FILL_2_BUFX2_insert679 (
);

FILL FILL_3__10637_ (
);

FILL FILL_1__11671_ (
);

FILL FILL_1__11251_ (
);

FILL FILL_0__15949_ (
);

FILL FILL_0__15529_ (
);

INVX1 _15814_ (
    .A(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_6275_)
);

FILL FILL_0__15109_ (
);

FILL FILL_2__8696_ (
);

FILL FILL_0__10664_ (
);

FILL FILL_2__8276_ (
);

FILL FILL_0__10244_ (
);

FILL FILL_5__13856_ (
);

FILL FILL_5__13436_ (
);

FILL FILL_3__14890_ (
);

FILL FILL_3__14470_ (
);

FILL FILL_5__13016_ (
);

INVX1 _7736_ (
    .A(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_436_)
);

FILL FILL_3__14050_ (
);

INVX1 _7316_ (
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_217_)
);

FILL FILL_4__9983_ (
);

FILL FILL_4__9143_ (
);

FILL FILL_4__12849_ (
);

FILL FILL_2__13883_ (
);

FILL FILL_4__12429_ (
);

FILL FILL_2__13463_ (
);

FILL FILL_4__12009_ (
);

FILL FILL_2__13043_ (
);

FILL FILL_1__12876_ (
);

FILL FILL_1__12456_ (
);

FILL SFILL78760x77050 (
);

FILL FILL_1__12036_ (
);

FILL FILL_6_CLKBUF1_insert121 (
);

FILL FILL_0__9883_ (
);

FILL FILL_3__7980_ (
);

FILL FILL_3__7560_ (
);

FILL FILL_0__9463_ (
);

FILL FILL_0__11869_ (
);

FILL FILL_0__9043_ (
);

AOI21X1 _11734_ (
    .A(_2168_),
    .B(_2478_),
    .C(_2830_),
    .Y(_2831_)
);

FILL FILL_0__11449_ (
);

FILL FILL_6_CLKBUF1_insert127 (
);

FILL FILL_0__11029_ (
);

INVX1 _11314_ (
    .A(_2224_),
    .Y(_2433_)
);

FILL FILL_5__7486_ (
);

FILL FILL_5__7066_ (
);

FILL FILL_4__16262_ (
);

FILL FILL_3__15675_ (
);

FILL FILL_3__15255_ (
);

FILL FILL_1__7478_ (
);

FILL FILL_1__7058_ (
);

FILL FILL_3__10390_ (
);

FILL FILL_2__14668_ (
);

FILL FILL_2__14248_ (
);

FILL FILL_0__15282_ (
);

FILL SFILL28760x2050 (
);

FILL FILL_1_BUFX2_insert690 (
);

FILL FILL_3__8765_ (
);

FILL FILL_1_BUFX2_insert691 (
);

FILL FILL_3__8345_ (
);

FILL FILL_1_BUFX2_insert692 (
);

DFFSR _12939_ (
    .Q(\datapath_1.a [20]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3555_[20])
);

OAI21X1 _12519_ (
    .A(_3411_),
    .B(vdd),
    .C(_3412_),
    .Y(_3360_[26])
);

FILL FILL_1_BUFX2_insert693 (
);

FILL FILL_1_BUFX2_insert694 (
);

FILL FILL_1_BUFX2_insert695 (
);

FILL FILL_1_BUFX2_insert696 (
);

FILL FILL_1__14602_ (
);

FILL FILL_1_BUFX2_insert697 (
);

FILL FILL_1_BUFX2_insert698 (
);

FILL FILL_6__11988_ (
);

FILL FILL_1_BUFX2_insert699 (
);

FILL SFILL24360x71050 (
);

FILL FILL_4__12182_ (
);

FILL FILL_5__9632_ (
);

FILL FILL_3__11595_ (
);

FILL FILL_5__9212_ (
);

FILL FILL_3__11175_ (
);

FILL FILL_0__16067_ (
);

NAND2X1 _16352_ (
    .A(gnd),
    .B(gnd),
    .Y(_6789_)
);

FILL FILL112360x44050 (
);

FILL FILL_2__10168_ (
);

FILL FILL_5__11922_ (
);

FILL FILL_1__9624_ (
);

FILL FILL_5__11502_ (
);

FILL FILL_4__10915_ (
);

FILL SFILL64040x53050 (
);

FILL FILL_5__14394_ (
);

FILL FILL_6__7555_ (
);

INVX1 _8694_ (
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_976_)
);

FILL FILL_1__15807_ (
);

OAI21X1 _8274_ (
    .A(_712_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .C(_713_),
    .Y(_653_[30])
);

FILL FILL_1__10942_ (
);

FILL FILL_4__13387_ (
);

FILL FILL_1__10522_ (
);

FILL FILL_1__10102_ (
);

FILL FILL_2__7967_ (
);

FILL FILL_2__7547_ (
);

BUFX2 BUFX2_insert360 (
    .A(_2470_),
    .Y(_2470__bF$buf3)
);

BUFX2 BUFX2_insert361 (
    .A(_2470_),
    .Y(_2470__bF$buf2)
);

BUFX2 BUFX2_insert362 (
    .A(_2470_),
    .Y(_2470__bF$buf1)
);

BUFX2 BUFX2_insert363 (
    .A(_2470_),
    .Y(_2470__bF$buf0)
);

BUFX2 BUFX2_insert364 (
    .A(_3998_),
    .Y(_3998__bF$buf3)
);

BUFX2 BUFX2_insert365 (
    .A(_3998_),
    .Y(_3998__bF$buf2)
);

BUFX2 BUFX2_insert366 (
    .A(_3998_),
    .Y(_3998__bF$buf1)
);

BUFX2 BUFX2_insert367 (
    .A(_3998_),
    .Y(_3998__bF$buf0)
);

BUFX2 BUFX2_insert368 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf7 )
);

DFFSR _12692_ (
    .Q(\datapath_1.Data [29]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3425_[29])
);

BUFX2 BUFX2_insert369 (
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf6 )
);

NAND3X1 _12272_ (
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [16]),
    .C(_3198__bF$buf2),
    .Y(_3243_)
);

FILL FILL_5__12707_ (
);

FILL FILL_3__13741_ (
);

FILL FILL_3__13321_ (
);

FILL FILL_6__16186_ (
);

FILL FILL_4__8834_ (
);

FILL FILL_2__12734_ (
);

FILL FILL_5__15599_ (
);

FILL FILL_5__15179_ (
);

FILL FILL_2__12314_ (
);

OAI21X1 _9899_ (
    .A(_1531_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .C(_1532_),
    .Y(_1498_[17])
);

OAI21X1 _9479_ (
    .A(_1312_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .C(_1313_),
    .Y(_1303_[5])
);

DFFSR _9059_ (
    .Q(\datapath_1.regfile_1.regOut[17] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_1043_[13])
);

FILL FILL_1__11727_ (
);

FILL FILL_1__11307_ (
);

FILL FILL_5__16120_ (
);

FILL FILL_0__8734_ (
);

FILL FILL_0__8314_ (
);

FILL FILL_1__14199_ (
);

FILL FILL_4__15953_ (
);

FILL FILL_4__15533_ (
);

FILL FILL_4__15113_ (
);

NAND3X1 _13897_ (
    .A(_4398_),
    .B(_4399_),
    .C(_4397_),
    .Y(_4400_)
);

INVX1 _13477_ (
    .A(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_3988_)
);

DFFSR _13057_ (
    .Q(_2_[10]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_3620_[10])
);

FILL FILL_3__14946_ (
);

FILL FILL_1__15980_ (
);

FILL FILL_3__14526_ (
);

FILL FILL_1__15560_ (
);

FILL FILL_3__14106_ (
);

FILL FILL_1__15140_ (
);

FILL FILL_4__9619_ (
);

FILL FILL_2__13939_ (
);

FILL FILL_0__14973_ (
);

FILL FILL_2__13519_ (
);

FILL FILL_0__14553_ (
);

FILL FILL_0__14133_ (
);

FILL FILL_5__11099_ (
);

FILL SFILL54040x51050 (
);

FILL FILL_0__9939_ (
);

FILL FILL_3__7616_ (
);

FILL FILL_0__9519_ (
);

FILL FILL_5__12880_ (
);

FILL FILL_5__12460_ (
);

FILL FILL_5__12040_ (
);

FILL FILL_4__16318_ (
);

FILL FILL_4__11873_ (
);

FILL FILL_6__10419_ (
);

FILL FILL_4__11453_ (
);

FILL FILL_4__11033_ (
);

FILL FILL_1__16345_ (
);

FILL FILL_5__8903_ (
);

FILL FILL_3__10446_ (
);

FILL FILL_3__10026_ (
);

FILL FILL_1__11480_ (
);

FILL FILL_1__11060_ (
);

FILL FILL_0__15758_ (
);

INVX1 _15623_ (
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_6089_)
);

FILL FILL_0__15338_ (
);

OAI21X1 _15203_ (
    .A(_4108_),
    .B(_5535__bF$buf0),
    .C(_5679_),
    .Y(_5680_)
);

FILL SFILL94520x16050 (
);

FILL FILL_0__10893_ (
);

FILL FILL_2__8085_ (
);

FILL FILL_0__10053_ (
);

FILL FILL_6__14672_ (
);

FILL FILL_6__14252_ (
);

FILL FILL_4__6900_ (
);

FILL FILL_5__13665_ (
);

FILL FILL_2__10800_ (
);

FILL FILL_5__13245_ (
);

INVX1 _7965_ (
    .A(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_548_)
);

INVX1 _7545_ (
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_329_)
);

OAI21X1 _7125_ (
    .A(_129_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_130_),
    .Y(_68_[31])
);

FILL FILL_4__9792_ (
);

FILL FILL_4__9372_ (
);

FILL FILL_4__12658_ (
);

FILL FILL_4__12238_ (
);

FILL FILL_2__13692_ (
);

FILL FILL_2__13272_ (
);

FILL FILL_1__12265_ (
);

INVX1 _16408_ (
    .A(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_6826_)
);

NAND2X1 _11963_ (
    .A(IorD_bF$buf6),
    .B(ALUOut[25]),
    .Y(_3017_)
);

FILL FILL_0__9272_ (
);

FILL FILL_0__11678_ (
);

NAND3X1 _11543_ (
    .A(_2462__bF$buf1),
    .B(_2652_),
    .C(_2632_),
    .Y(_2653_)
);

FILL FILL_0__11258_ (
);

INVX1 _11123_ (
    .A(\datapath_1.alu_1.ALUInA [19]),
    .Y(_2242_)
);

FILL FILL_5_CLKBUF1_insert111 (
);

FILL FILL_5_CLKBUF1_insert112 (
);

FILL FILL_5__7295_ (
);

FILL FILL_5_CLKBUF1_insert113 (
);

FILL FILL_5_CLKBUF1_insert114 (
);

FILL FILL_4__16071_ (
);

FILL FILL_5_CLKBUF1_insert115 (
);

FILL FILL_5_CLKBUF1_insert116 (
);

FILL FILL_5_CLKBUF1_insert117 (
);

FILL FILL_5_CLKBUF1_insert118 (
);

FILL FILL_5_CLKBUF1_insert119 (
);

FILL FILL_3__15484_ (
);

FILL FILL_3__15064_ (
);

FILL FILL_1__7287_ (
);

FILL SFILL23480x29050 (
);

FILL FILL_2__14897_ (
);

FILL FILL_2__14477_ (
);

FILL FILL_6_BUFX2_insert904 (
);

FILL FILL_2__14057_ (
);

FILL FILL_0__15091_ (
);

FILL FILL_5__15811_ (
);

FILL FILL_6_BUFX2_insert909 (
);

FILL FILL_4__14804_ (
);

FILL FILL_3__8994_ (
);

FILL FILL_3__8574_ (
);

OAI21X1 _12748_ (
    .A(_3523_),
    .B(IRWrite_bF$buf5),
    .C(_3524_),
    .Y(_3490_[17])
);

NAND3X1 _12328_ (
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf0),
    .Y(_3285_)
);

FILL FILL_1__14831_ (
);

FILL FILL_1__14411_ (
);

FILL FILL_0__13824_ (
);

FILL FILL_0__13404_ (
);

FILL FILL_3__16269_ (
);

FILL FILL_2__6991_ (
);

FILL FILL_5__9861_ (
);

FILL FILL_5__9021_ (
);

FILL FILL_0__16296_ (
);

NOR2X1 _16161_ (
    .A(_6611_),
    .B(_6613_),
    .Y(_6614_)
);

FILL FILL_2__10397_ (
);

FILL FILL_5__11731_ (
);

FILL FILL_1__9853_ (
);

FILL FILL_5__11311_ (
);

FILL FILL_1__9013_ (
);

FILL FILL_2__16203_ (
);

FILL FILL_3__9779_ (
);

FILL FILL_3__9359_ (
);

FILL FILL_4__10304_ (
);

FILL FILL_1__15616_ (
);

OAI21X1 _8083_ (
    .A(_605_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_606_),
    .Y(_588_[9])
);

FILL FILL_1__10751_ (
);

FILL FILL_0__14609_ (
);

FILL FILL_2__7356_ (
);

FILL FILL_3__12189_ (
);

FILL SFILL74120x43050 (
);

FILL SFILL13480x27050 (
);

AOI22X1 _12081_ (
    .A(\datapath_1.ALUResult [23]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3107_)
);

FILL FILL_5__12516_ (
);

FILL FILL_3__13970_ (
);

FILL FILL_3__13550_ (
);

FILL FILL_3__13130_ (
);

FILL FILL_4__8643_ (
);

FILL FILL_4__11929_ (
);

FILL FILL_5_BUFX2_insert920 (
);

FILL FILL_4__8223_ (
);

FILL FILL_5_BUFX2_insert921 (
);

FILL FILL_2__12963_ (
);

FILL FILL_4__11509_ (
);

FILL FILL_5_BUFX2_insert922 (
);

FILL FILL_5_BUFX2_insert923 (
);

FILL FILL_2__12123_ (
);

FILL FILL_5_BUFX2_insert924 (
);

NAND2X1 _9288_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1227_)
);

FILL FILL_5_BUFX2_insert925 (
);

FILL SFILL13800x39050 (
);

FILL FILL_5_BUFX2_insert926 (
);

FILL FILL_5_BUFX2_insert927 (
);

FILL FILL_1__11956_ (
);

FILL FILL_5_BUFX2_insert928 (
);

FILL FILL_5_BUFX2_insert929 (
);

FILL FILL_1__11536_ (
);

FILL FILL_1__11116_ (
);

FILL FILL_0__8963_ (
);

FILL FILL_0__10949_ (
);

FILL FILL_0__8123_ (
);

INVX1 _10814_ (
    .A(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_2000_)
);

FILL FILL_0__10529_ (
);

FILL FILL_0__10109_ (
);

FILL FILL_5__6986_ (
);

FILL FILL_6__14728_ (
);

FILL FILL_6__14308_ (
);

FILL FILL_4__15762_ (
);

FILL FILL_4__15342_ (
);

OR2X2 _13286_ (
    .A(_3796_),
    .B(_3824_),
    .Y(_3825_)
);

FILL FILL_2__9922_ (
);

FILL FILL_3__14755_ (
);

FILL FILL_2__9502_ (
);

FILL FILL_3__14335_ (
);

FILL FILL_1__6978_ (
);

FILL FILL_4__9848_ (
);

FILL FILL_4__9428_ (
);

FILL FILL_4__9008_ (
);

FILL FILL_2__13748_ (
);

FILL FILL_2__13328_ (
);

FILL FILL_0__14782_ (
);

FILL FILL_0__14362_ (
);

FILL FILL_3__7845_ (
);

FILL FILL_0__9748_ (
);

FILL FILL_3__7425_ (
);

FILL FILL_4__16127_ (
);

FILL FILL_4__11682_ (
);

FILL FILL_4__11262_ (
);

FILL FILL_1__16154_ (
);

FILL FILL_5__8712_ (
);

FILL FILL_3__10675_ (
);

FILL FILL_3__10255_ (
);

FILL FILL_0__15987_ (
);

FILL FILL_0__15567_ (
);

AOI21X1 _15852_ (
    .A(_6286_),
    .B(_6312_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [19])
);

FILL FILL_0__15147_ (
);

NOR2X1 _15432_ (
    .A(_5902_),
    .B(_5900_),
    .Y(_5903_)
);

NAND2X1 _15012_ (
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5492_)
);

FILL FILL_0__10282_ (
);

FILL FILL_3_BUFX2_insert1000 (
);

FILL FILL_1__8704_ (
);

FILL FILL_3_BUFX2_insert1001 (
);

FILL FILL_3_BUFX2_insert1002 (
);

FILL FILL_3_BUFX2_insert1003 (
);

FILL FILL_3_BUFX2_insert1004 (
);

FILL FILL_3_BUFX2_insert1005 (
);

FILL FILL_3_BUFX2_insert1006 (
);

FILL FILL_3_BUFX2_insert1007 (
);

FILL SFILL64040x48050 (
);

FILL FILL_3_BUFX2_insert1008 (
);

FILL FILL_5__13894_ (
);

FILL FILL_5__13474_ (
);

FILL FILL_3_BUFX2_insert1009 (
);

DFFSR _7774_ (
    .Q(\datapath_1.regfile_1.regOut[7] [8]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_393_[8])
);

OAI21X1 _7354_ (
    .A(_241_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .C(_242_),
    .Y(_198_[22])
);

FILL FILL_4__12887_ (
);

FILL FILL_4__12467_ (
);

FILL FILL_4__12047_ (
);

FILL FILL_2__13081_ (
);

FILL FILL_5__9917_ (
);

FILL FILL_1__12494_ (
);

FILL FILL_1__12074_ (
);

NOR3X1 _16217_ (
    .A(_6666_),
    .B(_6667_),
    .C(_5688_),
    .Y(_6668_)
);

FILL SFILL49560x70050 (
);

FILL FILL_2__9099_ (
);

NAND3X1 _11772_ (
    .A(_2859_),
    .B(_2860_),
    .C(_2866_),
    .Y(_2867_)
);

FILL FILL_0__9081_ (
);

FILL FILL_0__11487_ (
);

FILL FILL_0__11067_ (
);

INVX8 _11352_ (
    .A(_2458_),
    .Y(_2470_)
);

FILL FILL_1__9909_ (
);

FILL FILL_3__12401_ (
);

FILL FILL_2__11814_ (
);

FILL FILL_5__14679_ (
);

FILL FILL_5__14259_ (
);

OAI21X1 _8979_ (
    .A(_1060_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1061_),
    .Y(_1043_[9])
);

FILL FILL_3__15293_ (
);

DFFSR _8559_ (
    .Q(\datapath_1.regfile_1.regOut[13] [25]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_783_[25])
);

NAND2X1 _8139_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_644_)
);

FILL FILL_1__7096_ (
);

FILL FILL_1__10807_ (
);

FILL FILL_2__14286_ (
);

FILL FILL_5__15620_ (
);

FILL FILL_5__15200_ (
);

FILL FILL_0__7814_ (
);

OAI21X1 _9920_ (
    .A(_1545_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1546_),
    .Y(_1498_[24])
);

OAI21X1 _9500_ (
    .A(_1326_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .C(_1327_),
    .Y(_1303_[12])
);

FILL FILL_1__13699_ (
);

FILL FILL_1__13279_ (
);

FILL FILL_4__14613_ (
);

FILL FILL_3__8383_ (
);

OAI21X1 _12977_ (
    .A(_3635_),
    .B(vdd),
    .C(_3636_),
    .Y(_3620_[8])
);

DFFSR _12557_ (
    .Q(ALUOut[22]),
    .CLK(clk_bF$buf45),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3360_[22])
);

NAND2X1 _12137_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [7]),
    .Y(_3145_)
);

FILL FILL_3__13606_ (
);

FILL FILL_1__14640_ (
);

FILL FILL_1__14220_ (
);

FILL FILL_0__13633_ (
);

FILL FILL_0__13213_ (
);

FILL FILL_3__16078_ (
);

FILL SFILL54040x46050 (
);

FILL FILL_5__9670_ (
);

FILL FILL_5__10179_ (
);

FILL FILL_5__9250_ (
);

INVX1 _16390_ (
    .A(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_6814_)
);

FILL FILL_5__16405_ (
);

FILL FILL_5__11960_ (
);

FILL FILL_1__9662_ (
);

FILL FILL_5__11540_ (
);

FILL FILL_1__9242_ (
);

FILL FILL_5__11120_ (
);

FILL FILL_4__15818_ (
);

FILL FILL_2__16012_ (
);

FILL FILL_4__10953_ (
);

FILL FILL_3__9168_ (
);

FILL FILL_4__10533_ (
);

FILL FILL_4__10113_ (
);

FILL FILL_1__15845_ (
);

FILL FILL_1__15425_ (
);

FILL FILL_1__15005_ (
);

FILL FILL_1__10980_ (
);

FILL FILL_1__10560_ (
);

FILL FILL_1__10140_ (
);

FILL FILL_0__14838_ (
);

INVX1 _14703_ (
    .A(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_5189_)
);

FILL FILL_0__14418_ (
);

FILL FILL_2__7585_ (
);

BUFX2 BUFX2_insert740 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf1 )
);

BUFX2 BUFX2_insert741 (
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf0 )
);

FILL FILL_2__7165_ (
);

BUFX2 BUFX2_insert742 (
    .A(_5535_),
    .Y(_5535__bF$buf4)
);

BUFX2 BUFX2_insert743 (
    .A(_5535_),
    .Y(_5535__bF$buf3)
);

BUFX2 BUFX2_insert744 (
    .A(_5535_),
    .Y(_5535__bF$buf2)
);

BUFX2 BUFX2_insert745 (
    .A(_5535_),
    .Y(_5535__bF$buf1)
);

BUFX2 BUFX2_insert746 (
    .A(_5535_),
    .Y(_5535__bF$buf0)
);

BUFX2 BUFX2_insert747 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf7 )
);

BUFX2 BUFX2_insert748 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf6 )
);

BUFX2 BUFX2_insert749 (
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf5 )
);

FILL FILL_5__12745_ (
);

FILL FILL_5__12325_ (
);

FILL FILL_4__8872_ (
);

FILL FILL_4__8452_ (
);

FILL FILL_4__11738_ (
);

FILL FILL_2__12772_ (
);

FILL FILL_4__11318_ (
);

FILL FILL_2__12352_ (
);

NAND2X1 _9097_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1120_)
);

FILL FILL_1__11765_ (
);

FILL FILL_1__11345_ (
);

NOR2X1 _15908_ (
    .A(_6366_),
    .B(_6364_),
    .Y(_6367_)
);

FILL FILL_0__8772_ (
);

FILL FILL_0__8352_ (
);

FILL FILL_0__10758_ (
);

INVX1 _10623_ (
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_1893_)
);

DFFSR _10203_ (
    .Q(\datapath_1.regfile_1.regOut[26] [5]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_1628_[5])
);

FILL SFILL109400x76050 (
);

FILL FILL_4__15991_ (
);

FILL FILL_4__15571_ (
);

FILL SFILL44040x44050 (
);

FILL FILL_4__15151_ (
);

NAND2X1 _13095_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [5]),
    .Y(_3695_)
);

FILL FILL_3__14984_ (
);

FILL FILL_2__9731_ (
);

FILL FILL_3__14564_ (
);

FILL FILL_3__14144_ (
);

FILL FILL_4_BUFX2_insert580 (
);

FILL FILL_4_BUFX2_insert581 (
);

FILL FILL_4__9657_ (
);

FILL FILL_4_BUFX2_insert582 (
);

FILL FILL_4__9237_ (
);

FILL FILL_4_BUFX2_insert583 (
);

FILL FILL_2__13977_ (
);

FILL SFILL109000x62050 (
);

FILL FILL_4_BUFX2_insert584 (
);

FILL FILL_2__13557_ (
);

FILL FILL_0__14591_ (
);

FILL FILL_2__13137_ (
);

FILL FILL_4_BUFX2_insert585 (
);

FILL FILL_0__14171_ (
);

FILL FILL_4_BUFX2_insert586 (
);

FILL FILL_4_BUFX2_insert587 (
);

FILL FILL_4_BUFX2_insert588 (
);

FILL FILL_4_BUFX2_insert589 (
);

FILL FILL_0__9977_ (
);

FILL FILL_0__9557_ (
);

FILL FILL_0__9137_ (
);

NAND3X1 _11828_ (
    .A(_2914_),
    .B(_2915_),
    .C(_2917_),
    .Y(_2918_)
);

FILL FILL_3__7234_ (
);

INVX1 _11408_ (
    .A(_2283_),
    .Y(_2525_)
);

FILL SFILL8520x14050 (
);

FILL FILL_1__13911_ (
);

FILL FILL_4__16356_ (
);

FILL FILL_4__11491_ (
);

FILL FILL_4__11071_ (
);

FILL FILL_0__12904_ (
);

FILL FILL_3__15769_ (
);

FILL FILL_3__15349_ (
);

FILL FILL_1__16383_ (
);

FILL FILL_5__8521_ (
);

FILL FILL_3__10064_ (
);

FILL FILL_5__8101_ (
);

FILL FILL_0__15796_ (
);

FILL FILL_0__15376_ (
);

AOI22X1 _15661_ (
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_6126_)
);

NAND3X1 _15241_ (
    .A(_5707_),
    .B(_5716_),
    .C(_5710_),
    .Y(_5717_)
);

FILL FILL_5__10811_ (
);

FILL FILL_1__8513_ (
);

FILL SFILL109320x38050 (
);

FILL FILL_2__15703_ (
);

FILL FILL_3__8859_ (
);

FILL FILL_3__8439_ (
);

FILL FILL_3__8019_ (
);

FILL FILL_5__13283_ (
);

OAI21X1 _7583_ (
    .A(_353_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .C(_354_),
    .Y(_328_[13])
);

OAI21X1 _7163_ (
    .A(_134_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .C(_135_),
    .Y(_133_[1])
);

FILL SFILL99400x80050 (
);

FILL FILL_4__12696_ (
);

FILL FILL_4__12276_ (
);

FILL SFILL69160x55050 (
);

FILL FILL_3__9800_ (
);

FILL FILL_2__6856_ (
);

FILL FILL_3__11689_ (
);

FILL FILL_5__9726_ (
);

FILL FILL_3__11269_ (
);

FILL FILL_6__12603_ (
);

FILL SFILL74120x38050 (
);

DFFSR _16446_ (
    .Q(\datapath_1.regfile_1.regOut[0] [29]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_6769_[29])
);

OAI22X1 _16026_ (
    .A(_5480__bF$buf0),
    .B(_5086_),
    .C(_6481_),
    .D(_5499__bF$buf2),
    .Y(_6482_)
);

OAI21X1 _11581_ (
    .A(_2507_),
    .B(_2518_),
    .C(_2519_),
    .Y(_2688_)
);

FILL FILL_0__11296_ (
);

NOR2X1 _11161_ (
    .A(\datapath_1.alu_1.ALUInB [22]),
    .B(_2279_),
    .Y(_2280_)
);

FILL FILL_1__9718_ (
);

FILL FILL_3__12630_ (
);

FILL FILL_6__15495_ (
);

FILL FILL_3__12210_ (
);

FILL FILL_4__7723_ (
);

FILL FILL_4__7303_ (
);

FILL FILL_5__14488_ (
);

FILL FILL_2__11623_ (
);

FILL FILL_5__14068_ (
);

FILL FILL_2__11203_ (
);

NAND2X1 _8788_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_975_)
);

FILL FILL_6__7229_ (
);

NAND2X1 _8368_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_756_)
);

FILL FILL_1__10616_ (
);

FILL FILL_2__14095_ (
);

FILL FILL_0__7623_ (
);

FILL SFILL69160x10050 (
);

FILL FILL_0__7203_ (
);

FILL FILL_1__13088_ (
);

FILL FILL_4__14842_ (
);

FILL FILL_4__14422_ (
);

FILL FILL_4__14002_ (
);

NAND2X1 _12786_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[30]),
    .Y(_3550_)
);

FILL FILL_3__8192_ (
);

OAI21X1 _12366_ (
    .A(_3308_),
    .B(MemToReg_bF$buf7),
    .C(_3309_),
    .Y(\datapath_1.mux_wd3.dout [7])
);

FILL FILL_3__13835_ (
);

FILL FILL_3__13415_ (
);

FILL FILL_4__8508_ (
);

FILL FILL_2__12828_ (
);

FILL FILL_2__12408_ (
);

FILL FILL_0__13862_ (
);

FILL SFILL99320x42050 (
);

FILL FILL_0__13442_ (
);

FILL FILL_0__13022_ (
);

FILL FILL_3__6925_ (
);

FILL FILL_5__16214_ (
);

FILL FILL_0__8828_ (
);

FILL SFILL59160x53050 (
);

FILL FILL_1__9891_ (
);

FILL FILL_1__9471_ (
);

FILL FILL_4__15627_ (
);

FILL FILL_4__15207_ (
);

FILL FILL_2__16241_ (
);

FILL FILL_3__9397_ (
);

FILL FILL_4__10762_ (
);

FILL SFILL64120x36050 (
);

FILL FILL_1__15654_ (
);

FILL FILL_1__15234_ (
);

FILL FILL_0__14647_ (
);

INVX1 _14932_ (
    .A(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_5413_)
);

FILL FILL_0__14227_ (
);

NAND3X1 _14512_ (
    .A(_5000_),
    .B(_5001_),
    .C(_4997_),
    .Y(_5002_)
);

FILL SFILL68440x44050 (
);

FILL FILL_6__13981_ (
);

FILL FILL_6__13561_ (
);

FILL FILL_6__13141_ (
);

FILL FILL_5__12974_ (
);

FILL SFILL113880x47050 (
);

FILL FILL_5__12134_ (
);

BUFX2 _6854_ (
    .A(_1_[16]),
    .Y(memoryAddress[16])
);

FILL SFILL84200x3050 (
);

FILL FILL_4__11967_ (
);

FILL FILL_4__8261_ (
);

FILL FILL_4__11547_ (
);

FILL FILL_2__12581_ (
);

FILL FILL_4__11127_ (
);

FILL FILL_2__12161_ (
);

FILL FILL_1__16019_ (
);

FILL FILL_1__11994_ (
);

FILL FILL_1__11574_ (
);

FILL FILL_1__11154_ (
);

NOR2X1 _15717_ (
    .A(_6180_),
    .B(_5501_),
    .Y(_6181_)
);

FILL SFILL33960x80050 (
);

FILL FILL_2__8599_ (
);

FILL FILL_0__8581_ (
);

DFFSR _10852_ (
    .Q(\datapath_1.regfile_1.regOut[31] [14]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_1953_[14])
);

FILL FILL_0__10567_ (
);

OAI21X1 _10432_ (
    .A(_1805_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1806_),
    .Y(_1758_[24])
);

FILL FILL_0__10147_ (
);

FILL SFILL89320x40050 (
);

OAI21X1 _10012_ (
    .A(_1586_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .C(_1587_),
    .Y(_1563_[12])
);

FILL SFILL28680x24050 (
);

FILL FILL_3__11901_ (
);

FILL FILL_4__15380_ (
);

FILL FILL_5__13759_ (
);

FILL FILL_5__13339_ (
);

FILL FILL_3__14793_ (
);

FILL FILL_2__9540_ (
);

FILL FILL_2__9120_ (
);

FILL FILL_3__14373_ (
);

DFFSR _7639_ (
    .Q(\datapath_1.regfile_1.regOut[6] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_328_[1])
);

NAND2X1 _7219_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_173_)
);

FILL FILL_4__9886_ (
);

FILL FILL_4__9466_ (
);

FILL FILL_2__13786_ (
);

FILL FILL_2__13366_ (
);

FILL FILL_5__14700_ (
);

FILL SFILL54120x34050 (
);

FILL FILL_1__12779_ (
);

FILL FILL_1__12359_ (
);

FILL FILL_3__7883_ (
);

FILL FILL_0__9786_ (
);

FILL FILL_3__7463_ (
);

FILL FILL_0__9366_ (
);

FILL FILL_3__7043_ (
);

OAI21X1 _11637_ (
    .A(_2720_),
    .B(_2408_),
    .C(_2740_),
    .Y(_2741_)
);

NOR2X1 _11217_ (
    .A(gnd),
    .B(_2335_),
    .Y(_2336_)
);

FILL FILL_1__13720_ (
);

FILL FILL_1__13300_ (
);

FILL FILL_4__16165_ (
);

FILL FILL_3__15998_ (
);

FILL FILL_0__12713_ (
);

FILL FILL_3__15578_ (
);

FILL FILL_3__15158_ (
);

FILL FILL_1__16192_ (
);

FILL FILL_5__8750_ (
);

FILL FILL_3__10293_ (
);

FILL FILL_5__8330_ (
);

NOR3X1 _15890_ (
    .A(_6337_),
    .B(_6327_),
    .C(_6349_),
    .Y(_6350_)
);

FILL FILL_0__15185_ (
);

OAI22X1 _15470_ (
    .A(_4459_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf3),
    .D(_4456_),
    .Y(_5940_)
);

FILL FILL_5__15905_ (
);

NAND3X1 _15050_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5468_),
    .C(_5471__bF$buf5),
    .Y(_5530_)
);

FILL FILL_1__8742_ (
);

FILL FILL_5__10620_ (
);

FILL FILL_1__8322_ (
);

FILL FILL_2__15932_ (
);

FILL FILL_2__15512_ (
);

FILL FILL_3__8248_ (
);

FILL FILL_5__13092_ (
);

FILL FILL_1__14925_ (
);

FILL FILL_1__14505_ (
);

DFFSR _7392_ (
    .Q(\datapath_1.regfile_1.regOut[4] [10]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_198_[10])
);

FILL SFILL18680x22050 (
);

FILL FILL_4__12085_ (
);

FILL FILL_0__13918_ (
);

FILL FILL_5__9535_ (
);

FILL FILL_3__11498_ (
);

FILL FILL_5__9115_ (
);

FILL FILL_3__11078_ (
);

FILL FILL111960x51050 (
);

INVX1 _16255_ (
    .A(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_6705_)
);

AOI21X1 _11390_ (
    .A(_2496_),
    .B(_2502_),
    .C(_2506_),
    .Y(_2507_)
);

FILL FILL_5__11825_ (
);

FILL FILL_1__9527_ (
);

FILL FILL_5__11405_ (
);

FILL FILL_1__9107_ (
);

FILL SFILL79240x45050 (
);

FILL FILL_4__7952_ (
);

FILL FILL_4__7112_ (
);

FILL FILL_4__10818_ (
);

FILL FILL_2__11852_ (
);

FILL FILL_5__14297_ (
);

FILL FILL_2__11432_ (
);

FILL FILL_2__11012_ (
);

NAND2X1 _8597_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_868_)
);

DFFSR _8177_ (
    .Q(\datapath_1.regfile_1.regOut[10] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_588_[27])
);

FILL FILL_6__7038_ (
);

FILL FILL_1__10425_ (
);

FILL FILL_1__10005_ (
);

FILL FILL_0__7852_ (
);

FILL FILL_0__7432_ (
);

FILL SFILL44040x39050 (
);

FILL FILL_4__14651_ (
);

FILL FILL_4__14231_ (
);

FILL SFILL94360x5050 (
);

NAND2X1 _12595_ (
    .A(vdd),
    .B(memoryOutData[9]),
    .Y(_3443_)
);

INVX1 _12175_ (
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3170_)
);

FILL FILL_3__13644_ (
);

FILL FILL_3__13224_ (
);

FILL FILL_6__16089_ (
);

FILL FILL_4__8737_ (
);

FILL FILL_4__8317_ (
);

FILL FILL_2__12637_ (
);

FILL FILL_0__13671_ (
);

FILL FILL_2__12217_ (
);

FILL FILL_0__13251_ (
);

FILL FILL111880x13050 (
);

FILL FILL_0__8637_ (
);

FILL FILL_5__16023_ (
);

NOR2X1 _10908_ (
    .A(_2053_),
    .B(_2054_),
    .Y(ALUOp[1])
);

FILL FILL_0__8217_ (
);

FILL SFILL104520x8050 (
);

FILL FILL_1__9280_ (
);

FILL FILL_4__15856_ (
);

FILL FILL_4__15436_ (
);

FILL FILL_4__15016_ (
);

FILL FILL_2__16050_ (
);

FILL FILL_4__10991_ (
);

FILL FILL_4__10571_ (
);

FILL FILL_4__10151_ (
);

FILL FILL_3__14849_ (
);

FILL FILL_1__15883_ (
);

FILL FILL_3__14429_ (
);

FILL FILL_3__14009_ (
);

FILL FILL_1__15463_ (
);

FILL FILL_1__15043_ (
);

FILL FILL_5__7601_ (
);

FILL FILL_0__14876_ (
);

FILL SFILL69240x43050 (
);

FILL FILL_0__14456_ (
);

NOR2X1 _14741_ (
    .A(_5216_),
    .B(_5226_),
    .Y(_5227_)
);

FILL FILL_0__14036_ (
);

NOR2X1 _14321_ (
    .A(_4811_),
    .B(_4814_),
    .Y(_4815_)
);

FILL FILL_3__7939_ (
);

FILL FILL_5__12783_ (
);

FILL FILL_5__12363_ (
);

FILL SFILL99400x75050 (
);

FILL FILL_4__8490_ (
);

FILL FILL_4__11776_ (
);

FILL FILL_4__8070_ (
);

FILL FILL_4__11356_ (
);

FILL FILL_2__12390_ (
);

FILL FILL_1__16248_ (
);

FILL FILL_3__10769_ (
);

FILL FILL_1__11383_ (
);

OAI21X1 _15946_ (
    .A(_5524__bF$buf1),
    .B(_5007_),
    .C(_6403_),
    .Y(_6404_)
);

INVX1 _15526_ (
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_5995_)
);

OAI22X1 _15106_ (
    .A(_5530__bF$buf0),
    .B(_5584_),
    .C(_5532__bF$buf1),
    .D(_4019_),
    .Y(_5585_)
);

FILL FILL_0__8390_ (
);

FILL FILL_0__10796_ (
);

OAI21X1 _10661_ (
    .A(_1917_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .C(_1918_),
    .Y(_1888_[15])
);

FILL FILL_0__10376_ (
);

OAI21X1 _10241_ (
    .A(_1698_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1699_),
    .Y(_1693_[3])
);

FILL FILL_3__11710_ (
);

FILL FILL_6__14155_ (
);

FILL FILL_5__13988_ (
);

FILL FILL_2__10703_ (
);

FILL FILL_5__13568_ (
);

FILL FILL_5__13148_ (
);

NAND2X1 _7868_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_504_)
);

FILL FILL_3__14182_ (
);

NAND2X1 _7448_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_285_)
);

DFFSR _7028_ (
    .Q(\datapath_1.regfile_1.regOut[1] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_3_[30])
);

FILL FILL_4_BUFX2_insert960 (
);

FILL FILL_4_BUFX2_insert961 (
);

FILL FILL_4_BUFX2_insert962 (
);

FILL FILL_4__9275_ (
);

FILL FILL_4_BUFX2_insert963 (
);

FILL FILL_2__13595_ (
);

FILL FILL_4_BUFX2_insert964 (
);

FILL FILL_4_BUFX2_insert965 (
);

FILL FILL_4_BUFX2_insert966 (
);

FILL SFILL99400x30050 (
);

FILL FILL_4_BUFX2_insert967 (
);

FILL SFILL38760x14050 (
);

FILL FILL_4_BUFX2_insert968 (
);

FILL FILL_4_BUFX2_insert969 (
);

FILL FILL_1__12588_ (
);

FILL FILL_1__12168_ (
);

FILL FILL_4__13922_ (
);

FILL FILL_4__13502_ (
);

FILL FILL_3__7692_ (
);

FILL FILL_0__9595_ (
);

NOR2X1 _11866_ (
    .A(\datapath_1.ALUResult [28]),
    .B(\datapath_1.ALUResult [26]),
    .Y(_2953_)
);

NAND2X1 _11446_ (
    .A(_2559_),
    .B(_2561_),
    .Y(_2562_)
);

OAI22X1 _11026_ (
    .A(_2141_),
    .B(_2142_),
    .C(_2143_),
    .D(_2144_),
    .Y(_2145_)
);

FILL FILL_3__12915_ (
);

FILL FILL_4__16394_ (
);

FILL FILL_5__7198_ (
);

FILL FILL_2__11908_ (
);

FILL SFILL99320x37050 (
);

FILL FILL_3__15387_ (
);

FILL FILL_0__12522_ (
);

FILL FILL_0__12102_ (
);

FILL SFILL23800x9050 (
);

FILL FILL_5__15714_ (
);

FILL SFILL28760x57050 (
);

FILL SFILL59160x48050 (
);

FILL FILL_1__8971_ (
);

FILL FILL_1__8131_ (
);

FILL FILL_4__14707_ (
);

FILL FILL_2__15741_ (
);

FILL FILL_2__15321_ (
);

FILL FILL_3__8897_ (
);

FILL FILL_3__8477_ (
);

FILL FILL_3__8057_ (
);

FILL FILL_1__14734_ (
);

FILL FILL_1__14314_ (
);

FILL SFILL28360x43050 (
);

FILL FILL_0__13727_ (
);

FILL FILL_0__13307_ (
);

FILL FILL_2__6894_ (
);

FILL FILL_5__9764_ (
);

FILL FILL_5__9344_ (
);

FILL FILL_0__16199_ (
);

FILL FILL_0_BUFX2_insert1084 (
);

OAI22X1 _16064_ (
    .A(_6518_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf3),
    .D(_5150_),
    .Y(_6519_)
);

FILL FILL_0_BUFX2_insert1085 (
);

FILL FILL_0_BUFX2_insert1086 (
);

FILL FILL_0_BUFX2_insert1087 (
);

FILL FILL_0_BUFX2_insert1088 (
);

FILL FILL_0_BUFX2_insert1089 (
);

FILL FILL_1__9756_ (
);

FILL FILL_5__11634_ (
);

FILL FILL_1__9336_ (
);

FILL FILL_5__11214_ (
);

FILL FILL_3_BUFX2_insert980 (
);

FILL FILL_2__16106_ (
);

FILL FILL_4__7761_ (
);

FILL FILL_4__7341_ (
);

FILL FILL_3_BUFX2_insert981 (
);

FILL FILL_4__10627_ (
);

FILL FILL_3_BUFX2_insert982 (
);

FILL FILL_3_BUFX2_insert983 (
);

FILL FILL_2__11661_ (
);

FILL FILL_3_BUFX2_insert984 (
);

FILL FILL_2__11241_ (
);

FILL FILL_1__15939_ (
);

FILL FILL_3_BUFX2_insert985 (
);

FILL FILL_3_BUFX2_insert986 (
);

FILL FILL_1__15519_ (
);

FILL FILL_3_BUFX2_insert987 (
);

FILL FILL_3_BUFX2_insert988 (
);

FILL FILL_3_BUFX2_insert989 (
);

FILL FILL_1__10654_ (
);

FILL FILL_4__13099_ (
);

FILL FILL_1__10234_ (
);

FILL FILL_2__7679_ (
);

FILL FILL_0__7241_ (
);

FILL SFILL89320x35050 (
);

FILL SFILL28680x19050 (
);

FILL FILL_4__14880_ (
);

FILL FILL_4__14460_ (
);

FILL FILL_6__13006_ (
);

FILL FILL_4__14040_ (
);

FILL FILL_5__12839_ (
);

FILL FILL_3__13873_ (
);

FILL FILL_5__12419_ (
);

FILL FILL_2__8620_ (
);

FILL FILL_2__8200_ (
);

FILL FILL_3__13453_ (
);

FILL SFILL18760x55050 (
);

FILL FILL_3__13033_ (
);

FILL FILL_4__8966_ (
);

FILL FILL_4__8126_ (
);

FILL FILL_2__12866_ (
);

FILL FILL_2__12446_ (
);

FILL FILL_2__12026_ (
);

FILL FILL_0__13480_ (
);

FILL SFILL54120x29050 (
);

FILL FILL_1__11859_ (
);

FILL FILL_1__11439_ (
);

FILL FILL_1__11019_ (
);

FILL FILL_0__8866_ (
);

FILL FILL_5__16252_ (
);

FILL FILL_3__6963_ (
);

FILL FILL_0__8446_ (
);

DFFSR _10717_ (
    .Q(\datapath_1.regfile_1.regOut[30] [7]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1888_[7])
);

FILL SFILL79320x78050 (
);

FILL FILL_5__6889_ (
);

FILL FILL_4__15665_ (
);

FILL FILL_4__15245_ (
);

FILL FILL_4__10380_ (
);

DFFSR _13189_ (
    .Q(\datapath_1.mux_iord.din0 [14]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3685_[14])
);

FILL FILL_2__9405_ (
);

FILL FILL_3__14658_ (
);

FILL FILL_3__14238_ (
);

FILL FILL_1__15692_ (
);

FILL FILL_1__15272_ (
);

FILL FILL_5__7830_ (
);

FILL SFILL18760x10050 (
);

INVX1 _14970_ (
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_5451_)
);

FILL FILL_0__14685_ (
);

INVX1 _14550_ (
    .A(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_5039_)
);

FILL FILL_0__14265_ (
);

AOI22X1 _14130_ (
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .B(_4005__bF$buf2),
    .C(_3950__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_4628_)
);

FILL FILL_1__7822_ (
);

FILL FILL_3__7748_ (
);

FILL FILL_3__7328_ (
);

FILL FILL_5__12592_ (
);

FILL FILL_5__12172_ (
);

BUFX2 _6892_ (
    .A(_2_[22]),
    .Y(memoryWriteData[22])
);

FILL SFILL18680x17050 (
);

FILL SFILL59000x4050 (
);

FILL FILL_4__11585_ (
);

FILL FILL_4__11165_ (
);

FILL FILL_1__16057_ (
);

FILL FILL_3__10998_ (
);

FILL SFILL33640x5050 (
);

FILL FILL_5__8615_ (
);

FILL FILL_6_BUFX2_insert490 (
);

FILL FILL_3__10578_ (
);

FILL FILL111960x46050 (
);

FILL FILL_3__10158_ (
);

FILL FILL_1__11192_ (
);

INVX1 _15755_ (
    .A(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_6218_)
);

NOR2X1 _15335_ (
    .A(_5805_),
    .B(_5808_),
    .Y(_5809_)
);

FILL FILL_6_BUFX2_insert495 (
);

INVX1 _10890_ (
    .A(ALUOp[1]),
    .Y(_2036_)
);

DFFSR _10470_ (
    .Q(\datapath_1.regfile_1.regOut[28] [16]),
    .CLK(clk_bF$buf6),
    .R(rst_bF$buf89),
    .S(vdd),
    .D(_1758_[16])
);

FILL FILL_0__10185_ (
);

FILL FILL_5__10905_ (
);

NAND2X1 _10050_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1613_)
);

FILL FILL_1__8607_ (
);

FILL FILL_0__16411_ (
);

FILL FILL_2__10932_ (
);

FILL FILL_5__13797_ (
);

FILL FILL_2__10512_ (
);

FILL FILL_5__13377_ (
);

NAND2X1 _7677_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_397_)
);

DFFSR _7257_ (
    .Q(\datapath_1.regfile_1.regOut[3] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_133_[3])
);

FILL FILL_4__9084_ (
);

FILL FILL_0__6932_ (
);

FILL FILL_1__12397_ (
);

FILL FILL_4__13731_ (
);

FILL FILL_4__13311_ (
);

FILL FILL_3__7081_ (
);

INVX1 _11675_ (
    .A(_2776_),
    .Y(\datapath_1.ALUResult [14])
);

AOI21X1 _11255_ (
    .A(_2138_),
    .B(_2373_),
    .C(_2136_),
    .Y(_2374_)
);

FILL FILL_3__12724_ (
);

FILL FILL_3__12304_ (
);

FILL FILL_4__7817_ (
);

FILL FILL_2__11717_ (
);

FILL FILL_0__12751_ (
);

FILL FILL_3__15196_ (
);

FILL FILL_0__12331_ (
);

FILL FILL_2__14189_ (
);

FILL FILL_5__15943_ (
);

FILL FILL_5__15523_ (
);

FILL FILL_0__7717_ (
);

FILL FILL_5__15103_ (
);

DFFSR _9823_ (
    .Q(\datapath_1.regfile_1.regOut[23] [9]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_1433_[9])
);

INVX1 _9403_ (
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_1283_)
);

FILL FILL_1__8780_ (
);

FILL FILL_1__8360_ (
);

FILL FILL_4__14936_ (
);

FILL FILL_2__15970_ (
);

FILL FILL_4__14516_ (
);

FILL FILL_2__15550_ (
);

FILL FILL_2__15130_ (
);

FILL SFILL29160x42050 (
);

FILL FILL_3__13929_ (
);

FILL FILL_1__14963_ (
);

FILL FILL_3__13509_ (
);

FILL FILL_1__14543_ (
);

FILL FILL_1__14123_ (
);

FILL FILL_0__13956_ (
);

OAI22X1 _13821_ (
    .A(_4325_),
    .B(_3941_),
    .C(_3960_),
    .D(_4324_),
    .Y(_4326_)
);

FILL FILL_0__13536_ (
);

NAND3X1 _13401_ (
    .A(_3886_),
    .B(_3895_),
    .C(_3912_),
    .Y(_3913_)
);

FILL FILL_0__13116_ (
);

FILL FILL_5__9993_ (
);

FILL FILL_5__9153_ (
);

AOI22X1 _16293_ (
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [31]),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_6742_)
);

FILL FILL_5__16308_ (
);

FILL FILL_1__9985_ (
);

FILL FILL_5__11863_ (
);

FILL FILL_5__11443_ (
);

FILL FILL_1__9145_ (
);

FILL FILL_5__11023_ (
);

FILL FILL_4__7990_ (
);

FILL FILL_2__16335_ (
);

FILL FILL_4__7570_ (
);

FILL SFILL104760x77050 (
);

FILL FILL_4__10436_ (
);

FILL FILL_2__11890_ (
);

FILL FILL_4__10016_ (
);

FILL FILL_2__11470_ (
);

FILL FILL_2__11050_ (
);

FILL FILL_1__15748_ (
);

FILL FILL_1__15328_ (
);

FILL FILL_1__10883_ (
);

FILL FILL_1__10043_ (
);

AOI22X1 _14606_ (
    .A(\datapath_1.regfile_1.regOut[2] [24]),
    .B(_3998__bF$buf2),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_5094_)
);

FILL FILL_0__7890_ (
);

FILL FILL_2__7488_ (
);

FILL FILL_0__7470_ (
);

FILL FILL_0__7050_ (
);

FILL FILL_2__7068_ (
);

FILL SFILL43880x2050 (
);

FILL FILL_5__12648_ (
);

FILL FILL_3__13682_ (
);

FILL FILL_5__12228_ (
);

FILL FILL_3__13262_ (
);

NAND2X1 _6948_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_33_)
);

FILL FILL_4__8775_ (
);

FILL FILL_4__8355_ (
);

FILL SFILL8600x2050 (
);

FILL FILL_2__12255_ (
);

FILL FILL_1__11668_ (
);

FILL FILL_1__11248_ (
);

FILL FILL_5__16061_ (
);

FILL FILL_0__8255_ (
);

NAND2X1 _10946_ (
    .A(_2055_),
    .B(_2059_),
    .Y(_2079_)
);

NAND2X1 _10526_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1849_)
);

NAND2X1 _10106_ (
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1630_)
);

FILL FILL_4__15894_ (
);

FILL FILL_4__15474_ (
);

FILL FILL_4__15054_ (
);

FILL FILL_2__9634_ (
);

FILL FILL_3__14887_ (
);

FILL FILL_3__14467_ (
);

FILL FILL_2__9214_ (
);

FILL FILL_0__11602_ (
);

FILL FILL_3__14047_ (
);

FILL FILL_1__15081_ (
);

FILL FILL_0__14494_ (
);

FILL SFILL89400x68050 (
);

FILL FILL_0__14074_ (
);

FILL FILL_1__7631_ (
);

FILL SFILL104280x25050 (
);

FILL FILL_1__7211_ (
);

FILL FILL_2__14821_ (
);

FILL FILL_2__14401_ (
);

FILL FILL_3__7977_ (
);

FILL FILL_3__7557_ (
);

FILL FILL_1__13814_ (
);

FILL FILL_4__16259_ (
);

FILL FILL_4__11394_ (
);

FILL FILL_1__16286_ (
);

FILL FILL_5__8844_ (
);

FILL FILL_3__10387_ (
);

FILL FILL_5__8004_ (
);

NOR2X1 _15984_ (
    .A(_6440_),
    .B(_6433_),
    .Y(_6441_)
);

FILL FILL_0__15699_ (
);

NOR2X1 _15564_ (
    .A(_6030_),
    .B(_6031_),
    .Y(_6032_)
);

FILL FILL_0__15279_ (
);

NOR2X1 _15144_ (
    .A(_5621_),
    .B(_5614_),
    .Y(_5622_)
);

FILL FILL_1__8836_ (
);

FILL SFILL94280x74050 (
);

FILL FILL_2__15606_ (
);

FILL FILL_4__6841_ (
);

FILL FILL_0__16220_ (
);

FILL FILL_2__10321_ (
);

INVX1 _7486_ (
    .A(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_310_)
);

INVX1 _7066_ (
    .A(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_91_)
);

FILL FILL_4__12599_ (
);

FILL FILL_4__12179_ (
);

FILL FILL_5__9629_ (
);

FILL FILL_5__9209_ (
);

FILL FILL_4__13960_ (
);

FILL FILL_4__13540_ (
);

NAND2X1 _16349_ (
    .A(gnd),
    .B(gnd),
    .Y(_6787_)
);

FILL FILL_4__13120_ (
);

FILL FILL_0__11199_ (
);

OAI22X1 _11484_ (
    .A(_2286_),
    .B(_2346_),
    .C(_2347__bF$buf0),
    .D(_2285_),
    .Y(_2598_)
);

FILL FILL_5__11919_ (
);

INVX2 _11064_ (
    .A(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2183_)
);

FILL FILL_3__12953_ (
);

FILL FILL_2__7700_ (
);

FILL FILL_6__15398_ (
);

FILL FILL_3__12533_ (
);

FILL FILL_3__12113_ (
);

FILL FILL_4__7626_ (
);

FILL FILL_4__7206_ (
);

FILL FILL_2__11946_ (
);

FILL FILL_0__12980_ (
);

FILL FILL_2__11526_ (
);

FILL FILL_2__11106_ (
);

FILL FILL_0__12140_ (
);

FILL FILL_1__10939_ (
);

FILL FILL_1__10519_ (
);

FILL FILL_5__15752_ (
);

FILL FILL_0__7946_ (
);

FILL FILL_5__15332_ (
);

FILL FILL_6__8913_ (
);

INVX1 _9632_ (
    .A(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_1395_)
);

FILL FILL_0__7106_ (
);

INVX1 _9212_ (
    .A(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_1176_)
);

FILL FILL_4__14745_ (
);

FILL FILL_4__14325_ (
);

DFFSR _12689_ (
    .Q(\datapath_1.Data [26]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_3425_[26])
);

FILL FILL_3__8095_ (
);

AOI22X1 _12269_ (
    .A(_2_[13]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump [13]),
    .Y(_3241_)
);

FILL FILL_2__8905_ (
);

FILL FILL_3__13738_ (
);

FILL FILL_3__13318_ (
);

FILL FILL_1__14772_ (
);

FILL FILL_1__14352_ (
);

FILL FILL_5__6910_ (
);

FILL FILL_0__13765_ (
);

FILL FILL_0__13345_ (
);

OAI22X1 _13630_ (
    .A(_4137_),
    .B(_3925_),
    .C(_3881_),
    .D(_4138_),
    .Y(_4139_)
);

NAND2X1 _13210_ (
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_3753_)
);

FILL FILL_5__9382_ (
);

FILL FILL_1__6902_ (
);

FILL FILL_5__16117_ (
);

FILL FILL_1__9794_ (
);

FILL FILL_5__11672_ (
);

FILL FILL_5__11252_ (
);

FILL FILL_1__9374_ (
);

FILL SFILL79320x28050 (
);

FILL FILL_2__16144_ (
);

FILL FILL_4__10665_ (
);

FILL FILL_4__10245_ (
);

FILL FILL_1__15977_ (
);

FILL FILL_1__15557_ (
);

FILL FILL_1__15137_ (
);

FILL FILL_1__10692_ (
);

FILL SFILL84200x70050 (
);

FILL FILL_1__10272_ (
);

FILL SFILL105160x62050 (
);

AOI22X1 _14835_ (
    .A(\datapath_1.regfile_1.regOut[3] [29]),
    .B(_3942__bF$buf1),
    .C(_3891__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_5318_)
);

INVX1 _14415_ (
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_4907_)
);

FILL FILL_2__7297_ (
);

FILL FILL_6__13884_ (
);

FILL FILL_6__13464_ (
);

FILL FILL_0__15911_ (
);

FILL FILL_5__12877_ (
);

FILL FILL_5__12457_ (
);

FILL FILL_5__12037_ (
);

FILL FILL_3__13491_ (
);

FILL FILL_4__8584_ (
);

FILL FILL_2__12484_ (
);

FILL SFILL114440x53050 (
);

FILL FILL_2__12064_ (
);

FILL FILL_2_BUFX2_insert1010 (
);

FILL FILL_2_BUFX2_insert1011 (
);

FILL FILL_1__11897_ (
);

FILL FILL_2_BUFX2_insert1012 (
);

FILL FILL_2_BUFX2_insert1013 (
);

FILL FILL_1__11477_ (
);

FILL FILL_2_BUFX2_insert1014 (
);

FILL FILL_1__11057_ (
);

FILL FILL_2_BUFX2_insert1015 (
);

FILL FILL_2_BUFX2_insert1016 (
);

FILL FILL_2_BUFX2_insert1017 (
);

FILL FILL_2_BUFX2_insert1018 (
);

FILL FILL_5__16290_ (
);

FILL FILL_0__8484_ (
);

FILL FILL_2_BUFX2_insert1019 (
);

FILL SFILL74280x70050 (
);

FILL FILL_0__8064_ (
);

NAND2X1 _10755_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1961_)
);

DFFSR _10335_ (
    .Q(\datapath_1.regfile_1.regOut[27] [9]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_1693_[9])
);

FILL FILL_3__11804_ (
);

FILL FILL_4__15283_ (
);

FILL FILL_2__9863_ (
);

FILL FILL_3__14696_ (
);

FILL FILL_0__11831_ (
);

FILL FILL_2__9023_ (
);

FILL FILL_3__14276_ (
);

FILL FILL_0__11411_ (
);

FILL FILL_4__9789_ (
);

FILL FILL_4__9369_ (
);

FILL FILL_2__13689_ (
);

FILL FILL_2__13269_ (
);

FILL SFILL69320x26050 (
);

FILL FILL_5__14603_ (
);

INVX1 _8903_ (
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_1031_)
);

FILL FILL_1__7860_ (
);

FILL FILL_1__7440_ (
);

FILL FILL_2__14630_ (
);

FILL FILL_2__14210_ (
);

FILL FILL_0__9269_ (
);

FILL FILL_3__7366_ (
);

FILL FILL_1__13623_ (
);

FILL FILL_4__16068_ (
);

FILL FILL_1_BUFX2_insert310 (
);

FILL FILL_1_BUFX2_insert311 (
);

FILL FILL_0__12616_ (
);

INVX1 _12901_ (
    .A(\datapath_1.a [26]),
    .Y(_3606_)
);

FILL FILL_1_BUFX2_insert312 (
);

FILL FILL_1_BUFX2_insert313 (
);

FILL FILL_1__16095_ (
);

FILL FILL_1_BUFX2_insert314 (
);

FILL FILL_1_BUFX2_insert315 (
);

FILL FILL_5__8653_ (
);

FILL FILL_1_BUFX2_insert316 (
);

FILL FILL_1_BUFX2_insert317 (
);

FILL FILL_3__10196_ (
);

FILL FILL_5__8233_ (
);

FILL FILL_1_BUFX2_insert318 (
);

FILL FILL_1_BUFX2_insert319 (
);

FILL FILL_6_BUFX2_insert874 (
);

NOR2X1 _15793_ (
    .A(_6252_),
    .B(_6254_),
    .Y(_6255_)
);

AOI21X1 _15373_ (
    .A(_5845_),
    .B(_5828_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [7])
);

FILL FILL_0__15088_ (
);

FILL FILL_5__15808_ (
);

FILL FILL_3__16002_ (
);

FILL FILL_6_BUFX2_insert879 (
);

FILL FILL_5__10943_ (
);

FILL FILL_1__8645_ (
);

FILL FILL_5__10523_ (
);

FILL FILL_1__8225_ (
);

FILL FILL_5__10103_ (
);

FILL FILL_2__15835_ (
);

FILL FILL_2__15415_ (
);

FILL FILL_2__10970_ (
);

FILL FILL_2__10550_ (
);

FILL FILL_6__6996_ (
);

FILL FILL_2__10130_ (
);

FILL FILL_1__14828_ (
);

INVX1 _7295_ (
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_203_)
);

FILL FILL_1__14408_ (
);

FILL SFILL59720x38050 (
);

FILL FILL_3__9932_ (
);

FILL FILL_3__9512_ (
);

FILL FILL_2__6988_ (
);

FILL FILL_0__6970_ (
);

FILL SFILL104360x58050 (
);

FILL FILL_5__9858_ (
);

FILL FILL_5__9018_ (
);

OAI22X1 _16158_ (
    .A(_6610_),
    .B(_5548__bF$buf4),
    .C(_5534__bF$buf3),
    .D(_5241_),
    .Y(_6611_)
);

NOR2X1 _11293_ (
    .A(_2410_),
    .B(_2411_),
    .Y(_2412_)
);

FILL FILL_5__11728_ (
);

FILL FILL_3__12762_ (
);

FILL FILL_5__11308_ (
);

FILL FILL_3__12342_ (
);

FILL SFILL108680x66050 (
);

FILL FILL_4__7855_ (
);

FILL FILL_4__7435_ (
);

FILL FILL_2__11755_ (
);

FILL FILL_2__11335_ (
);

FILL FILL_1__10748_ (
);

FILL FILL_5__15981_ (
);

FILL FILL_5__15561_ (
);

FILL FILL_0__7755_ (
);

FILL FILL_5__15141_ (
);

FILL SFILL43640x46050 (
);

FILL FILL112440x64050 (
);

FILL FILL_0__7335_ (
);

INVX1 _9861_ (
    .A(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_1507_)
);

DFFSR _9441_ (
    .Q(\datapath_1.regfile_1.regOut[20] [11]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1238_[11])
);

OAI21X1 _9021_ (
    .A(_1088_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1089_),
    .Y(_1043_[23])
);

FILL FILL_4__14974_ (
);

FILL FILL_4__14554_ (
);

FILL FILL_4__14134_ (
);

OAI21X1 _12498_ (
    .A(_3397_),
    .B(vdd),
    .C(_3398_),
    .Y(_3360_[19])
);

NAND3X1 _12078_ (
    .A(_3102_),
    .B(_3103_),
    .C(_3104_),
    .Y(\datapath_1.mux_pcsrc.dout [22])
);

FILL FILL_2__8714_ (
);

FILL FILL_3__13967_ (
);

FILL FILL_3__13547_ (
);

FILL FILL_1__14581_ (
);

FILL FILL_3__13127_ (
);

FILL FILL_1__14161_ (
);

FILL FILL_5_BUFX2_insert890 (
);

FILL FILL_5_BUFX2_insert891 (
);

FILL FILL_5_BUFX2_insert892 (
);

FILL FILL_0__13994_ (
);

FILL FILL_5_BUFX2_insert893 (
);

FILL FILL_0__13574_ (
);

FILL FILL_5_BUFX2_insert894 (
);

FILL FILL_0__13154_ (
);

FILL FILL_5_BUFX2_insert895 (
);

FILL FILL_5_BUFX2_insert896 (
);

FILL FILL_5_BUFX2_insert897 (
);

FILL FILL_5_BUFX2_insert898 (
);

FILL FILL_5_BUFX2_insert899 (
);

FILL FILL_2__13901_ (
);

FILL FILL_5__16346_ (
);

FILL FILL_6__9927_ (
);

FILL FILL_5__11481_ (
);

FILL FILL_5__11061_ (
);

FILL FILL_4__15759_ (
);

FILL FILL_4__15339_ (
);

FILL FILL_2__16373_ (
);

FILL FILL_4__10894_ (
);

FILL FILL_2__9919_ (
);

FILL FILL_4__10054_ (
);

FILL FILL_0__9901_ (
);

FILL FILL_1__15786_ (
);

FILL FILL_1__15366_ (
);

FILL FILL_5__7504_ (
);

FILL FILL_6__10801_ (
);

FILL FILL_0__14779_ (
);

NOR2X1 _14644_ (
    .A(_5131_),
    .B(_5128_),
    .Y(_5132_)
);

FILL FILL_0__14359_ (
);

NOR2X1 _14224_ (
    .A(_4719_),
    .B(_4716_),
    .Y(_4720_)
);

FILL SFILL89400x18050 (
);

FILL FILL_0__15720_ (
);

FILL FILL_0__15300_ (
);

FILL FILL_5__12266_ (
);

INVX1 _6986_ (
    .A(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_58_)
);

FILL FILL_4__8393_ (
);

FILL FILL_4__11679_ (
);

FILL FILL_4__11259_ (
);

FILL FILL_2__12293_ (
);

FILL FILL_5__8709_ (
);

FILL SFILL23720x80050 (
);

FILL FILL_1__11286_ (
);

NOR2X1 _15849_ (
    .A(_6309_),
    .B(_6306_),
    .Y(_6310_)
);

FILL FILL_4__12620_ (
);

OAI22X1 _15429_ (
    .A(_5526__bF$buf1),
    .B(_4426_),
    .C(_4407_),
    .D(_5527__bF$buf2),
    .Y(_5900_)
);

NAND3X1 _15009_ (
    .A(_5459__bF$buf1),
    .B(_5468_),
    .C(_5471__bF$buf3),
    .Y(_5489_)
);

FILL FILL_4__12200_ (
);

DFFSR _10984_ (
    .Q(\control_1.reg_state.dout [0]),
    .CLK(clk_bF$buf36),
    .R(rst_bF$buf100),
    .S(vdd),
    .D(_2098_[0])
);

FILL FILL_0__10699_ (
);

FILL FILL_0__10279_ (
);

INVX1 _10564_ (
    .A(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_1874_)
);

FILL FILL_6__9260_ (
);

INVX1 _10144_ (
    .A(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_1655_)
);

FILL FILL_3__11613_ (
);

FILL FILL_6__14058_ (
);

FILL FILL_4__15092_ (
);

FILL FILL_2__9672_ (
);

FILL FILL_2__9252_ (
);

FILL FILL_0__11640_ (
);

FILL FILL_0__11220_ (
);

FILL FILL_3__14085_ (
);

FILL FILL_4__9598_ (
);

FILL FILL_2__13498_ (
);

FILL FILL_5__14832_ (
);

FILL FILL_5__14412_ (
);

INVX1 _8712_ (
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_924_)
);

FILL FILL_4__13825_ (
);

FILL FILL_4__13405_ (
);

FILL FILL_0__9498_ (
);

FILL FILL_3__7595_ (
);

FILL FILL_0__9078_ (
);

OAI21X1 _11769_ (
    .A(_2863_),
    .B(_2139_),
    .C(_2861_),
    .Y(_2864_)
);

FILL FILL_3__7175_ (
);

OAI22X1 _11349_ (
    .A(_2115_),
    .B(_2347__bF$buf2),
    .C(_2350_),
    .D(_2346_),
    .Y(_2467_)
);

FILL FILL_1__13852_ (
);

FILL FILL_1__13432_ (
);

FILL FILL_4__16297_ (
);

FILL SFILL98920x44050 (
);

FILL FILL_1__13012_ (
);

FILL FILL_6__10398_ (
);

FILL SFILL84280x67050 (
);

FILL FILL_0__12845_ (
);

INVX1 _12710_ (
    .A(\aluControl_1.inst [5]),
    .Y(_3499_)
);

FILL FILL_0__12425_ (
);

FILL FILL_0__12005_ (
);

FILL FILL_5__8882_ (
);

FILL FILL_5__8462_ (
);

OAI22X1 _15182_ (
    .A(_4124_),
    .B(_5548__bF$buf0),
    .C(_5495__bF$buf1),
    .D(_5658_),
    .Y(_5659_)
);

FILL FILL_5__15617_ (
);

OAI21X1 _9917_ (
    .A(_1543_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1544_),
    .Y(_1498_[23])
);

FILL FILL_3__16231_ (
);

FILL FILL_5__10752_ (
);

FILL FILL_1__8874_ (
);

FILL FILL_1__8454_ (
);

FILL SFILL8680x41050 (
);

FILL FILL_2__15644_ (
);

FILL SFILL84680x36050 (
);

FILL FILL_2__15224_ (
);

FILL FILL_1__14637_ (
);

FILL FILL_1__14217_ (
);

FILL SFILL69400x59050 (
);

FILL SFILL84200x65050 (
);

FILL FILL_3__9741_ (
);

INVX1 _13915_ (
    .A(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_4418_)
);

FILL FILL_5__9667_ (
);

FILL FILL_5__9247_ (
);

INVX1 _16387_ (
    .A(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_6812_)
);

FILL FILL_5__11957_ (
);

FILL FILL_1__9659_ (
);

FILL FILL_3__12991_ (
);

FILL FILL_5__11537_ (
);

FILL FILL_3__12571_ (
);

FILL FILL_1__9239_ (
);

FILL FILL_5__11117_ (
);

FILL FILL_3__12151_ (
);

FILL FILL_2__16009_ (
);

FILL FILL_4__7244_ (
);

FILL FILL_2__11984_ (
);

FILL SFILL114440x48050 (
);

FILL FILL_2__11564_ (
);

FILL FILL_2__11144_ (
);

FILL FILL_1__10977_ (
);

FILL FILL_1__10557_ (
);

FILL FILL_1__10137_ (
);

FILL FILL_5__15790_ (
);

FILL SFILL84200x20050 (
);

FILL FILL_5__15370_ (
);

FILL FILL_0__7984_ (
);

FILL SFILL74280x65050 (
);

FILL FILL_0__7564_ (
);

FILL FILL_6__8951_ (
);

FILL FILL_6__8531_ (
);

OAI21X1 _9670_ (
    .A(_1419_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1420_),
    .Y(_1368_[26])
);

OAI21X1 _9250_ (
    .A(_1200_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .C(_1201_),
    .Y(_1173_[14])
);

FILL SFILL99160x50 (
);

FILL FILL_4__14783_ (
);

FILL FILL_4__14363_ (
);

FILL SFILL13640x40050 (
);

FILL FILL_0__10911_ (
);

FILL FILL_3__13776_ (
);

FILL FILL_2__8523_ (
);

FILL FILL_3__13356_ (
);

FILL FILL_2__8103_ (
);

FILL SFILL27880x12050 (
);

FILL FILL_1__14390_ (
);

FILL FILL_4__8869_ (
);

FILL FILL_4__8449_ (
);

FILL FILL_2__12769_ (
);

FILL FILL_2__12349_ (
);

FILL FILL_0__13383_ (
);

FILL FILL_1__6940_ (
);

FILL FILL_4__9810_ (
);

FILL FILL_2__13710_ (
);

FILL SFILL74200x63050 (
);

FILL FILL_3__6866_ (
);

FILL FILL_5__16155_ (
);

FILL FILL_0__8769_ (
);

FILL FILL_6__9736_ (
);

FILL FILL_0__8349_ (
);

FILL FILL_5__11290_ (
);

FILL FILL_4__15988_ (
);

FILL SFILL74280x20050 (
);

FILL FILL_1__12703_ (
);

FILL FILL_4__15568_ (
);

FILL FILL_4__15148_ (
);

FILL FILL_2__16182_ (
);

FILL FILL_4__10283_ (
);

FILL SFILL19240x68050 (
);

FILL FILL_2__9728_ (
);

FILL FILL_1__15595_ (
);

FILL FILL_1__15175_ (
);

FILL FILL_5__7733_ (
);

FILL FILL_5__7313_ (
);

INVX1 _14873_ (
    .A(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_5356_)
);

FILL FILL_0__14588_ (
);

OAI22X1 _14453_ (
    .A(_4942_),
    .B(_3982__bF$buf3),
    .C(_3978_),
    .D(_4943_),
    .Y(_4944_)
);

FILL FILL_0__14168_ (
);

INVX1 _14033_ (
    .A(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_4533_)
);

FILL FILL_3__15922_ (
);

FILL FILL_3__15502_ (
);

FILL FILL_1__7725_ (
);

FILL FILL_1__7305_ (
);

FILL FILL_2__14915_ (
);

FILL FILL_5__12495_ (
);

FILL FILL112120x83050 (
);

FILL FILL_5__12075_ (
);

FILL FILL_1__13908_ (
);

FILL SFILL64280x63050 (
);

FILL FILL_4__11488_ (
);

FILL FILL_4__11068_ (
);

FILL FILL_5__8518_ (
);

FILL FILL_1__11095_ (
);

NOR3X1 _15658_ (
    .A(_6119_),
    .B(_6121_),
    .C(_6122_),
    .Y(_6123_)
);

INVX1 _15238_ (
    .A(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_5714_)
);

INVX1 _10793_ (
    .A(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_1986_)
);

INVX1 _10373_ (
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_1767_)
);

FILL FILL_5__10808_ (
);

FILL FILL_3__11842_ (
);

FILL FILL_3__11422_ (
);

FILL FILL_3__11002_ (
);

FILL FILL_4__6935_ (
);

FILL FILL_0__16314_ (
);

FILL FILL_2__10835_ (
);

FILL FILL_2__9481_ (
);

FILL FILL_2__10415_ (
);

FILL SFILL33800x70050 (
);

FILL FILL_5__14641_ (
);

FILL FILL112440x59050 (
);

FILL FILL_5__14221_ (
);

DFFSR _8941_ (
    .Q(\datapath_1.regfile_1.regOut[16] [23]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_978_[23])
);

OAI21X1 _8521_ (
    .A(_836_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_837_),
    .Y(_783_[27])
);

OAI21X1 _8101_ (
    .A(_617_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .C(_618_),
    .Y(_588_[15])
);

FILL FILL_4__13634_ (
);

FILL FILL_4__13214_ (
);

NAND3X1 _11998_ (
    .A(_3042_),
    .B(_3043_),
    .C(_3044_),
    .Y(\datapath_1.mux_pcsrc.dout [2])
);

OAI21X1 _11578_ (
    .A(_2684_),
    .B(_2685_),
    .C(_2683_),
    .Y(_2686_)
);

OAI21X1 _11158_ (
    .A(_2229_),
    .B(_2230_),
    .C(_2276_),
    .Y(_2277_)
);

FILL FILL_3__12627_ (
);

FILL FILL_1__13661_ (
);

FILL FILL_3__12207_ (
);

FILL FILL_1__13241_ (
);

FILL FILL_0__12654_ (
);

FILL FILL_0__12234_ (
);

FILL FILL_3__15099_ (
);

FILL FILL_5__8271_ (
);

FILL FILL_5__15846_ (
);

FILL FILL_5__15426_ (
);

FILL FILL_5__15006_ (
);

FILL FILL_3__16040_ (
);

OAI21X1 _9726_ (
    .A(_1436_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .C(_1437_),
    .Y(_1433_[2])
);

FILL FILL_5__10981_ (
);

DFFSR _9306_ (
    .Q(\datapath_1.regfile_1.regOut[19] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_1173_[4])
);

FILL FILL_5__10561_ (
);

FILL FILL_1__8263_ (
);

FILL FILL_5__10141_ (
);

FILL FILL112440x14050 (
);

FILL FILL_4__14839_ (
);

FILL FILL_4__14419_ (
);

FILL FILL_2__15873_ (
);

FILL FILL_2__15453_ (
);

FILL FILL_2__15033_ (
);

FILL FILL_3__8189_ (
);

FILL FILL_1__14866_ (
);

FILL FILL_1__14446_ (
);

FILL FILL_1__14026_ (
);

FILL FILL_3__9550_ (
);

FILL FILL_0__13859_ (
);

FILL FILL_0__13439_ (
);

FILL FILL_3__9130_ (
);

INVX1 _13724_ (
    .A(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_4231_)
);

NOR2X1 _13304_ (
    .A(_3794_),
    .B(_3838_),
    .Y(_3839_)
);

FILL FILL_0__13019_ (
);

FILL FILL_5__9896_ (
);

FILL FILL_5__9476_ (
);

OAI22X1 _16196_ (
    .A(_5495__bF$buf1),
    .B(_5289_),
    .C(_5288_),
    .D(_5534__bF$buf2),
    .Y(_6648_)
);

FILL FILL_0__14800_ (
);

FILL FILL_1__9888_ (
);

FILL FILL_5__11766_ (
);

FILL FILL_5__11346_ (
);

FILL FILL_1__9468_ (
);

FILL FILL_3__12380_ (
);

FILL FILL_2__16238_ (
);

FILL FILL_4__7893_ (
);

FILL FILL_4__7473_ (
);

FILL FILL_4__7053_ (
);

FILL FILL_4__10759_ (
);

FILL FILL_2__11793_ (
);

FILL FILL_2__11373_ (
);

FILL SFILL23720x75050 (
);

FILL FILL_1__10786_ (
);

FILL FILL_1__10366_ (
);

AOI21X1 _14929_ (
    .A(_5410_),
    .B(_5389_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [30])
);

NOR2X1 _14509_ (
    .A(_4998_),
    .B(_3944__bF$buf3),
    .Y(_4999_)
);

FILL FILL_4__11700_ (
);

FILL FILL_0__7373_ (
);

FILL FILL_6__8340_ (
);

FILL FILL_4__14592_ (
);

FILL FILL_4__14172_ (
);

FILL SFILL58440x74050 (
);

FILL SFILL94280x19050 (
);

FILL FILL_2__8752_ (
);

FILL FILL_2__8332_ (
);

FILL FILL_3__13585_ (
);

FILL FILL_0__10300_ (
);

FILL FILL_3__13165_ (
);

FILL FILL_4__8258_ (
);

FILL FILL_2__12998_ (
);

FILL FILL_2__12578_ (
);

FILL FILL_2__12158_ (
);

FILL FILL_5_BUFX2_insert0 (
);

FILL FILL_5_BUFX2_insert1 (
);

FILL FILL_5_BUFX2_insert2 (
);

FILL FILL_5__13912_ (
);

FILL FILL_5_BUFX2_insert3 (
);

FILL FILL_5_BUFX2_insert4 (
);

FILL FILL_5_BUFX2_insert5 (
);

FILL FILL_5_BUFX2_insert6 (
);

FILL FILL_5_BUFX2_insert7 (
);

FILL FILL_5_BUFX2_insert8 (
);

FILL FILL_5_BUFX2_insert9 (
);

FILL FILL_4__12905_ (
);

FILL SFILL23720x30050 (
);

FILL FILL_0__8998_ (
);

FILL FILL_5__16384_ (
);

FILL FILL_0__8578_ (
);

DFFSR _10849_ (
    .Q(\datapath_1.regfile_1.regOut[31] [11]),
    .CLK(clk_bF$buf79),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_1953_[11])
);

OAI21X1 _10429_ (
    .A(_1803_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .C(_1804_),
    .Y(_1758_[23])
);

OAI21X1 _10009_ (
    .A(_1584_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1585_),
    .Y(_1563_[11])
);

FILL FILL_4__15797_ (
);

FILL FILL_4__15377_ (
);

FILL FILL_1__12512_ (
);

FILL FILL_0__11925_ (
);

FILL FILL_2__9537_ (
);

FILL FILL_0__11505_ (
);

FILL FILL_2__9117_ (
);

FILL FILL_5__7962_ (
);

FILL FILL_5__7542_ (
);

FILL FILL_5__7122_ (
);

FILL FILL_0__14397_ (
);

INVX1 _14682_ (
    .A(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_5169_)
);

AOI22X1 _14262_ (
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .B(_4102_),
    .C(_4090_),
    .D(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_4758_)
);

FILL SFILL8600x79050 (
);

FILL FILL_3__15731_ (
);

FILL FILL_3__15311_ (
);

FILL FILL_1__7954_ (
);

FILL FILL_1__7114_ (
);

FILL SFILL8680x36050 (
);

FILL SFILL13720x73050 (
);

FILL FILL_2__14724_ (
);

FILL FILL_2__14304_ (
);

FILL SFILL27960x45050 (
);

FILL FILL_1__13717_ (
);

FILL FILL_4__11297_ (
);

FILL FILL_3__8401_ (
);

FILL FILL_1__16189_ (
);

FILL FILL_5__8747_ (
);

FILL FILL_5__8327_ (
);

OAI22X1 _15887_ (
    .A(_5480__bF$buf2),
    .B(_6345_),
    .C(_5523_),
    .D(_6346_),
    .Y(_6347_)
);

AOI22X1 _15467_ (
    .A(\datapath_1.regfile_1.regOut[1] [10]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_5937_)
);

NAND3X1 _15047_ (
    .A(_5459__bF$buf2),
    .B(_5465_),
    .C(_5476_),
    .Y(_5527_)
);

OAI21X1 _10182_ (
    .A(_1679_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1680_),
    .Y(_1628_[26])
);

FILL FILL_1__8739_ (
);

FILL FILL_5__10617_ (
);

FILL FILL_1__8319_ (
);

FILL FILL_3__11651_ (
);

FILL FILL_3__11231_ (
);

FILL FILL_2__15929_ (
);

FILL FILL_2__15509_ (
);

FILL FILL_0__16123_ (
);

FILL FILL_2__10644_ (
);

FILL FILL_5__13089_ (
);

FILL FILL_2__9290_ (
);

DFFSR _7389_ (
    .Q(\datapath_1.regfile_1.regOut[4] [7]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_198_[7])
);

FILL FILL_3__9606_ (
);

FILL SFILL84200x15050 (
);

FILL FILL_5__14870_ (
);

FILL FILL_5__14450_ (
);

FILL FILL_5__14030_ (
);

FILL FILL_3_BUFX2_insert225 (
);

FILL FILL_6__7611_ (
);

OAI21X1 _8750_ (
    .A(_948_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .C(_949_),
    .Y(_913_[18])
);

FILL FILL_3_BUFX2_insert226 (
);

OAI21X1 _8330_ (
    .A(_729_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_730_),
    .Y(_718_[6])
);

FILL FILL_3_BUFX2_insert227 (
);

FILL FILL_3_BUFX2_insert228 (
);

FILL FILL_3_BUFX2_insert229 (
);

FILL FILL_4__13863_ (
);

FILL FILL_4__13443_ (
);

FILL FILL_4__13023_ (
);

FILL SFILL13640x35050 (
);

OAI21X1 _11387_ (
    .A(_2385_),
    .B(_2386_),
    .C(_2503_),
    .Y(_2504_)
);

FILL SFILL88520x23050 (
);

FILL FILL_3__12856_ (
);

FILL FILL_2__7603_ (
);

FILL FILL_3__12436_ (
);

FILL FILL_1__13890_ (
);

FILL SFILL109480x15050 (
);

FILL FILL_3__12016_ (
);

FILL FILL_1__13470_ (
);

FILL FILL_4__7949_ (
);

FILL FILL_4__7109_ (
);

FILL FILL_2__11849_ (
);

FILL FILL_0__12883_ (
);

FILL FILL_2__11429_ (
);

FILL FILL_0__12463_ (
);

FILL FILL_2__11009_ (
);

FILL FILL_0__12043_ (
);

FILL FILL_6__16242_ (
);

FILL FILL_5__8080_ (
);

FILL FILL_5__15655_ (
);

FILL FILL_5__15235_ (
);

FILL FILL_0__7849_ (
);

FILL FILL_0__7429_ (
);

DFFSR _9955_ (
    .Q(\datapath_1.regfile_1.regOut[24] [13]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_1498_[13])
);

NAND2X1 _9535_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1351_)
);

FILL FILL_5__10790_ (
);

NAND2X1 _9115_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1132_)
);

FILL FILL_5__10370_ (
);

FILL FILL_1__8492_ (
);

FILL SFILL74280x15050 (
);

FILL FILL_1__8072_ (
);

FILL FILL_4__14648_ (
);

FILL FILL_2__15682_ (
);

FILL FILL_4__14228_ (
);

FILL FILL_2__15262_ (
);

FILL FILL112200x71050 (
);

FILL FILL_1__14675_ (
);

FILL SFILL99480x64050 (
);

FILL FILL_1__14255_ (
);

FILL FILL_0_BUFX2_insert350 (
);

FILL FILL_0_BUFX2_insert351 (
);

FILL FILL_0_BUFX2_insert352 (
);

FILL FILL_0_BUFX2_insert353 (
);

FILL FILL_0_BUFX2_insert354 (
);

FILL FILL_0__13668_ (
);

NOR2X1 _13953_ (
    .A(_4444_),
    .B(_4454_),
    .Y(_4455_)
);

FILL FILL_0__13248_ (
);

FILL FILL_0_BUFX2_insert355 (
);

AOI21X1 _13533_ (
    .A(_4043_),
    .B(_4015_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [1])
);

FILL FILL_0_BUFX2_insert356 (
);

NAND2X1 _13113_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_pcsrc.dout [11]),
    .Y(_3707_)
);

FILL FILL_0_BUFX2_insert357 (
);

FILL FILL_0_BUFX2_insert358 (
);

FILL FILL_5__9285_ (
);

FILL FILL_0_BUFX2_insert359 (
);

FILL FILL_6__12162_ (
);

FILL FILL_5__11995_ (
);

FILL FILL112120x78050 (
);

FILL FILL_5__11575_ (
);

FILL SFILL74200x13050 (
);

FILL FILL_1__9277_ (
);

FILL FILL_5__11155_ (
);

FILL FILL_2__16047_ (
);

FILL FILL_4__10988_ (
);

FILL FILL_4__10568_ (
);

FILL FILL_4__10148_ (
);

FILL FILL_2__11182_ (
);

FILL FILL_1__10175_ (
);

AOI22X1 _14738_ (
    .A(_3891__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [26]),
    .C(\datapath_1.regfile_1.regOut[8] [26]),
    .D(_4090_),
    .Y(_5224_)
);

INVX1 _14318_ (
    .A(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_4812_)
);

FILL FILL_0__7182_ (
);

FILL FILL_2_BUFX2_insert30 (
);

FILL SFILL28840x82050 (
);

FILL FILL_2_BUFX2_insert31 (
);

FILL FILL_1__16401_ (
);

FILL FILL_2_BUFX2_insert32 (
);

FILL FILL_3__10922_ (
);

FILL FILL_6__13787_ (
);

FILL FILL_2_BUFX2_insert33 (
);

FILL FILL_2_BUFX2_insert34 (
);

FILL FILL_6__13367_ (
);

FILL FILL_3__10502_ (
);

FILL FILL_2_BUFX2_insert35 (
);

FILL FILL_2_BUFX2_insert36 (
);

FILL FILL_0__15814_ (
);

FILL FILL_2_BUFX2_insert37 (
);

FILL FILL_2_BUFX2_insert38 (
);

FILL FILL_2_BUFX2_insert39 (
);

FILL SFILL68920x78050 (
);

FILL FILL_2__8981_ (
);

FILL SFILL33800x65050 (
);

FILL SFILL64200x56050 (
);

FILL FILL_2__8141_ (
);

FILL FILL_3__13394_ (
);

FILL FILL112120x33050 (
);

FILL FILL_4__8487_ (
);

FILL FILL_4__8067_ (
);

FILL FILL_2__12387_ (
);

FILL SFILL68760x6050 (
);

FILL FILL_5__13721_ (
);

FILL FILL_5__13301_ (
);

OAI21X1 _7601_ (
    .A(_365_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .C(_366_),
    .Y(_328_[19])
);

FILL FILL_0_CLKBUF1_insert1074 (
);

FILL FILL_0_CLKBUF1_insert1075 (
);

FILL FILL_4__12714_ (
);

FILL FILL_0_CLKBUF1_insert1076 (
);

FILL FILL_0_CLKBUF1_insert1077 (
);

FILL FILL_0_CLKBUF1_insert1078 (
);

FILL FILL_5__16193_ (
);

FILL FILL_0_CLKBUF1_insert1079 (
);

FILL FILL_0__8387_ (
);

OAI21X1 _10658_ (
    .A(_1915_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .C(_1916_),
    .Y(_1888_[14])
);

OAI21X1 _10238_ (
    .A(_1696_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1697_),
    .Y(_1693_[2])
);

FILL FILL_3__11707_ (
);

FILL FILL_1__12741_ (
);

FILL FILL_4__15186_ (
);

FILL FILL_1__12321_ (
);

FILL FILL_2__9766_ (
);

FILL FILL_3__14599_ (
);

FILL FILL_2__9346_ (
);

FILL FILL_0__11734_ (
);

FILL FILL_3__14179_ (
);

FILL FILL_0__11314_ (
);

FILL FILL_5__7351_ (
);

FILL SFILL64200x11050 (
);

INVX1 _14491_ (
    .A(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_4982_)
);

OAI22X1 _14071_ (
    .A(_4569_),
    .B(_3893__bF$buf0),
    .C(_3971__bF$buf3),
    .D(_4570_),
    .Y(_4571_)
);

FILL FILL_5__14926_ (
);

FILL FILL_3__15960_ (
);

FILL FILL_5__14506_ (
);

FILL FILL_3__15540_ (
);

DFFSR _8806_ (
    .Q(\datapath_1.regfile_1.regOut[15] [16]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_913_[16])
);

FILL FILL_3__15120_ (
);

FILL FILL_1__7763_ (
);

FILL FILL_1__7343_ (
);

FILL FILL_4__13919_ (
);

FILL FILL_2__14953_ (
);

FILL FILL_2__14533_ (
);

FILL FILL_3__7689_ (
);

FILL FILL_2__14113_ (
);

FILL FILL_1__13946_ (
);

FILL FILL_1__13526_ (
);

FILL FILL_1__13106_ (
);

FILL FILL_3__8630_ (
);

DFFSR _12804_ (
    .Q(\datapath_1.PCJump [15]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3490_[13])
);

FILL FILL_0__12519_ (
);

FILL FILL_3__8210_ (
);

FILL FILL_5__8976_ (
);

FILL SFILL58920x76050 (
);

FILL FILL_5__8136_ (
);

AOI22X1 _15696_ (
    .A(_5562_),
    .B(\datapath_1.regfile_1.regOut[25] [16]),
    .C(\datapath_1.regfile_1.regOut[22] [16]),
    .D(_5650_),
    .Y(_6160_)
);

NOR3X1 _15276_ (
    .A(_5515__bF$buf2),
    .B(_5750_),
    .C(_5521__bF$buf1),
    .Y(_5751_)
);

FILL FILL_3__16325_ (
);

FILL FILL_1__8968_ (
);

FILL FILL_3__11880_ (
);

FILL FILL_5__10426_ (
);

FILL FILL_1__8128_ (
);

FILL FILL_3__11460_ (
);

FILL FILL_5__10006_ (
);

FILL FILL_3__11040_ (
);

FILL FILL_2__15738_ (
);

FILL FILL_4__6973_ (
);

FILL FILL_2__15318_ (
);

FILL FILL_0__16352_ (
);

FILL FILL_2__10873_ (
);

FILL FILL_2__10453_ (
);

FILL FILL_2__10033_ (
);

FILL FILL_6__6899_ (
);

NAND2X1 _7198_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_159_)
);

FILL FILL_3__9415_ (
);

FILL FILL_0__6873_ (
);

FILL FILL_4__13672_ (
);

FILL FILL_6__12218_ (
);

FILL FILL_4__13252_ (
);

OAI21X1 _11196_ (
    .A(_2311_),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .C(_2314_),
    .Y(_2315_)
);

FILL FILL_2__7832_ (
);

FILL FILL_3__12245_ (
);

FILL FILL_4__7758_ (
);

FILL FILL_4__7338_ (
);

FILL FILL_2__11658_ (
);

FILL FILL_2__11238_ (
);

FILL SFILL39480x3050 (
);

FILL FILL_0__12272_ (
);

FILL SFILL109240x72050 (
);

FILL SFILL74120x4050 (
);

FILL SFILL23720x25050 (
);

FILL FILL_5__15884_ (
);

FILL FILL_5__15464_ (
);

FILL FILL_5__15044_ (
);

NAND2X1 _9764_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1463_)
);

FILL FILL_0__7238_ (
);

NAND2X1 _9344_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_1244_)
);

FILL FILL_4__14877_ (
);

FILL FILL_4__14457_ (
);

FILL FILL_4__14037_ (
);

FILL FILL_2__15491_ (
);

FILL FILL_2__15071_ (
);

FILL FILL_2__8617_ (
);

FILL FILL_1__14484_ (
);

FILL FILL_1__14064_ (
);

FILL FILL_0__13897_ (
);

INVX1 _13762_ (
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_4268_)
);

FILL FILL_0__13477_ (
);

NAND3X1 _13342_ (
    .A(_3783_),
    .B(_3826_),
    .C(_3861_),
    .Y(_3863_)
);

FILL FILL_3__14811_ (
);

FILL FILL_5__9094_ (
);

FILL FILL_4__9904_ (
);

FILL FILL_2__13804_ (
);

FILL FILL_5__16249_ (
);

FILL SFILL109560x48050 (
);

FILL FILL_5__11384_ (
);

FILL FILL_1__9086_ (
);

FILL FILL_2__16276_ (
);

FILL FILL_4__10797_ (
);

FILL FILL_4__7091_ (
);

FILL FILL_4__10377_ (
);

FILL FILL_0__9804_ (
);

FILL FILL_1__15689_ (
);

FILL FILL_1__15269_ (
);

FILL FILL_5__7827_ (
);

NOR2X1 _14967_ (
    .A(_5447_),
    .B(_3935__bF$buf2),
    .Y(_5448_)
);

NAND3X1 _14547_ (
    .A(_5028_),
    .B(_5029_),
    .C(_5036_),
    .Y(_5037_)
);

INVX1 _14127_ (
    .A(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_4625_)
);

FILL FILL_1__16210_ (
);

FILL FILL_1__7819_ (
);

FILL SFILL8600x29050 (
);

FILL FILL_3__10311_ (
);

FILL FILL_0__15623_ (
);

FILL FILL_0__15203_ (
);

FILL SFILL13720x23050 (
);

FILL FILL_5__12589_ (
);

FILL FILL_5__12169_ (
);

FILL FILL_2__8370_ (
);

BUFX2 _6889_ (
    .A(_2_[19]),
    .Y(memoryWriteData[19])
);

FILL FILL_2__12196_ (
);

FILL SFILL38920x72050 (
);

FILL FILL_5__13950_ (
);

FILL FILL_5__13530_ (
);

FILL FILL_5__13110_ (
);

OAI21X1 _7830_ (
    .A(_477_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .C(_478_),
    .Y(_458_[10])
);

DFFSR _7410_ (
    .Q(\datapath_1.regfile_1.regOut[4] [28]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_198_[28])
);

FILL FILL_1__11189_ (
);

FILL FILL_4__12523_ (
);

FILL FILL_4__12103_ (
);

FILL FILL_0__8196_ (
);

OAI21X1 _10887_ (
    .A(_2022_),
    .B(_2033_),
    .C(_2031_),
    .Y(_2034_)
);

DFFSR _10467_ (
    .Q(\datapath_1.regfile_1.regOut[28] [13]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_1758_[13])
);

NAND2X1 _10047_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1611_)
);

FILL FILL_3__11936_ (
);

FILL FILL_3__11516_ (
);

FILL FILL_1__12970_ (
);

FILL FILL_1__12130_ (
);

FILL FILL_0__16408_ (
);

FILL SFILL38840x79050 (
);

FILL FILL_2__9995_ (
);

FILL FILL_2__10929_ (
);

FILL FILL_2__10509_ (
);

FILL FILL_0__11963_ (
);

FILL SFILL34120x57050 (
);

FILL FILL_2__9155_ (
);

FILL FILL_0__11543_ (
);

FILL FILL_0__11123_ (
);

FILL FILL_5__7580_ (
);

FILL FILL_5__7160_ (
);

FILL SFILL3560x71050 (
);

FILL FILL_5__14735_ (
);

FILL FILL_5__14315_ (
);

FILL FILL_0__6929_ (
);

NAND2X1 _8615_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_880_)
);

FILL FILL_1__7992_ (
);

FILL FILL_1__7572_ (
);

FILL FILL_4__13728_ (
);

FILL FILL_4__13308_ (
);

FILL FILL_2__14762_ (
);

FILL FILL_2__14342_ (
);

FILL FILL_3__7498_ (
);

FILL FILL_3__7078_ (
);

FILL FILL112200x66050 (
);

FILL SFILL99480x59050 (
);

FILL FILL_1__13755_ (
);

FILL FILL_1__13335_ (
);

FILL SFILL44040x8050 (
);

FILL FILL_0__12748_ (
);

NAND2X1 _12613_ (
    .A(vdd),
    .B(memoryOutData[15]),
    .Y(_3455_)
);

FILL FILL_0__12328_ (
);

FILL SFILL38840x34050 (
);

FILL FILL_5__8785_ (
);

FILL FILL_5__8365_ (
);

NAND3X1 _15085_ (
    .A(_5561_),
    .B(_5563_),
    .C(_5559_),
    .Y(_5564_)
);

FILL FILL_3__16134_ (
);

FILL SFILL28920x70050 (
);

FILL FILL_1__8777_ (
);

FILL FILL_5__10655_ (
);

FILL FILL_1__8357_ (
);

FILL FILL_5__10235_ (
);

FILL FILL_2__15967_ (
);

FILL FILL_2__15547_ (
);

FILL FILL_2__15127_ (
);

FILL FILL_0__16161_ (
);

FILL FILL_2__10682_ (
);

FILL FILL_2__10262_ (
);

FILL FILL112200x21050 (
);

FILL SFILL99480x14050 (
);

FILL FILL_3_BUFX2_insert600 (
);

FILL FILL_3__9644_ (
);

AOI22X1 _13818_ (
    .A(_3891__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [7]),
    .C(\datapath_1.regfile_1.regOut[8] [7]),
    .D(_4090_),
    .Y(_4323_)
);

FILL FILL_3__9224_ (
);

FILL FILL_3_BUFX2_insert601 (
);

FILL FILL_3_BUFX2_insert602 (
);

FILL FILL_3_BUFX2_insert603 (
);

FILL FILL_3_BUFX2_insert604 (
);

FILL SFILL28840x77050 (
);

FILL FILL_3_BUFX2_insert605 (
);

FILL FILL_1__15901_ (
);

FILL FILL_3_BUFX2_insert606 (
);

FILL FILL_3_BUFX2_insert607 (
);

FILL FILL_3_BUFX2_insert608 (
);

FILL FILL_6__12867_ (
);

FILL FILL_3_BUFX2_insert609 (
);

FILL FILL_4__13481_ (
);

FILL FILL_3__12894_ (
);

FILL FILL_2__7221_ (
);

FILL FILL_3__12474_ (
);

FILL FILL_3__12054_ (
);

FILL FILL112120x28050 (
);

FILL FILL_4__7987_ (
);

FILL FILL_4__7567_ (
);

FILL FILL_2__11887_ (
);

FILL FILL_2__11467_ (
);

FILL FILL_2__11047_ (
);

FILL FILL_0__12081_ (
);

FILL FILL_5__15693_ (
);

FILL FILL_0__7887_ (
);

FILL FILL_5__15273_ (
);

NAND2X1 _9993_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1575_)
);

FILL FILL_0__7467_ (
);

DFFSR _9573_ (
    .Q(\datapath_1.regfile_1.regOut[21] [15]),
    .CLK(clk_bF$buf32),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_1303_[15])
);

FILL FILL_0__7047_ (
);

FILL FILL_6__8014_ (
);

INVX1 _9153_ (
    .A(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_1157_)
);

FILL FILL_1__11821_ (
);

FILL FILL_4__14686_ (
);

FILL SFILL28840x32050 (
);

FILL FILL_4__14266_ (
);

FILL FILL_1__11401_ (
);

FILL FILL_2__8846_ (
);

FILL FILL_0__10814_ (
);

FILL FILL_3__13679_ (
);

FILL FILL_3__13259_ (
);

FILL FILL_2__8006_ (
);

FILL FILL_1__14293_ (
);

FILL SFILL33800x15050 (
);

FILL FILL_0_BUFX2_insert730 (
);

FILL FILL_5__6851_ (
);

FILL FILL_0_BUFX2_insert731 (
);

FILL FILL_0_BUFX2_insert732 (
);

FILL FILL_0_BUFX2_insert733 (
);

INVX1 _13991_ (
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_4492_)
);

FILL FILL_0_BUFX2_insert734 (
);

FILL FILL_0__13286_ (
);

FILL FILL_0_BUFX2_insert735 (
);

NAND3X1 _13571_ (
    .A(_4078_),
    .B(_4080_),
    .C(_4077_),
    .Y(_4081_)
);

INVX1 _13151_ (
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3732_)
);

FILL FILL_0_BUFX2_insert736 (
);

FILL FILL_0_BUFX2_insert737 (
);

FILL FILL_3__14620_ (
);

FILL FILL_0_BUFX2_insert738 (
);

FILL FILL_3__14200_ (
);

FILL FILL_0_BUFX2_insert739 (
);

FILL FILL_1__6843_ (
);

FILL FILL_2__13613_ (
);

FILL FILL_5__16058_ (
);

FILL FILL_6__9219_ (
);

FILL FILL_5__11193_ (
);

FILL FILL_1__12606_ (
);

FILL SFILL18840x75050 (
);

FILL FILL_2__16085_ (
);

FILL FILL_4__10186_ (
);

FILL FILL_0__9613_ (
);

FILL FILL_3__7710_ (
);

FILL FILL_1__15498_ (
);

FILL FILL_1__15078_ (
);

FILL FILL_5__7636_ (
);

FILL FILL_5__7216_ (
);

FILL FILL_4__16412_ (
);

INVX1 _14776_ (
    .A(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_5261_)
);

NOR2X1 _14356_ (
    .A(_4849_),
    .B(_4839_),
    .Y(_4850_)
);

FILL FILL_3__15825_ (
);

FILL FILL_3__15405_ (
);

FILL FILL_3__10960_ (
);

FILL FILL_1__7628_ (
);

FILL FILL_1__7208_ (
);

FILL FILL_3__10540_ (
);

FILL FILL_3__10120_ (
);

FILL FILL_2__14818_ (
);

FILL FILL_0__15852_ (
);

FILL FILL_0__15432_ (
);

FILL FILL_0__15012_ (
);

FILL FILL_5__12398_ (
);

FILL FILL_3__8915_ (
);

FILL SFILL18840x30050 (
);

FILL FILL_4__12752_ (
);

FILL FILL_4__12332_ (
);

NAND2X1 _10696_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1942_)
);

FILL SFILL103560x46050 (
);

NAND2X1 _10276_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1723_)
);

FILL FILL_2__6912_ (
);

FILL FILL_3__11745_ (
);

FILL FILL_3__11325_ (
);

FILL FILL_4__6838_ (
);

FILL FILL_0__16217_ (
);

FILL FILL_2__10318_ (
);

FILL FILL_2__9384_ (
);

FILL FILL_0__11772_ (
);

FILL FILL_0__11352_ (
);

FILL FILL_6__15971_ (
);

FILL FILL_5__14964_ (
);

FILL FILL_5__14544_ (
);

FILL FILL_5__14124_ (
);

NAND2X1 _8844_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_992_)
);

FILL FILL_6__7705_ (
);

DFFSR _8424_ (
    .Q(\datapath_1.regfile_1.regOut[12] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_718_[18])
);

INVX1 _8004_ (
    .A(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_574_)
);

FILL FILL_1__7381_ (
);

FILL FILL_4__13957_ (
);

FILL SFILL48920x69050 (
);

FILL FILL_2__14991_ (
);

FILL FILL_4__13537_ (
);

FILL FILL_2__14571_ (
);

FILL FILL_4__13117_ (
);

FILL FILL_2__14151_ (
);

FILL FILL_1__13984_ (
);

FILL FILL_1__13564_ (
);

FILL FILL_1__13144_ (
);

FILL FILL_0__12977_ (
);

NAND2X1 _12842_ (
    .A(vdd),
    .B(\datapath_1.rd1 [6]),
    .Y(_3567_)
);

NAND2X1 _12422_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [26]),
    .Y(_3347_)
);

FILL FILL_0__12137_ (
);

NAND3X1 _12002_ (
    .A(_3045_),
    .B(_3046_),
    .C(_3047_),
    .Y(\datapath_1.mux_pcsrc.dout [3])
);

FILL FILL_5__8594_ (
);

FILL FILL_6__11891_ (
);

FILL FILL_6__11471_ (
);

FILL FILL_5__15749_ (
);

FILL FILL_5__15329_ (
);

FILL FILL_3__16363_ (
);

FILL SFILL69000x82050 (
);

INVX1 _9629_ (
    .A(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_1393_)
);

FILL FILL_5__10884_ (
);

INVX1 _9209_ (
    .A(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_1174_)
);

FILL FILL_1__8586_ (
);

FILL FILL_5__10044_ (
);

FILL FILL_2__15776_ (
);

FILL FILL_2__15356_ (
);

FILL FILL_0__16390_ (
);

FILL SFILL48920x24050 (
);

FILL FILL_2__10491_ (
);

FILL FILL_1__14769_ (
);

FILL FILL_1__14349_ (
);

FILL FILL_5__6907_ (
);

FILL FILL_3__9873_ (
);

AOI22X1 _13627_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [3]),
    .C(\datapath_1.regfile_1.regOut[18] [3]),
    .D(_4135_),
    .Y(_4136_)
);

FILL FILL_3__9033_ (
);

INVX4 _13207_ (
    .A(\datapath_1.a3 [4]),
    .Y(_3750_)
);

FILL FILL_5__9799_ (
);

FILL FILL_5__9379_ (
);

FILL FILL_1__15710_ (
);

FILL FILL_4__13290_ (
);

OAI22X1 _16099_ (
    .A(_5182_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf3),
    .D(_5210_),
    .Y(_6553_)
);

FILL FILL_0__14703_ (
);

FILL SFILL13720x18050 (
);

FILL FILL_2__7870_ (
);

FILL FILL_5__11669_ (
);

FILL FILL_2__7450_ (
);

FILL FILL_5__11249_ (
);

FILL FILL_2__7030_ (
);

FILL FILL_3__12283_ (
);

FILL SFILL59080x82050 (
);

FILL FILL_4__7376_ (
);

FILL FILL_2__11696_ (
);

FILL FILL_2__11276_ (
);

FILL FILL_5__12610_ (
);

OAI21X1 _6910_ (
    .A(_6_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .C(_7_),
    .Y(_3_[2])
);

FILL FILL_2_BUFX2_insert260 (
);

FILL FILL_1__10689_ (
);

FILL FILL_2_BUFX2_insert261 (
);

FILL FILL_1__10269_ (
);

FILL FILL_2_BUFX2_insert262 (
);

FILL FILL_2_BUFX2_insert263 (
);

FILL FILL_2_BUFX2_insert264 (
);

FILL FILL_4__11603_ (
);

FILL FILL_2_BUFX2_insert265 (
);

FILL FILL_0__7696_ (
);

FILL FILL_5__15082_ (
);

FILL FILL_2_BUFX2_insert266 (
);

FILL FILL_2_BUFX2_insert267 (
);

INVX1 _9382_ (
    .A(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_1269_)
);

FILL FILL_2_BUFX2_insert268 (
);

FILL FILL_2_BUFX2_insert269 (
);

FILL FILL_4__14495_ (
);

FILL FILL_1__11630_ (
);

FILL FILL_4__14075_ (
);

FILL FILL_1__11210_ (
);

FILL FILL_0__15908_ (
);

FILL FILL_2__8655_ (
);

FILL FILL_0__10623_ (
);

FILL FILL_2__8235_ (
);

FILL FILL_3__13488_ (
);

NOR2X1 _13380_ (
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3892_)
);

FILL FILL_0__13095_ (
);

FILL FILL_5__13815_ (
);

FILL SFILL38920x22050 (
);

FILL FILL_4__9522_ (
);

FILL FILL_4__9102_ (
);

FILL FILL_2__13842_ (
);

FILL FILL_2__13422_ (
);

FILL FILL_5__16287_ (
);

FILL FILL_2__13002_ (
);

FILL FILL_1__12835_ (
);

FILL FILL_1__12415_ (
);

FILL FILL_0__9422_ (
);

FILL FILL_0__11828_ (
);

FILL FILL_0__9002_ (
);

FILL FILL_0__11408_ (
);

FILL SFILL38840x29050 (
);

FILL FILL_5__7865_ (
);

FILL FILL_5__7445_ (
);

FILL FILL_4__16221_ (
);

INVX1 _14585_ (
    .A(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_5074_)
);

INVX1 _14165_ (
    .A(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_4663_)
);

FILL FILL_3__15634_ (
);

FILL FILL_3__15214_ (
);

FILL SFILL3560x21050 (
);

FILL FILL_1__7857_ (
);

FILL FILL_1__7437_ (
);

FILL SFILL38440x15050 (
);

FILL FILL_2__14627_ (
);

FILL FILL_0__15661_ (
);

FILL FILL_2__14207_ (
);

FILL FILL_0__15241_ (
);

FILL FILL112200x16050 (
);

FILL FILL_1_BUFX2_insert280 (
);

FILL FILL_1_BUFX2_insert281 (
);

FILL FILL_3__8724_ (
);

FILL FILL_1_BUFX2_insert282 (
);

FILL FILL_1_BUFX2_insert283 (
);

FILL FILL_1_BUFX2_insert284 (
);

FILL FILL_1_BUFX2_insert285 (
);

FILL SFILL3480x28050 (
);

FILL FILL_1_BUFX2_insert286 (
);

FILL FILL_1_BUFX2_insert287 (
);

FILL FILL_1_BUFX2_insert288 (
);

FILL FILL_6__11947_ (
);

FILL FILL_1_BUFX2_insert289 (
);

FILL FILL_4__12981_ (
);

FILL FILL_4__12141_ (
);

DFFSR _10085_ (
    .Q(\datapath_1.regfile_1.regOut[25] [15]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_1563_[15])
);

FILL FILL_3__11974_ (
);

FILL FILL_3__11554_ (
);

FILL FILL_3__11134_ (
);

FILL FILL_0__16026_ (
);

OAI22X1 _16311_ (
    .A(_5518__bF$buf0),
    .B(_5454_),
    .C(_5503__bF$buf1),
    .D(_6759_),
    .Y(_6760_)
);

FILL FILL_2__10967_ (
);

FILL FILL_2__10547_ (
);

FILL FILL_2__10127_ (
);

FILL FILL_0__11581_ (
);

FILL FILL_0__11161_ (
);

FILL SFILL115000x49050 (
);

FILL FILL_3__9929_ (
);

FILL FILL_3__9509_ (
);

FILL FILL_5__14773_ (
);

FILL FILL_0__6967_ (
);

FILL FILL_5__14353_ (
);

INVX1 _8653_ (
    .A(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_905_)
);

INVX1 _8233_ (
    .A(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_686_)
);

FILL FILL_1__7190_ (
);

FILL SFILL28840x27050 (
);

FILL FILL_1__10901_ (
);

FILL FILL_4__13766_ (
);

FILL FILL_4__13346_ (
);

FILL FILL_2__14380_ (
);

FILL FILL_2__7926_ (
);

FILL FILL_3__12759_ (
);

FILL FILL_2__7506_ (
);

FILL FILL_1__13793_ (
);

FILL FILL_3__12339_ (
);

FILL FILL_1__13373_ (
);

FILL SFILL18920x63050 (
);

FILL FILL_0__12786_ (
);

INVX1 _12651_ (
    .A(\datapath_1.Data [28]),
    .Y(_3480_)
);

FILL FILL_0__12366_ (
);

NAND3X1 _12231_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3212_)
);

FILL FILL_3__13700_ (
);

FILL FILL_6__16145_ (
);

FILL FILL_5__15978_ (
);

FILL FILL_5__15558_ (
);

FILL FILL_5__15138_ (
);

INVX1 _9858_ (
    .A(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_1505_)
);

FILL FILL_3__16172_ (
);

DFFSR _9438_ (
    .Q(\datapath_1.regfile_1.regOut[20] [8]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_1238_[8])
);

FILL FILL_5__10693_ (
);

OAI21X1 _9018_ (
    .A(_1086_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .C(_1087_),
    .Y(_1043_[22])
);

FILL FILL_1__8395_ (
);

FILL FILL_5__10273_ (
);

FILL FILL_2__15585_ (
);

FILL FILL_2__15165_ (
);

FILL FILL_1__14998_ (
);

FILL FILL_1__14578_ (
);

FILL FILL_1__14158_ (
);

FILL FILL_4__15912_ (
);

FILL FILL_3__9682_ (
);

INVX1 _13856_ (
    .A(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_4360_)
);

FILL FILL_3__9262_ (
);

INVX8 _13436_ (
    .A(_3947__bF$buf2),
    .Y(_3948_)
);

OAI21X1 _13016_ (
    .A(_3661_),
    .B(vdd),
    .C(_3662_),
    .Y(_3620_[21])
);

FILL FILL_3__14905_ (
);

FILL FILL_6__12065_ (
);

FILL FILL_0__14932_ (
);

FILL FILL_0__14512_ (
);

FILL FILL_5__11898_ (
);

FILL FILL_5__11478_ (
);

FILL FILL_5__11058_ (
);

FILL FILL_3__12092_ (
);

FILL FILL_4__7185_ (
);

FILL FILL_2__11085_ (
);

FILL FILL_1__10498_ (
);

FILL FILL_4__11832_ (
);

FILL FILL_4__11412_ (
);

FILL FILL_0__7085_ (
);

FILL FILL_1__16304_ (
);

DFFSR _9191_ (
    .Q(\datapath_1.regfile_1.regOut[18] [17]),
    .CLK(clk_bF$buf107),
    .R(rst_bF$buf31),
    .S(vdd),
    .D(_1108_[17])
);

FILL FILL_3__10825_ (
);

FILL FILL_3__10405_ (
);

FILL FILL_0__15717_ (
);

FILL FILL_2__8884_ (
);

FILL FILL_2__8464_ (
);

FILL FILL_3__13297_ (
);

FILL FILL_0__10432_ (
);

FILL FILL_0__10012_ (
);

FILL FILL_6__14631_ (
);

FILL FILL_6__14211_ (
);

FILL FILL_5__13624_ (
);

DFFSR _7924_ (
    .Q(\datapath_1.regfile_1.regOut[8] [30]),
    .CLK(clk_bF$buf106),
    .R(rst_bF$buf108),
    .S(vdd),
    .D(_458_[30])
);

INVX1 _7504_ (
    .A(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_322_)
);

FILL FILL_1__6881_ (
);

FILL FILL_4__9751_ (
);

FILL FILL_4__12617_ (
);

FILL FILL_2__13651_ (
);

FILL FILL_2__13231_ (
);

FILL FILL_5__16096_ (
);

FILL FILL_1__12644_ (
);

FILL FILL_1__12224_ (
);

FILL FILL_4__15089_ (
);

FILL FILL_2__9669_ (
);

FILL FILL_0__9651_ (
);

FILL FILL_0__9231_ (
);

FILL FILL_2__9249_ (
);

OAI21X1 _11922_ (
    .A(_2988_),
    .B(IorD_bF$buf4),
    .C(_2989_),
    .Y(_1_[11])
);

FILL FILL_0__11637_ (
);

FILL SFILL114520x73050 (
);

FILL FILL_0__11217_ (
);

NOR2X1 _11502_ (
    .A(_2614_),
    .B(_2574_),
    .Y(_2615_)
);

FILL SFILL53880x63050 (
);

FILL FILL_5__7674_ (
);

FILL FILL_4__16450_ (
);

FILL FILL_4__16030_ (
);

FILL FILL_6__10971_ (
);

INVX1 _14394_ (
    .A(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_4887_)
);

FILL FILL_5__14829_ (
);

FILL FILL_5__14409_ (
);

FILL FILL_3__15863_ (
);

FILL FILL_3__15443_ (
);

FILL FILL_3__15023_ (
);

INVX1 _8709_ (
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_922_)
);

FILL FILL_1__7246_ (
);

FILL SFILL94600x7050 (
);

FILL SFILL69080x34050 (
);

FILL FILL_2__14856_ (
);

FILL FILL_0__15890_ (
);

FILL FILL_2__14436_ (
);

FILL FILL_2__14016_ (
);

FILL FILL_0__15470_ (
);

FILL FILL_0__15050_ (
);

FILL FILL_1__13849_ (
);

FILL FILL_1__13429_ (
);

FILL FILL_1__13009_ (
);

FILL FILL_3__8953_ (
);

FILL FILL_3__8533_ (
);

INVX1 _12707_ (
    .A(\aluControl_1.inst [4]),
    .Y(_3497_)
);

FILL FILL_3__8113_ (
);

FILL FILL_5__8879_ (
);

FILL FILL_5__8459_ (
);

FILL FILL_4__12790_ (
);

OAI22X1 _15599_ (
    .A(_4602_),
    .B(_5539__bF$buf0),
    .C(_5526__bF$buf4),
    .D(_4606_),
    .Y(_6066_)
);

INVX1 _15179_ (
    .A(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_5656_)
);

FILL FILL_4__12370_ (
);

FILL FILL_3__16228_ (
);

FILL FILL_2__6950_ (
);

FILL FILL_5__10749_ (
);

FILL FILL_3__11783_ (
);

FILL FILL_5__9400_ (
);

FILL FILL_3__11363_ (
);

FILL SFILL59080x77050 (
);

FILL FILL_4__6876_ (
);

FILL FILL_0__16255_ (
);

OAI22X1 _16120_ (
    .A(_5463__bF$buf1),
    .B(_6573_),
    .C(_6572_),
    .D(_5504__bF$buf3),
    .Y(_6574_)
);

FILL FILL_2__10776_ (
);

FILL FILL_0__11390_ (
);

FILL FILL_1__9812_ (
);

FILL FILL_3__9738_ (
);

FILL SFILL3640x54050 (
);

FILL FILL_5__14582_ (
);

FILL FILL_5__14162_ (
);

INVX1 _8882_ (
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_1017_)
);

INVX1 _8462_ (
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_798_)
);

DFFSR _8042_ (
    .Q(\datapath_1.regfile_1.regOut[9] [20]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_523_[20])
);

FILL SFILL104520x71050 (
);

FILL SFILL43880x61050 (
);

FILL FILL_4__13995_ (
);

FILL FILL_4__13575_ (
);

FILL FILL_4__13155_ (
);

NAND2X1 _11099_ (
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2218_)
);

FILL FILL_2__7735_ (
);

FILL FILL_3__12988_ (
);

FILL FILL_3__12568_ (
);

FILL FILL_2__7315_ (
);

FILL FILL_3__12148_ (
);

FILL SFILL59000x75050 (
);

FILL SFILL59080x32050 (
);

FILL FILL_0__12595_ (
);

INVX1 _12880_ (
    .A(\datapath_1.a [19]),
    .Y(_3592_)
);

INVX1 _12460_ (
    .A(ALUOut[7]),
    .Y(_3373_)
);

FILL FILL_0__12175_ (
);

NAND3X1 _12040_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [13]),
    .C(_3034__bF$buf3),
    .Y(_3076_)
);

FILL SFILL104440x78050 (
);

FILL FILL_4__8602_ (
);

FILL FILL_5_BUFX2_insert510 (
);

FILL FILL_5_BUFX2_insert511 (
);

FILL FILL_5__15787_ (
);

FILL FILL_5__15367_ (
);

FILL FILL_2__12502_ (
);

FILL FILL_5_BUFX2_insert512 (
);

FILL FILL_5_BUFX2_insert513 (
);

FILL FILL_5_BUFX2_insert514 (
);

OAI21X1 _9667_ (
    .A(_1417_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .C(_1418_),
    .Y(_1368_[25])
);

FILL FILL_5_BUFX2_insert515 (
);

OAI21X1 _9247_ (
    .A(_1198_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1199_),
    .Y(_1173_[13])
);

FILL FILL_6__8108_ (
);

FILL FILL_5_BUFX2_insert516 (
);

FILL FILL_5_BUFX2_insert517 (
);

FILL FILL_5_BUFX2_insert518 (
);

FILL FILL_1__11915_ (
);

FILL FILL_5_BUFX2_insert519 (
);

FILL FILL_2__15394_ (
);

FILL FILL_0__8502_ (
);

FILL FILL_0__10908_ (
);

FILL FILL_1__14387_ (
);

FILL FILL_5__6945_ (
);

FILL FILL_4__15721_ (
);

FILL FILL_1_BUFX2_insert1040 (
);

FILL FILL_4__15301_ (
);

FILL FILL_1_BUFX2_insert1041 (
);

FILL FILL_1_BUFX2_insert1042 (
);

FILL SFILL59000x30050 (
);

FILL FILL_1_BUFX2_insert1043 (
);

FILL FILL_3__9491_ (
);

FILL SFILL49080x75050 (
);

FILL FILL_1_BUFX2_insert1044 (
);

AOI22X1 _13665_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [4]),
    .C(\datapath_1.regfile_1.regOut[6] [4]),
    .D(_4001__bF$buf0),
    .Y(_4173_)
);

AND2X2 _13245_ (
    .A(_3787_),
    .B(_3785_),
    .Y(_3788_)
);

FILL FILL_1_BUFX2_insert1045 (
);

FILL FILL_1_BUFX2_insert1046 (
);

FILL FILL_1_BUFX2_insert1047 (
);

FILL FILL_3__14714_ (
);

FILL FILL_1_BUFX2_insert1048 (
);

FILL SFILL3560x16050 (
);

FILL FILL_1_BUFX2_insert1049 (
);

FILL FILL_1__6937_ (
);

FILL FILL_4__9807_ (
);

FILL SFILL104440x33050 (
);

FILL FILL_2__13707_ (
);

FILL FILL_0__14741_ (
);

FILL FILL_0__14321_ (
);

FILL FILL_5__11287_ (
);

FILL FILL_2__16179_ (
);

FILL FILL_3__7804_ (
);

FILL SFILL108760x41050 (
);

FILL FILL_2_BUFX2_insert640 (
);

FILL FILL_2_BUFX2_insert641 (
);

FILL FILL_2_BUFX2_insert642 (
);

FILL SFILL49000x73050 (
);

FILL FILL_2_BUFX2_insert643 (
);

FILL FILL_2_BUFX2_insert644 (
);

FILL FILL_4__11641_ (
);

FILL FILL_2_BUFX2_insert645 (
);

FILL FILL_4__11221_ (
);

FILL FILL_3__15919_ (
);

FILL FILL_2_BUFX2_insert646 (
);

FILL FILL_2_BUFX2_insert647 (
);

FILL FILL_2_BUFX2_insert648 (
);

FILL SFILL49080x30050 (
);

FILL FILL_2_BUFX2_insert649 (
);

FILL FILL_1__16113_ (
);

FILL FILL_3__10634_ (
);

FILL FILL_6__13079_ (
);

FILL SFILL28920x15050 (
);

FILL FILL_0__15946_ (
);

FILL FILL_0__15526_ (
);

NOR3X1 _15811_ (
    .A(_6262_),
    .B(_6250_),
    .C(_6272_),
    .Y(_6273_)
);

FILL FILL_0__15106_ (
);

FILL FILL_0__10661_ (
);

FILL FILL_2__8273_ (
);

FILL FILL_0__10241_ (
);

FILL FILL_4__8199_ (
);

FILL FILL_2__12099_ (
);

FILL FILL_5__13853_ (
);

FILL FILL_5__13433_ (
);

FILL FILL_5__13013_ (
);

INVX1 _7733_ (
    .A(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_434_)
);

INVX1 _7313_ (
    .A(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_215_)
);

FILL FILL_4__9980_ (
);

FILL FILL_4__12846_ (
);

FILL FILL_4__9140_ (
);

FILL FILL_2__13880_ (
);

FILL FILL_4__12426_ (
);

FILL FILL_2__13460_ (
);

FILL FILL_4__12006_ (
);

FILL FILL_2__13040_ (
);

FILL FILL_0__8099_ (
);

FILL SFILL114600x6050 (
);

FILL FILL_3__11839_ (
);

FILL FILL_1__12873_ (
);

FILL FILL_3__11419_ (
);

FILL FILL_1__12453_ (
);

FILL FILL_1__12033_ (
);

FILL FILL_0__9880_ (
);

FILL FILL_2__9898_ (
);

FILL SFILL79160x69050 (
);

FILL FILL_0__11866_ (
);

FILL FILL_2__9478_ (
);

FILL FILL_0__9040_ (
);

FILL FILL_0__11446_ (
);

OAI21X1 _11731_ (
    .A(_2826_),
    .B(_2168_),
    .C(_2470__bF$buf1),
    .Y(_2828_)
);

FILL FILL_0__11026_ (
);

INVX2 _11311_ (
    .A(_2234_),
    .Y(_2430_)
);

FILL FILL_5__7483_ (
);

FILL FILL_5__7063_ (
);

FILL FILL_5__14638_ (
);

FILL FILL_5__14218_ (
);

FILL FILL_3__15672_ (
);

FILL FILL_3__15252_ (
);

DFFSR _8938_ (
    .Q(\datapath_1.regfile_1.regOut[16] [20]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_978_[20])
);

OAI21X1 _8518_ (
    .A(_834_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .C(_835_),
    .Y(_783_[26])
);

FILL FILL_1__7475_ (
);

FILL FILL_1__7055_ (
);

FILL FILL_2__14665_ (
);

FILL FILL111800x73050 (
);

FILL FILL_2__14245_ (
);

FILL SFILL63960x53050 (
);

FILL SFILL39000x71050 (
);

FILL SFILL94360x44050 (
);

FILL FILL_1__13658_ (
);

FILL FILL_1__13238_ (
);

FILL FILL_1_BUFX2_insert660 (
);

FILL FILL_3__8762_ (
);

FILL FILL_1_BUFX2_insert661 (
);

DFFSR _12936_ (
    .Q(\datapath_1.a [17]),
    .CLK(clk_bF$buf2),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_3555_[17])
);

FILL FILL_1_BUFX2_insert662 (
);

FILL FILL_3__8342_ (
);

OAI21X1 _12516_ (
    .A(_3409_),
    .B(vdd),
    .C(_3410_),
    .Y(_3360_[25])
);

FILL FILL_1_BUFX2_insert663 (
);

FILL FILL_1_BUFX2_insert664 (
);

FILL FILL_1_BUFX2_insert665 (
);

FILL SFILL98680x52050 (
);

FILL FILL_1_BUFX2_insert666 (
);

FILL SFILL79160x24050 (
);

FILL FILL_5__8268_ (
);

FILL FILL_1_BUFX2_insert667 (
);

FILL FILL_1_BUFX2_insert668 (
);

FILL FILL_1_BUFX2_insert669 (
);

FILL FILL_3__16037_ (
);

FILL SFILL103640x29050 (
);

FILL FILL_5__10978_ (
);

FILL FILL_5__10558_ (
);

FILL FILL_5__10138_ (
);

FILL FILL_3__11592_ (
);

FILL FILL_3__11172_ (
);

FILL FILL_0__16064_ (
);

FILL FILL_2__10165_ (
);

FILL FILL_1__9621_ (
);

FILL FILL_3__9547_ (
);

FILL FILL_4__10912_ (
);

FILL FILL_3__9127_ (
);

FILL FILL_5__14391_ (
);

DFFSR _8691_ (
    .Q(\datapath_1.regfile_1.regOut[14] [29]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_848_[29])
);

FILL FILL_1__15804_ (
);

OAI21X1 _8271_ (
    .A(_710_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .C(_711_),
    .Y(_653_[29])
);

FILL FILL_4__13384_ (
);

FILL SFILL8760x61050 (
);

FILL FILL_2__7964_ (
);

FILL FILL_2__7544_ (
);

BUFX2 BUFX2_insert330 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf3 )
);

FILL FILL_3__12377_ (
);

FILL FILL_2__7124_ (
);

BUFX2 BUFX2_insert331 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf2 )
);

BUFX2 BUFX2_insert332 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf1 )
);

BUFX2 BUFX2_insert333 (
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf0 )
);

BUFX2 BUFX2_insert334 (
    .A(_4005_),
    .Y(_4005__bF$buf3)
);

BUFX2 BUFX2_insert335 (
    .A(_4005_),
    .Y(_4005__bF$buf2)
);

BUFX2 BUFX2_insert336 (
    .A(_4005_),
    .Y(_4005__bF$buf1)
);

BUFX2 BUFX2_insert337 (
    .A(_4005_),
    .Y(_4005__bF$buf0)
);

BUFX2 BUFX2_insert338 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf3 )
);

BUFX2 BUFX2_insert339 (
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf2 )
);

FILL SFILL114600x61050 (
);

FILL SFILL99400x9050 (
);

FILL FILL_5__12704_ (
);

FILL SFILL53960x51050 (
);

FILL FILL_4__8831_ (
);

FILL FILL_2__12731_ (
);

FILL FILL_5__15596_ (
);

FILL FILL_5__15176_ (
);

FILL FILL_2__12311_ (
);

OAI21X1 _9896_ (
    .A(_1529_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1530_),
    .Y(_1498_[16])
);

OAI21X1 _9476_ (
    .A(_1310_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .C(_1311_),
    .Y(_1303_[4])
);

DFFSR _9056_ (
    .Q(\datapath_1.regfile_1.regOut[17] [10]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_1043_[10])
);

FILL FILL_4__14589_ (
);

FILL FILL_1__11724_ (
);

FILL FILL_4__14169_ (
);

FILL FILL_1__11304_ (
);

FILL FILL_0__8731_ (
);

FILL FILL_2__8749_ (
);

FILL SFILL114520x68050 (
);

FILL FILL_2__8329_ (
);

FILL FILL_0__8311_ (
);

FILL FILL_1__14196_ (
);

FILL FILL_4__15950_ (
);

FILL FILL_4__15530_ (
);

FILL FILL_4__15110_ (
);

NOR2X1 _13894_ (
    .A(_4396_),
    .B(_4393_),
    .Y(_4397_)
);

NAND2X1 _13474_ (
    .A(_3974_),
    .B(_3985_),
    .Y(_3986_)
);

DFFSR _13054_ (
    .Q(_2_[7]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3620_[7])
);

FILL FILL_5__13909_ (
);

FILL FILL_3__14943_ (
);

FILL FILL_3__14523_ (
);

FILL FILL_3__14103_ (
);

FILL FILL_4__9616_ (
);

FILL SFILL69080x29050 (
);

FILL FILL_2__13936_ (
);

FILL FILL_0__14970_ (
);

FILL FILL_2__13516_ (
);

FILL FILL_0__14550_ (
);

FILL FILL_0__14130_ (
);

FILL FILL_5__11096_ (
);

FILL FILL_1__12509_ (
);

FILL FILL_0__9936_ (
);

FILL FILL_3__7613_ (
);

FILL FILL_0__9516_ (
);

FILL FILL_5__7959_ (
);

FILL SFILL114520x23050 (
);

FILL FILL_5__7119_ (
);

FILL FILL_4__16315_ (
);

FILL FILL_4__11870_ (
);

NOR2X1 _14679_ (
    .A(_5165_),
    .B(_5162_),
    .Y(_5166_)
);

OAI22X1 _14259_ (
    .A(_3983__bF$buf0),
    .B(_4753_),
    .C(_3977__bF$buf1),
    .D(_4754_),
    .Y(_4755_)
);

FILL FILL_4__11450_ (
);

FILL FILL_4__11030_ (
);

FILL SFILL3720x42050 (
);

FILL FILL_3__15728_ (
);

FILL FILL_3__15308_ (
);

FILL FILL_1__16342_ (
);

FILL FILL_5__8900_ (
);

FILL FILL_3__10443_ (
);

FILL FILL_3__10023_ (
);

FILL FILL_0__15755_ (
);

AOI22X1 _15620_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [14]),
    .C(\datapath_1.regfile_1.regOut[22] [14]),
    .D(_5650_),
    .Y(_6086_)
);

FILL FILL_0__15335_ (
);

OAI22X1 _15200_ (
    .A(_5499__bF$buf2),
    .B(_5676_),
    .C(_5532__bF$buf3),
    .D(_5675_),
    .Y(_5677_)
);

FILL FILL_0__10890_ (
);

FILL FILL_2__8082_ (
);

FILL FILL_0__10050_ (
);

FILL SFILL3640x49050 (
);

FILL FILL_5__13662_ (
);

FILL FILL_5__13242_ (
);

INVX1 _7962_ (
    .A(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_546_)
);

INVX1 _7542_ (
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_391_)
);

FILL SFILL104520x66050 (
);

OAI21X1 _7122_ (
    .A(_127_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .C(_128_),
    .Y(_68_[30])
);

FILL FILL_4__12655_ (
);

FILL FILL_4__12235_ (
);

DFFSR _10599_ (
    .Q(\datapath_1.regfile_1.regOut[29] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_1823_[17])
);

OAI21X1 _10179_ (
    .A(_1677_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .C(_1678_),
    .Y(_1628_[25])
);

FILL FILL_3__11648_ (
);

FILL FILL_3__11228_ (
);

FILL FILL_1__12262_ (
);

INVX1 _16405_ (
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_6824_)
);

FILL SFILL59080x27050 (
);

FILL FILL112280x60050 (
);

NAND2X1 _11960_ (
    .A(IorD_bF$buf2),
    .B(ALUOut[24]),
    .Y(_3015_)
);

FILL FILL_2__9287_ (
);

FILL FILL_0__11675_ (
);

FILL FILL_0__11255_ (
);

NAND3X1 _11540_ (
    .A(_2470__bF$buf0),
    .B(_2646_),
    .C(_2650_),
    .Y(_2651_)
);

NOR2X1 _11120_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2239_)
);

FILL FILL_6__15874_ (
);

FILL FILL_6__15454_ (
);

FILL FILL_5__7292_ (
);

FILL FILL_5__14867_ (
);

FILL FILL_5__14447_ (
);

FILL FILL_5__14027_ (
);

FILL FILL_3__15481_ (
);

FILL FILL_3__15061_ (
);

OAI21X1 _8747_ (
    .A(_946_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .C(_947_),
    .Y(_913_[17])
);

OAI21X1 _8327_ (
    .A(_727_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .C(_728_),
    .Y(_718_[5])
);

FILL FILL_2__14894_ (
);

FILL FILL_2__14474_ (
);

FILL SFILL104520x21050 (
);

FILL FILL_2__14054_ (
);

FILL SFILL43880x11050 (
);

FILL FILL_1__13887_ (
);

FILL FILL_1__13467_ (
);

FILL FILL_4__14801_ (
);

FILL SFILL59000x25050 (
);

FILL FILL_3__8991_ (
);

FILL FILL_3__8571_ (
);

OAI21X1 _12745_ (
    .A(_3521_),
    .B(IRWrite_bF$buf1),
    .C(_3522_),
    .Y(_3490_[16])
);

AOI22X1 _12325_ (
    .A(_2_[27]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3283_)
);

FILL FILL_5__8497_ (
);

FILL FILL_5__8077_ (
);

FILL FILL_6__11794_ (
);

FILL FILL_6__11374_ (
);

FILL SFILL104440x28050 (
);

FILL FILL_0__13821_ (
);

FILL FILL_0__13401_ (
);

FILL FILL_3__16266_ (
);

FILL FILL_5__10787_ (
);

FILL FILL_5__10367_ (
);

FILL FILL_1__8489_ (
);

FILL FILL_1__8069_ (
);

FILL FILL_2__15679_ (
);

FILL FILL_2__15259_ (
);

FILL FILL_0__16293_ (
);

FILL SFILL33880x54050 (
);

FILL FILL_2__10394_ (
);

FILL FILL_1__9850_ (
);

FILL FILL_1__9010_ (
);

FILL FILL_2__16200_ (
);

FILL FILL_3__9776_ (
);

FILL FILL_3__9356_ (
);

FILL SFILL113720x19050 (
);

FILL FILL_4__10301_ (
);

FILL SFILL49080x25050 (
);

FILL FILL_1__15613_ (
);

OAI21X1 _8080_ (
    .A(_603_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .C(_604_),
    .Y(_588_[8])
);

FILL SFILL94440x77050 (
);

FILL FILL_0__14606_ (
);

FILL FILL_2__7353_ (
);

FILL FILL_3__12186_ (
);

FILL FILL_6__13940_ (
);

FILL FILL_4__7699_ (
);

FILL FILL_6__13100_ (
);

FILL FILL_2__11599_ (
);

FILL FILL_2__11179_ (
);

FILL FILL_5__12513_ (
);

FILL FILL_4__8640_ (
);

FILL FILL_4__8220_ (
);

FILL FILL_4__11926_ (
);

FILL FILL_2__12960_ (
);

FILL FILL_4__11506_ (
);

FILL FILL_6__8986_ (
);

FILL FILL_0__7599_ (
);

FILL FILL_2__12120_ (
);

FILL SFILL49000x23050 (
);

FILL FILL_0__7179_ (
);

NAND2X1 _9285_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1225_)
);

FILL FILL_3__10919_ (
);

FILL FILL_1__11953_ (
);

FILL FILL_4__14398_ (
);

FILL FILL_1__11533_ (
);

FILL FILL_1__11113_ (
);

FILL FILL_0__8960_ (
);

FILL FILL_2__8978_ (
);

FILL SFILL94440x32050 (
);

FILL FILL_0__10946_ (
);

INVX1 _10811_ (
    .A(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_1998_)
);

FILL FILL_0__8120_ (
);

FILL FILL_2__8138_ (
);

FILL FILL_0__10526_ (
);

FILL FILL_0__10106_ (
);

FILL FILL_5__6983_ (
);

NOR2X1 _13283_ (
    .A(_3812_),
    .B(_3773_),
    .Y(_3822_)
);

FILL FILL_5__13718_ (
);

FILL SFILL23880x52050 (
);

FILL FILL_3__14752_ (
);

FILL FILL_3__14332_ (
);

FILL FILL_1__6975_ (
);

FILL FILL_4__9425_ (
);

FILL FILL_4__9005_ (
);

FILL FILL_2__13745_ (
);

FILL FILL_2__13325_ (
);

FILL SFILL39000x66050 (
);

FILL SFILL94360x39050 (
);

FILL FILL_1__12738_ (
);

FILL FILL_1__12318_ (
);

FILL FILL_3__7842_ (
);

FILL FILL_0__9745_ (
);

FILL FILL_3__7422_ (
);

FILL SFILL63560x34050 (
);

FILL FILL_5__7348_ (
);

FILL FILL_4__16124_ (
);

INVX1 _14488_ (
    .A(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_4979_)
);

OAI22X1 _14068_ (
    .A(_4566_),
    .B(_3936__bF$buf3),
    .C(_3902__bF$buf2),
    .D(_4567_),
    .Y(_4568_)
);

FILL FILL_3__15957_ (
);

FILL FILL_3__15537_ (
);

FILL FILL_3__15117_ (
);

FILL FILL_1__16151_ (
);

FILL FILL_3__10672_ (
);

FILL FILL_3__10252_ (
);

FILL FILL_0__15984_ (
);

FILL FILL_0__15564_ (
);

FILL FILL_0__15144_ (
);

FILL SFILL79160x9050 (
);

FILL SFILL39000x21050 (
);

FILL FILL_1__8701_ (
);

FILL SFILL4440x48050 (
);

FILL FILL_3__8627_ (
);

FILL FILL_3__8207_ (
);

FILL FILL_5__13891_ (
);

FILL FILL_5__13471_ (
);

DFFSR _7771_ (
    .Q(\datapath_1.regfile_1.regOut[7] [5]),
    .CLK(clk_bF$buf60),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_393_[5])
);

FILL SFILL78520x6050 (
);

OAI21X1 _7351_ (
    .A(_239_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_240_),
    .Y(_198_[21])
);

FILL FILL_4__12884_ (
);

FILL FILL_4__12464_ (
);

FILL SFILL8760x56050 (
);

FILL FILL_4__12044_ (
);

FILL FILL_3__11877_ (
);

FILL FILL_5__9914_ (
);

FILL FILL_3__11457_ (
);

FILL FILL_1__12491_ (
);

FILL FILL_3__11037_ (
);

FILL FILL_1__12071_ (
);

FILL FILL_0__16349_ (
);

AND2X2 _16214_ (
    .A(_5494_),
    .B(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_6665_)
);

FILL FILL_2__9096_ (
);

FILL FILL_0__11484_ (
);

FILL FILL_0__11064_ (
);

FILL SFILL53960x46050 (
);

FILL FILL_1__9906_ (
);

FILL SFILL29000x64050 (
);

FILL SFILL84360x37050 (
);

FILL FILL_2__11811_ (
);

FILL FILL_5__14676_ (
);

FILL FILL_5__14256_ (
);

OAI21X1 _8976_ (
    .A(_1058_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .C(_1059_),
    .Y(_1043_[8])
);

FILL FILL_3__15290_ (
);

DFFSR _8556_ (
    .Q(\datapath_1.regfile_1.regOut[13] [22]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_783_[22])
);

NAND2X1 _8136_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_642_)
);

FILL FILL_1__7093_ (
);

FILL FILL_4__13669_ (
);

FILL FILL_1__10804_ (
);

FILL FILL_4__13249_ (
);

FILL FILL_2__14283_ (
);

FILL FILL_0__7811_ (
);

FILL FILL_2__7829_ (
);

FILL FILL_1__13696_ (
);

FILL FILL_1__13276_ (
);

FILL SFILL78760x81050 (
);

FILL FILL_4__14610_ (
);

FILL FILL_3__8380_ (
);

OAI21X1 _12974_ (
    .A(_3633_),
    .B(vdd),
    .C(_3634_),
    .Y(_3620_[7])
);

DFFSR _12554_ (
    .Q(ALUOut[19]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3360_[19])
);

FILL FILL_0__12269_ (
);

NAND2X1 _12134_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.a [6]),
    .Y(_3143_)
);

FILL FILL_3__13603_ (
);

FILL FILL_6__16048_ (
);

FILL FILL_0__13630_ (
);

FILL FILL_0__13210_ (
);

FILL FILL_3__16075_ (
);

FILL FILL_5__10176_ (
);

FILL FILL_2__15488_ (
);

FILL FILL_2__15068_ (
);

FILL FILL_5__16402_ (
);

FILL FILL_4__15815_ (
);

FILL FILL_4__10950_ (
);

FILL FILL_3__9165_ (
);

NOR2X1 _13759_ (
    .A(_4261_),
    .B(_4264_),
    .Y(_4265_)
);

NAND2X1 _13339_ (
    .A(\datapath_1.a3 [4]),
    .B(_3822_),
    .Y(_3861_)
);

FILL FILL_4__10530_ (
);

FILL FILL_4__10110_ (
);

FILL FILL_3__14808_ (
);

FILL FILL_1__15842_ (
);

FILL FILL_1__15422_ (
);

FILL FILL_1__15002_ (
);

FILL SFILL43960x44050 (
);

FILL FILL_0__14835_ (
);

OAI22X1 _14700_ (
    .A(_3947__bF$buf0),
    .B(_5185_),
    .C(_3935__bF$buf1),
    .D(_5184_),
    .Y(_5186_)
);

FILL FILL_0__14415_ (
);

BUFX2 BUFX2_insert710 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf1 )
);

FILL FILL_2__7582_ (
);

BUFX2 BUFX2_insert711 (
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf0 )
);

FILL FILL_2__7162_ (
);

BUFX2 BUFX2_insert712 (
    .A(_5503_),
    .Y(_5503__bF$buf3)
);

BUFX2 BUFX2_insert713 (
    .A(_5503_),
    .Y(_5503__bF$buf2)
);

BUFX2 BUFX2_insert714 (
    .A(_5503_),
    .Y(_5503__bF$buf1)
);

BUFX2 BUFX2_insert715 (
    .A(_5503_),
    .Y(_5503__bF$buf0)
);

FILL SFILL108920x62050 (
);

BUFX2 BUFX2_insert716 (
    .A(_3930_),
    .Y(_3930__bF$buf3)
);

FILL FILL_4__7088_ (
);

FILL SFILL38200x17050 (
);

BUFX2 BUFX2_insert717 (
    .A(_3930_),
    .Y(_3930__bF$buf2)
);

BUFX2 BUFX2_insert718 (
    .A(_3930_),
    .Y(_3930__bF$buf1)
);

BUFX2 BUFX2_insert719 (
    .A(_3930_),
    .Y(_3930__bF$buf0)
);

FILL FILL_5__12742_ (
);

FILL FILL_5__12322_ (
);

FILL SFILL48920x6050 (
);

FILL FILL_4__11735_ (
);

FILL FILL_4__11315_ (
);

FILL SFILL23880x4050 (
);

FILL FILL_1__16207_ (
);

NAND2X1 _9094_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1118_)
);

FILL FILL_3__10308_ (
);

FILL FILL_1__11762_ (
);

FILL FILL_1__11342_ (
);

OAI22X1 _15905_ (
    .A(_5526__bF$buf0),
    .B(_4976_),
    .C(_4979_),
    .D(_5527__bF$buf0),
    .Y(_6364_)
);

FILL FILL112280x55050 (
);

FILL FILL_2__8787_ (
);

FILL FILL_0__10755_ (
);

FILL FILL_2__8367_ (
);

INVX1 _10620_ (
    .A(\datapath_1.regfile_1.regOut[30] [2]),
    .Y(_1891_)
);

DFFSR _10200_ (
    .Q(\datapath_1.regfile_1.regOut[26] [2]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1628_[2])
);

FILL FILL_6__14114_ (
);

NAND2X1 _13092_ (
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [4]),
    .Y(_3693_)
);

FILL FILL_5__13947_ (
);

FILL FILL_5__13527_ (
);

FILL FILL_3__14981_ (
);

FILL FILL_3__14561_ (
);

FILL FILL_5__13107_ (
);

FILL FILL_3__14141_ (
);

OAI21X1 _7827_ (
    .A(_475_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_476_),
    .Y(_458_[9])
);

DFFSR _7407_ (
    .Q(\datapath_1.regfile_1.regOut[4] [25]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_198_[25])
);

FILL FILL_4_BUFX2_insert550 (
);

FILL FILL_4__9654_ (
);

FILL FILL_4_BUFX2_insert551 (
);

FILL FILL_4_BUFX2_insert552 (
);

FILL FILL_4__9234_ (
);

FILL FILL_4_BUFX2_insert553 (
);

FILL FILL_2__13974_ (
);

FILL SFILL104520x16050 (
);

FILL FILL_4_BUFX2_insert554 (
);

FILL FILL_2__13554_ (
);

FILL FILL_2__13134_ (
);

FILL FILL_4_BUFX2_insert555 (
);

FILL FILL_4_BUFX2_insert556 (
);

FILL FILL_4_BUFX2_insert557 (
);

FILL FILL_4_BUFX2_insert558 (
);

FILL FILL_4_BUFX2_insert559 (
);

FILL FILL_1__12967_ (
);

FILL FILL_1__12127_ (
);

FILL SFILL28600x29050 (
);

FILL FILL_0__9974_ (
);

FILL FILL_0__9554_ (
);

FILL FILL_3__7231_ (
);

FILL FILL_0__9134_ (
);

AOI22X1 _11825_ (
    .A(_2351_),
    .B(_2481__bF$buf1),
    .C(_2620_),
    .D(_2133_),
    .Y(_2915_)
);

OAI21X1 _11405_ (
    .A(_2507_),
    .B(_2518_),
    .C(_2521_),
    .Y(_2522_)
);

FILL FILL112280x10050 (
);

FILL FILL_5__7997_ (
);

FILL FILL_5__7577_ (
);

FILL FILL_4__16353_ (
);

FILL FILL_6__10874_ (
);

NOR2X1 _14297_ (
    .A(_4788_),
    .B(_4791_),
    .Y(_4792_)
);

FILL FILL_0__12901_ (
);

FILL FILL_3__15766_ (
);

FILL FILL_3__15346_ (
);

FILL FILL_1__16380_ (
);

FILL SFILL33080x66050 (
);

FILL FILL_1__7989_ (
);

FILL FILL_1__7569_ (
);

FILL FILL_3__10061_ (
);

FILL FILL_2__14759_ (
);

FILL SFILL94520x65050 (
);

FILL FILL_0__15793_ (
);

FILL FILL_2__14339_ (
);

FILL SFILL33880x49050 (
);

FILL FILL_0__15373_ (
);

FILL FILL_1__8510_ (
);

FILL FILL_2__15700_ (
);

FILL FILL_3__8856_ (
);

FILL FILL_3__8016_ (
);

FILL FILL_5__13280_ (
);

OAI21X1 _7580_ (
    .A(_351_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .C(_352_),
    .Y(_328_[12])
);

OAI21X1 _7160_ (
    .A(_196_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .C(_197_),
    .Y(_133_[0])
);

FILL FILL_4__12273_ (
);

FILL FILL_2__6853_ (
);

FILL FILL_5__9723_ (
);

FILL FILL_3__11686_ (
);

FILL FILL_3__11266_ (
);

DFFSR _16443_ (
    .Q(\datapath_1.regfile_1.regOut[0] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_6769_[26])
);

FILL FILL_0__16158_ (
);

INVX1 _16023_ (
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_6479_)
);

FILL FILL_2__10679_ (
);

FILL FILL_2__10259_ (
);

FILL FILL_0__11293_ (
);

FILL FILL_4__7720_ (
);

FILL FILL_3_BUFX2_insert570 (
);

FILL FILL_4__7300_ (
);

FILL FILL_3_BUFX2_insert571 (
);

FILL FILL_3_BUFX2_insert572 (
);

FILL SFILL18600x27050 (
);

FILL FILL_5__14485_ (
);

FILL FILL_3_BUFX2_insert573 (
);

FILL FILL_2__11620_ (
);

FILL SFILL49000x18050 (
);

FILL FILL_5__14065_ (
);

FILL FILL_2__11200_ (
);

FILL FILL_3_BUFX2_insert574 (
);

FILL FILL_3_BUFX2_insert575 (
);

NAND2X1 _8785_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_973_)
);

NAND2X1 _8365_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_754_)
);

FILL FILL_3_BUFX2_insert576 (
);

FILL FILL_3_BUFX2_insert577 (
);

FILL FILL_3_BUFX2_insert578 (
);

FILL FILL_3_BUFX2_insert579 (
);

FILL FILL_4__13898_ (
);

FILL FILL_4__13478_ (
);

FILL FILL_2__14092_ (
);

FILL SFILL94440x27050 (
);

FILL FILL_0__7620_ (
);

FILL FILL_0__7200_ (
);

FILL FILL_2__7218_ (
);

FILL FILL_1__13085_ (
);

NAND2X1 _12783_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[29]),
    .Y(_3548_)
);

FILL FILL_0__12498_ (
);

FILL SFILL84520x63050 (
);

OAI21X1 _12363_ (
    .A(_3306_),
    .B(MemToReg_bF$buf1),
    .C(_3307_),
    .Y(\datapath_1.mux_wd3.dout [6])
);

FILL FILL_0__12078_ (
);

FILL SFILL23880x47050 (
);

FILL FILL_3__13832_ (
);

FILL FILL_3__13412_ (
);

FILL FILL_4__8505_ (
);

FILL FILL_2__12825_ (
);

FILL FILL_2__12405_ (
);

FILL FILL_1__11818_ (
);

FILL SFILL23480x33050 (
);

FILL FILL_2__15297_ (
);

FILL FILL_5__16211_ (
);

FILL FILL_3__6922_ (
);

FILL FILL_0__8825_ (
);

FILL FILL_0__8405_ (
);

FILL FILL_5__6848_ (
);

FILL FILL_4__15624_ (
);

FILL FILL_4__15204_ (
);

AOI22X1 _13988_ (
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .B(_4005__bF$buf2),
    .C(_4001__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_4489_)
);

FILL FILL_3__9394_ (
);

AOI22X1 _13568_ (
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .C(\datapath_1.regfile_1.regOut[31] [2]),
    .D(_3995__bF$buf0),
    .Y(_4078_)
);

FILL SFILL23800x45050 (
);

INVX1 _13148_ (
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3730_)
);

FILL FILL_3__14617_ (
);

FILL FILL_1__15651_ (
);

FILL FILL_1__15231_ (
);

FILL FILL_0__14644_ (
);

FILL FILL_0__14224_ (
);

FILL SFILL39000x16050 (
);

FILL FILL_3__7707_ (
);

FILL FILL_5__12971_ (
);

FILL FILL_5__12131_ (
);

BUFX2 _6851_ (
    .A(_1_[13]),
    .Y(memoryAddress[13])
);

FILL FILL_4__16409_ (
);

FILL FILL_4__11964_ (
);

FILL FILL_4__11544_ (
);

FILL FILL_4__11124_ (
);

FILL FILL_1__16016_ (
);

FILL FILL_3__10957_ (
);

FILL FILL_1__11991_ (
);

FILL FILL_3__10537_ (
);

FILL FILL_1__11571_ (
);

FILL FILL_3__10117_ (
);

FILL FILL_1__11151_ (
);

FILL FILL_0__15849_ (
);

NOR2X1 _15714_ (
    .A(_6175_),
    .B(_6177_),
    .Y(_6178_)
);

FILL FILL_0__15429_ (
);

FILL FILL_0__15009_ (
);

FILL FILL_2__8596_ (
);

FILL FILL_0__10564_ (
);

FILL FILL_0__10144_ (
);

FILL FILL_5__13756_ (
);

FILL FILL_5__13336_ (
);

FILL FILL_3__14790_ (
);

FILL FILL_3__14370_ (
);

NAND2X1 _7636_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_390_)
);

NAND2X1 _7216_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_171_)
);

FILL FILL_4__9883_ (
);

FILL FILL_4__9463_ (
);

FILL FILL_4__12749_ (
);

FILL FILL_4__9043_ (
);

FILL FILL_2__13783_ (
);

FILL FILL_4__12329_ (
);

FILL FILL_2__13363_ (
);

FILL FILL_6__9389_ (
);

FILL FILL_2__6909_ (
);

FILL FILL_1__12776_ (
);

FILL FILL_1__12356_ (
);

FILL FILL_0__9783_ (
);

FILL FILL_3__7880_ (
);

FILL FILL_3__7460_ (
);

FILL FILL_0__11769_ (
);

FILL FILL_0__9363_ (
);

FILL FILL_3__7040_ (
);

FILL FILL_0__11349_ (
);

OAI21X1 _11634_ (
    .A(_2253_),
    .B(_2346_),
    .C(_2737_),
    .Y(_2738_)
);

INVX2 _11214_ (
    .A(ALUControl[1]),
    .Y(_2333_)
);

FILL FILL_4__16162_ (
);

FILL FILL_3__15995_ (
);

FILL FILL_0__12710_ (
);

FILL FILL_3__15575_ (
);

FILL FILL_3__15155_ (
);

FILL FILL_1__7798_ (
);

FILL FILL_1__7378_ (
);

FILL FILL_3__10290_ (
);

FILL FILL_2__14988_ (
);

FILL FILL_2__14568_ (
);

FILL FILL_2__14148_ (
);

FILL FILL_0__15182_ (
);

FILL FILL_5__15902_ (
);

FILL SFILL28760x1050 (
);

FILL SFILL28680x6050 (
);

FILL FILL_3__8245_ (
);

NAND2X1 _12839_ (
    .A(vdd),
    .B(\datapath_1.rd1 [5]),
    .Y(_3565_)
);

NAND2X1 _12419_ (
    .A(MemToReg_bF$buf0),
    .B(\datapath_1.Data [25]),
    .Y(_3345_)
);

FILL FILL_1__14922_ (
);

FILL FILL_1__14502_ (
);

FILL SFILL43960x39050 (
);

FILL FILL_4__12082_ (
);

FILL FILL_0__13915_ (
);

FILL FILL_5__9532_ (
);

FILL FILL_3__11495_ (
);

FILL FILL_5__9112_ (
);

FILL FILL_3__11075_ (
);

FILL FILL_0__16387_ (
);

AOI22X1 _16252_ (
    .A(\datapath_1.regfile_1.regOut[1] [30]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_6702_)
);

FILL FILL112360x43050 (
);

FILL FILL_2__10488_ (
);

FILL FILL_2__10068_ (
);

FILL FILL_5__11822_ (
);

FILL FILL_1__9524_ (
);

FILL FILL_5__11402_ (
);

FILL FILL_1__9104_ (
);

FILL FILL_4__10815_ (
);

FILL SFILL64040x52050 (
);

FILL FILL_5__14294_ (
);

FILL FILL_6__7875_ (
);

FILL FILL_1__15707_ (
);

NAND2X1 _8594_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_866_)
);

DFFSR _8174_ (
    .Q(\datapath_1.regfile_1.regOut[10] [24]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_588_[24])
);

FILL FILL_1__10422_ (
);

FILL FILL_4__13287_ (
);

FILL FILL_1__10002_ (
);

FILL FILL_2__7867_ (
);

FILL FILL_2__7447_ (
);

NAND2X1 _12592_ (
    .A(vdd),
    .B(memoryOutData[8]),
    .Y(_3441_)
);

INVX1 _12172_ (
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3168_)
);

FILL FILL_5__12607_ (
);

FILL FILL_3__13641_ (
);

FILL FILL_3__13221_ (
);

OAI21X1 _6907_ (
    .A(_4_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .C(_5_),
    .Y(_3_[1])
);

FILL FILL_4__8734_ (
);

FILL FILL_4__8314_ (
);

FILL FILL_2__12634_ (
);

FILL FILL_5__15499_ (
);

FILL FILL_2__12214_ (
);

FILL FILL_5__15079_ (
);

INVX1 _9799_ (
    .A(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_1486_)
);

INVX1 _9379_ (
    .A(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_1267_)
);

FILL SFILL54840x78050 (
);

FILL FILL_1__11627_ (
);

FILL FILL_1__11207_ (
);

FILL FILL_5__16020_ (
);

FILL FILL_0__8634_ (
);

INVX2 _10905_ (
    .A(\control_1.reg_state.dout [3]),
    .Y(_2052_)
);

FILL FILL_0__8214_ (
);

FILL FILL_1__14099_ (
);

FILL FILL_4__15853_ (
);

FILL FILL_4__15433_ (
);

FILL FILL_4__15013_ (
);

INVX1 _13797_ (
    .A(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_4302_)
);

NOR3X1 _13377_ (
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(\datapath_1.PCJump [19]),
    .C(\datapath_1.PCJump [18]),
    .Y(_3889_)
);

FILL FILL_3__14846_ (
);

FILL FILL_3__14426_ (
);

FILL FILL_1__15880_ (
);

FILL FILL_3__14006_ (
);

FILL FILL_1__15460_ (
);

FILL FILL_1__15040_ (
);

FILL FILL_4__9939_ (
);

FILL FILL_4__9519_ (
);

FILL FILL_2__13839_ (
);

FILL FILL_0__14873_ (
);

FILL FILL_2__13419_ (
);

FILL FILL_0__14453_ (
);

FILL FILL_0__14033_ (
);

FILL FILL_3__7936_ (
);

FILL FILL_0__9419_ (
);

FILL FILL_5__12780_ (
);

FILL FILL_5__12360_ (
);

FILL FILL_4__16218_ (
);

FILL FILL_4__11773_ (
);

FILL FILL_4__11353_ (
);

FILL SFILL58680x79050 (
);

FILL FILL_1__16245_ (
);

FILL FILL_3__10766_ (
);

FILL FILL_1__11380_ (
);

FILL FILL_0__15658_ (
);

NOR2X1 _15943_ (
    .A(_6394_),
    .B(_6400_),
    .Y(_6401_)
);

FILL FILL_0__15238_ (
);

NAND2X1 _15523_ (
    .A(_5987_),
    .B(_5991_),
    .Y(_5992_)
);

NOR3X1 _15103_ (
    .A(_5581_),
    .B(_5573_),
    .C(_5564_),
    .Y(_5582_)
);

FILL FILL_0__10793_ (
);

FILL FILL_0__10373_ (
);

FILL FILL_5__13985_ (
);

FILL FILL_2__10700_ (
);

FILL FILL_5__13565_ (
);

FILL FILL_5__13145_ (
);

FILL SFILL54360x26050 (
);

NAND2X1 _7865_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_502_)
);

NAND2X1 _7445_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_283_)
);

FILL FILL_4_BUFX2_insert930 (
);

DFFSR _7025_ (
    .Q(\datapath_1.regfile_1.regOut[1] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_3_[27])
);

FILL FILL_4_BUFX2_insert931 (
);

FILL FILL_4__9272_ (
);

FILL FILL_4_BUFX2_insert932 (
);

FILL FILL_4__12978_ (
);

FILL FILL_4_BUFX2_insert933 (
);

FILL FILL_2__13592_ (
);

FILL FILL_4__12138_ (
);

FILL FILL_4_BUFX2_insert934 (
);

FILL FILL_4_BUFX2_insert935 (
);

FILL FILL_2__13172_ (
);

FILL FILL_4_BUFX2_insert936 (
);

FILL FILL_4_BUFX2_insert937 (
);

FILL FILL_4_BUFX2_insert938 (
);

FILL FILL_4_BUFX2_insert939 (
);

FILL FILL_1__12585_ (
);

FILL FILL_1__12165_ (
);

FILL SFILL23080x59050 (
);

NAND2X1 _16308_ (
    .A(_6751_),
    .B(_6756_),
    .Y(_6757_)
);

FILL FILL_0__11998_ (
);

FILL FILL_0__9592_ (
);

NOR3X1 _11863_ (
    .A(_2946_),
    .B(_2949_),
    .C(_2947_),
    .Y(_2950_)
);

FILL FILL_0__9172_ (
);

FILL FILL_0__11578_ (
);

NOR2X1 _11443_ (
    .A(_2154_),
    .B(_2558_),
    .Y(_2559_)
);

FILL FILL_0__11158_ (
);

NOR2X1 _11023_ (
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2142_)
);

FILL FILL_3__12912_ (
);

FILL FILL_6__15777_ (
);

FILL SFILL109400x80050 (
);

FILL FILL_6__15357_ (
);

FILL FILL_5__7195_ (
);

FILL FILL_4__16391_ (
);

FILL FILL_6__10492_ (
);

FILL FILL_2__11905_ (
);

FILL FILL_3__15384_ (
);

FILL FILL_1__7187_ (
);

FILL FILL_2__14797_ (
);

FILL FILL_2__14377_ (
);

FILL FILL_5__15711_ (
);

FILL FILL_4__14704_ (
);

FILL FILL_3__8894_ (
);

FILL FILL_3__8474_ (
);

INVX1 _12648_ (
    .A(\datapath_1.Data [27]),
    .Y(_3478_)
);

FILL FILL_3__8054_ (
);

NAND3X1 _12228_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [3]),
    .C(_3198__bF$buf4),
    .Y(_3210_)
);

FILL FILL_1__14731_ (
);

FILL FILL_1__14311_ (
);

FILL FILL_6__11697_ (
);

FILL FILL_6__11277_ (
);

FILL FILL_0__13724_ (
);

FILL FILL_0__13304_ (
);

FILL FILL_3__16169_ (
);

FILL FILL_2__6891_ (
);

FILL FILL_5__9761_ (
);

FILL SFILL23400x26050 (
);

FILL FILL_5__9341_ (
);

FILL FILL_0_BUFX2_insert1050 (
);

FILL FILL_0_BUFX2_insert1051 (
);

FILL FILL_0_BUFX2_insert1052 (
);

FILL FILL_0__16196_ (
);

FILL FILL_0_BUFX2_insert1053 (
);

FILL FILL_0_BUFX2_insert1054 (
);

AOI22X1 _16061_ (
    .A(_5565__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [25]),
    .C(\datapath_1.regfile_1.regOut[5] [25]),
    .D(_5700_),
    .Y(_6516_)
);

FILL FILL_0_BUFX2_insert1055 (
);

FILL FILL_0_BUFX2_insert1056 (
);

FILL FILL_2__10297_ (
);

FILL FILL_0_BUFX2_insert1057 (
);

FILL FILL_0_BUFX2_insert1058 (
);

FILL FILL_1__9753_ (
);

FILL FILL_0_BUFX2_insert1059 (
);

FILL FILL_5__11631_ (
);

FILL FILL_5__11211_ (
);

FILL FILL_4__15909_ (
);

FILL FILL_3__9679_ (
);

FILL FILL_2__16103_ (
);

FILL FILL_3_BUFX2_insert950 (
);

FILL FILL_3_BUFX2_insert951 (
);

FILL FILL_3__9259_ (
);

FILL FILL_4__10624_ (
);

FILL FILL_3_BUFX2_insert952 (
);

FILL FILL_3_BUFX2_insert953 (
);

FILL FILL_3_BUFX2_insert954 (
);

FILL FILL_3_BUFX2_insert955 (
);

FILL FILL_6__7684_ (
);

FILL FILL_1__15936_ (
);

FILL FILL_3_BUFX2_insert956 (
);

FILL FILL_1__15516_ (
);

FILL SFILL74520x56050 (
);

FILL FILL_3_BUFX2_insert957 (
);

FILL FILL_3_BUFX2_insert958 (
);

FILL FILL_3_BUFX2_insert959 (
);

FILL FILL_1__10651_ (
);

FILL FILL_1__10231_ (
);

FILL FILL_4__13096_ (
);

FILL FILL_0__14929_ (
);

FILL FILL_0__14509_ (
);

FILL FILL_2__7676_ (
);

FILL FILL_3__12089_ (
);

FILL FILL_6__13843_ (
);

FILL FILL_6__13423_ (
);

FILL SFILL74120x42050 (
);

FILL FILL_5__12836_ (
);

FILL FILL_5__12416_ (
);

FILL FILL_3__13870_ (
);

FILL FILL_3__13450_ (
);

FILL FILL_3__13030_ (
);

FILL FILL_4__8963_ (
);

FILL FILL_4__8123_ (
);

FILL FILL_4__11829_ (
);

FILL FILL_2__12863_ (
);

FILL FILL_4__11409_ (
);

FILL FILL_2__12443_ (
);

FILL FILL_2__12023_ (
);

DFFSR _9188_ (
    .Q(\datapath_1.regfile_1.regOut[18] [14]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_1108_[14])
);

FILL SFILL13800x38050 (
);

FILL FILL_1__11856_ (
);

FILL FILL_1__11436_ (
);

FILL FILL_1__11016_ (
);

FILL FILL_3__6960_ (
);

FILL FILL_0__8863_ (
);

FILL FILL_0__8443_ (
);

FILL FILL_0__10429_ (
);

DFFSR _10714_ (
    .Q(\datapath_1.regfile_1.regOut[30] [4]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_1888_[4])
);

FILL FILL_6__9410_ (
);

FILL FILL_0__10009_ (
);

FILL FILL_5__6886_ (
);

FILL FILL_4__15662_ (
);

FILL FILL_4__15242_ (
);

DFFSR _13186_ (
    .Q(\datapath_1.mux_iord.din0 [11]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3685_[11])
);

FILL FILL_2__9402_ (
);

FILL FILL_3__14655_ (
);

FILL FILL_3__14235_ (
);

FILL FILL_1__6878_ (
);

FILL FILL_4__9748_ (
);

FILL FILL_2__13648_ (
);

FILL FILL_2__13228_ (
);

FILL FILL_0__14682_ (
);

FILL FILL_0__14262_ (
);

FILL FILL_0__9648_ (
);

FILL FILL_3__7745_ (
);

FILL FILL_0__9228_ (
);

OAI21X1 _11919_ (
    .A(_2986_),
    .B(IorD_bF$buf3),
    .C(_2987_),
    .Y(_1_[10])
);

FILL FILL_3__7325_ (
);

FILL FILL_4__16027_ (
);

FILL FILL_6__10548_ (
);

FILL FILL_4__11582_ (
);

FILL FILL_4__11162_ (
);

FILL SFILL64120x40050 (
);

FILL FILL_1__16054_ (
);

FILL FILL_3__10995_ (
);

FILL FILL_3__10575_ (
);

FILL FILL_5__8612_ (
);

FILL FILL_3__10155_ (
);

FILL FILL_0__15887_ (
);

OAI22X1 _15752_ (
    .A(_5478__bF$buf2),
    .B(_6214_),
    .C(_5552__bF$buf3),
    .D(_4779_),
    .Y(_6215_)
);

FILL FILL_0__15467_ (
);

FILL FILL_6_BUFX2_insert464 (
);

INVX1 _15332_ (
    .A(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_5806_)
);

FILL FILL_0__15047_ (
);

FILL FILL112360x38050 (
);

FILL FILL_0__10182_ (
);

FILL FILL_6_BUFX2_insert469 (
);

FILL FILL_5__10902_ (
);

FILL FILL_1__8604_ (
);

FILL SFILL68760x69050 (
);

FILL SFILL64040x47050 (
);

FILL FILL_5__13794_ (
);

FILL FILL_5__13374_ (
);

FILL FILL_6__6955_ (
);

NAND2X1 _7674_ (
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_395_)
);

DFFSR _7254_ (
    .Q(\datapath_1.regfile_1.regOut[3] [0]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_133_[0])
);

FILL FILL_4__12787_ (
);

FILL FILL_4__9081_ (
);

FILL FILL_4__12367_ (
);

FILL SFILL54120x83050 (
);

FILL FILL_2__6947_ (
);

FILL FILL_1__12394_ (
);

OAI22X1 _16117_ (
    .A(_5193_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf3),
    .D(_5190_),
    .Y(_6571_)
);

FILL FILL_0__11387_ (
);

OAI21X1 _11672_ (
    .A(_2758_),
    .B(_2752_),
    .C(_2470__bF$buf1),
    .Y(_2774_)
);

INVX1 _11252_ (
    .A(_2142_),
    .Y(_2371_)
);

FILL FILL_1__9809_ (
);

FILL FILL_3__12721_ (
);

FILL FILL_3__12301_ (
);

FILL FILL_4__7814_ (
);

FILL FILL_5__14999_ (
);

FILL SFILL80040x3050 (
);

FILL FILL_5__14579_ (
);

FILL FILL_2__11714_ (
);

FILL FILL_5__14159_ (
);

FILL FILL_3__15193_ (
);

INVX1 _8879_ (
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_1015_)
);

INVX1 _8459_ (
    .A(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_796_)
);

DFFSR _8039_ (
    .Q(\datapath_1.regfile_1.regOut[9] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_523_[17])
);

FILL FILL_1__10707_ (
);

FILL FILL_2__14186_ (
);

FILL FILL_5__15940_ (
);

FILL FILL_5__15520_ (
);

FILL FILL_5__15100_ (
);

FILL FILL_0__7714_ (
);

DFFSR _9820_ (
    .Q(\datapath_1.regfile_1.regOut[23] [6]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_1433_[6])
);

FILL SFILL89240x51050 (
);

FILL FILL_1__13599_ (
);

INVX1 _9400_ (
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_1281_)
);

FILL FILL_4__14933_ (
);

FILL FILL_4__14513_ (
);

INVX1 _12877_ (
    .A(\datapath_1.a [18]),
    .Y(_3590_)
);

INVX1 _12457_ (
    .A(ALUOut[6]),
    .Y(_3371_)
);

AOI22X1 _12037_ (
    .A(\datapath_1.ALUResult [12]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3074_)
);

FILL FILL_3__13926_ (
);

FILL FILL_1__14960_ (
);

FILL FILL_3__13506_ (
);

FILL SFILL18680x71050 (
);

FILL FILL_1__14540_ (
);

FILL FILL_1__14120_ (
);

FILL FILL_5_BUFX2_insert480 (
);

FILL FILL_5_BUFX2_insert481 (
);

FILL FILL_5_BUFX2_insert482 (
);

FILL FILL_0__13953_ (
);

FILL FILL_5_BUFX2_insert483 (
);

FILL FILL_0__13533_ (
);

FILL FILL_3__16398_ (
);

FILL FILL_0__13113_ (
);

FILL FILL_5_BUFX2_insert484 (
);

FILL FILL_5_BUFX2_insert485 (
);

FILL FILL_5__10499_ (
);

FILL FILL_5_BUFX2_insert486 (
);

FILL FILL_5__9990_ (
);

FILL SFILL54040x45050 (
);

FILL FILL_5_BUFX2_insert487 (
);

FILL FILL_5__9150_ (
);

FILL FILL_5_BUFX2_insert488 (
);

FILL FILL_5_BUFX2_insert489 (
);

NAND3X1 _16290_ (
    .A(_6736_),
    .B(_6737_),
    .C(_6738_),
    .Y(_6739_)
);

FILL FILL_5__16305_ (
);

FILL FILL_5__11860_ (
);

FILL FILL_1__9982_ (
);

FILL FILL_5__11440_ (
);

FILL FILL_1__9142_ (
);

FILL FILL_5__11020_ (
);

FILL FILL_4__15718_ (
);

FILL FILL_2__16332_ (
);

FILL FILL_3__9488_ (
);

FILL FILL_4__10433_ (
);

FILL FILL_4__10013_ (
);

FILL FILL_1__15745_ (
);

FILL FILL_1__15325_ (
);

FILL FILL_1__10880_ (
);

FILL FILL_1__10040_ (
);

FILL FILL_0__14738_ (
);

OAI22X1 _14603_ (
    .A(_5089_),
    .B(_3936__bF$buf2),
    .C(_3935__bF$buf3),
    .D(_5090_),
    .Y(_5091_)
);

FILL FILL_0__14318_ (
);

FILL FILL_2__7485_ (
);

FILL FILL_2__7065_ (
);

FILL FILL_5__12645_ (
);

FILL FILL_5__12225_ (
);

NAND2X1 _6945_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_31_)
);

FILL FILL_4__8772_ (
);

FILL FILL_4__8352_ (
);

FILL FILL_4__11638_ (
);

FILL FILL_4__11218_ (
);

FILL FILL_2__12252_ (
);

FILL FILL111880x62050 (
);

FILL FILL_1__11665_ (
);

FILL FILL_1__11245_ (
);

OAI22X1 _15808_ (
    .A(_5485__bF$buf4),
    .B(_6268_),
    .C(_6269_),
    .D(_5549__bF$buf3),
    .Y(_6270_)
);

NAND3X1 _10943_ (
    .A(_2071_),
    .B(_2076_),
    .C(_2072_),
    .Y(_2077_)
);

FILL FILL_0__8252_ (
);

FILL FILL_0__10658_ (
);

NAND2X1 _10523_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1847_)
);

FILL FILL_0__10238_ (
);

NAND2X1 _10103_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .Y(_1692_)
);

FILL SFILL109400x75050 (
);

FILL FILL_4__15891_ (
);

FILL FILL_6__14017_ (
);

FILL FILL_4__15471_ (
);

FILL SFILL44040x43050 (
);

FILL FILL_4__15051_ (
);

FILL FILL_3__14884_ (
);

FILL FILL_2__9631_ (
);

FILL FILL_3__14464_ (
);

FILL FILL_2__9211_ (
);

FILL FILL_3__14044_ (
);

FILL FILL_4__9977_ (
);

FILL FILL112200x3050 (
);

FILL FILL_4__9557_ (
);

FILL FILL_4__9137_ (
);

FILL FILL_2__13877_ (
);

FILL FILL_2__13457_ (
);

FILL FILL_0__14491_ (
);

FILL FILL_2__13037_ (
);

FILL FILL_0__14071_ (
);

FILL SFILL109800x44050 (
);

FILL FILL_3__7974_ (
);

FILL FILL_0__9877_ (
);

FILL FILL_3__7554_ (
);

FILL SFILL79960x3050 (
);

FILL FILL_0__9037_ (
);

OAI21X1 _11728_ (
    .A(_2563_),
    .B(_2375_),
    .C(_2169_),
    .Y(_2825_)
);

OAI21X1 _11308_ (
    .A(_2416_),
    .B(_2424_),
    .C(_2426_),
    .Y(_2427_)
);

FILL FILL_1__13811_ (
);

FILL FILL_4__16256_ (
);

FILL FILL_4__11391_ (
);

FILL FILL_3__15669_ (
);

FILL FILL_3__15249_ (
);

FILL FILL_1__16283_ (
);

FILL FILL_5__8841_ (
);

FILL FILL_3__10384_ (
);

FILL FILL_5__8001_ (
);

OAI22X1 _15981_ (
    .A(_5052_),
    .B(_5548__bF$buf3),
    .C(_5504__bF$buf1),
    .D(_5081_),
    .Y(_6438_)
);

FILL FILL_0__15696_ (
);

INVX1 _15561_ (
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_6029_)
);

FILL FILL_0__15276_ (
);

OAI22X1 _15141_ (
    .A(_5618_),
    .B(_5548__bF$buf4),
    .C(_5504__bF$buf0),
    .D(_4055_),
    .Y(_5619_)
);

FILL FILL_1__8833_ (
);

FILL SFILL69560x68050 (
);

FILL FILL_2__15603_ (
);

FILL FILL_3__8759_ (
);

FILL FILL_3__8339_ (
);

INVX1 _7483_ (
    .A(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_308_)
);

INVX1 _7063_ (
    .A(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_89_)
);

FILL FILL_4__12596_ (
);

FILL FILL_4__12176_ (
);

FILL SFILL69160x54050 (
);

FILL FILL_5__9626_ (
);

FILL FILL_3__11589_ (
);

FILL FILL_5__9206_ (
);

FILL FILL_3__11169_ (
);

FILL SFILL74120x37050 (
);

NAND2X1 _16346_ (
    .A(gnd),
    .B(gnd),
    .Y(_6785_)
);

FILL FILL_0__11196_ (
);

NAND3X1 _11481_ (
    .A(_2462__bF$buf2),
    .B(_2594_),
    .C(_2575_),
    .Y(_2595_)
);

FILL FILL_5__11916_ (
);

OAI21X1 _11061_ (
    .A(_2178_),
    .B(_2179_),
    .C(_2177_),
    .Y(_2180_)
);

FILL FILL_1__9618_ (
);

FILL FILL_3__12530_ (
);

FILL FILL_3__12110_ (
);

FILL FILL_4__7623_ (
);

FILL FILL_4__7203_ (
);

FILL FILL_4__10909_ (
);

FILL FILL_2__11943_ (
);

FILL FILL_5__14388_ (
);

FILL FILL_2__11523_ (
);

FILL FILL_2__11103_ (
);

DFFSR _8688_ (
    .Q(\datapath_1.regfile_1.regOut[14] [26]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_848_[26])
);

OAI21X1 _8268_ (
    .A(_708_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .C(_709_),
    .Y(_653_[28])
);

FILL FILL_1__10936_ (
);

FILL FILL_1__10516_ (
);

FILL FILL_0__7943_ (
);

FILL FILL_0__7103_ (
);

FILL FILL_4__14742_ (
);

FILL FILL_4__14322_ (
);

FILL FILL_3__8092_ (
);

DFFSR _12686_ (
    .Q(\datapath_1.Data [23]),
    .CLK(clk_bF$buf43),
    .R(rst_bF$buf37),
    .S(vdd),
    .D(_3425_[23])
);

NAND3X1 _12266_ (
    .A(_3236_),
    .B(_3237_),
    .C(_3238_),
    .Y(\datapath_1.alu_1.ALUInB [12])
);

FILL FILL_2__8902_ (
);

FILL FILL_3__13735_ (
);

FILL FILL_3__13315_ (
);

FILL FILL_4__8828_ (
);

FILL FILL_2__12728_ (
);

FILL FILL_0__13762_ (
);

FILL FILL_2__12308_ (
);

FILL SFILL99320x41050 (
);

FILL FILL_0__13342_ (
);

FILL FILL_0__8728_ (
);

FILL FILL_5__16114_ (
);

FILL SFILL59160x52050 (
);

FILL FILL_1__9791_ (
);

FILL FILL_1__9371_ (
);

FILL FILL_4__15947_ (
);

FILL FILL_4__15527_ (
);

FILL FILL_4__15107_ (
);

FILL FILL_2__16141_ (
);

FILL FILL_3__9297_ (
);

FILL FILL_4__10662_ (
);

FILL FILL_4__10242_ (
);

FILL SFILL64120x35050 (
);

FILL FILL_1__15974_ (
);

FILL SFILL84920x9050 (
);

FILL FILL_1__15554_ (
);

FILL FILL_1__15134_ (
);

FILL FILL_0__14967_ (
);

NAND3X1 _14832_ (
    .A(_5307_),
    .B(_5308_),
    .C(_5315_),
    .Y(_5316_)
);

FILL FILL_0__14547_ (
);

FILL FILL_0__14127_ (
);

NAND3X1 _14412_ (
    .A(_4895_),
    .B(_4896_),
    .C(_4903_),
    .Y(_4904_)
);

FILL SFILL28680x68050 (
);

FILL FILL_2__7294_ (
);

FILL FILL_5__12874_ (
);

FILL FILL_5__12454_ (
);

FILL FILL_5__12034_ (
);

FILL SFILL84200x2050 (
);

FILL FILL_4__8581_ (
);

FILL FILL_4__11867_ (
);

FILL FILL_4__11447_ (
);

FILL SFILL89720x53050 (
);

FILL FILL_2__12481_ (
);

FILL FILL_4__11027_ (
);

FILL FILL_2__12061_ (
);

FILL FILL_1__16339_ (
);

FILL FILL_6__8087_ (
);

FILL FILL_1__11894_ (
);

FILL SFILL9320x57050 (
);

FILL FILL_1__11474_ (
);

FILL FILL_1__11054_ (
);

AOI22X1 _15617_ (
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .B(_5577_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_6083_)
);

FILL FILL_0__8481_ (
);

FILL FILL_0__10887_ (
);

FILL FILL_2__8499_ (
);

FILL FILL_2__8079_ (
);

NAND2X1 _10752_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_1959_)
);

FILL FILL_0__8061_ (
);

DFFSR _10332_ (
    .Q(\datapath_1.regfile_1.regOut[27] [6]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_1693_[6])
);

FILL FILL_0__10047_ (
);

FILL FILL_3__11801_ (
);

FILL FILL_4__15280_ (
);

FILL FILL_2__9860_ (
);

FILL FILL_5__13659_ (
);

FILL SFILL113800x44050 (
);

FILL FILL_5__13239_ (
);

FILL FILL_3__14693_ (
);

FILL FILL_2__9020_ (
);

INVX1 _7959_ (
    .A(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_544_)
);

FILL FILL_3__14273_ (
);

DFFSR _7539_ (
    .Q(\datapath_1.regfile_1.regOut[5] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_263_[29])
);

OAI21X1 _7119_ (
    .A(_125_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_126_),
    .Y(_68_[29])
);

FILL SFILL49160x50050 (
);

FILL FILL_4__9786_ (
);

FILL FILL_4__9366_ (
);

FILL FILL_2__13686_ (
);

FILL FILL_2__13266_ (
);

FILL FILL_5__14600_ (
);

FILL SFILL89240x46050 (
);

INVX1 _8900_ (
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_1029_)
);

FILL SFILL54120x33050 (
);

FILL FILL_1__12259_ (
);

NAND2X1 _11957_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[23]),
    .Y(_3013_)
);

FILL FILL_0__9266_ (
);

FILL FILL_3__7363_ (
);

OAI21X1 _11537_ (
    .A(_2647_),
    .B(_2427_),
    .C(_2414_),
    .Y(_2648_)
);

NOR2X1 _11117_ (
    .A(_2235_),
    .B(_2234_),
    .Y(_2236_)
);

FILL SFILL79320x82050 (
);

FILL FILL_1__13620_ (
);

FILL FILL_5__7289_ (
);

FILL FILL_4__16065_ (
);

FILL FILL_3__15898_ (
);

FILL FILL_0__12613_ (
);

FILL FILL_3__15478_ (
);

FILL FILL_3__15058_ (
);

FILL FILL_1__16092_ (
);

FILL FILL_5__8650_ (
);

FILL FILL_5__8230_ (
);

FILL FILL_3__10193_ (
);

FILL FILL_6_BUFX2_insert843 (
);

OAI21X1 _15790_ (
    .A(_5524__bF$buf0),
    .B(_4820_),
    .C(_6251_),
    .Y(_6252_)
);

NOR2X1 _15370_ (
    .A(_5841_),
    .B(_5842_),
    .Y(_5843_)
);

FILL FILL_0__15085_ (
);

FILL FILL_5__15805_ (
);

FILL FILL_6_BUFX2_insert848 (
);

FILL FILL_5__10940_ (
);

FILL FILL_5__10520_ (
);

FILL FILL_1__8642_ (
);

FILL FILL_1__8222_ (
);

FILL FILL_2__15832_ (
);

FILL FILL_2__15412_ (
);

FILL FILL_3__8988_ (
);

FILL FILL_3__8568_ (
);

FILL FILL_3__8148_ (
);

FILL FILL_1__14825_ (
);

FILL FILL_1__14405_ (
);

INVX1 _7292_ (
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_201_)
);

FILL SFILL18680x21050 (
);

FILL FILL_0__13818_ (
);

FILL FILL_2__6985_ (
);

FILL FILL_5__9855_ (
);

FILL FILL_3__11398_ (
);

FILL FILL_5__9015_ (
);

OAI22X1 _16155_ (
    .A(_5527__bF$buf3),
    .B(_5236_),
    .C(_5243_),
    .D(_5532__bF$buf2),
    .Y(_6608_)
);

INVX1 _11290_ (
    .A(_2217_),
    .Y(_2409_)
);

FILL FILL_1__9847_ (
);

FILL FILL_5__11725_ (
);

FILL FILL_1__9427_ (
);

FILL FILL_5__11305_ (
);

FILL FILL_1__9007_ (
);

FILL SFILL79240x44050 (
);

FILL FILL_4__7852_ (
);

FILL FILL_4__7432_ (
);

FILL FILL_2__11752_ (
);

FILL FILL_5__14197_ (
);

FILL FILL_2__11332_ (
);

FILL FILL_6__7358_ (
);

OAI21X1 _8497_ (
    .A(_820_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .C(_821_),
    .Y(_783_[19])
);

OAI21X1 _8077_ (
    .A(_601_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .C(_602_),
    .Y(_588_[7])
);

FILL FILL_1__10745_ (
);

FILL FILL_1__10325_ (
);

FILL FILL_0__7752_ (
);

FILL FILL_0__7332_ (
);

FILL FILL_4__14971_ (
);

FILL SFILL44040x38050 (
);

FILL SFILL54120x6050 (
);

FILL FILL_4__14551_ (
);

FILL FILL_4__14131_ (
);

FILL SFILL94360x4050 (
);

OAI21X1 _12495_ (
    .A(_3395_),
    .B(vdd),
    .C(_3396_),
    .Y(_3360_[18])
);

NAND3X1 _12075_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[22]),
    .C(_3032__bF$buf4),
    .Y(_3102_)
);

FILL FILL_3__13964_ (
);

FILL FILL_2__8711_ (
);

FILL SFILL94280x9050 (
);

FILL FILL_3__13544_ (
);

FILL FILL_3__13124_ (
);

FILL FILL_4__8637_ (
);

FILL FILL_5_BUFX2_insert860 (
);

FILL FILL_4__8217_ (
);

FILL FILL_2__12957_ (
);

FILL FILL_5_BUFX2_insert861 (
);

FILL FILL_5_BUFX2_insert862 (
);

FILL FILL_0__13991_ (
);

FILL FILL_5_BUFX2_insert863 (
);

FILL FILL_2__12117_ (
);

FILL FILL_0__13571_ (
);

FILL FILL_0__13151_ (
);

FILL FILL_5_BUFX2_insert864 (
);

FILL FILL_5_BUFX2_insert865 (
);

FILL FILL_5_BUFX2_insert866 (
);

FILL FILL_5_BUFX2_insert867 (
);

FILL FILL_5_BUFX2_insert868 (
);

FILL FILL_5_BUFX2_insert869 (
);

FILL FILL111880x12050 (
);

FILL FILL_5__16343_ (
);

FILL FILL_0__8957_ (
);

FILL FILL_0__8117_ (
);

INVX1 _10808_ (
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_1996_)
);

FILL SFILL104520x7050 (
);

FILL FILL_4__15756_ (
);

FILL FILL_4__15336_ (
);

FILL FILL_2__16370_ (
);

FILL FILL_4__10891_ (
);

FILL FILL_2__9916_ (
);

FILL FILL_4__10051_ (
);

FILL FILL_3__14749_ (
);

FILL FILL_1__15783_ (
);

FILL FILL_3__14329_ (
);

FILL FILL_1__15363_ (
);

FILL FILL_5__7501_ (
);

FILL FILL_0__14776_ (
);

FILL SFILL69240x42050 (
);

INVX1 _14641_ (
    .A(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_5129_)
);

FILL FILL_0__14356_ (
);

INVX1 _14221_ (
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_4717_)
);

FILL FILL_6__13270_ (
);

FILL FILL_3__7839_ (
);

FILL FILL_3__7419_ (
);

FILL FILL_5__12263_ (
);

INVX1 _6983_ (
    .A(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_56_)
);

FILL FILL_2_BUFX2_insert990 (
);

FILL FILL_2_BUFX2_insert991 (
);

FILL FILL_2_BUFX2_insert992 (
);

FILL FILL_2_BUFX2_insert993 (
);

FILL FILL_4__8390_ (
);

FILL SFILL38760x58050 (
);

FILL FILL_2_BUFX2_insert994 (
);

FILL FILL_4__11676_ (
);

FILL SFILL69160x49050 (
);

FILL FILL_2_BUFX2_insert995 (
);

FILL FILL_4__11256_ (
);

FILL FILL_2_BUFX2_insert996 (
);

FILL FILL_2__12290_ (
);

FILL FILL_2_BUFX2_insert997 (
);

FILL FILL_2_BUFX2_insert998 (
);

FILL FILL_2_BUFX2_insert999 (
);

FILL FILL_1__16148_ (
);

FILL FILL_5__8706_ (
);

FILL FILL_3__10669_ (
);

FILL FILL_3__10249_ (
);

FILL FILL_1__11283_ (
);

INVX1 _15846_ (
    .A(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_6307_)
);

NAND3X1 _15426_ (
    .A(_5886_),
    .B(_5896_),
    .C(_5892_),
    .Y(_5897_)
);

INVX4 _15006_ (
    .A(_5485__bF$buf1),
    .Y(_5486_)
);

INVX1 _10981_ (
    .A(\control_1.reg_state.dout [3]),
    .Y(_2105_)
);

FILL FILL_0__10696_ (
);

FILL FILL_0__10276_ (
);

INVX1 _10561_ (
    .A(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_1872_)
);

INVX1 _10141_ (
    .A(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_1653_)
);

FILL FILL_3__11610_ (
);

FILL FILL_5__13888_ (
);

FILL FILL_5__13468_ (
);

FILL FILL_3__14082_ (
);

DFFSR _7768_ (
    .Q(\datapath_1.regfile_1.regOut[7] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_393_[2])
);

OAI21X1 _7348_ (
    .A(_237_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .C(_238_),
    .Y(_198_[20])
);

FILL FILL_4__9595_ (
);

FILL SFILL59640x54050 (
);

FILL FILL_2__13495_ (
);

FILL FILL_1__12488_ (
);

FILL FILL_1__12068_ (
);

FILL FILL_4__13822_ (
);

FILL FILL_4__13402_ (
);

FILL FILL_3__7592_ (
);

FILL FILL_0__9495_ (
);

FILL FILL_3__7172_ (
);

INVX1 _11766_ (
    .A(_2138_),
    .Y(_2861_)
);

AOI21X1 _11346_ (
    .A(_2116_),
    .B(_2461_),
    .C(_2463_),
    .Y(_2464_)
);

FILL FILL_5__7098_ (
);

FILL FILL_4__16294_ (
);

FILL FILL_2__11808_ (
);

FILL FILL_0__12842_ (
);

FILL FILL_0__12422_ (
);

FILL FILL_3__15287_ (
);

FILL FILL_0__12002_ (
);

FILL SFILL23800x8050 (
);

FILL FILL_6__16201_ (
);

FILL SFILL89400x72050 (
);

FILL FILL_5__15614_ (
);

FILL FILL_0__7808_ (
);

FILL SFILL59160x47050 (
);

OAI21X1 _9914_ (
    .A(_1541_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1542_),
    .Y(_1498_[22])
);

FILL FILL_1__8871_ (
);

FILL FILL_1__8451_ (
);

FILL SFILL3720x4050 (
);

FILL FILL_4__14607_ (
);

FILL FILL_2__15641_ (
);

FILL FILL_2__15221_ (
);

FILL FILL_3__8377_ (
);

FILL SFILL3640x9050 (
);

FILL FILL_1__14634_ (
);

FILL FILL_1__14214_ (
);

FILL FILL_0__13627_ (
);

INVX1 _13912_ (
    .A(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_4415_)
);

FILL FILL_0__13207_ (
);

FILL FILL_5__9664_ (
);

FILL FILL_5__9244_ (
);

INVX1 _16384_ (
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .Y(_6810_)
);

FILL FILL_6__12121_ (
);

FILL FILL_0__16099_ (
);

FILL FILL_5__11954_ (
);

FILL FILL_1__9656_ (
);

FILL FILL_5__11534_ (
);

FILL SFILL114360x3050 (
);

FILL FILL_5__11114_ (
);

FILL FILL_1__9236_ (
);

FILL SFILL28760x11050 (
);

FILL FILL_2__16006_ (
);

FILL FILL_4__10947_ (
);

FILL FILL_4__7241_ (
);

FILL FILL_2__11981_ (
);

FILL FILL_4__10527_ (
);

FILL FILL_2__11561_ (
);

FILL FILL_4__10107_ (
);

FILL FILL_2__11141_ (
);

FILL FILL_1__15839_ (
);

FILL FILL_6__7167_ (
);

FILL FILL_1__15419_ (
);

FILL FILL_1__10974_ (
);

FILL FILL_1__10554_ (
);

FILL FILL_1__10134_ (
);

FILL SFILL33960x74050 (
);

FILL FILL_2__7999_ (
);

FILL FILL_0__7981_ (
);

FILL FILL_0__7561_ (
);

BUFX2 BUFX2_insert680 (
    .A(_5485_),
    .Y(_5485__bF$buf3)
);

FILL FILL_2__7579_ (
);

FILL FILL_2__7159_ (
);

BUFX2 BUFX2_insert681 (
    .A(_5485_),
    .Y(_5485__bF$buf2)
);

FILL SFILL89320x34050 (
);

BUFX2 BUFX2_insert682 (
    .A(_5485_),
    .Y(_5485__bF$buf1)
);

BUFX2 BUFX2_insert683 (
    .A(_5485_),
    .Y(_5485__bF$buf0)
);

FILL FILL_6__13746_ (
);

BUFX2 BUFX2_insert684 (
    .A(_3971_),
    .Y(_3971__bF$buf4)
);

FILL FILL_6__13326_ (
);

BUFX2 BUFX2_insert685 (
    .A(_3971_),
    .Y(_3971__bF$buf3)
);

FILL FILL_4__14780_ (
);

BUFX2 BUFX2_insert686 (
    .A(_3971_),
    .Y(_3971__bF$buf2)
);

FILL FILL_4__14360_ (
);

BUFX2 BUFX2_insert687 (
    .A(_3971_),
    .Y(_3971__bF$buf1)
);

BUFX2 BUFX2_insert688 (
    .A(_3971_),
    .Y(_3971__bF$buf0)
);

BUFX2 BUFX2_insert689 (
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf7 )
);

FILL FILL_5__12739_ (
);

FILL FILL_3__13773_ (
);

FILL FILL_2__8520_ (
);

FILL FILL_5__12319_ (
);

FILL FILL_2__8100_ (
);

FILL FILL_3__13353_ (
);

FILL SFILL18760x54050 (
);

FILL SFILL33560x60050 (
);

FILL FILL_4__8866_ (
);

FILL FILL_4__8446_ (
);

FILL FILL_2__12766_ (
);

FILL FILL_2__12346_ (
);

FILL FILL_0__13380_ (
);

FILL SFILL94440x50 (
);

FILL FILL_1__11759_ (
);

FILL FILL_1__11339_ (
);

FILL FILL_0__8766_ (
);

FILL FILL_3__6863_ (
);

FILL FILL_5__16152_ (
);

FILL FILL_0__8346_ (
);

INVX1 _10617_ (
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_1889_)
);

FILL FILL_4__15985_ (
);

FILL FILL_1__12700_ (
);

FILL FILL_4__15565_ (
);

FILL FILL_4__15145_ (
);

NAND2X1 _13089_ (
    .A(PCEn_bF$buf6),
    .B(\datapath_1.mux_pcsrc.dout [3]),
    .Y(_3691_)
);

FILL FILL_4__10280_ (
);

FILL FILL_3__14978_ (
);

FILL FILL_2__9725_ (
);

FILL FILL_3__14558_ (
);

FILL FILL_3__14138_ (
);

FILL FILL_1__15592_ (
);

FILL FILL_1__15172_ (
);

FILL FILL_5__7730_ (
);

FILL FILL_5__7310_ (
);

INVX1 _14870_ (
    .A(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_5353_)
);

FILL FILL_0__14585_ (
);

FILL FILL_0__14165_ (
);

AOI21X1 _14450_ (
    .A(_4941_),
    .B(_4915_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [20])
);

OAI22X1 _14030_ (
    .A(_3982__bF$buf2),
    .B(_4529_),
    .C(_3966__bF$buf2),
    .D(_4528_),
    .Y(_4530_)
);

FILL FILL_1__7722_ (
);

FILL FILL_1__7302_ (
);

FILL FILL_2__14912_ (
);

FILL FILL_3__7228_ (
);

FILL FILL_5__12492_ (
);

FILL FILL_5__12072_ (
);

FILL FILL_1__13905_ (
);

FILL SFILL79320x32050 (
);

FILL SFILL18680x16050 (
);

FILL SFILL59000x3050 (
);

FILL FILL_4__11485_ (
);

FILL FILL_4__11065_ (
);

FILL FILL_1__16377_ (
);

FILL FILL_3__10898_ (
);

FILL FILL_5__8515_ (
);

FILL FILL_3__10058_ (
);

FILL FILL_1__11092_ (
);

INVX1 _15655_ (
    .A(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_6120_)
);

INVX1 _15235_ (
    .A(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_5711_)
);

INVX1 _10790_ (
    .A(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_1984_)
);

INVX1 _10370_ (
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_1765_)
);

FILL FILL_5__10805_ (
);

FILL FILL_1__8507_ (
);

FILL FILL_4__6932_ (
);

FILL FILL_0__16311_ (
);

FILL FILL_2__10832_ (
);

FILL FILL_5__13697_ (
);

FILL FILL_5__13277_ (
);

FILL FILL_2__10412_ (
);

OAI21X1 _7997_ (
    .A(_568_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_569_),
    .Y(_523_[23])
);

FILL FILL_6__6858_ (
);

OAI21X1 _7577_ (
    .A(_349_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .C(_350_),
    .Y(_328_[11])
);

DFFSR _7157_ (
    .Q(\datapath_1.regfile_1.regOut[2] [31]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf91),
    .S(vdd),
    .D(_68_[31])
);

FILL FILL_1__12297_ (
);

FILL FILL_4__13631_ (
);

FILL FILL_4__13211_ (
);

NAND3X1 _11995_ (
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[2]),
    .C(_3032__bF$buf2),
    .Y(_3042_)
);

AOI21X1 _11575_ (
    .A(_2669_),
    .B(_2620_),
    .C(_2682_),
    .Y(_2683_)
);

AOI21X1 _11155_ (
    .A(_2272_),
    .B(_2248_),
    .C(_2273_),
    .Y(_2274_)
);

FILL FILL_3__12624_ (
);

FILL FILL_3__12204_ (
);

FILL FILL_4__7717_ (
);

FILL FILL_2__11617_ (
);

FILL FILL_0__12651_ (
);

FILL FILL_0__12231_ (
);

FILL FILL_3__15096_ (
);

FILL FILL_2__14089_ (
);

FILL FILL_5__15843_ (
);

FILL FILL_5__15423_ (
);

FILL FILL_5__15003_ (
);

FILL FILL_0__7617_ (
);

OAI21X1 _9723_ (
    .A(_1434_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1435_),
    .Y(_1433_[1])
);

DFFSR _9303_ (
    .Q(\datapath_1.regfile_1.regOut[19] [1]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_1173_[1])
);

FILL FILL_1__8260_ (
);

FILL FILL_4__14836_ (
);

FILL FILL_2__15870_ (
);

FILL FILL_4__14416_ (
);

FILL FILL_2__15450_ (
);

FILL FILL_2__15030_ (
);

FILL FILL_3__8186_ (
);

FILL FILL_3__13829_ (
);

FILL FILL_1__14863_ (
);

FILL FILL_3__13409_ (
);

FILL FILL_1__14443_ (
);

FILL FILL_1__14023_ (
);

FILL SFILL69240x37050 (
);

FILL FILL_0__13856_ (
);

FILL FILL_0__13436_ (
);

INVX1 _13721_ (
    .A(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_4228_)
);

NOR2X1 _13301_ (
    .A(_3781_),
    .B(_3836_),
    .Y(\datapath_1.regfile_1.regEn [8])
);

FILL FILL_0__13016_ (
);

FILL FILL_5__9893_ (
);

FILL FILL_5__9473_ (
);

NAND3X1 _16193_ (
    .A(\datapath_1.regfile_1.regOut[24] [28]),
    .B(_5465_),
    .C(_5531__bF$buf4),
    .Y(_6645_)
);

FILL FILL_5__16208_ (
);

FILL FILL_3__6919_ (
);

FILL FILL_5__11763_ (
);

FILL FILL_1__9885_ (
);

FILL FILL_1__9465_ (
);

FILL FILL_5__11343_ (
);

FILL FILL_1__9045_ (
);

FILL SFILL99400x69050 (
);

FILL FILL_2__16235_ (
);

FILL FILL_4__7890_ (
);

FILL FILL_4__7470_ (
);

FILL FILL_4__7050_ (
);

FILL FILL_4__10756_ (
);

FILL FILL_2__11790_ (
);

FILL FILL_2__11370_ (
);

FILL FILL_1__15648_ (
);

FILL FILL_1__15228_ (
);

FILL FILL_1__10783_ (
);

FILL FILL_1__10363_ (
);

AOI22X1 _14926_ (
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .B(_4005__bF$buf2),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_5408_)
);

OAI22X1 _14506_ (
    .A(_3884__bF$buf2),
    .B(_4994_),
    .C(_3955__bF$buf4),
    .D(_4995_),
    .Y(_4996_)
);

FILL FILL_0__7370_ (
);

FILL SFILL69160x5050 (
);

FILL FILL_5__12968_ (
);

FILL FILL_5__12128_ (
);

FILL FILL_3__13582_ (
);

BUFX2 _6848_ (
    .A(_1_[10]),
    .Y(memoryAddress[10])
);

FILL FILL_3__13162_ (
);

FILL FILL_4__8255_ (
);

FILL SFILL8600x1050 (
);

FILL FILL_2__12995_ (
);

FILL FILL_2__12575_ (
);

FILL FILL_2__12155_ (
);

FILL SFILL99400x24050 (
);

FILL FILL_1__11988_ (
);

FILL FILL_1__11568_ (
);

FILL FILL_1__11148_ (
);

FILL FILL_4__12902_ (
);

FILL FILL_0__8995_ (
);

FILL FILL_5__16381_ (
);

FILL FILL_0__8575_ (
);

DFFSR _10846_ (
    .Q(\datapath_1.regfile_1.regOut[31] [8]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf72),
    .S(vdd),
    .D(_1953_[8])
);

OAI21X1 _10426_ (
    .A(_1801_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .C(_1802_),
    .Y(_1758_[22])
);

OAI21X1 _10006_ (
    .A(_1582_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .C(_1583_),
    .Y(_1563_[10])
);

FILL FILL_4__15794_ (
);

FILL FILL_4__15374_ (
);

FILL FILL_2__9534_ (
);

FILL FILL_0__11922_ (
);

FILL FILL_3__14787_ (
);

FILL FILL_2__9114_ (
);

FILL FILL_3__14367_ (
);

FILL FILL_0__11502_ (
);

FILL FILL_0__14394_ (
);

FILL SFILL89400x67050 (
);

FILL FILL_1__7951_ (
);

FILL FILL_1__7111_ (
);

FILL FILL_2__14721_ (
);

FILL FILL_3__7877_ (
);

FILL FILL_2__14301_ (
);

FILL FILL_3__7457_ (
);

FILL FILL_3__7037_ (
);

FILL FILL_1__13714_ (
);

FILL FILL_4__16159_ (
);

FILL FILL_4__11294_ (
);

FILL FILL_0__12707_ (
);

FILL FILL_1__16186_ (
);

FILL FILL_5__8744_ (
);

FILL FILL_5__8324_ (
);

FILL FILL_3__10287_ (
);

OAI22X1 _15884_ (
    .A(_5534__bF$buf1),
    .B(_4919_),
    .C(_6343_),
    .D(_5549__bF$buf0),
    .Y(_6344_)
);

FILL FILL_0__15599_ (
);

FILL FILL_0__15179_ (
);

OAI22X1 _15464_ (
    .A(_5472__bF$buf0),
    .B(_4437_),
    .C(_4470_),
    .D(_5552__bF$buf1),
    .Y(_5934_)
);

NAND3X1 _15044_ (
    .A(_5459__bF$buf3),
    .B(_5461_),
    .C(_5471__bF$buf5),
    .Y(_5524_)
);

FILL SFILL89400x22050 (
);

FILL FILL_1__8736_ (
);

FILL FILL_5__10614_ (
);

FILL FILL_1__8316_ (
);

FILL SFILL94280x73050 (
);

FILL FILL_2__15926_ (
);

FILL FILL_2__15506_ (
);

FILL FILL_0__16120_ (
);

FILL FILL_2__10641_ (
);

FILL FILL_5__13086_ (
);

FILL FILL_1__14919_ (
);

DFFSR _7386_ (
    .Q(\datapath_1.regfile_1.regOut[4] [4]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_198_[4])
);

FILL FILL_4__12499_ (
);

FILL FILL_4__12079_ (
);

FILL FILL_3__9603_ (
);

FILL SFILL33960x69050 (
);

FILL FILL_5__9529_ (
);

FILL FILL_5__9109_ (
);

FILL FILL_6__12826_ (
);

FILL FILL_4__13860_ (
);

FILL FILL_4__13440_ (
);

NOR2X1 _16249_ (
    .A(_6698_),
    .B(_6697_),
    .Y(_6699_)
);

FILL FILL_4__13020_ (
);

OAI21X1 _11384_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2157_),
    .C(_2500_),
    .Y(_2501_)
);

FILL FILL_0__11099_ (
);

FILL FILL_5__11819_ (
);

FILL FILL_2__7600_ (
);

FILL FILL_3__12853_ (
);

FILL SFILL18760x49050 (
);

FILL FILL_3__12433_ (
);

FILL SFILL33560x55050 (
);

FILL FILL_3__12013_ (
);

FILL FILL_4__7946_ (
);

FILL FILL_4__7106_ (
);

FILL FILL_2__11846_ (
);

FILL FILL_0__12880_ (
);

FILL FILL_2__11426_ (
);

FILL FILL_0__12460_ (
);

FILL FILL_2__11006_ (
);

FILL FILL_0__12040_ (
);

FILL FILL_1__10419_ (
);

FILL FILL_5__15652_ (
);

FILL FILL_0__7846_ (
);

FILL FILL_5__15232_ (
);

FILL FILL_0__7426_ (
);

DFFSR _9952_ (
    .Q(\datapath_1.regfile_1.regOut[24] [10]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_1498_[10])
);

NAND2X1 _9532_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1349_)
);

NAND2X1 _9112_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1130_)
);

FILL SFILL33960x24050 (
);

FILL FILL_4__14645_ (
);

FILL FILL_4__14225_ (
);

NAND2X1 _12589_ (
    .A(vdd),
    .B(memoryOutData[7]),
    .Y(_3439_)
);

INVX1 _12169_ (
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3166_)
);

FILL FILL_3__13638_ (
);

FILL FILL_3__13218_ (
);

FILL FILL_1__14672_ (
);

FILL FILL_1__14252_ (
);

FILL FILL_0_BUFX2_insert320 (
);

FILL SFILL79400x20050 (
);

FILL FILL_0_BUFX2_insert321 (
);

FILL FILL_0_BUFX2_insert322 (
);

FILL FILL_0_BUFX2_insert323 (
);

FILL FILL_0__13665_ (
);

FILL FILL_0_BUFX2_insert324 (
);

AOI22X1 _13950_ (
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .B(_4246_),
    .C(_4129_),
    .D(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_4452_)
);

FILL FILL_0__13245_ (
);

FILL FILL_0_BUFX2_insert325 (
);

AOI22X1 _13530_ (
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .B(_3885_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_4041_)
);

FILL FILL_0_BUFX2_insert326 (
);

NAND2X1 _13110_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_pcsrc.dout [10]),
    .Y(_3705_)
);

FILL FILL_0_BUFX2_insert327 (
);

FILL FILL_0_BUFX2_insert328 (
);

FILL FILL_0_BUFX2_insert329 (
);

FILL FILL_5__9282_ (
);

FILL FILL_5__16017_ (
);

FILL FILL_5__11992_ (
);

FILL FILL_5__11572_ (
);

FILL FILL_1__9274_ (
);

FILL FILL_5__11152_ (
);

FILL SFILL79320x27050 (
);

FILL FILL_2__16044_ (
);

FILL FILL_4__10565_ (
);

FILL FILL_4__10145_ (
);

FILL FILL_1__15877_ (
);

FILL FILL_1__15457_ (
);

FILL FILL_1__15037_ (
);

FILL FILL_1__10172_ (
);

INVX1 _14735_ (
    .A(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_5221_)
);

INVX1 _14315_ (
    .A(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_4809_)
);

FILL FILL_2__7197_ (
);

FILL FILL_0__15811_ (
);

FILL FILL_5__12777_ (
);

FILL FILL_5__12357_ (
);

FILL FILL_3__13391_ (
);

FILL FILL_4__8484_ (
);

FILL FILL_4__8064_ (
);

FILL FILL_2__12384_ (
);

FILL SFILL114440x52050 (
);

FILL FILL_1__11797_ (
);

FILL FILL_1__11377_ (
);

FILL FILL_4__12711_ (
);

FILL FILL_5__16190_ (
);

FILL FILL_0__8384_ (
);

OAI21X1 _10655_ (
    .A(_1913_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1914_),
    .Y(_1888_[13])
);

OAI21X1 _10235_ (
    .A(_1694_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .C(_1695_),
    .Y(_1693_[1])
);

FILL FILL_6__14989_ (
);

FILL FILL_6__14569_ (
);

FILL FILL_3__11704_ (
);

FILL FILL_4__15183_ (
);

FILL FILL_2__9763_ (
);

FILL FILL_2__9343_ (
);

FILL FILL_3__14596_ (
);

FILL FILL_0__11731_ (
);

FILL FILL_3__14176_ (
);

FILL FILL_0__11311_ (
);

FILL FILL_6__15930_ (
);

FILL FILL_4__9269_ (
);

FILL FILL_2__13589_ (
);

FILL FILL_2__13169_ (
);

FILL FILL_5__14923_ (
);

FILL FILL_5__14503_ (
);

DFFSR _8803_ (
    .Q(\datapath_1.regfile_1.regOut[15] [13]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_913_[13])
);

FILL FILL_1__7760_ (
);

FILL FILL_1__7340_ (
);

FILL FILL_4__13916_ (
);

FILL FILL_2__14950_ (
);

FILL FILL_2__14530_ (
);

FILL FILL_3__7686_ (
);

FILL FILL_2__14110_ (
);

FILL FILL_0__9169_ (
);

FILL FILL_3__12909_ (
);

FILL FILL_1__13943_ (
);

FILL FILL_4__16388_ (
);

FILL FILL_1__13523_ (
);

FILL FILL_1__13103_ (
);

DFFSR _12801_ (
    .Q(\datapath_1.PCJump [12]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf99),
    .S(vdd),
    .D(_3490_[10])
);

FILL FILL_0__12516_ (
);

FILL FILL_5__8973_ (
);

FILL FILL_5__8133_ (
);

FILL FILL_6__11850_ (
);

OAI22X1 _15693_ (
    .A(_5549__bF$buf4),
    .B(_4732_),
    .C(_5532__bF$buf0),
    .D(_4731_),
    .Y(_6157_)
);

NAND3X1 _15273_ (
    .A(_5741_),
    .B(_5742_),
    .C(_5747_),
    .Y(_5748_)
);

FILL FILL_5__15708_ (
);

FILL FILL_3__16322_ (
);

FILL FILL_1__8965_ (
);

FILL FILL_5__10423_ (
);

FILL FILL_1__8125_ (
);

FILL FILL_5__10003_ (
);

FILL FILL_2__15735_ (
);

FILL FILL_2__15315_ (
);

FILL FILL_4__6970_ (
);

FILL FILL_2__10870_ (
);

FILL FILL_2__10450_ (
);

FILL FILL_2__10030_ (
);

FILL FILL_1__14728_ (
);

NAND2X1 _7195_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_157_)
);

FILL FILL_1__14308_ (
);

FILL FILL_3__9412_ (
);

FILL FILL_0__6870_ (
);

FILL FILL_2__6888_ (
);

FILL FILL_5__9758_ (
);

FILL FILL_5__9338_ (
);

NOR2X1 _16058_ (
    .A(_6511_),
    .B(_6512_),
    .Y(_6513_)
);

INVX1 _11193_ (
    .A(\datapath_1.alu_1.ALUInA [26]),
    .Y(_2312_)
);

FILL FILL_5__11628_ (
);

FILL FILL_3__12662_ (
);

FILL FILL_5__11208_ (
);

FILL FILL_3__12242_ (
);

FILL FILL_4__7755_ (
);

FILL FILL_4__7335_ (
);

FILL FILL_2__11655_ (
);

FILL SFILL99400x19050 (
);

FILL FILL_2__11235_ (
);

FILL FILL_1__10648_ (
);

FILL FILL_5__15881_ (
);

FILL FILL_5__15461_ (
);

FILL FILL_5__15041_ (
);

FILL FILL112440x63050 (
);

NAND2X1 _9761_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1461_)
);

FILL FILL_0__7235_ (
);

NAND2X1 _9341_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1242_)
);

FILL FILL_4__14874_ (
);

FILL SFILL104360x12050 (
);

FILL FILL_4__14454_ (
);

FILL FILL_4__14034_ (
);

NAND2X1 _12398_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [18]),
    .Y(_3331_)
);

FILL FILL_3__13867_ (
);

FILL FILL_2__8614_ (
);

FILL FILL_3__13447_ (
);

FILL SFILL108600x63050 (
);

FILL FILL_1__14481_ (
);

FILL FILL_3__13027_ (
);

FILL FILL_1__14061_ (
);

FILL FILL_0__13894_ (
);

FILL FILL_0__13474_ (
);

FILL FILL_5__9091_ (
);

FILL SFILL104280x19050 (
);

FILL FILL_4__9901_ (
);

FILL FILL_2__13801_ (
);

FILL FILL_3__6957_ (
);

FILL FILL_5__16246_ (
);

FILL FILL_5__11381_ (
);

FILL FILL_1__9083_ (
);

FILL FILL_4__15659_ (
);

FILL FILL_4__15239_ (
);

FILL FILL_2__16273_ (
);

FILL FILL_4__10794_ (
);

FILL FILL_4__10374_ (
);

FILL FILL_0__9801_ (
);

FILL FILL_1__15686_ (
);

FILL FILL_1__15266_ (
);

FILL FILL_5__7824_ (
);

NAND3X1 _14964_ (
    .A(_5436_),
    .B(_5437_),
    .C(_5444_),
    .Y(_5445_)
);

FILL FILL_0__14679_ (
);

FILL FILL_0__14259_ (
);

INVX1 _14544_ (
    .A(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_5034_)
);

INVX1 _14124_ (
    .A(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_4622_)
);

FILL SFILL89400x17050 (
);

FILL FILL_1__7816_ (
);

FILL FILL_0__15620_ (
);

FILL FILL_0__15200_ (
);

FILL FILL_5__12586_ (
);

FILL FILL_5__12166_ (
);

BUFX2 _6886_ (
    .A(_2_[16]),
    .Y(memoryWriteData[16])
);

FILL SFILL49240x28050 (
);

FILL FILL_4__11999_ (
);

FILL FILL_4__11579_ (
);

FILL FILL_4__11159_ (
);

FILL FILL_2__12193_ (
);

FILL FILL_5__8609_ (
);

FILL FILL_1__11186_ (
);

FILL FILL_6__11906_ (
);

INVX1 _15749_ (
    .A(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_6212_)
);

NOR2X1 _15329_ (
    .A(_5802_),
    .B(_5800_),
    .Y(_5803_)
);

FILL FILL_4__12520_ (
);

FILL FILL_4__12100_ (
);

FILL FILL_0__8193_ (
);

NOR2X1 _10884_ (
    .A(\aluControl_1.inst [0]),
    .B(_2030_),
    .Y(_2031_)
);

FILL FILL_0__10179_ (
);

DFFSR _10464_ (
    .Q(\datapath_1.regfile_1.regOut[28] [10]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_1758_[10])
);

NAND2X1 _10044_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1609_)
);

FILL FILL_3__11933_ (
);

FILL FILL_3__11513_ (
);

FILL FILL_0__16405_ (
);

FILL SFILL94280x23050 (
);

FILL FILL_2__10926_ (
);

FILL FILL_2__9992_ (
);

FILL FILL_0__11960_ (
);

FILL FILL_2__10506_ (
);

FILL FILL_2__9152_ (
);

FILL FILL_0__11540_ (
);

FILL FILL_0__11120_ (
);

FILL FILL_4__9498_ (
);

FILL SFILL98520x74050 (
);

FILL FILL_4__9078_ (
);

FILL FILL_2__13398_ (
);

FILL FILL_5__14732_ (
);

FILL FILL_0__6926_ (
);

FILL FILL_5__14312_ (
);

NAND2X1 _8612_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_878_)
);

FILL SFILL33960x19050 (
);

FILL FILL_4__13725_ (
);

FILL FILL_4__13305_ (
);

FILL SFILL23240x72050 (
);

FILL FILL_0__9398_ (
);

FILL FILL_3__7495_ (
);

FILL FILL_3__7075_ (
);

OAI21X1 _11669_ (
    .A(_2179_),
    .B(_2347__bF$buf3),
    .C(_2770_),
    .Y(_2771_)
);

XOR2X1 _11249_ (
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2368_)
);

FILL FILL_3__12718_ (
);

FILL FILL_1__13752_ (
);

FILL FILL_1__13332_ (
);

FILL FILL_4__16197_ (
);

FILL SFILL84280x66050 (
);

FILL FILL_0__12745_ (
);

NAND2X1 _12610_ (
    .A(vdd),
    .B(memoryOutData[14]),
    .Y(_3453_)
);

FILL FILL_0__12325_ (
);

FILL FILL_5__8782_ (
);

FILL FILL_6__16104_ (
);

FILL FILL_5__8362_ (
);

FILL FILL_5__15937_ (
);

NAND2X1 _15082_ (
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .B(_5560_),
    .Y(_5561_)
);

FILL FILL_5__15517_ (
);

FILL SFILL8600x83050 (
);

DFFSR _9817_ (
    .Q(\datapath_1.regfile_1.regOut[23] [3]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_1433_[3])
);

FILL FILL_3__16131_ (
);

FILL FILL_1__8774_ (
);

FILL FILL_5__10652_ (
);

FILL FILL_1__8354_ (
);

FILL FILL_5__10232_ (
);

FILL FILL_2__15964_ (
);

FILL SFILL8680x40050 (
);

FILL FILL_2__15544_ (
);

FILL SFILL29320x62050 (
);

FILL SFILL84680x35050 (
);

FILL FILL_2__15124_ (
);

FILL FILL_1__14957_ (
);

FILL FILL_1__14537_ (
);

FILL FILL_1__14117_ (
);

FILL SFILL84200x64050 (
);

FILL FILL_3__9641_ (
);

NAND3X1 _13815_ (
    .A(_4311_),
    .B(_4312_),
    .C(_4319_),
    .Y(_4320_)
);

FILL FILL_3__9221_ (
);

FILL FILL_5__9987_ (
);

FILL FILL_5__9147_ (
);

FILL FILL_6__12024_ (
);

NAND2X1 _16287_ (
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .B(_5579_),
    .Y(_6736_)
);

FILL SFILL109480x64050 (
);

FILL FILL_5__11857_ (
);

FILL FILL_1__9979_ (
);

FILL FILL_3__12891_ (
);

FILL FILL_5__11437_ (
);

FILL FILL_3__12471_ (
);

FILL FILL_1__9139_ (
);

FILL FILL_5__11017_ (
);

FILL FILL_3__12051_ (
);

FILL FILL_4__7984_ (
);

FILL FILL_2__16329_ (
);

FILL FILL_4__7564_ (
);

FILL FILL_2__11884_ (
);

FILL FILL_2__11464_ (
);

FILL FILL_2__11044_ (
);

FILL FILL_1__10877_ (
);

FILL FILL_1__10037_ (
);

FILL FILL_5__15690_ (
);

FILL FILL_0__7884_ (
);

FILL FILL_5__15270_ (
);

FILL SFILL74280x64050 (
);

FILL FILL_0__7464_ (
);

NAND2X1 _9990_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1573_)
);

FILL FILL_0__7044_ (
);

DFFSR _9570_ (
    .Q(\datapath_1.regfile_1.regOut[21] [12]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_1303_[12])
);

INVX1 _9150_ (
    .A(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_1155_)
);

FILL FILL_6__13229_ (
);

FILL FILL_4__14683_ (
);

FILL FILL_4__14263_ (
);

FILL FILL_2__8843_ (
);

FILL FILL_0__10811_ (
);

FILL FILL_3__13676_ (
);

FILL FILL_3__13256_ (
);

FILL FILL_2__8003_ (
);

FILL FILL_1__14290_ (
);

FILL FILL_4__8769_ (
);

FILL FILL_0_BUFX2_insert700 (
);

FILL FILL_0_BUFX2_insert701 (
);

FILL FILL_4__8349_ (
);

FILL FILL_0_BUFX2_insert702 (
);

FILL FILL_0_BUFX2_insert703 (
);

FILL FILL_0_BUFX2_insert704 (
);

FILL FILL_2__12249_ (
);

FILL FILL_0__13283_ (
);

FILL FILL_0_BUFX2_insert705 (
);

FILL FILL_0_BUFX2_insert706 (
);

FILL FILL_0_BUFX2_insert707 (
);

FILL FILL_0_BUFX2_insert708 (
);

FILL FILL_0_BUFX2_insert709 (
);

FILL FILL_1__6840_ (
);

FILL FILL_2__13610_ (
);

FILL FILL_5__16055_ (
);

FILL FILL_0__8249_ (
);

FILL FILL_5__11190_ (
);

FILL FILL_4__15888_ (
);

FILL FILL_1__12603_ (
);

FILL FILL_4__15468_ (
);

FILL FILL_4__15048_ (
);

FILL FILL_2__16082_ (
);

FILL FILL_4__10183_ (
);

FILL FILL_0__9610_ (
);

FILL FILL_2__9628_ (
);

FILL FILL_2__9208_ (
);

FILL FILL_1__15495_ (
);

FILL FILL_1__15075_ (
);

FILL FILL_5__7633_ (
);

FILL FILL_5__7213_ (
);

FILL FILL_6__10930_ (
);

FILL FILL_0__14488_ (
);

AOI22X1 _14773_ (
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .B(_3891__bF$buf2),
    .C(_3998__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_5258_)
);

FILL FILL_0__14068_ (
);

AOI22X1 _14353_ (
    .A(_3891__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[4] [18]),
    .C(\datapath_1.regfile_1.regOut[8] [18]),
    .D(_4090_),
    .Y(_4847_)
);

FILL FILL_3__15822_ (
);

FILL FILL_3__15402_ (
);

FILL FILL_1__7625_ (
);

FILL FILL_1__7205_ (
);

FILL FILL_2__14815_ (
);

FILL FILL_5__12395_ (
);

FILL FILL_1__13808_ (
);

FILL FILL_4__11388_ (
);

FILL FILL_3__8912_ (
);

FILL FILL_5__8838_ (
);

AOI22X1 _15978_ (
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_6435_)
);

OAI22X1 _15558_ (
    .A(_5472__bF$buf3),
    .B(_4550_),
    .C(_4533_),
    .D(_5483__bF$buf1),
    .Y(_6026_)
);

AOI22X1 _15138_ (
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_5616_)
);

NAND2X1 _10693_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1940_)
);

NAND2X1 _10273_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1721_)
);

FILL FILL_5__10708_ (
);

FILL FILL_3__11742_ (
);

FILL FILL_3__11322_ (
);

FILL FILL_0__16214_ (
);

FILL SFILL68920x82050 (
);

FILL FILL_2__10315_ (
);

FILL FILL_2__9381_ (
);

FILL FILL_5__14961_ (
);

FILL FILL_5__14541_ (
);

FILL FILL112440x58050 (
);

FILL FILL_5__14121_ (
);

NAND2X1 _8841_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_990_)
);

DFFSR _8421_ (
    .Q(\datapath_1.regfile_1.regOut[12] [15]),
    .CLK(clk_bF$buf110),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_718_[15])
);

INVX1 _8001_ (
    .A(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_572_)
);

FILL FILL_4__13954_ (
);

FILL FILL_4__13534_ (
);

FILL FILL_4__13114_ (
);

OAI21X1 _11898_ (
    .A(_2972_),
    .B(IorD_bF$buf2),
    .C(_2973_),
    .Y(_1_[3])
);

NAND3X1 _11478_ (
    .A(_2470__bF$buf3),
    .B(_2588_),
    .C(_2592_),
    .Y(_2593_)
);

FILL SFILL33720x76050 (
);

XNOR2X1 _11058_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2177_)
);

FILL FILL_3__12527_ (
);

FILL FILL_1__13981_ (
);

FILL FILL_3__12107_ (
);

FILL FILL_1__13561_ (
);

FILL FILL_1__13141_ (
);

FILL FILL112040x44050 (
);

FILL SFILL89640x8050 (
);

FILL FILL_0__12974_ (
);

FILL FILL_0__12134_ (
);

FILL FILL_5__8591_ (
);

FILL FILL_5_BUFX2_insert100 (
);

FILL FILL_5_BUFX2_insert101 (
);

FILL FILL_5__15746_ (
);

FILL FILL_5__15326_ (
);

FILL FILL_5_BUFX2_insert102 (
);

FILL FILL_5_BUFX2_insert103 (
);

FILL FILL_3__16360_ (
);

FILL FILL_5_BUFX2_insert104 (
);

INVX1 _9626_ (
    .A(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_1391_)
);

FILL FILL_5_BUFX2_insert105 (
);

INVX1 _9206_ (
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_1236_)
);

FILL FILL_5__10881_ (
);

FILL FILL_5_BUFX2_insert106 (
);

FILL FILL_1__8583_ (
);

FILL FILL_5_BUFX2_insert107 (
);

FILL FILL_5__10041_ (
);

FILL FILL112440x13050 (
);

FILL FILL_5_BUFX2_insert108 (
);

FILL FILL_4__14739_ (
);

FILL FILL_5_BUFX2_insert109 (
);

FILL FILL_4__14319_ (
);

FILL FILL_2__15773_ (
);

FILL FILL_2__15353_ (
);

FILL FILL_3__8089_ (
);

FILL FILL_1__14766_ (
);

FILL FILL_1__14346_ (
);

FILL FILL_5__6904_ (
);

FILL FILL_3__9870_ (
);

FILL FILL_0__13759_ (
);

FILL FILL_0__13339_ (
);

NOR2X1 _13624_ (
    .A(_4132_),
    .B(_3983__bF$buf0),
    .Y(_4133_)
);

FILL FILL_3__9030_ (
);

DFFSR _13204_ (
    .Q(\datapath_1.PCJump [29]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3685_[29])
);

FILL FILL_5__9796_ (
);

FILL FILL_5__9376_ (
);

AOI22X1 _16096_ (
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_6550_)
);

FILL FILL_0__14700_ (
);

FILL FILL_1__9788_ (
);

FILL FILL_5__11666_ (
);

FILL FILL_1__9368_ (
);

FILL FILL_5__11246_ (
);

FILL FILL_3__12280_ (
);

FILL FILL_2__16138_ (
);

FILL FILL_4__7373_ (
);

FILL FILL_4__10659_ (
);

FILL FILL_4__10239_ (
);

FILL FILL_2__11693_ (
);

FILL FILL_2__11273_ (
);

FILL SFILL23720x74050 (
);

FILL FILL_1__10686_ (
);

FILL FILL_2_BUFX2_insert230 (
);

FILL FILL_1__10266_ (
);

FILL FILL_2_BUFX2_insert231 (
);

FILL FILL_2_BUFX2_insert232 (
);

INVX1 _14829_ (
    .A(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_5313_)
);

FILL FILL_2_BUFX2_insert233 (
);

INVX1 _14409_ (
    .A(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_4901_)
);

FILL FILL_2_BUFX2_insert234 (
);

FILL FILL_4__11600_ (
);

FILL FILL_2_BUFX2_insert235 (
);

FILL FILL_0__7693_ (
);

FILL FILL_2_BUFX2_insert236 (
);

FILL FILL_6__8660_ (
);

FILL FILL_2_BUFX2_insert237 (
);

FILL FILL_2_BUFX2_insert238 (
);

FILL FILL_2_BUFX2_insert239 (
);

FILL FILL_4__14492_ (
);

FILL FILL_4__14072_ (
);

FILL FILL_0__15905_ (
);

FILL FILL_2__8652_ (
);

FILL FILL_2__8232_ (
);

FILL FILL_3__13485_ (
);

FILL FILL_0__10620_ (
);

FILL FILL_4__8998_ (
);

FILL FILL_4__8578_ (
);

FILL FILL_2__12898_ (
);

FILL FILL_2__12478_ (
);

FILL FILL_2__12058_ (
);

FILL FILL_0__13092_ (
);

FILL FILL_5__13812_ (
);

FILL FILL_3__6995_ (
);

FILL FILL_5__16284_ (
);

FILL FILL_0__8898_ (
);

FILL FILL_6__9865_ (
);

FILL FILL_0__8478_ (
);

NAND2X1 _10749_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1957_)
);

FILL FILL_0__8058_ (
);

DFFSR _10329_ (
    .Q(\datapath_1.regfile_1.regOut[27] [3]),
    .CLK(clk_bF$buf0),
    .R(rst_bF$buf15),
    .S(vdd),
    .D(_1693_[3])
);

FILL FILL_4__15697_ (
);

FILL FILL_1__12832_ (
);

FILL FILL_1__12412_ (
);

FILL FILL_4__15277_ (
);

FILL FILL_2__9857_ (
);

FILL FILL_0__11825_ (
);

FILL FILL_2__9017_ (
);

FILL FILL_0__11405_ (
);

FILL FILL_5__7862_ (
);

FILL FILL_5__7442_ (
);

INVX1 _14582_ (
    .A(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_5071_)
);

FILL FILL_0__14297_ (
);

INVX1 _14162_ (
    .A(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_4660_)
);

FILL SFILL8600x78050 (
);

FILL FILL_3__15631_ (
);

FILL FILL_3__15211_ (
);

FILL FILL_1__7854_ (
);

FILL FILL_1__7434_ (
);

FILL SFILL8680x35050 (
);

FILL SFILL13720x72050 (
);

FILL FILL_2__14624_ (
);

FILL FILL_2__14204_ (
);

FILL FILL_1__13617_ (
);

FILL SFILL84200x59050 (
);

FILL FILL_1_BUFX2_insert250 (
);

FILL FILL_4__11197_ (
);

FILL FILL_1_BUFX2_insert251 (
);

FILL FILL_3__8721_ (
);

FILL SFILL99480x4050 (
);

FILL FILL_1_BUFX2_insert252 (
);

FILL SFILL48440x71050 (
);

FILL FILL_1_BUFX2_insert253 (
);

FILL SFILL84280x16050 (
);

FILL FILL_1_BUFX2_insert254 (
);

FILL FILL_1__16089_ (
);

FILL FILL_1_BUFX2_insert255 (
);

FILL FILL_1_BUFX2_insert256 (
);

FILL FILL_5__8647_ (
);

FILL FILL_5__8227_ (
);

FILL FILL_1_BUFX2_insert257 (
);

FILL FILL_1_BUFX2_insert258 (
);

FILL FILL_1_BUFX2_insert259 (
);

INVX1 _15787_ (
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_6249_)
);

NOR2X1 _15367_ (
    .A(_5839_),
    .B(_5836_),
    .Y(_5840_)
);

FILL SFILL69000x39050 (
);

FILL SFILL109480x59050 (
);

FILL FILL_3__16416_ (
);

FILL FILL_5__10937_ (
);

DFFSR _10082_ (
    .Q(\datapath_1.regfile_1.regOut[25] [12]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_1563_[12])
);

FILL FILL_1__8639_ (
);

FILL FILL_3__11971_ (
);

FILL FILL_5__10517_ (
);

FILL FILL_1__8219_ (
);

FILL FILL_3__11551_ (
);

FILL SFILL8600x33050 (
);

FILL FILL_3__11131_ (
);

FILL FILL_2__15829_ (
);

FILL FILL_2__15409_ (
);

FILL FILL_0__16023_ (
);

FILL FILL_2__10964_ (
);

FILL FILL_2__10544_ (
);

FILL FILL_2__10124_ (
);

INVX1 _7289_ (
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_199_)
);

FILL FILL_3__9926_ (
);

FILL FILL_3__9506_ (
);

FILL SFILL109880x28050 (
);

FILL SFILL84200x14050 (
);

FILL FILL_5__14770_ (
);

FILL SFILL74280x59050 (
);

FILL FILL_5__14350_ (
);

FILL FILL_0__6964_ (
);

INVX1 _8650_ (
    .A(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_903_)
);

INVX1 _8230_ (
    .A(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_684_)
);

FILL FILL_4__13763_ (
);

FILL FILL_4__13343_ (
);

FILL SFILL13640x34050 (
);

OAI21X1 _11287_ (
    .A(_2377_),
    .B(_2400_),
    .C(_2405_),
    .Y(_2406_)
);

FILL FILL_2__7503_ (
);

FILL FILL_3__12756_ (
);

FILL FILL_1__13790_ (
);

FILL FILL_3__12336_ (
);

FILL FILL_1__13370_ (
);

FILL FILL_4__7849_ (
);

FILL FILL_4__7429_ (
);

FILL FILL_2__11749_ (
);

FILL SFILL38840x83050 (
);

FILL FILL_0__12783_ (
);

FILL FILL_2__11329_ (
);

FILL FILL_0__12363_ (
);

FILL FILL_5__15975_ (
);

FILL SFILL74200x57050 (
);

FILL FILL_5__15555_ (
);

FILL FILL_0__7749_ (
);

FILL FILL_5__15135_ (
);

INVX1 _9855_ (
    .A(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_1503_)
);

FILL FILL_0__7329_ (
);

DFFSR _9435_ (
    .Q(\datapath_1.regfile_1.regOut[20] [5]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_1238_[5])
);

OAI21X1 _9015_ (
    .A(_1084_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1085_),
    .Y(_1043_[21])
);

FILL FILL_5__10690_ (
);

FILL FILL_1__8392_ (
);

FILL FILL_5__10270_ (
);

FILL SFILL74280x14050 (
);

FILL FILL_4__14968_ (
);

FILL FILL_4__14548_ (
);

FILL FILL_4__14128_ (
);

FILL FILL_2__15582_ (
);

FILL FILL_2__15162_ (
);

FILL FILL_2__8708_ (
);

FILL FILL_1__14995_ (
);

FILL FILL_1__14575_ (
);

FILL SFILL99480x63050 (
);

FILL FILL_1__14155_ (
);

FILL FILL_0__13988_ (
);

AOI22X1 _13853_ (
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .B(_4115_),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_4357_)
);

FILL FILL_0__13568_ (
);

FILL FILL_0__13148_ (
);

NOR2X1 _13433_ (
    .A(_3943_),
    .B(_3944__bF$buf0),
    .Y(_3945_)
);

OAI21X1 _13013_ (
    .A(_3659_),
    .B(vdd),
    .C(_3660_),
    .Y(_3620_[20])
);

FILL FILL_3__14902_ (
);

FILL FILL_5__11895_ (
);

FILL SFILL43800x21050 (
);

FILL FILL_5__11475_ (
);

FILL FILL_1__9597_ (
);

FILL SFILL74200x12050 (
);

FILL FILL_5__11055_ (
);

FILL FILL_2__16367_ (
);

FILL FILL_4__7182_ (
);

FILL FILL_4__10888_ (
);

FILL FILL_4__10048_ (
);

FILL FILL_2__11082_ (
);

FILL FILL_1__10495_ (
);

INVX1 _14638_ (
    .A(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_5126_)
);

INVX1 _14218_ (
    .A(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_4714_)
);

FILL FILL_0__7082_ (
);

FILL SFILL28840x81050 (
);

FILL FILL_1__16301_ (
);

FILL FILL_3__10822_ (
);

FILL FILL_3__10402_ (
);

FILL FILL_0__15714_ (
);

FILL FILL_2__8881_ (
);

FILL SFILL33800x64050 (
);

FILL FILL_2__8461_ (
);

FILL FILL_3__13294_ (
);

FILL FILL_4__8387_ (
);

FILL FILL_2__12287_ (
);

FILL FILL_5__13621_ (
);

DFFSR _7921_ (
    .Q(\datapath_1.regfile_1.regOut[8] [27]),
    .CLK(clk_bF$buf73),
    .R(rst_bF$buf98),
    .S(vdd),
    .D(_458_[27])
);

INVX1 _7501_ (
    .A(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_320_)
);

FILL FILL_4__12614_ (
);

FILL FILL_5__16093_ (
);

INVX1 _10978_ (
    .A(\control_1.reg_state.dout [2]),
    .Y(_2103_)
);

INVX1 _10558_ (
    .A(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_1870_)
);

INVX1 _10138_ (
    .A(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_1651_)
);

FILL FILL_3__11607_ (
);

FILL FILL_1__12641_ (
);

FILL FILL_4__15086_ (
);

FILL FILL_1__12221_ (
);

FILL FILL_2__9666_ (
);

FILL FILL_3__14499_ (
);

FILL FILL_0__11634_ (
);

FILL FILL_2__9246_ (
);

FILL FILL_0__11214_ (
);

FILL FILL_3__14079_ (
);

FILL FILL_6__15833_ (
);

FILL FILL_6__15413_ (
);

FILL FILL_5__7671_ (
);

FILL FILL_5__7251_ (
);

FILL SFILL64200x10050 (
);

INVX1 _14391_ (
    .A(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_4884_)
);

FILL FILL_5__14826_ (
);

FILL FILL_3__15860_ (
);

FILL FILL_5__14406_ (
);

FILL FILL_3__15440_ (
);

INVX1 _8706_ (
    .A(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_920_)
);

FILL FILL_3__15020_ (
);

FILL FILL_1__7243_ (
);

FILL FILL_4__13819_ (
);

FILL FILL_2__14853_ (
);

FILL FILL_2__14433_ (
);

FILL FILL_3__7589_ (
);

FILL FILL_2__14013_ (
);

FILL FILL_3__7169_ (
);

FILL FILL_1__13846_ (
);

FILL FILL_1__13426_ (
);

FILL FILL_1__13006_ (
);

FILL FILL_3__8950_ (
);

FILL FILL_3__8530_ (
);

FILL FILL_0__12839_ (
);

INVX1 _12704_ (
    .A(\aluControl_1.inst [3]),
    .Y(_3495_)
);

FILL FILL_0__12419_ (
);

FILL FILL_3__8110_ (
);

FILL FILL_5__8876_ (
);

FILL FILL_5__8456_ (
);

FILL SFILL54200x53050 (
);

FILL FILL_6__11753_ (
);

FILL FILL_6__11333_ (
);

OAI22X1 _15596_ (
    .A(_5485__bF$buf2),
    .B(_4588_),
    .C(_5483__bF$buf0),
    .D(_4580_),
    .Y(_6063_)
);

NAND3X1 _15176_ (
    .A(_5651_),
    .B(_5652_),
    .C(_5648_),
    .Y(_5653_)
);

FILL FILL_3__16225_ (
);

FILL FILL_1__8868_ (
);

FILL FILL_5__10746_ (
);

FILL FILL_1__8448_ (
);

FILL FILL_3__11780_ (
);

FILL FILL_3__11360_ (
);

FILL FILL_2__15638_ (
);

FILL FILL_4__6873_ (
);

FILL FILL_2__15218_ (
);

FILL SFILL58520x61050 (
);

FILL FILL_0__16252_ (
);

FILL FILL_2__10773_ (
);

OAI21X1 _7098_ (
    .A(_111_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_112_),
    .Y(_68_[22])
);

FILL SFILL23720x69050 (
);

FILL FILL_3__9735_ (
);

AOI22X1 _13909_ (
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .B(_4102_),
    .C(_4001__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_4412_)
);

FILL FILL_6__7740_ (
);

FILL FILL_4__13992_ (
);

FILL FILL_4__13572_ (
);

FILL FILL_4__13152_ (
);

OAI21X1 _11096_ (
    .A(_2209_),
    .B(_2180_),
    .C(_2214_),
    .Y(_2215_)
);

FILL FILL_3__12985_ (
);

FILL FILL_2__7732_ (
);

FILL FILL_2__7312_ (
);

FILL FILL_3__12145_ (
);

FILL FILL_4__7238_ (
);

FILL FILL_2__11978_ (
);

FILL FILL_2__11558_ (
);

FILL FILL_0__12592_ (
);

FILL FILL_2__11138_ (
);

FILL FILL_0__12172_ (
);

FILL SFILL74120x3050 (
);

FILL SFILL23720x24050 (
);

FILL FILL_5__15784_ (
);

FILL FILL_5__15364_ (
);

FILL FILL_0__7978_ (
);

FILL FILL_0__7558_ (
);

OAI21X1 _9664_ (
    .A(_1415_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .C(_1416_),
    .Y(_1368_[24])
);

OAI21X1 _9244_ (
    .A(_1196_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1197_),
    .Y(_1173_[12])
);

FILL FILL_1__11912_ (
);

FILL FILL_4__14777_ (
);

FILL FILL_4__14357_ (
);

FILL SFILL48920x73050 (
);

FILL FILL_2__15391_ (
);

FILL FILL_0__10905_ (
);

FILL FILL_2__8517_ (
);

FILL FILL_1__14384_ (
);

FILL FILL_5__6942_ (
);

FILL FILL_1_BUFX2_insert1010 (
);

FILL FILL_1_BUFX2_insert1011 (
);

FILL FILL_1_BUFX2_insert1012 (
);

FILL FILL_0__13797_ (
);

FILL FILL_1_BUFX2_insert1013 (
);

NOR2X1 _13662_ (
    .A(_4169_),
    .B(_4166_),
    .Y(_4170_)
);

FILL FILL_1_BUFX2_insert1014 (
);

FILL FILL_0__13377_ (
);

AOI21X1 _13242_ (
    .A(_3750_),
    .B(_3782_),
    .C(_3784_),
    .Y(_3785_)
);

FILL FILL_1_BUFX2_insert1015 (
);

FILL FILL_1_BUFX2_insert1016 (
);

FILL FILL_1_BUFX2_insert1017 (
);

FILL FILL_3__14711_ (
);

FILL FILL_1_BUFX2_insert1018 (
);

FILL FILL_1_BUFX2_insert1019 (
);

FILL FILL_1__6934_ (
);

FILL FILL_4__9804_ (
);

FILL SFILL13720x67050 (
);

FILL FILL_2__13704_ (
);

FILL FILL_5__16149_ (
);

FILL SFILL109560x47050 (
);

FILL FILL_5__11284_ (
);

FILL FILL_2__16176_ (
);

FILL FILL_4__10697_ (
);

FILL FILL_4__10277_ (
);

FILL FILL_3__7801_ (
);

FILL FILL_1__15589_ (
);

FILL FILL_1__15169_ (
);

FILL FILL_5__7727_ (
);

FILL FILL_5__7307_ (
);

FILL FILL_2_BUFX2_insert610 (
);

FILL FILL_2_BUFX2_insert611 (
);

FILL FILL_2_BUFX2_insert612 (
);

AOI22X1 _14867_ (
    .A(\datapath_1.regfile_1.regOut[23] [29]),
    .B(_4038__bF$buf2),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_5350_)
);

FILL FILL_2_BUFX2_insert613 (
);

FILL FILL_2_BUFX2_insert614 (
);

AOI22X1 _14447_ (
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .B(_4135_),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_4939_)
);

FILL FILL_2_BUFX2_insert615 (
);

OAI22X1 _14027_ (
    .A(_4525_),
    .B(_3925_),
    .C(_3977__bF$buf4),
    .D(_4526_),
    .Y(_4527_)
);

FILL FILL_3__15916_ (
);

FILL FILL_2_BUFX2_insert616 (
);

FILL FILL_2_BUFX2_insert617 (
);

FILL FILL_2_BUFX2_insert618 (
);

FILL FILL_1__16110_ (
);

FILL FILL_2_BUFX2_insert619 (
);

FILL FILL_1__7719_ (
);

FILL SFILL8600x28050 (
);

FILL FILL_3__10631_ (
);

FILL FILL_2__14909_ (
);

FILL FILL_0__15943_ (
);

FILL FILL_0__15523_ (
);

FILL FILL_0__15103_ (
);

FILL SFILL13720x22050 (
);

FILL FILL_5__12489_ (
);

FILL FILL_2__8270_ (
);

FILL FILL_5__12069_ (
);

FILL FILL_4__8196_ (
);

FILL FILL_2__12096_ (
);

FILL SFILL38920x71050 (
);

FILL FILL_5__13850_ (
);

FILL FILL_5__13430_ (
);

FILL FILL_5__13010_ (
);

INVX1 _7730_ (
    .A(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_432_)
);

INVX1 _7310_ (
    .A(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_213_)
);

FILL FILL_1__11089_ (
);

FILL FILL_6__11809_ (
);

FILL FILL_4__12843_ (
);

FILL FILL_4__12423_ (
);

FILL FILL_4__12003_ (
);

FILL SFILL13640x29050 (
);

FILL FILL_6__9483_ (
);

INVX1 _10787_ (
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_1982_)
);

FILL FILL_0__8096_ (
);

INVX1 _10367_ (
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .Y(_1763_)
);

FILL FILL_3__11836_ (
);

FILL FILL_1__12870_ (
);

FILL FILL_3__11416_ (
);

FILL FILL_1__12450_ (
);

FILL FILL_1__12030_ (
);

FILL FILL_4__6929_ (
);

FILL FILL_0__16308_ (
);

FILL FILL_2__10829_ (
);

FILL FILL_2__9895_ (
);

FILL FILL_2__9475_ (
);

FILL FILL_2__10409_ (
);

FILL FILL_0__11863_ (
);

FILL FILL_0__11443_ (
);

FILL FILL_0__11023_ (
);

FILL FILL_5__7480_ (
);

FILL FILL_5__7060_ (
);

FILL SFILL3560x70050 (
);

FILL FILL_5__14635_ (
);

FILL FILL_5__14215_ (
);

DFFSR _8935_ (
    .Q(\datapath_1.regfile_1.regOut[16] [17]),
    .CLK(clk_bF$buf96),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_978_[17])
);

OAI21X1 _8515_ (
    .A(_832_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_833_),
    .Y(_783_[25])
);

FILL FILL_1__7892_ (
);

FILL FILL_1__7472_ (
);

FILL FILL_1__7052_ (
);

FILL FILL_4__13628_ (
);

FILL FILL_4__13208_ (
);

FILL FILL_2__14662_ (
);

FILL FILL_2__14242_ (
);

FILL FILL112200x65050 (
);

FILL FILL_3_BUFX2_insert70 (
);

FILL SFILL99480x58050 (
);

FILL FILL_1__13655_ (
);

FILL FILL_3_BUFX2_insert71 (
);

FILL FILL_1__13235_ (
);

FILL FILL_3_BUFX2_insert72 (
);

FILL FILL_3_BUFX2_insert73 (
);

FILL FILL_3_BUFX2_insert74 (
);

FILL SFILL44040x7050 (
);

FILL FILL_3_BUFX2_insert75 (
);

FILL FILL_3_BUFX2_insert76 (
);

FILL FILL_1_BUFX2_insert630 (
);

FILL FILL_3_BUFX2_insert77 (
);

FILL FILL_1_BUFX2_insert631 (
);

FILL FILL_0__12648_ (
);

FILL FILL_1_BUFX2_insert632 (
);

FILL FILL_3_BUFX2_insert78 (
);

DFFSR _12933_ (
    .Q(\datapath_1.a [14]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3555_[14])
);

FILL FILL_1_BUFX2_insert633 (
);

OAI21X1 _12513_ (
    .A(_3407_),
    .B(vdd),
    .C(_3408_),
    .Y(_3360_[24])
);

FILL FILL_3_BUFX2_insert79 (
);

FILL FILL_0__12228_ (
);

FILL FILL_1_BUFX2_insert634 (
);

FILL FILL_1_BUFX2_insert635 (
);

FILL SFILL38840x33050 (
);

FILL FILL_1_BUFX2_insert636 (
);

FILL FILL_6__16007_ (
);

FILL FILL_1_BUFX2_insert637 (
);

FILL FILL_5__8265_ (
);

FILL FILL_1_BUFX2_insert638 (
);

FILL FILL_1_BUFX2_insert639 (
);

FILL SFILL23800x50 (
);

FILL FILL_3__16034_ (
);

FILL FILL_5__10975_ (
);

FILL FILL_5__10555_ (
);

FILL FILL_5__10135_ (
);

FILL FILL_1__8257_ (
);

FILL FILL_2__15867_ (
);

FILL FILL_2__15447_ (
);

FILL FILL_2__15027_ (
);

FILL FILL_0__16061_ (
);

FILL FILL_2__10162_ (
);

FILL FILL112200x20050 (
);

FILL SFILL99480x13050 (
);

FILL FILL_3__9544_ (
);

FILL FILL_3__9124_ (
);

AND2X2 _13718_ (
    .A(_3917_),
    .B(_3888_),
    .Y(_4225_)
);

FILL SFILL28840x76050 (
);

FILL FILL_1__15801_ (
);

FILL FILL_4__13381_ (
);

FILL SFILL33800x59050 (
);

FILL FILL_2__7961_ (
);

BUFX2 BUFX2_insert300 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf3 )
);

BUFX2 BUFX2_insert301 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf2 )
);

FILL FILL_3__12374_ (
);

FILL FILL_2__7121_ (
);

BUFX2 BUFX2_insert302 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf1 )
);

BUFX2 BUFX2_insert303 (
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf0 )
);

FILL FILL112120x27050 (
);

FILL FILL_4__7887_ (
);

BUFX2 BUFX2_insert304 (
    .A(_3032_),
    .Y(_3032__bF$buf4)
);

BUFX2 BUFX2_insert305 (
    .A(_3032_),
    .Y(_3032__bF$buf3)
);

FILL FILL_4__7467_ (
);

BUFX2 BUFX2_insert306 (
    .A(_3032_),
    .Y(_3032__bF$buf2)
);

FILL FILL_4__7047_ (
);

BUFX2 BUFX2_insert307 (
    .A(_3032_),
    .Y(_3032__bF$buf1)
);

FILL FILL_2__11787_ (
);

BUFX2 BUFX2_insert308 (
    .A(_3032_),
    .Y(_3032__bF$buf0)
);

FILL FILL_2__11367_ (
);

BUFX2 BUFX2_insert309 (
    .A(_2341_),
    .Y(_2341__bF$buf3)
);

FILL FILL_5__12701_ (
);

FILL FILL_5__15593_ (
);

FILL FILL_5__15173_ (
);

OAI21X1 _9893_ (
    .A(_1527_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1528_),
    .Y(_1498_[15])
);

FILL FILL_0__7367_ (
);

FILL FILL_6__8754_ (
);

OAI21X1 _9473_ (
    .A(_1308_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .C(_1309_),
    .Y(_1303_[3])
);

DFFSR _9053_ (
    .Q(\datapath_1.regfile_1.regOut[17] [7]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_1043_[7])
);

FILL FILL_4__14586_ (
);

FILL FILL_1__11721_ (
);

FILL SFILL28840x31050 (
);

FILL FILL_4__14166_ (
);

FILL FILL_1__11301_ (
);

FILL FILL_3__13999_ (
);

FILL FILL_2__8746_ (
);

FILL FILL_3__13579_ (
);

FILL FILL_2__8326_ (
);

FILL FILL_3__13159_ (
);

FILL FILL_1__14193_ (
);

INVX1 _13891_ (
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_4394_)
);

NAND3X1 _13471_ (
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3904_),
    .C(_3879_),
    .Y(_3983_)
);

DFFSR _13051_ (
    .Q(_2_[4]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_3620_[4])
);

FILL FILL_5__13906_ (
);

FILL FILL_3__14940_ (
);

FILL FILL_3__14520_ (
);

FILL FILL_3__14100_ (
);

FILL FILL_4__9613_ (
);

FILL FILL_2__13933_ (
);

FILL FILL_5__16378_ (
);

FILL FILL_2__13513_ (
);

FILL FILL_6__9539_ (
);

FILL FILL_5__11093_ (
);

FILL FILL_1__12506_ (
);

FILL SFILL18840x74050 (
);

FILL FILL_0__9933_ (
);

FILL FILL_3__7610_ (
);

FILL FILL_0__11919_ (
);

FILL FILL_0__9513_ (
);

FILL FILL_1__15398_ (
);

FILL FILL_5__7956_ (
);

FILL FILL_5__7116_ (
);

FILL FILL_4__16312_ (
);

FILL FILL_6__10413_ (
);

INVX1 _14676_ (
    .A(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_5163_)
);

FILL SFILL13800x4050 (
);

OAI22X1 _14256_ (
    .A(_3902__bF$buf1),
    .B(_4751_),
    .C(_4750_),
    .D(_3944__bF$buf2),
    .Y(_4752_)
);

FILL FILL_3__15725_ (
);

FILL FILL_3__15305_ (
);

FILL SFILL13720x9050 (
);

FILL FILL_1__7948_ (
);

FILL FILL_1__7108_ (
);

FILL FILL_3__10440_ (
);

FILL FILL_3__10020_ (
);

FILL FILL_2__14718_ (
);

FILL FILL_0__15752_ (
);

FILL FILL_0__15332_ (
);

FILL FILL_5__12298_ (
);

FILL FILL_4__12652_ (
);

FILL FILL_4__12232_ (
);

DFFSR _10596_ (
    .Q(\datapath_1.regfile_1.regOut[29] [14]),
    .CLK(clk_bF$buf11),
    .R(rst_bF$buf3),
    .S(vdd),
    .D(_1823_[14])
);

OAI21X1 _10176_ (
    .A(_1675_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1676_),
    .Y(_1628_[24])
);

FILL FILL_3__11645_ (
);

FILL FILL_3__11225_ (
);

FILL FILL_0__16117_ (
);

INVX1 _16402_ (
    .A(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_6822_)
);

FILL FILL_2__10638_ (
);

FILL FILL_2__9284_ (
);

FILL FILL_0__11672_ (
);

FILL FILL_0__11252_ (
);

FILL SFILL23720x19050 (
);

FILL FILL_5__14864_ (
);

FILL FILL_5__14444_ (
);

FILL FILL_5__14024_ (
);

OAI21X1 _8744_ (
    .A(_944_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_945_),
    .Y(_913_[16])
);

FILL SFILL69080x83050 (
);

OAI21X1 _8324_ (
    .A(_725_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_726_),
    .Y(_718_[4])
);

FILL FILL_4__13857_ (
);

FILL FILL_4__13437_ (
);

FILL FILL_2__14891_ (
);

FILL FILL_2__14471_ (
);

FILL FILL_4__13017_ (
);

FILL FILL_2__14051_ (
);

FILL FILL_1__13884_ (
);

FILL FILL_1__13464_ (
);

FILL FILL_1__13044_ (
);

FILL FILL_0__12877_ (
);

OAI21X1 _12742_ (
    .A(_3519_),
    .B(IRWrite_bF$buf0),
    .C(_3520_),
    .Y(_3490_[15])
);

FILL FILL_0__12457_ (
);

FILL FILL_0__12037_ (
);

NAND3X1 _12322_ (
    .A(_3278_),
    .B(_3279_),
    .C(_3280_),
    .Y(\datapath_1.alu_1.ALUInB [26])
);

FILL FILL_5__8494_ (
);

FILL FILL_5__8074_ (
);

FILL FILL_5__15649_ (
);

FILL FILL_5__15229_ (
);

DFFSR _9949_ (
    .Q(\datapath_1.regfile_1.regOut[24] [7]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_1498_[7])
);

FILL FILL_3__16263_ (
);

NAND2X1 _9529_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1347_)
);

FILL FILL_5__10784_ (
);

NAND2X1 _9109_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1128_)
);

FILL FILL_1__8486_ (
);

FILL FILL_5__10364_ (
);

FILL FILL_1__8066_ (
);

FILL FILL_2__15676_ (
);

FILL FILL_2__15256_ (
);

FILL FILL_0__16290_ (
);

FILL SFILL48920x23050 (
);

FILL FILL_2__10391_ (
);

FILL FILL_1__14669_ (
);

FILL FILL_1__14249_ (
);

FILL FILL_0_BUFX2_insert290 (
);

FILL FILL_0_BUFX2_insert291 (
);

FILL FILL_0_BUFX2_insert292 (
);

FILL FILL_0_BUFX2_insert293 (
);

FILL FILL_3__9773_ (
);

FILL FILL_3__9353_ (
);

FILL FILL_0_BUFX2_insert294 (
);

INVX1 _13947_ (
    .A(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_4449_)
);

FILL FILL_0_BUFX2_insert295 (
);

INVX8 _13527_ (
    .A(_3916_),
    .Y(_4038_)
);

FILL FILL_0_BUFX2_insert296 (
);

NAND2X1 _13107_ (
    .A(PCEn_bF$buf2),
    .B(\datapath_1.mux_pcsrc.dout [9]),
    .Y(_3703_)
);

FILL FILL_0_BUFX2_insert297 (
);

FILL FILL_0_BUFX2_insert298 (
);

FILL FILL_5__9279_ (
);

FILL FILL_0_BUFX2_insert299 (
);

FILL FILL_1__15610_ (
);

FILL FILL_6__12996_ (
);

FILL FILL_0__14603_ (
);

FILL SFILL13720x17050 (
);

FILL FILL_5__11989_ (
);

FILL FILL_5__11569_ (
);

FILL FILL_2__7350_ (
);

FILL FILL_5__11149_ (
);

FILL FILL_3__12183_ (
);

FILL SFILL59080x81050 (
);

FILL FILL_4__7696_ (
);

FILL FILL_2__11596_ (
);

FILL SFILL38920x66050 (
);

FILL FILL_2__11176_ (
);

FILL FILL_5__12510_ (
);

FILL FILL_1__10169_ (
);

FILL FILL_4__11923_ (
);

FILL FILL_4__11503_ (
);

FILL FILL_0__7596_ (
);

FILL FILL_0__7176_ (
);

FILL FILL_6__8143_ (
);

NAND2X1 _9282_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1223_)
);

FILL FILL_3__10916_ (
);

FILL FILL_1__11950_ (
);

FILL FILL_4__14395_ (
);

FILL FILL_1__11530_ (
);

FILL FILL_1__11110_ (
);

FILL FILL_0__15808_ (
);

FILL FILL_2__8975_ (
);

FILL FILL_0__10943_ (
);

FILL FILL_3__13388_ (
);

FILL FILL_0__10523_ (
);

FILL FILL_2__8135_ (
);

FILL FILL_0__10103_ (
);

FILL FILL_5__6980_ (
);

FILL SFILL3560x65050 (
);

NOR2X1 _13280_ (
    .A(_3781_),
    .B(_3819_),
    .Y(\datapath_1.regfile_1.regEn [4])
);

FILL FILL_5__13715_ (
);

FILL SFILL38920x21050 (
);

FILL SFILL104440x82050 (
);

FILL FILL_1__6972_ (
);

FILL FILL_4__9422_ (
);

FILL FILL_4__12708_ (
);

FILL FILL_4__9002_ (
);

FILL FILL_2__13742_ (
);

FILL FILL_2__13322_ (
);

FILL FILL_5__16187_ (
);

FILL FILL_3__6898_ (
);

FILL FILL_6__9348_ (
);

FILL FILL_1__12735_ (
);

FILL FILL_1__12315_ (
);

FILL SFILL38040x45050 (
);

FILL FILL_0__9742_ (
);

FILL FILL_0__11728_ (
);

FILL FILL_0__11308_ (
);

FILL SFILL38840x28050 (
);

FILL FILL_5__7765_ (
);

FILL FILL_5__7345_ (
);

FILL FILL_4__16121_ (
);

FILL SFILL83480x54050 (
);

INVX1 _14485_ (
    .A(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_4976_)
);

AOI22X1 _14065_ (
    .A(\datapath_1.regfile_1.regOut[11] [12]),
    .B(_3950__bF$buf3),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_4565_)
);

FILL FILL_3__15954_ (
);

FILL FILL_3__15534_ (
);

FILL FILL_3__15114_ (
);

FILL SFILL28920x64050 (
);

FILL SFILL3560x20050 (
);

FILL FILL_1__7757_ (
);

FILL FILL_1__7337_ (
);

FILL FILL_2__14947_ (
);

FILL FILL_0__15981_ (
);

FILL FILL_2__14527_ (
);

FILL FILL_0__15561_ (
);

FILL FILL_2__14107_ (
);

FILL FILL_0__15141_ (
);

FILL SFILL28520x50050 (
);

FILL FILL_3__8624_ (
);

FILL FILL_3__8204_ (
);

FILL FILL_4__12881_ (
);

FILL FILL_4__12461_ (
);

FILL FILL_4__12041_ (
);

FILL FILL_3__16319_ (
);

FILL FILL_5__9911_ (
);

FILL FILL_3__11874_ (
);

FILL FILL_3__11454_ (
);

FILL FILL_3__11034_ (
);

FILL FILL_4__6967_ (
);

FILL FILL_0__16346_ (
);

NAND2X1 _16211_ (
    .A(\datapath_1.regfile_1.regOut[2] [29]),
    .B(_5479_),
    .Y(_6662_)
);

FILL FILL_2__10447_ (
);

FILL FILL_2__10027_ (
);

FILL FILL_0__11481_ (
);

FILL FILL_2__9093_ (
);

FILL FILL_0__11061_ (
);

FILL FILL_1__9903_ (
);

FILL FILL_6__15260_ (
);

FILL FILL_3__9409_ (
);

FILL FILL_5__14673_ (
);

FILL FILL_0__6867_ (
);

FILL FILL_5__14253_ (
);

OAI21X1 _8973_ (
    .A(_1056_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1057_),
    .Y(_1043_[7])
);

FILL FILL_6__7834_ (
);

DFFSR _8553_ (
    .Q(\datapath_1.regfile_1.regOut[13] [19]),
    .CLK(clk_bF$buf72),
    .R(rst_bF$buf36),
    .S(vdd),
    .D(_783_[19])
);

NAND2X1 _8133_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_640_)
);

FILL FILL_1__7090_ (
);

FILL SFILL28840x26050 (
);

FILL FILL_4__13666_ (
);

FILL FILL_1__10801_ (
);

FILL FILL_4__13246_ (
);

FILL FILL_2__14280_ (
);

FILL FILL_2__7826_ (
);

FILL FILL_3__12659_ (
);

FILL FILL_3__12239_ (
);

FILL FILL_1__13693_ (
);

FILL FILL_1__13273_ (
);

OAI21X1 _12971_ (
    .A(_3631_),
    .B(vdd),
    .C(_3632_),
    .Y(_3620_[6])
);

DFFSR _12551_ (
    .Q(ALUOut[16]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[16])
);

FILL FILL_0__12266_ (
);

NAND2X1 _12131_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.a [5]),
    .Y(_3141_)
);

FILL FILL_3__13600_ (
);

FILL FILL_6__11180_ (
);

FILL FILL_5__15878_ (
);

FILL FILL_5__15458_ (
);

FILL FILL_5__15038_ (
);

FILL FILL_6__8619_ (
);

FILL FILL_3__16072_ (
);

NAND2X1 _9758_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1459_)
);

NAND2X1 _9338_ (
    .A(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1240_)
);

FILL FILL_5__10173_ (
);

FILL FILL_2__15485_ (
);

FILL FILL_2__15065_ (
);

FILL FILL_1__14898_ (
);

FILL FILL_1__14478_ (
);

FILL FILL_1__14058_ (
);

FILL FILL_4__15812_ (
);

INVX1 _13756_ (
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_4262_)
);

FILL FILL_3__9162_ (
);

AOI21X1 _13336_ (
    .A(_3751_),
    .B(_3772_),
    .C(_3820_),
    .Y(_3859_)
);

FILL FILL_3__14805_ (
);

FILL FILL_5__9088_ (
);

FILL FILL_0__14832_ (
);

FILL FILL_0__14412_ (
);

FILL FILL_5__11798_ (
);

FILL FILL_5__11378_ (
);

FILL FILL_4__7085_ (
);

FILL SFILL18840x24050 (
);

FILL FILL_1__10398_ (
);

FILL FILL_4__11732_ (
);

FILL FILL_4__11312_ (
);

NAND2X1 _9091_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1116_)
);

FILL FILL_1__16204_ (
);

FILL FILL_3__10305_ (
);

NAND3X1 _15902_ (
    .A(_6351_),
    .B(_6360_),
    .C(_6355_),
    .Y(_6361_)
);

FILL FILL_0__15617_ (
);

FILL FILL_2__8784_ (
);

FILL FILL_0__10752_ (
);

FILL FILL_2__8364_ (
);

FILL FILL_5__13944_ (
);

FILL FILL_5__13524_ (
);

FILL FILL_5__13104_ (
);

OAI21X1 _7824_ (
    .A(_473_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_474_),
    .Y(_458_[8])
);

DFFSR _7404_ (
    .Q(\datapath_1.regfile_1.regOut[4] [22]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf17),
    .S(vdd),
    .D(_198_[22])
);

FILL FILL_4_BUFX2_insert520 (
);

FILL FILL_4_BUFX2_insert521 (
);

FILL FILL_4__9651_ (
);

FILL FILL_4__9231_ (
);

FILL FILL_4_BUFX2_insert522 (
);

FILL FILL_4_BUFX2_insert523 (
);

FILL FILL_4__12517_ (
);

FILL FILL_2__13971_ (
);

FILL FILL_4_BUFX2_insert524 (
);

FILL FILL_2__13551_ (
);

FILL FILL_2__13131_ (
);

FILL FILL_4_BUFX2_insert525 (
);

FILL FILL_4_BUFX2_insert526 (
);

FILL FILL_4_BUFX2_insert527 (
);

FILL FILL_4_BUFX2_insert528 (
);

FILL FILL_4_BUFX2_insert529 (
);

FILL FILL_1__12964_ (
);

FILL FILL_1__12124_ (
);

FILL FILL_2__9989_ (
);

FILL FILL_0__9551_ (
);

FILL FILL_0__11957_ (
);

FILL FILL_2__9149_ (
);

FILL FILL_0__9131_ (
);

OAI21X1 _11822_ (
    .A(_2911_),
    .B(_2541_),
    .C(_2462__bF$buf0),
    .Y(_2912_)
);

FILL FILL_0__11537_ (
);

FILL SFILL114520x72050 (
);

FILL FILL_0__11117_ (
);

INVX1 _11402_ (
    .A(_2258_),
    .Y(_2519_)
);

FILL FILL_5__7994_ (
);

FILL FILL_6__15736_ (
);

FILL FILL_6__15316_ (
);

FILL FILL_5__7574_ (
);

FILL FILL_4__16350_ (
);

FILL FILL_6__10031_ (
);

INVX1 _14294_ (
    .A(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_4789_)
);

FILL FILL_5__14729_ (
);

FILL FILL_3__15763_ (
);

FILL FILL_5__14309_ (
);

FILL FILL_3__15343_ (
);

NAND2X1 _8609_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_876_)
);

FILL FILL_1__7986_ (
);

FILL FILL_1__7566_ (
);

FILL SFILL69080x33050 (
);

FILL FILL_2__14756_ (
);

FILL FILL_0__15790_ (
);

FILL FILL_2__14336_ (
);

FILL FILL_0__15370_ (
);

FILL SFILL48920x18050 (
);

FILL FILL_1__13749_ (
);

FILL FILL_1__13329_ (
);

FILL FILL_3__8853_ (
);

FILL FILL_3__8013_ (
);

NAND2X1 _12607_ (
    .A(vdd),
    .B(memoryOutData[13]),
    .Y(_3451_)
);

FILL FILL_5__8779_ (
);

FILL FILL_5__8359_ (
);

FILL SFILL114040x65050 (
);

FILL FILL_6__11656_ (
);

OAI22X1 _15499_ (
    .A(_4492_),
    .B(_5539__bF$buf3),
    .C(_5552__bF$buf0),
    .D(_4491_),
    .Y(_5968_)
);

FILL FILL_6__11236_ (
);

FILL FILL_4__12270_ (
);

INVX1 _15079_ (
    .A(_5549__bF$buf1),
    .Y(_5558_)
);

FILL FILL_3__16128_ (
);

FILL FILL_5__10649_ (
);

FILL FILL_2__6850_ (
);

FILL FILL_5__9720_ (
);

FILL FILL_3__11683_ (
);

FILL FILL_5__9300_ (
);

FILL FILL_3__11263_ (
);

DFFSR _16440_ (
    .Q(\datapath_1.regfile_1.regOut[0] [23]),
    .CLK(clk_bF$buf75),
    .R(rst_bF$buf0),
    .S(vdd),
    .D(_6769_[23])
);

FILL FILL_0__16155_ (
);

NAND3X1 _16020_ (
    .A(_6469_),
    .B(_6470_),
    .C(_6475_),
    .Y(_6476_)
);

FILL FILL_2__10676_ (
);

FILL FILL_2__10256_ (
);

FILL FILL_0__11290_ (
);

FILL FILL_3__9638_ (
);

FILL FILL_3_BUFX2_insert540 (
);

FILL FILL_3__9218_ (
);

FILL FILL_3_BUFX2_insert541 (
);

FILL FILL_3_BUFX2_insert542 (
);

FILL SFILL3640x53050 (
);

FILL FILL_5__14482_ (
);

FILL FILL_3_BUFX2_insert543 (
);

FILL FILL_3_BUFX2_insert544 (
);

FILL FILL_5__14062_ (
);

NAND2X1 _8782_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_971_)
);

FILL FILL_3_BUFX2_insert545 (
);

FILL FILL_3_BUFX2_insert546 (
);

NAND2X1 _8362_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_752_)
);

FILL FILL_3_BUFX2_insert547 (
);

FILL SFILL104520x70050 (
);

FILL FILL_3_BUFX2_insert548 (
);

FILL SFILL43880x60050 (
);

FILL FILL_3_BUFX2_insert549 (
);

FILL FILL_4__13895_ (
);

FILL FILL_4__13475_ (
);

FILL FILL_3__12888_ (
);

FILL FILL_2__7635_ (
);

FILL FILL_3__12468_ (
);

FILL FILL_2__7215_ (
);

FILL FILL_3__12048_ (
);

FILL FILL_1__13082_ (
);

FILL FILL_6__13802_ (
);

FILL SFILL59080x31050 (
);

NAND2X1 _12780_ (
    .A(IRWrite_bF$buf7),
    .B(memoryOutData[28]),
    .Y(_3546_)
);

FILL FILL_0__12495_ (
);

FILL FILL_0__12075_ (
);

OAI21X1 _12360_ (
    .A(_3304_),
    .B(MemToReg_bF$buf4),
    .C(_3305_),
    .Y(\datapath_1.mux_wd3.dout [5])
);

FILL SFILL38920x16050 (
);

FILL FILL_4__8502_ (
);

FILL FILL_5__15687_ (
);

FILL FILL_2__12402_ (
);

FILL FILL_5__15267_ (
);

NAND2X1 _9987_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1571_)
);

DFFSR _9567_ (
    .Q(\datapath_1.regfile_1.regOut[21] [9]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf6),
    .S(vdd),
    .D(_1303_[9])
);

INVX1 _9147_ (
    .A(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_1153_)
);

FILL FILL_1__11815_ (
);

FILL FILL_2__15294_ (
);

FILL FILL_0__8822_ (
);

FILL FILL_0__10808_ (
);

FILL FILL_0__8402_ (
);

FILL FILL_1__14287_ (
);

FILL FILL_5__6845_ (
);

FILL FILL_0_BUFX2_insert670 (
);

FILL FILL_0_BUFX2_insert671 (
);

FILL FILL_4__15621_ (
);

FILL FILL_4__15201_ (
);

FILL FILL_0_BUFX2_insert672 (
);

FILL FILL_0_BUFX2_insert673 (
);

OAI22X1 _13985_ (
    .A(_4485_),
    .B(_3916_),
    .C(_3881_),
    .D(_4484_),
    .Y(_4486_)
);

FILL FILL_0_BUFX2_insert674 (
);

FILL FILL_3__9391_ (
);

FILL FILL_0_BUFX2_insert675 (
);

INVX1 _13565_ (
    .A(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_4075_)
);

INVX1 _13145_ (
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3728_)
);

FILL FILL_0_BUFX2_insert676 (
);

FILL FILL_0_BUFX2_insert677 (
);

FILL FILL_3__14614_ (
);

FILL FILL_0_BUFX2_insert678 (
);

FILL SFILL28920x59050 (
);

FILL FILL_0_BUFX2_insert679 (
);

FILL SFILL3560x15050 (
);

FILL FILL_1__6837_ (
);

FILL SFILL104440x32050 (
);

FILL FILL_2__13607_ (
);

FILL FILL_0__14641_ (
);

FILL FILL_0__14221_ (
);

FILL FILL_5__11187_ (
);

FILL FILL_2__16079_ (
);

FILL FILL_3__7704_ (
);

FILL FILL_0__9607_ (
);

FILL SFILL64600x5050 (
);

FILL FILL_4__16406_ (
);

FILL SFILL49000x72050 (
);

FILL FILL_6__10507_ (
);

FILL FILL_4__11961_ (
);

FILL FILL_4__11541_ (
);

FILL FILL_4__11121_ (
);

FILL FILL_3__15819_ (
);

FILL FILL_1__16013_ (
);

FILL FILL_3__10954_ (
);

FILL FILL_3__10534_ (
);

FILL FILL_3__10114_ (
);

FILL SFILL94440x81050 (
);

FILL FILL_0__15846_ (
);

OAI22X1 _15711_ (
    .A(_6173_),
    .B(_5548__bF$buf0),
    .C(_5489__bF$buf1),
    .D(_6174_),
    .Y(_6175_)
);

FILL FILL_0__15426_ (
);

FILL FILL_0__15006_ (
);

FILL FILL_0__10981_ (
);

FILL FILL_2__8593_ (
);

FILL FILL_0__10561_ (
);

FILL FILL_0__10141_ (
);

FILL FILL_4__8099_ (
);

FILL FILL_3__8909_ (
);

FILL FILL_5__13753_ (
);

FILL FILL_5__13333_ (
);

FILL FILL_6__6914_ (
);

NAND2X1 _7633_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_388_)
);

NAND2X1 _7213_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_169_)
);

FILL FILL_4__9880_ (
);

FILL FILL_4__12746_ (
);

FILL FILL_4__9040_ (
);

FILL FILL_2__13780_ (
);

FILL FILL_4__12326_ (
);

FILL FILL_2__13360_ (
);

FILL FILL_2__6906_ (
);

FILL FILL_3__11739_ (
);

FILL FILL_1__12773_ (
);

FILL FILL_3__11319_ (
);

FILL FILL_1__12353_ (
);

FILL FILL_2__9798_ (
);

FILL FILL_0__9780_ (
);

FILL FILL_0__9360_ (
);

FILL FILL_2__9378_ (
);

FILL FILL_0__11766_ (
);

FILL FILL_0__11346_ (
);

NAND3X1 _11631_ (
    .A(_2462__bF$buf0),
    .B(_2728_),
    .C(_2734_),
    .Y(_2735_)
);

OAI21X1 _11211_ (
    .A(_2317_),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .C(_2329_),
    .Y(_2330_)
);

FILL FILL_5__14958_ (
);

FILL FILL_3__15992_ (
);

FILL FILL_5__14538_ (
);

FILL FILL_3__15572_ (
);

FILL FILL_5__14118_ (
);

FILL FILL_3__15152_ (
);

NAND2X1 _8838_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_988_)
);

DFFSR _8418_ (
    .Q(\datapath_1.regfile_1.regOut[12] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_718_[12])
);

FILL FILL_1__7375_ (
);

FILL FILL_2__14985_ (
);

FILL FILL_2__14565_ (
);

FILL FILL_2__14145_ (
);

FILL SFILL39000x70050 (
);

FILL SFILL94360x43050 (
);

FILL FILL_1__13978_ (
);

FILL FILL_1__13558_ (
);

FILL FILL_1__13138_ (
);

NAND2X1 _12836_ (
    .A(vdd),
    .B(\datapath_1.rd1 [4]),
    .Y(_3563_)
);

FILL FILL_3__8242_ (
);

NAND2X1 _12416_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [24]),
    .Y(_3343_)
);

FILL FILL_5__8588_ (
);

FILL FILL_0__13912_ (
);

FILL FILL_3__16357_ (
);

FILL FILL_5__10878_ (
);

FILL FILL_5__10038_ (
);

FILL FILL_3__11492_ (
);

FILL FILL_3__11072_ (
);

FILL FILL_0__16384_ (
);

FILL SFILL18840x19050 (
);

FILL FILL_2__10065_ (
);

FILL FILL_1__9941_ (
);

FILL FILL_1__9521_ (
);

FILL FILL_1__9101_ (
);

FILL FILL_3__9867_ (
);

FILL FILL_4__10812_ (
);

FILL FILL_3__9027_ (
);

FILL FILL_5__14291_ (
);

NAND2X1 _8591_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_864_)
);

FILL FILL_1__15704_ (
);

DFFSR _8171_ (
    .Q(\datapath_1.regfile_1.regOut[10] [21]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf97),
    .S(vdd),
    .D(_588_[21])
);

FILL FILL_4__13284_ (
);

FILL SFILL8760x60050 (
);

FILL FILL111880x6050 (
);

FILL FILL_2__7864_ (
);

FILL FILL_3__12697_ (
);

FILL FILL_2__7444_ (
);

FILL FILL_3__12277_ (
);

FILL SFILL114600x60050 (
);

FILL FILL_5__12604_ (
);

FILL SFILL53960x50050 (
);

FILL SFILL84360x41050 (
);

OAI21X1 _6904_ (
    .A(_66_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .C(_67_),
    .Y(_3_[0])
);

FILL FILL_4__8731_ (
);

FILL FILL_4__8311_ (
);

FILL FILL_2__12631_ (
);

FILL FILL_5__15496_ (
);

FILL FILL_5__15076_ (
);

FILL FILL_2__12211_ (
);

INVX1 _9796_ (
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .Y(_1484_)
);

INVX1 _9376_ (
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_1265_)
);

FILL FILL_6__8237_ (
);

FILL FILL_4__14489_ (
);

FILL FILL_1__11624_ (
);

FILL FILL_4__14069_ (
);

FILL FILL_1__11204_ (
);

FILL FILL_0__8631_ (
);

FILL FILL_2__8649_ (
);

FILL SFILL114520x67050 (
);

FILL FILL_2__8229_ (
);

INVX1 _10902_ (
    .A(\control_1.reg_state.dout [0]),
    .Y(_2050_)
);

FILL FILL_0__10617_ (
);

FILL FILL_0__8211_ (
);

FILL FILL_1__14096_ (
);

FILL FILL_4__15850_ (
);

FILL FILL_4__15430_ (
);

FILL FILL_4__15010_ (
);

INVX1 _13794_ (
    .A(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_4299_)
);

FILL FILL_0__13089_ (
);

AOI22X1 _13374_ (
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .B(_3885_),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_3886_)
);

FILL FILL_5__13809_ (
);

FILL FILL_3__14843_ (
);

FILL FILL_3__14423_ (
);

FILL FILL_3__14003_ (
);

FILL FILL_4__9936_ (
);

FILL FILL_4__9516_ (
);

FILL SFILL69080x28050 (
);

FILL FILL_2__13836_ (
);

FILL FILL_0__14870_ (
);

FILL FILL_2__13416_ (
);

FILL FILL_0__14450_ (
);

FILL FILL_0__14030_ (
);

FILL FILL_1__12829_ (
);

FILL FILL_1__12409_ (
);

CLKBUF1 CLKBUF1_insert220 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert221 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert222 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert223 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf1)
);

FILL FILL_3__7933_ (
);

CLKBUF1 CLKBUF1_insert224 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf0)
);

FILL FILL_0__9416_ (
);

FILL FILL_5__7859_ (
);

FILL FILL_5__7439_ (
);

FILL SFILL114520x22050 (
);

FILL FILL_4__16215_ (
);

INVX4 _14999_ (
    .A(_5478__bF$buf3),
    .Y(_5479_)
);

NOR2X1 _14579_ (
    .A(_5067_),
    .B(_5064_),
    .Y(_5068_)
);

FILL FILL_4__11770_ (
);

INVX1 _14159_ (
    .A(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_4657_)
);

FILL FILL_4__11350_ (
);

FILL SFILL3720x41050 (
);

FILL FILL_3__15628_ (
);

FILL FILL_3__15208_ (
);

FILL FILL_1__16242_ (
);

FILL FILL_3__10763_ (
);

FILL FILL_0__15655_ (
);

NOR2X1 _15940_ (
    .A(_5004_),
    .B(_5539__bF$buf0),
    .Y(_6398_)
);

FILL FILL_0__15235_ (
);

OAI21X1 _15520_ (
    .A(_4510_),
    .B(_5535__bF$buf4),
    .C(_5988_),
    .Y(_5989_)
);

INVX4 _15100_ (
    .A(_5548__bF$buf3),
    .Y(_5579_)
);

FILL FILL_0__10790_ (
);

FILL FILL_0__10370_ (
);

FILL FILL_3__8718_ (
);

FILL FILL_5__13982_ (
);

FILL FILL_5__13562_ (
);

FILL FILL_5__13142_ (
);

NAND2X1 _7862_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_500_)
);

NAND2X1 _7442_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_281_)
);

FILL SFILL104520x65050 (
);

DFFSR _7022_ (
    .Q(\datapath_1.regfile_1.regOut[1] [24]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_3_[24])
);

FILL FILL_4_BUFX2_insert900 (
);

FILL SFILL43880x55050 (
);

FILL FILL_4_BUFX2_insert901 (
);

FILL FILL_4__12975_ (
);

FILL FILL_4_BUFX2_insert902 (
);

FILL FILL_4_BUFX2_insert903 (
);

FILL FILL_4_BUFX2_insert904 (
);

FILL FILL_4__12135_ (
);

FILL FILL_4_BUFX2_insert905 (
);

FILL FILL_4_BUFX2_insert906 (
);

FILL FILL_4_BUFX2_insert907 (
);

NAND2X1 _10499_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1831_)
);

FILL FILL_4_BUFX2_insert908 (
);

DFFSR _10079_ (
    .Q(\datapath_1.regfile_1.regOut[25] [9]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_1563_[9])
);

FILL FILL_4_BUFX2_insert909 (
);

FILL FILL_3__11968_ (
);

FILL FILL_3__11548_ (
);

FILL SFILL59000x69050 (
);

FILL FILL_1__12582_ (
);

FILL FILL_3__11128_ (
);

FILL FILL_1__12162_ (
);

INVX1 _16305_ (
    .A(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_6754_)
);

FILL SFILL59080x26050 (
);

FILL FILL_0__11995_ (
);

NAND2X1 _11860_ (
    .A(_2687_),
    .B(_2718_),
    .Y(_2947_)
);

FILL FILL_0__11575_ (
);

INVX1 _11440_ (
    .A(_2449_),
    .Y(_2556_)
);

FILL FILL_0__11155_ (
);

NOR2X1 _11020_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2139_)
);

FILL FILL_5__7192_ (
);

FILL FILL_2__11902_ (
);

FILL FILL_5__14767_ (
);

FILL FILL_5__14347_ (
);

FILL FILL_3__15381_ (
);

FILL FILL_6__7508_ (
);

INVX1 _8647_ (
    .A(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_901_)
);

INVX1 _8227_ (
    .A(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_682_)
);

FILL FILL_1__7184_ (
);

FILL FILL_2__14794_ (
);

FILL FILL_2__14374_ (
);

FILL SFILL104520x20050 (
);

FILL SFILL43880x10050 (
);

FILL FILL_1__13787_ (
);

FILL FILL_1__13367_ (
);

FILL FILL_4__14701_ (
);

FILL SFILL59000x24050 (
);

FILL FILL_3__8891_ (
);

FILL SFILL49080x69050 (
);

FILL FILL_3__8471_ (
);

INVX1 _12645_ (
    .A(\datapath_1.Data [26]),
    .Y(_3476_)
);

AOI22X1 _12225_ (
    .A(_2_[2]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf3),
    .D(\aluControl_1.inst [0]),
    .Y(_3208_)
);

FILL FILL_5__8397_ (
);

FILL FILL_0__13721_ (
);

FILL FILL_0__13301_ (
);

FILL FILL_3__16166_ (
);

FILL FILL_5__10687_ (
);

FILL FILL_1__8389_ (
);

FILL FILL_5__10267_ (
);

FILL FILL_2__15999_ (
);

FILL FILL_0_BUFX2_insert1020 (
);

FILL FILL_0_BUFX2_insert1021 (
);

FILL FILL_2__15579_ (
);

FILL FILL_0_BUFX2_insert1022 (
);

FILL FILL_2__15159_ (
);

FILL FILL_0__16193_ (
);

FILL FILL_0_BUFX2_insert1023 (
);

FILL SFILL33880x53050 (
);

FILL FILL_0_BUFX2_insert1024 (
);

FILL FILL_0_BUFX2_insert1025 (
);

FILL FILL_2__10294_ (
);

FILL FILL_0_BUFX2_insert1026 (
);

FILL FILL_0_BUFX2_insert1027 (
);

FILL SFILL104040x13050 (
);

FILL FILL_0_BUFX2_insert1028 (
);

FILL FILL_0_BUFX2_insert1029 (
);

FILL FILL_1__9750_ (
);

FILL FILL_4__15906_ (
);

FILL SFILL49000x67050 (
);

FILL FILL_3__9676_ (
);

FILL FILL_2__16100_ (
);

FILL FILL_3_BUFX2_insert920 (
);

FILL FILL_3__9256_ (
);

FILL FILL_3_BUFX2_insert921 (
);

FILL FILL_3_BUFX2_insert922 (
);

FILL FILL_4__10621_ (
);

FILL FILL_3_BUFX2_insert923 (
);

FILL FILL_3_BUFX2_insert924 (
);

FILL FILL_1__15933_ (
);

FILL FILL_3_BUFX2_insert925 (
);

FILL FILL_1__15513_ (
);

FILL FILL_3_BUFX2_insert926 (
);

FILL FILL_3_BUFX2_insert927 (
);

FILL FILL_3_BUFX2_insert928 (
);

FILL FILL_6__12479_ (
);

FILL FILL_3_BUFX2_insert929 (
);

FILL SFILL94440x76050 (
);

FILL FILL_4__13093_ (
);

FILL FILL_0__14926_ (
);

FILL FILL_0__14506_ (
);

FILL FILL_2__7673_ (
);

FILL FILL_2__7253_ (
);

FILL FILL_3__12086_ (
);

FILL FILL_4__7599_ (
);

FILL FILL_4__7179_ (
);

FILL FILL_2__11499_ (
);

FILL FILL_2__11079_ (
);

FILL FILL_5__12833_ (
);

FILL FILL_5__12413_ (
);

FILL FILL_4__8960_ (
);

FILL FILL_4__8120_ (
);

FILL FILL_4__11826_ (
);

FILL FILL_2__12860_ (
);

FILL FILL_4__11406_ (
);

FILL FILL_2__12440_ (
);

FILL SFILL18120x69050 (
);

FILL FILL_0__7499_ (
);

FILL FILL_2__12020_ (
);

FILL SFILL49000x22050 (
);

FILL FILL_0__7079_ (
);

FILL SFILL39080x67050 (
);

DFFSR _9185_ (
    .Q(\datapath_1.regfile_1.regOut[18] [11]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf69),
    .S(vdd),
    .D(_1108_[11])
);

FILL FILL_3__10819_ (
);

FILL FILL_1__11853_ (
);

FILL FILL_4__14298_ (
);

FILL FILL_1__11433_ (
);

FILL FILL_1__11013_ (
);

FILL FILL_0__8860_ (
);

FILL FILL_2__8878_ (
);

FILL FILL_2__8458_ (
);

FILL FILL_0__8440_ (
);

FILL FILL_0__8020_ (
);

FILL FILL_0__10426_ (
);

DFFSR _10711_ (
    .Q(\datapath_1.regfile_1.regOut[30] [1]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_1888_[1])
);

FILL FILL_0__10006_ (
);

FILL FILL_5__6883_ (
);

DFFSR _13183_ (
    .Q(\datapath_1.mux_iord.din0 [8]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3685_[8])
);

FILL FILL_5__13618_ (
);

FILL FILL_3__14652_ (
);

FILL SFILL54280x42050 (
);

DFFSR _7918_ (
    .Q(\datapath_1.regfile_1.regOut[8] [24]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_458_[24])
);

FILL FILL_3__14232_ (
);

FILL FILL_1__6875_ (
);

FILL FILL_4__9745_ (
);

FILL FILL_2__13645_ (
);

FILL FILL_2__13225_ (
);

FILL SFILL39000x65050 (
);

FILL SFILL94360x38050 (
);

FILL FILL_1__12638_ (
);

FILL FILL_1__12218_ (
);

FILL FILL_3__7742_ (
);

FILL FILL_0__9645_ (
);

FILL SFILL84440x74050 (
);

FILL FILL_0__9225_ (
);

OAI21X1 _11916_ (
    .A(_2984_),
    .B(IorD_bF$buf4),
    .C(_2985_),
    .Y(_1_[9])
);

FILL FILL_3__7322_ (
);

FILL SFILL79160x18050 (
);

FILL FILL_5__7248_ (
);

FILL FILL_4__16024_ (
);

AOI22X1 _14388_ (
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .B(_4135_),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_4881_)
);

FILL FILL_3__15857_ (
);

FILL FILL_3__15437_ (
);

FILL FILL_3__15017_ (
);

FILL FILL_1__16051_ (
);

FILL FILL_3__10992_ (
);

FILL FILL_3__10572_ (
);

FILL FILL_3__10152_ (
);

FILL FILL_0__15884_ (
);

FILL FILL_6_BUFX2_insert434 (
);

FILL FILL_0__15464_ (
);

FILL FILL_0__15044_ (
);

FILL FILL111800x22050 (
);

FILL FILL_6_BUFX2_insert439 (
);

FILL FILL_1__8601_ (
);

FILL SFILL53880x4050 (
);

FILL FILL_3__8527_ (
);

FILL FILL_3__8107_ (
);

FILL FILL_5__13791_ (
);

FILL FILL_5__13371_ (
);

NAND2X1 _7671_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .Y(_457_)
);

INVX1 _7251_ (
    .A(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_194_)
);

FILL FILL_4__12784_ (
);

FILL FILL_4__12364_ (
);

FILL FILL_2__6944_ (
);

FILL FILL_3__11777_ (
);

FILL FILL_3__11357_ (
);

FILL FILL_1__12391_ (
);

FILL FILL_0__16249_ (
);

INVX1 _16114_ (
    .A(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_6568_)
);

FILL FILL_0__11384_ (
);

FILL SFILL53960x45050 (
);

FILL FILL_1__9806_ (
);

FILL FILL_6__15163_ (
);

FILL FILL_4__7811_ (
);

FILL FILL_5__14996_ (
);

FILL FILL_5__14576_ (
);

FILL FILL_2__11711_ (
);

FILL FILL_5__14156_ (
);

FILL FILL_3__15190_ (
);

INVX1 _8876_ (
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_1013_)
);

INVX1 _8456_ (
    .A(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_794_)
);

FILL FILL_6__7317_ (
);

DFFSR _8036_ (
    .Q(\datapath_1.regfile_1.regOut[9] [14]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_523_[14])
);

FILL FILL_4__13989_ (
);

FILL FILL_4__13569_ (
);

FILL FILL_1__10704_ (
);

FILL SFILL53560x31050 (
);

FILL FILL_4__13149_ (
);

FILL FILL_2__14183_ (
);

FILL FILL_2__7729_ (
);

FILL FILL_0__7711_ (
);

FILL SFILL8760x10050 (
);

FILL FILL_2__7309_ (
);

FILL FILL_1__13596_ (
);

FILL FILL_4__14930_ (
);

FILL FILL_4__14510_ (
);

FILL FILL_0__12589_ (
);

INVX1 _12874_ (
    .A(\datapath_1.a [17]),
    .Y(_3588_)
);

INVX1 _12454_ (
    .A(ALUOut[5]),
    .Y(_3369_)
);

FILL FILL_0__12169_ (
);

NAND3X1 _12034_ (
    .A(_3069_),
    .B(_3070_),
    .C(_3071_),
    .Y(\datapath_1.mux_pcsrc.dout [11])
);

FILL FILL_3__13923_ (
);

FILL FILL_3__13503_ (
);

FILL SFILL114600x10050 (
);

FILL FILL_5_BUFX2_insert450 (
);

FILL FILL_6__11083_ (
);

FILL FILL_5_BUFX2_insert451 (
);

FILL FILL_2__12916_ (
);

FILL FILL_5_BUFX2_insert452 (
);

FILL FILL_0__13950_ (
);

FILL FILL_3__16395_ (
);

FILL FILL_5_BUFX2_insert453 (
);

FILL FILL_0__13530_ (
);

FILL FILL_5_BUFX2_insert454 (
);

FILL FILL_0__13110_ (
);

FILL FILL_5_BUFX2_insert455 (
);

FILL FILL_5__10496_ (
);

FILL FILL_5_BUFX2_insert456 (
);

FILL FILL_5_BUFX2_insert457 (
);

FILL FILL_1__8198_ (
);

FILL FILL_1__11909_ (
);

FILL FILL_5_BUFX2_insert458 (
);

FILL FILL_5_BUFX2_insert459 (
);

FILL FILL_2__15388_ (
);

FILL FILL_5__16302_ (
);

FILL FILL_0__8916_ (
);

FILL FILL_5__6939_ (
);

FILL SFILL114520x17050 (
);

FILL FILL_4__15715_ (
);

FILL FILL_3__9485_ (
);

INVX1 _13659_ (
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_4167_)
);

NOR2X1 _13239_ (
    .A(_3759_),
    .B(_3753_),
    .Y(_3782_)
);

FILL FILL_4__10430_ (
);

FILL SFILL3720x36050 (
);

FILL FILL_4__10010_ (
);

FILL FILL_3__14708_ (
);

FILL FILL_1__15742_ (
);

FILL FILL_1__15322_ (
);

FILL SFILL43960x43050 (
);

FILL FILL_0__14735_ (
);

OAI22X1 _14600_ (
    .A(_5086_),
    .B(_3884__bF$buf1),
    .C(_3881_),
    .D(_5087_),
    .Y(_5088_)
);

FILL FILL_0__14315_ (
);

FILL FILL_2__7482_ (
);

FILL FILL_2__7062_ (
);

FILL SFILL49560x8050 (
);

FILL FILL_5__12642_ (
);

FILL FILL_5__12222_ (
);

NAND2X1 _6942_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_29_)
);

FILL FILL_2_BUFX2_insert580 (
);

FILL FILL_2_BUFX2_insert581 (
);

FILL FILL_2_BUFX2_insert582 (
);

FILL FILL_2_BUFX2_insert583 (
);

FILL FILL_2_BUFX2_insert584 (
);

FILL FILL_4__11635_ (
);

FILL FILL_2_BUFX2_insert585 (
);

FILL FILL_4__11215_ (
);

FILL FILL_2_BUFX2_insert586 (
);

FILL SFILL23880x3050 (
);

FILL FILL_2_BUFX2_insert587 (
);

FILL FILL_2_BUFX2_insert588 (
);

FILL FILL_2_BUFX2_insert589 (
);

FILL FILL_1__16107_ (
);

FILL FILL_3__10628_ (
);

FILL FILL_1__11662_ (
);

FILL FILL_1__11242_ (
);

OAI22X1 _15805_ (
    .A(_6266_),
    .B(_5548__bF$buf2),
    .C(_5534__bF$buf4),
    .D(_4831_),
    .Y(_6267_)
);

FILL FILL112280x54050 (
);

NAND2X1 _10940_ (
    .A(\control_1.op [5]),
    .B(_2073_),
    .Y(_2074_)
);

FILL FILL_2__8267_ (
);

FILL FILL_0__10655_ (
);

NAND2X1 _10520_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1845_)
);

FILL FILL_0__10235_ (
);

DFFSR _10100_ (
    .Q(\datapath_1.regfile_1.regOut[25] [30]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1563_[30])
);

FILL FILL_5__13847_ (
);

FILL FILL_3__14881_ (
);

FILL FILL_5__13427_ (
);

FILL FILL_3__14461_ (
);

FILL FILL_5__13007_ (
);

FILL FILL_3__14041_ (
);

INVX1 _7727_ (
    .A(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_430_)
);

INVX1 _7307_ (
    .A(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_211_)
);

FILL FILL_4__9974_ (
);

FILL FILL_4__9554_ (
);

FILL FILL_4__9134_ (
);

FILL FILL_2__13874_ (
);

FILL SFILL104520x15050 (
);

FILL FILL_2__13454_ (
);

FILL FILL_2__13034_ (
);

FILL FILL_1__12867_ (
);

FILL FILL_1__12447_ (
);

FILL FILL_1__12027_ (
);

FILL SFILL59000x19050 (
);

FILL FILL_3__7971_ (
);

FILL FILL_0__9874_ (
);

FILL FILL_3__7551_ (
);

FILL FILL_0__9034_ (
);

AOI21X1 _11725_ (
    .A(_2172_),
    .B(_2811_),
    .C(_2458_),
    .Y(_2823_)
);

INVX2 _11305_ (
    .A(_2423_),
    .Y(_2424_)
);

FILL FILL_6__15639_ (
);

FILL FILL_5__7477_ (
);

FILL FILL_6__15219_ (
);

FILL FILL_4__16253_ (
);

FILL FILL_5__7057_ (
);

AOI22X1 _14197_ (
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .B(_4135_),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_4694_)
);

FILL FILL_3__15666_ (
);

FILL FILL_3__15246_ (
);

FILL FILL_1__16280_ (
);

FILL FILL_1__7889_ (
);

FILL FILL_1__7469_ (
);

FILL FILL_3__10381_ (
);

FILL FILL_1__7049_ (
);

FILL FILL_2__14659_ (
);

FILL FILL_2__14239_ (
);

FILL FILL_0__15693_ (
);

FILL SFILL33880x48050 (
);

FILL FILL_0__15273_ (
);

FILL FILL_1__8830_ (
);

FILL FILL_2__15600_ (
);

FILL FILL_3__8756_ (
);

FILL FILL_3__8336_ (
);

FILL SFILL98840x72050 (
);

INVX1 _7480_ (
    .A(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_306_)
);

INVX1 _7060_ (
    .A(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_87_)
);

FILL FILL_4__12593_ (
);

FILL FILL_6__11139_ (
);

FILL FILL_4__12173_ (
);

FILL FILL_5__9623_ (
);

FILL FILL_3__11586_ (
);

FILL FILL_3__11166_ (
);

FILL FILL_6__12500_ (
);

NAND2X1 _16343_ (
    .A(gnd),
    .B(gnd),
    .Y(_6783_)
);

FILL FILL_0__16058_ (
);

FILL FILL_2__10999_ (
);

FILL FILL_2__10579_ (
);

FILL FILL_2__10159_ (
);

FILL FILL_0__11193_ (
);

FILL FILL_5__11913_ (
);

FILL FILL_1__9615_ (
);

FILL FILL_4__7620_ (
);

FILL FILL_4__10906_ (
);

FILL FILL_4__7200_ (
);

FILL FILL_2__11940_ (
);

FILL FILL_5__14385_ (
);

FILL FILL_2__11520_ (
);

FILL SFILL49000x17050 (
);

FILL FILL_2__11100_ (
);

DFFSR _8685_ (
    .Q(\datapath_1.regfile_1.regOut[14] [23]),
    .CLK(clk_bF$buf82),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_848_[23])
);

OAI21X1 _8265_ (
    .A(_706_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_707_),
    .Y(_653_[27])
);

FILL FILL_1__10933_ (
);

FILL FILL_4__13798_ (
);

FILL FILL_4__13378_ (
);

FILL FILL_1__10513_ (
);

FILL SFILL94440x26050 (
);

FILL FILL_0__7940_ (
);

FILL FILL_2__7958_ (
);

BUFX2 BUFX2_insert270 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf6 )
);

FILL FILL_0__7100_ (
);

FILL FILL_2__7118_ (
);

BUFX2 BUFX2_insert271 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf5 )
);

BUFX2 BUFX2_insert272 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf4 )
);

BUFX2 BUFX2_insert273 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf3 )
);

FILL SFILL18840x9050 (
);

BUFX2 BUFX2_insert274 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf2 )
);

FILL FILL_6__13705_ (
);

BUFX2 BUFX2_insert275 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf1 )
);

BUFX2 BUFX2_insert276 (
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf0 )
);

BUFX2 BUFX2_insert277 (
    .A(_3931_),
    .Y(_3931__bF$buf3)
);

BUFX2 BUFX2_insert278 (
    .A(_3931_),
    .Y(_3931__bF$buf2)
);

FILL FILL_0__12398_ (
);

DFFSR _12683_ (
    .Q(\datapath_1.Data [20]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3425_[20])
);

BUFX2 BUFX2_insert279 (
    .A(_3931_),
    .Y(_3931__bF$buf1)
);

NAND3X1 _12263_ (
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3236_)
);

FILL FILL_3__13732_ (
);

FILL FILL_3__13312_ (
);

FILL FILL_4__8825_ (
);

FILL FILL_4__8405_ (
);

FILL FILL_2__12725_ (
);

FILL FILL_2__12305_ (
);

FILL FILL_1__11718_ (
);

FILL FILL_2__15197_ (
);

FILL FILL_5__16111_ (
);

FILL FILL_0__8725_ (
);

FILL FILL_4__15944_ (
);

FILL FILL_4__15524_ (
);

FILL FILL_4__15104_ (
);

FILL FILL_3__9294_ (
);

INVX1 _13888_ (
    .A(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_4391_)
);

INVX1 _13468_ (
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_3980_)
);

DFFSR _13048_ (
    .Q(_2_[1]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_3620_[1])
);

FILL FILL_3__14937_ (
);

FILL FILL_1__15971_ (
);

FILL FILL_3__14517_ (
);

FILL FILL_1__15551_ (
);

FILL FILL_1__15131_ (
);

FILL FILL_0__14964_ (
);

FILL FILL_0__14544_ (
);

FILL FILL_0__14124_ (
);

FILL FILL_2__7291_ (
);

FILL FILL_3__7607_ (
);

FILL FILL_5__12871_ (
);

FILL FILL_5__12451_ (
);

FILL FILL_5__12031_ (
);

FILL FILL_4__16309_ (
);

FILL FILL_4__11864_ (
);

FILL FILL_4__11444_ (
);

FILL FILL_4__11024_ (
);

FILL FILL_1__16336_ (
);

FILL FILL_3__10437_ (
);

FILL FILL_1__11891_ (
);

FILL FILL_3__10017_ (
);

FILL FILL_1__11471_ (
);

FILL FILL_1__11051_ (
);

FILL FILL_0__15749_ (
);

FILL SFILL84040x10050 (
);

FILL FILL_0__15329_ (
);

OAI22X1 _15614_ (
    .A(_5569_),
    .B(_6078_),
    .C(_5523_),
    .D(_6079_),
    .Y(_6080_)
);

FILL FILL_0__10884_ (
);

FILL FILL_2__8496_ (
);

FILL FILL_2__8076_ (
);

FILL FILL_0__10044_ (
);

FILL FILL_5__13656_ (
);

FILL FILL_5__13236_ (
);

FILL FILL_3__14690_ (
);

FILL FILL_3__14270_ (
);

INVX1 _7956_ (
    .A(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_542_)
);

DFFSR _7536_ (
    .Q(\datapath_1.regfile_1.regOut[5] [26]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_263_[26])
);

OAI21X1 _7116_ (
    .A(_123_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .C(_124_),
    .Y(_68_[28])
);

FILL FILL_4__9783_ (
);

FILL FILL_4__9363_ (
);

FILL FILL_4__12649_ (
);

FILL FILL_2__13683_ (
);

FILL FILL_4__12229_ (
);

FILL FILL_2__13263_ (
);

FILL FILL_1__12256_ (
);

FILL FILL_0__9683_ (
);

FILL FILL_3__7360_ (
);

NAND2X1 _11954_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[22]),
    .Y(_3011_)
);

FILL FILL_0__9263_ (
);

FILL FILL_0__11669_ (
);

FILL FILL_0__11249_ (
);

OAI21X1 _11534_ (
    .A(_2644_),
    .B(_2431_),
    .C(_2220_),
    .Y(_2645_)
);

INVX1 _11114_ (
    .A(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2233_)
);

FILL SFILL74840x36050 (
);

FILL FILL_5__7286_ (
);

FILL FILL_4__16062_ (
);

FILL FILL_3__15895_ (
);

FILL FILL_0__12610_ (
);

FILL FILL_3__15475_ (
);

FILL FILL_3__15055_ (
);

FILL FILL_1__7698_ (
);

FILL FILL_3__10190_ (
);

FILL FILL_2__14888_ (
);

FILL FILL_6_BUFX2_insert812 (
);

FILL FILL_2__14468_ (
);

FILL FILL_2__14048_ (
);

FILL FILL_0__15082_ (
);

FILL FILL_5__15802_ (
);

FILL FILL_6_BUFX2_insert817 (
);

FILL FILL_3__8985_ (
);

OAI21X1 _12739_ (
    .A(_3517_),
    .B(IRWrite_bF$buf6),
    .C(_3518_),
    .Y(_3490_[14])
);

FILL FILL_3__8145_ (
);

NAND3X1 _12319_ (
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3278_)
);

FILL FILL_1__14822_ (
);

FILL FILL_1__14402_ (
);

FILL SFILL43960x38050 (
);

FILL SFILL74360x29050 (
);

FILL FILL_0__13815_ (
);

FILL FILL_2__6982_ (
);

FILL FILL_5__9852_ (
);

FILL FILL_3__11395_ (
);

FILL FILL_5__9012_ (
);

FILL FILL_0__16287_ (
);

NOR2X1 _16152_ (
    .A(_6602_),
    .B(_6604_),
    .Y(_6605_)
);

FILL FILL112360x42050 (
);

FILL FILL_2__10388_ (
);

FILL FILL_5__11722_ (
);

FILL FILL_1__9424_ (
);

FILL FILL_5__11302_ (
);

FILL FILL_1__9004_ (
);

FILL SFILL64040x51050 (
);

FILL FILL_5__14194_ (
);

OAI21X1 _8494_ (
    .A(_818_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_819_),
    .Y(_783_[18])
);

FILL FILL_1__15607_ (
);

OAI21X1 _8074_ (
    .A(_599_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .C(_600_),
    .Y(_588_[6])
);

FILL FILL_1__10742_ (
);

FILL FILL_1__10322_ (
);

FILL FILL112280x49050 (
);

FILL FILL_2__7347_ (
);

OAI21X1 _12492_ (
    .A(_3393_),
    .B(vdd),
    .C(_3394_),
    .Y(_3360_[17])
);

NAND3X1 _12072_ (
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [21]),
    .C(_3034__bF$buf2),
    .Y(_3100_)
);

FILL FILL_5__12507_ (
);

FILL FILL_3__13961_ (
);

FILL FILL_3__13541_ (
);

FILL FILL_3__13121_ (
);

FILL FILL_4__8634_ (
);

FILL FILL_5_BUFX2_insert830 (
);

FILL FILL_4__8214_ (
);

FILL FILL_5_BUFX2_insert831 (
);

FILL FILL_2__12954_ (
);

FILL FILL_5__15399_ (
);

FILL FILL_5_BUFX2_insert832 (
);

FILL FILL_2__12534_ (
);

FILL FILL_2__12114_ (
);

FILL FILL_5_BUFX2_insert833 (
);

FILL FILL_5_BUFX2_insert834 (
);

DFFSR _9699_ (
    .Q(\datapath_1.regfile_1.regOut[22] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_1368_[13])
);

NAND2X1 _9279_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1221_)
);

FILL FILL_5_BUFX2_insert835 (
);

FILL FILL_5_BUFX2_insert836 (
);

FILL FILL_5_BUFX2_insert837 (
);

FILL FILL_5_BUFX2_insert838 (
);

FILL FILL_1__11947_ (
);

FILL FILL_5_BUFX2_insert839 (
);

FILL FILL_1__11527_ (
);

FILL FILL_1__11107_ (
);

FILL FILL_5__16340_ (
);

FILL FILL_0__8954_ (
);

FILL FILL_6__9921_ (
);

INVX1 _10805_ (
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_1994_)
);

FILL FILL_0__8114_ (
);

FILL FILL_5__6977_ (
);

FILL FILL_4__15753_ (
);

FILL FILL_4__15333_ (
);

NOR2X1 _13697_ (
    .A(_4200_),
    .B(_4203_),
    .Y(_4204_)
);

NOR2X1 _13277_ (
    .A(_3797_),
    .B(_3804_),
    .Y(_3817_)
);

FILL FILL_2__9913_ (
);

FILL FILL_3__14746_ (
);

FILL FILL_1__15780_ (
);

FILL FILL_3__14326_ (
);

FILL FILL_1__15360_ (
);

FILL FILL_1__6969_ (
);

FILL FILL_4__9419_ (
);

FILL SFILL94520x59050 (
);

FILL FILL_2__13739_ (
);

FILL FILL_2__13319_ (
);

FILL FILL_0__14773_ (
);

FILL FILL_0__14353_ (
);

FILL FILL_0__9739_ (
);

FILL FILL_3__7836_ (
);

FILL FILL_3__7416_ (
);

FILL FILL_5__12260_ (
);

INVX1 _6980_ (
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_54_)
);

FILL FILL_2_BUFX2_insert960 (
);

FILL FILL_4__16118_ (
);

FILL FILL_2_BUFX2_insert961 (
);

FILL FILL_2_BUFX2_insert962 (
);

FILL FILL_2_BUFX2_insert963 (
);

FILL FILL_2_BUFX2_insert964 (
);

FILL FILL_4__11673_ (
);

FILL FILL_2_BUFX2_insert965 (
);

FILL FILL_4__11253_ (
);

FILL FILL_2_BUFX2_insert966 (
);

FILL FILL_2_BUFX2_insert967 (
);

FILL FILL_2_BUFX2_insert968 (
);

FILL FILL_2_BUFX2_insert969 (
);

FILL FILL_1__16145_ (
);

FILL FILL_5__8703_ (
);

FILL FILL_3__10666_ (
);

FILL FILL_3__10246_ (
);

FILL FILL_1__11280_ (
);

FILL FILL_0__15978_ (
);

FILL FILL_0__15558_ (
);

NOR2X1 _15843_ (
    .A(_6303_),
    .B(_6302_),
    .Y(_6304_)
);

OAI22X1 _15423_ (
    .A(_5530__bF$buf1),
    .B(_5893_),
    .C(_5532__bF$buf2),
    .D(_4391_),
    .Y(_5894_)
);

FILL FILL_0__15138_ (
);

NAND3X1 _15003_ (
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5465_),
    .C(_5476_),
    .Y(_5483_)
);

FILL FILL_0__10693_ (
);

FILL FILL_0__10273_ (
);

FILL FILL_6__14892_ (
);

FILL FILL_6__14472_ (
);

FILL FILL_5__13885_ (
);

FILL FILL_5__13465_ (
);

FILL FILL_5__13045_ (
);

OAI21X1 _7765_ (
    .A(_454_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_455_),
    .Y(_393_[31])
);

OAI21X1 _7345_ (
    .A(_235_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .C(_236_),
    .Y(_198_[19])
);

FILL FILL_4__9592_ (
);

FILL FILL_4__12878_ (
);

FILL FILL_4__9172_ (
);

FILL FILL_4__12458_ (
);

FILL FILL_4__12038_ (
);

FILL FILL_2__13492_ (
);

FILL FILL_5__9908_ (
);

FILL FILL_1__12485_ (
);

FILL FILL_1__12065_ (
);

OAI22X1 _16208_ (
    .A(_6658_),
    .B(_5469__bF$buf0),
    .C(_5472__bF$buf1),
    .D(_5323_),
    .Y(_6659_)
);

FILL FILL_0__11898_ (
);

FILL FILL_0__9492_ (
);

AOI21X1 _11763_ (
    .A(_2364_),
    .B(_2853_),
    .C(_2857_),
    .Y(_2858_)
);

FILL FILL_0__11478_ (
);

NOR2X1 _11343_ (
    .A(_2330_),
    .B(_2326_),
    .Y(_2461_)
);

FILL FILL_0__11058_ (
);

FILL FILL_5__7095_ (
);

FILL FILL_4__16291_ (
);

FILL FILL_2__11805_ (
);

FILL FILL_3__15284_ (
);

FILL FILL_1__7087_ (
);

FILL FILL_2__14697_ (
);

FILL FILL_2__14277_ (
);

FILL FILL_5__15611_ (
);

FILL FILL_0__7805_ (
);

OAI21X1 _9911_ (
    .A(_1539_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1540_),
    .Y(_1498_[21])
);

FILL FILL_4__14604_ (
);

FILL FILL_1_BUFX2_insert980 (
);

FILL FILL_1_BUFX2_insert981 (
);

FILL FILL_3__8374_ (
);

FILL FILL_1_BUFX2_insert982 (
);

OAI21X1 _12968_ (
    .A(_3629_),
    .B(vdd),
    .C(_3630_),
    .Y(_3620_[5])
);

FILL SFILL23800x39050 (
);

FILL FILL_1_BUFX2_insert983 (
);

DFFSR _12548_ (
    .Q(ALUOut[13]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[13])
);

NAND2X1 _12128_ (
    .A(ALUSrcA_bF$buf4),
    .B(\datapath_1.a [4]),
    .Y(_3139_)
);

FILL FILL_1_BUFX2_insert984 (
);

FILL FILL_1_BUFX2_insert985 (
);

FILL FILL_1_BUFX2_insert986 (
);

FILL FILL_1__14631_ (
);

FILL FILL_1_BUFX2_insert987 (
);

FILL FILL_1_BUFX2_insert988 (
);

FILL FILL_1__14211_ (
);

FILL FILL_1_BUFX2_insert989 (
);

FILL FILL_0__13624_ (
);

FILL FILL_3__16069_ (
);

FILL FILL_5__9661_ (
);

FILL FILL_5__9241_ (
);

FILL FILL_0__16096_ (
);

INVX1 _16381_ (
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_6808_)
);

FILL FILL_2__10197_ (
);

FILL FILL_5__11951_ (
);

FILL FILL_1__9653_ (
);

FILL FILL_5__11531_ (
);

FILL FILL_5__11111_ (
);

FILL FILL_1__9233_ (
);

FILL FILL_4__15809_ (
);

FILL FILL_3__9999_ (
);

FILL FILL_2__16003_ (
);

FILL FILL_4__10944_ (
);

FILL FILL_3__9159_ (
);

FILL FILL_4__10524_ (
);

FILL FILL_4__10104_ (
);

FILL FILL_1__15836_ (
);

FILL FILL_1__15416_ (
);

FILL FILL_1__10971_ (
);

FILL FILL_1__10551_ (
);

FILL FILL_1__10131_ (
);

FILL FILL_0__14829_ (
);

FILL FILL_0__14409_ (
);

FILL FILL_2__7996_ (
);

BUFX2 BUFX2_insert650 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf1)
);

FILL FILL_2__7576_ (
);

BUFX2 BUFX2_insert651 (
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf0)
);

FILL SFILL13400x68050 (
);

BUFX2 BUFX2_insert652 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf4 )
);

BUFX2 BUFX2_insert653 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf3 )
);

BUFX2 BUFX2_insert654 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf2 )
);

BUFX2 BUFX2_insert655 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf1 )
);

BUFX2 BUFX2_insert656 (
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf0 )
);

FILL SFILL74120x41050 (
);

BUFX2 BUFX2_insert657 (
    .A(_3037_),
    .Y(_3037__bF$buf4)
);

BUFX2 BUFX2_insert658 (
    .A(_3037_),
    .Y(_3037__bF$buf3)
);

BUFX2 BUFX2_insert659 (
    .A(_3037_),
    .Y(_3037__bF$buf2)
);

FILL FILL_5__12736_ (
);

FILL FILL_3__13770_ (
);

FILL FILL_5__12316_ (
);

FILL FILL_3__13350_ (
);

FILL FILL_4__8863_ (
);

FILL FILL_4__8443_ (
);

FILL FILL_4__11729_ (
);

FILL FILL_2__12763_ (
);

FILL FILL_4__11309_ (
);

FILL FILL_2__12343_ (
);

FILL FILL_6__8789_ (
);

NAND2X1 _9088_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1114_)
);

FILL SFILL13800x37050 (
);

FILL FILL_1__11756_ (
);

FILL FILL_1__11336_ (
);

FILL SFILL74040x48050 (
);

FILL FILL_0__8763_ (
);

FILL FILL_3__6860_ (
);

FILL FILL_0__8343_ (
);

FILL FILL_0__10749_ (
);

INVX1 _10614_ (
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .Y(_1951_)
);

FILL FILL_6__14948_ (
);

FILL FILL_4__15982_ (
);

FILL FILL_6__14528_ (
);

FILL FILL_4__15562_ (
);

FILL FILL_4__15142_ (
);

NAND2X1 _13086_ (
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [2]),
    .Y(_3689_)
);

FILL FILL_3__14975_ (
);

FILL FILL_2__9722_ (
);

FILL FILL_3__14555_ (
);

FILL FILL_3__14135_ (
);

FILL FILL_4_BUFX2_insert490 (
);

FILL FILL_4__9648_ (
);

FILL FILL_4_BUFX2_insert491 (
);

FILL FILL_4__9228_ (
);

FILL FILL_4_BUFX2_insert492 (
);

FILL FILL_4_BUFX2_insert493 (
);

FILL FILL_2__13968_ (
);

FILL FILL_4_BUFX2_insert494 (
);

FILL FILL_2__13548_ (
);

FILL FILL_0__14582_ (
);

FILL FILL_2__13128_ (
);

FILL FILL_4_BUFX2_insert495 (
);

FILL FILL_4_BUFX2_insert496 (
);

FILL FILL_0__14162_ (
);

FILL FILL_4_BUFX2_insert497 (
);

FILL FILL_4_BUFX2_insert498 (
);

FILL FILL_4_BUFX2_insert499 (
);

FILL FILL_0__9548_ (
);

FILL FILL_0__9128_ (
);

FILL FILL_3__7225_ (
);

AND2X2 _11819_ (
    .A(_2909_),
    .B(_2906_),
    .Y(_2910_)
);

FILL FILL_1__13902_ (
);

FILL FILL_4__16347_ (
);

FILL FILL_4__11482_ (
);

FILL FILL_4__11062_ (
);

FILL FILL_1__16374_ (
);

FILL FILL_3__10895_ (
);

FILL FILL_5__8512_ (
);

FILL FILL_3__10055_ (
);

FILL FILL_0__15787_ (
);

AOI22X1 _15652_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [15]),
    .C(\datapath_1.regfile_1.regOut[22] [15]),
    .D(_5650_),
    .Y(_6117_)
);

FILL FILL_0__15367_ (
);

INVX1 _15232_ (
    .A(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_5708_)
);

FILL FILL112360x37050 (
);

FILL FILL_5__10802_ (
);

FILL FILL_1__8504_ (
);

FILL SFILL64040x46050 (
);

FILL FILL_5__13694_ (
);

FILL FILL_5__13274_ (
);

OAI21X1 _7994_ (
    .A(_566_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_567_),
    .Y(_523_[22])
);

OAI21X1 _7574_ (
    .A(_347_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_348_),
    .Y(_328_[10])
);

DFFSR _7154_ (
    .Q(\datapath_1.regfile_1.regOut[2] [28]),
    .CLK(clk_bF$buf34),
    .R(rst_bF$buf96),
    .S(vdd),
    .D(_68_[28])
);

FILL FILL_4__12267_ (
);

FILL SFILL54120x82050 (
);

FILL FILL_2__6847_ (
);

FILL FILL_1__12294_ (
);

DFFSR _16437_ (
    .Q(\datapath_1.regfile_1.regOut[0] [20]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_6769_[20])
);

INVX1 _16017_ (
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_6473_)
);

NAND3X1 _11992_ (
    .A(PCSource_1_bF$buf4),
    .B(gnd),
    .C(_3034__bF$buf1),
    .Y(_3040_)
);

AOI21X1 _11572_ (
    .A(_2236_),
    .B(_2678_),
    .C(_2679_),
    .Y(_2680_)
);

FILL FILL_0__11287_ (
);

INVX1 _11152_ (
    .A(\datapath_1.alu_1.ALUInA [18]),
    .Y(_2271_)
);

FILL FILL_3__12621_ (
);

FILL FILL_6__15066_ (
);

FILL FILL_3__12201_ (
);

FILL FILL_4__7714_ (
);

FILL FILL_5__14899_ (
);

FILL FILL_5__14479_ (
);

FILL FILL_2__11614_ (
);

FILL FILL_5__14059_ (
);

NAND2X1 _8779_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_969_)
);

FILL FILL_3__15093_ (
);

FILL SFILL68760x23050 (
);

NAND2X1 _8359_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_750_)
);

FILL FILL_2__14086_ (
);

FILL FILL_5__15840_ (
);

FILL FILL_5__15420_ (
);

FILL FILL_0__7614_ (
);

FILL FILL_5__15000_ (
);

OAI21X1 _9720_ (
    .A(_1496_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1497_),
    .Y(_1433_[0])
);

FILL SFILL89240x50050 (
);

NAND2X1 _9300_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_1235_)
);

FILL FILL_1__13499_ (
);

FILL FILL_1__13079_ (
);

FILL FILL_4__14833_ (
);

FILL FILL_4__14413_ (
);

NAND2X1 _12777_ (
    .A(IRWrite_bF$buf7),
    .B(memoryOutData[27]),
    .Y(_3544_)
);

FILL FILL_3__8183_ (
);

OAI21X1 _12357_ (
    .A(_3302_),
    .B(MemToReg_bF$buf3),
    .C(_3303_),
    .Y(\datapath_1.mux_wd3.dout [4])
);

FILL FILL_3__13826_ (
);

FILL FILL_1__14860_ (
);

FILL FILL_3__13406_ (
);

FILL FILL_1__14440_ (
);

FILL FILL_1__14020_ (
);

FILL FILL_0__13853_ (
);

FILL FILL_0__13433_ (
);

FILL FILL_3__16298_ (
);

FILL FILL_0__13013_ (
);

FILL FILL_5__9890_ (
);

FILL FILL_5__10399_ (
);

FILL SFILL54040x44050 (
);

FILL FILL_5__9470_ (
);

NAND2X1 _16190_ (
    .A(_6641_),
    .B(_6636_),
    .Y(_6642_)
);

FILL FILL_5__16205_ (
);

FILL FILL_3__6916_ (
);

FILL FILL_1__9882_ (
);

FILL FILL_5__11760_ (
);

FILL FILL_1__9462_ (
);

FILL FILL_5__11340_ (
);

FILL FILL_1__9042_ (
);

FILL FILL_4__15618_ (
);

FILL FILL_2__16232_ (
);

FILL FILL_3__9388_ (
);

FILL FILL_4__10753_ (
);

FILL FILL_1__15645_ (
);

FILL FILL_1__15225_ (
);

FILL FILL_1__10780_ (
);

FILL FILL_1__10360_ (
);

FILL FILL_0__14638_ (
);

OAI22X1 _14923_ (
    .A(_3983__bF$buf1),
    .B(_5403_),
    .C(_3971__bF$buf0),
    .D(_5404_),
    .Y(_5405_)
);

FILL FILL_0__14218_ (
);

OAI22X1 _14503_ (
    .A(_3947__bF$buf1),
    .B(_4992_),
    .C(_3909_),
    .D(_4991_),
    .Y(_4993_)
);

FILL FILL_5__12965_ (
);

FILL FILL_5__12125_ (
);

BUFX2 _6845_ (
    .A(_1_[7]),
    .Y(memoryAddress[7])
);

FILL FILL_4__8252_ (
);

FILL FILL_4__11958_ (
);

FILL FILL_2__12992_ (
);

FILL FILL_4__11538_ (
);

FILL FILL_2__12572_ (
);

FILL FILL_4__11118_ (
);

FILL FILL_2__12152_ (
);

FILL FILL_1__11985_ (
);

FILL FILL111880x61050 (
);

FILL FILL_1__11565_ (
);

FILL FILL_1__11145_ (
);

NOR3X1 _15708_ (
    .A(_5515__bF$buf3),
    .B(_6171_),
    .C(_5521__bF$buf3),
    .Y(_6172_)
);

FILL FILL_0__8992_ (
);

FILL FILL_0__10978_ (
);

FILL FILL_0__8572_ (
);

FILL FILL_0__10558_ (
);

DFFSR _10843_ (
    .Q(\datapath_1.regfile_1.regOut[31] [5]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_1953_[5])
);

FILL FILL_0__10138_ (
);

OAI21X1 _10423_ (
    .A(_1799_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .C(_1800_),
    .Y(_1758_[21])
);

OAI21X1 _10003_ (
    .A(_1580_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1581_),
    .Y(_1563_[9])
);

FILL SFILL109400x74050 (
);

FILL FILL_4__15791_ (
);

FILL FILL_4__15371_ (
);

FILL FILL_2__9531_ (
);

FILL FILL_3__14784_ (
);

FILL FILL_2__9111_ (
);

FILL FILL_3__14364_ (
);

FILL FILL_4__9877_ (
);

FILL FILL_4__9037_ (
);

FILL FILL_2__13777_ (
);

FILL FILL_2__13357_ (
);

FILL SFILL8920x26050 (
);

FILL FILL_0__14391_ (
);

FILL FILL112120x7050 (
);

FILL FILL_0__9777_ (
);

FILL FILL_3__7874_ (
);

FILL FILL_0__9357_ (
);

FILL FILL_3__7454_ (
);

AOI21X1 _11628_ (
    .A(_2723_),
    .B(_2724_),
    .C(_2732_),
    .Y(_2733_)
);

FILL FILL_3__7034_ (
);

INVX1 _11208_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .Y(_2327_)
);

FILL FILL_1__13711_ (
);

FILL FILL_4__16156_ (
);

FILL FILL_6__10677_ (
);

FILL FILL_4__11291_ (
);

FILL FILL_3__15989_ (
);

FILL FILL_0__12704_ (
);

FILL FILL_3__15569_ (
);

FILL FILL_3__15149_ (
);

FILL FILL_1__16183_ (
);

FILL FILL_5__8741_ (
);

FILL FILL_5__8321_ (
);

FILL FILL_3__10284_ (
);

OAI22X1 _15881_ (
    .A(_5518__bF$buf3),
    .B(_4935_),
    .C(_5503__bF$buf2),
    .D(_6340_),
    .Y(_6341_)
);

FILL FILL_0__15596_ (
);

FILL FILL_0__15176_ (
);

NOR2X1 _15461_ (
    .A(_4449_),
    .B(_5549__bF$buf0),
    .Y(_5931_)
);

OR2X2 _15041_ (
    .A(_5520_),
    .B(_5517_),
    .Y(_5521_)
);

FILL FILL_1__8733_ (
);

FILL FILL_1__8313_ (
);

FILL FILL_2__15923_ (
);

FILL SFILL109320x36050 (
);

FILL FILL_2__15503_ (
);

FILL FILL_3__8659_ (
);

FILL FILL_3__8239_ (
);

FILL FILL_5__13083_ (
);

FILL FILL_1__14916_ (
);

DFFSR _7383_ (
    .Q(\datapath_1.regfile_1.regOut[4] [1]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_198_[1])
);

FILL FILL_4__12496_ (
);

FILL FILL_4__12076_ (
);

FILL SFILL69160x53050 (
);

FILL FILL_3__9600_ (
);

FILL FILL_0__13909_ (
);

FILL FILL_5__9526_ (
);

FILL FILL_3__11489_ (
);

FILL FILL_5__9106_ (
);

FILL FILL_3__11069_ (
);

FILL FILL_6__12403_ (
);

INVX1 _16246_ (
    .A(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_6696_)
);

OAI21X1 _11381_ (
    .A(_2141_),
    .B(_2142_),
    .C(_2152_),
    .Y(_2498_)
);

FILL FILL_0__11096_ (
);

FILL FILL_1__9938_ (
);

FILL FILL_5__11816_ (
);

FILL FILL_1__9518_ (
);

FILL FILL_3__12850_ (
);

FILL FILL_3__12430_ (
);

FILL FILL_3__12010_ (
);

FILL FILL_4__7943_ (
);

FILL FILL_4__7103_ (
);

FILL FILL_4__10809_ (
);

FILL FILL_2__11843_ (
);

FILL FILL_5__14288_ (
);

FILL FILL_2__11423_ (
);

FILL FILL_2__11003_ (
);

NAND2X1 _8588_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_862_)
);

DFFSR _8168_ (
    .Q(\datapath_1.regfile_1.regOut[10] [18]),
    .CLK(clk_bF$buf113),
    .R(rst_bF$buf22),
    .S(vdd),
    .D(_588_[18])
);

FILL FILL_1__10836_ (
);

FILL FILL_1__10416_ (
);

FILL FILL_0__7843_ (
);

FILL FILL_0__7423_ (
);

FILL FILL_6__13608_ (
);

FILL FILL_4__14642_ (
);

FILL SFILL64120x79050 (
);

FILL FILL_4__14222_ (
);

NAND2X1 _12586_ (
    .A(vdd),
    .B(memoryOutData[6]),
    .Y(_3437_)
);

INVX1 _12166_ (
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3164_)
);

FILL FILL_3__13635_ (
);

FILL FILL_3__13215_ (
);

FILL FILL_4__8728_ (
);

FILL FILL_2__12628_ (
);

FILL FILL_0__13662_ (
);

FILL FILL_2__12208_ (
);

FILL SFILL99320x40050 (
);

FILL FILL_0__13242_ (
);

FILL FILL_5__16014_ (
);

FILL FILL_0__8628_ (
);

FILL SFILL28760x60050 (
);

FILL FILL_0__8208_ (
);

FILL SFILL59160x51050 (
);

FILL FILL_1__9271_ (
);

FILL FILL_4__15847_ (
);

FILL FILL_4__15427_ (
);

FILL FILL_4__15007_ (
);

FILL FILL_2__16041_ (
);

FILL FILL_4__10982_ (
);

FILL FILL_4__10562_ (
);

FILL SFILL99240x47050 (
);

FILL FILL_4__10142_ (
);

FILL FILL_1__15874_ (
);

FILL FILL_1__15454_ (
);

FILL FILL_1__15034_ (
);

FILL FILL_0__14867_ (
);

INVX1 _14732_ (
    .A(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_5218_)
);

FILL FILL_0__14447_ (
);

FILL SFILL89320x83050 (
);

FILL FILL_0__14027_ (
);

AOI21X1 _14312_ (
    .A(_4806_),
    .B(_4783_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [17])
);

FILL FILL_2__7194_ (
);

FILL FILL_6__13781_ (
);

CLKBUF1 CLKBUF1_insert190 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert191 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert192 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert193 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert194 (
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert195 (
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf29)
);

FILL FILL_5__12774_ (
);

CLKBUF1 CLKBUF1_insert196 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf28)
);

FILL FILL_5__12354_ (
);

CLKBUF1 CLKBUF1_insert197 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert198 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert199 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf25)
);

FILL SFILL84200x1050 (
);

FILL FILL_4__8481_ (
);

FILL FILL_4__11767_ (
);

FILL FILL_4__8061_ (
);

FILL FILL_4__11347_ (
);

FILL FILL_2__12381_ (
);

FILL SFILL54120x77050 (
);

FILL FILL_1__16239_ (
);

FILL FILL_1__11794_ (
);

FILL FILL_1__11374_ (
);

OAI22X1 _15937_ (
    .A(_5472__bF$buf3),
    .B(_5013_),
    .C(_4995_),
    .D(_5552__bF$buf2),
    .Y(_6395_)
);

OAI22X1 _15517_ (
    .A(_5480__bF$buf3),
    .B(_5984_),
    .C(_5985_),
    .D(_5499__bF$buf1),
    .Y(_5986_)
);

FILL FILL_0__10787_ (
);

FILL FILL_0__8381_ (
);

FILL FILL_2__8399_ (
);

FILL FILL_0__10367_ (
);

OAI21X1 _10652_ (
    .A(_1911_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .C(_1912_),
    .Y(_1888_[12])
);

OAI21X1 _10232_ (
    .A(_1756_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1757_),
    .Y(_1693_[0])
);

FILL FILL_3__11701_ (
);

FILL FILL_4__15180_ (
);

FILL FILL_5__13979_ (
);

FILL FILL_2__9760_ (
);

FILL FILL_5__13559_ (
);

FILL FILL_3__14593_ (
);

FILL FILL_5__13139_ (
);

FILL FILL_2__9340_ (
);

FILL FILL_3__14173_ (
);

NAND2X1 _7859_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_498_)
);

NAND2X1 _7439_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_279_)
);

DFFSR _7019_ (
    .Q(\datapath_1.regfile_1.regOut[1] [21]),
    .CLK(clk_bF$buf9),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_3_[21])
);

FILL FILL_4_BUFX2_insert870 (
);

FILL FILL_4_BUFX2_insert871 (
);

FILL FILL_4_BUFX2_insert872 (
);

FILL FILL_4__9266_ (
);

FILL FILL_4_BUFX2_insert873 (
);

FILL FILL_2__13586_ (
);

FILL FILL_4_BUFX2_insert874 (
);

FILL FILL_2__13166_ (
);

FILL FILL_4_BUFX2_insert875 (
);

FILL FILL_4_BUFX2_insert876 (
);

FILL FILL_4_BUFX2_insert877 (
);

FILL FILL_5__14920_ (
);

FILL FILL_5__14500_ (
);

FILL FILL_4_BUFX2_insert878 (
);

FILL FILL_4_BUFX2_insert879 (
);

FILL SFILL89240x45050 (
);

FILL FILL_1__12999_ (
);

DFFSR _8800_ (
    .Q(\datapath_1.regfile_1.regOut[15] [10]),
    .CLK(clk_bF$buf42),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_913_[10])
);

FILL SFILL54120x32050 (
);

FILL FILL_1__12579_ (
);

FILL FILL_1__12159_ (
);

FILL FILL_4__13913_ (
);

FILL FILL_3__7683_ (
);

FILL FILL_0__9166_ (
);

NAND3X1 _11857_ (
    .A(_2943_),
    .B(_2675_),
    .C(_2776_),
    .Y(_2944_)
);

OAI21X1 _11437_ (
    .A(_2552_),
    .B(_2550_),
    .C(_2434_),
    .Y(_2553_)
);

AND2X2 _11017_ (
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2136_)
);

FILL FILL_3__12906_ (
);

FILL SFILL18680x65050 (
);

FILL FILL_1__13940_ (
);

FILL FILL_4__16385_ (
);

FILL FILL_1__13520_ (
);

FILL FILL_5__7189_ (
);

FILL FILL_1__13100_ (
);

FILL FILL_6__10486_ (
);

FILL FILL_3__15798_ (
);

FILL FILL_3__15378_ (
);

FILL FILL_0__12513_ (
);

FILL FILL_5__8970_ (
);

FILL FILL_5__8130_ (
);

NOR2X1 _15690_ (
    .A(_6144_),
    .B(_6154_),
    .Y(_6155_)
);

INVX1 _15270_ (
    .A(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_5745_)
);

FILL FILL_5__15705_ (
);

FILL FILL_1__8962_ (
);

FILL FILL_5__10420_ (
);

FILL FILL_1__8122_ (
);

FILL FILL_5__10000_ (
);

FILL FILL_2__15732_ (
);

FILL FILL_2__15312_ (
);

FILL FILL_3__8888_ (
);

FILL FILL_3__8468_ (
);

FILL FILL_1__14725_ (
);

NAND2X1 _7192_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_155_)
);

FILL FILL_1__14305_ (
);

FILL SFILL18680x20050 (
);

FILL FILL_0__13718_ (
);

FILL FILL_2__6885_ (
);

FILL FILL_5__9755_ (
);

FILL FILL_5__9335_ (
);

FILL FILL_3__11298_ (
);

INVX1 _16055_ (
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_6510_)
);

INVX2 _11190_ (
    .A(_2308_),
    .Y(_2309_)
);

FILL FILL_1__9747_ (
);

FILL FILL_5__11625_ (
);

FILL FILL_5__11205_ (
);

FILL SFILL79240x43050 (
);

FILL FILL_3_BUFX2_insert890 (
);

FILL FILL_4__7752_ (
);

FILL FILL_3_BUFX2_insert891 (
);

FILL FILL_4__7332_ (
);

FILL FILL_3_BUFX2_insert892 (
);

FILL FILL_4__10618_ (
);

FILL FILL_3_BUFX2_insert893 (
);

FILL FILL_2__11652_ (
);

FILL FILL_3_BUFX2_insert894 (
);

FILL FILL_2__11232_ (
);

FILL FILL_5__14097_ (
);

FILL FILL_3_BUFX2_insert895 (
);

INVX1 _8397_ (
    .A(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_775_)
);

FILL FILL_3_BUFX2_insert896 (
);

FILL SFILL95080x1050 (
);

FILL FILL_3_BUFX2_insert897 (
);

FILL FILL_3_BUFX2_insert898 (
);

FILL FILL_3_BUFX2_insert899 (
);

FILL FILL_1__10645_ (
);

FILL FILL_0__7232_ (
);

FILL SFILL109400x69050 (
);

FILL FILL_4__14871_ (
);

FILL SFILL44040x37050 (
);

FILL SFILL54120x5050 (
);

FILL FILL_4__14451_ (
);

FILL FILL_4__14031_ (
);

FILL SFILL94360x3050 (
);

NAND2X1 _12395_ (
    .A(MemToReg_bF$buf4),
    .B(\datapath_1.Data [17]),
    .Y(_3329_)
);

FILL FILL_3__13864_ (
);

FILL FILL_2__8611_ (
);

FILL SFILL94280x8050 (
);

FILL FILL_3__13444_ (
);

FILL FILL_3__13024_ (
);

FILL FILL_4__8957_ (
);

FILL FILL_4__8117_ (
);

FILL FILL_2__12857_ (
);

FILL FILL_2__12437_ (
);

FILL FILL_0__13891_ (
);

FILL FILL_2__12017_ (
);

FILL FILL_0__13471_ (
);

FILL FILL111880x11050 (
);

FILL FILL_5__16243_ (
);

FILL FILL_0__8857_ (
);

FILL FILL_3__6954_ (
);

NAND2X1 _10708_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1950_)
);

FILL FILL_0__8017_ (
);

FILL SFILL104520x6050 (
);

FILL FILL_1__9080_ (
);

FILL FILL_4__15656_ (
);

FILL FILL_4__15236_ (
);

FILL FILL_2__16270_ (
);

FILL FILL_4__10791_ (
);

FILL FILL_4__10371_ (
);

FILL FILL_3__14649_ (
);

FILL FILL_3__14229_ (
);

FILL FILL_1__15683_ (
);

FILL FILL_1__15263_ (
);

FILL FILL_5__7821_ (
);

INVX1 _14961_ (
    .A(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_5442_)
);

FILL FILL_0__14676_ (
);

FILL FILL_0__14256_ (
);

INVX1 _14541_ (
    .A(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_5031_)
);

NOR2X1 _14121_ (
    .A(_4605_),
    .B(_4619_),
    .Y(_4620_)
);

FILL FILL_1__7813_ (
);

FILL FILL_3__7739_ (
);

FILL FILL_3__7319_ (
);

FILL FILL_5__12583_ (
);

FILL FILL_5__12163_ (
);

BUFX2 _6883_ (
    .A(_2_[13]),
    .Y(memoryWriteData[13])
);

FILL SFILL99400x73050 (
);

FILL FILL_4__11996_ (
);

FILL FILL_4__11576_ (
);

FILL SFILL69160x48050 (
);

FILL FILL_4__11156_ (
);

FILL FILL_2__12190_ (
);

FILL FILL_1__16048_ (
);

FILL FILL_3__10989_ (
);

FILL FILL_3__10569_ (
);

FILL FILL_5__8606_ (
);

FILL FILL_3__10149_ (
);

FILL FILL_1__11183_ (
);

NOR3X1 _15746_ (
    .A(_6208_),
    .B(_6203_),
    .C(_6199_),
    .Y(_6209_)
);

OAI22X1 _15326_ (
    .A(_4273_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf0),
    .D(_4250_),
    .Y(_5800_)
);

NAND2X1 _10881_ (
    .A(_2024_),
    .B(_2028_),
    .Y(_2029_)
);

FILL FILL_0__8190_ (
);

DFFSR _10461_ (
    .Q(\datapath_1.regfile_1.regOut[28] [7]),
    .CLK(clk_bF$buf33),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_1758_[7])
);

FILL FILL_0__10176_ (
);

NAND2X1 _10041_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1607_)
);

FILL FILL_3__11930_ (
);

FILL FILL_6__14375_ (
);

FILL FILL_3__11510_ (
);

FILL FILL_0__16402_ (
);

FILL FILL_2__10923_ (
);

FILL FILL_5__13788_ (
);

FILL FILL_5__13368_ (
);

FILL FILL_2__10503_ (
);

DFFSR _7668_ (
    .Q(\datapath_1.regfile_1.regOut[6] [30]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_328_[30])
);

INVX1 _7248_ (
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_192_)
);

FILL FILL_4__9495_ (
);

FILL FILL_2__13395_ (
);

FILL FILL_0__6923_ (
);

FILL FILL_1__12388_ (
);

FILL FILL_4__13722_ (
);

FILL FILL_4__13302_ (
);

FILL FILL_3__7492_ (
);

FILL FILL_0__9395_ (
);

FILL FILL_3__7072_ (
);

NAND2X1 _11666_ (
    .A(_2179_),
    .B(_2341__bF$buf1),
    .Y(_2768_)
);

XOR2X1 _11246_ (
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2365_)
);

FILL FILL_3__12715_ (
);

FILL FILL_4__16194_ (
);

FILL FILL_4__7808_ (
);

FILL FILL_6__10295_ (
);

FILL FILL_2__11708_ (
);

FILL SFILL99320x35050 (
);

FILL FILL_0__12742_ (
);

FILL FILL_3__15187_ (
);

FILL FILL_0__12322_ (
);

FILL SFILL23800x7050 (
);

FILL FILL_5__15934_ (
);

FILL SFILL89400x71050 (
);

FILL FILL_5__15514_ (
);

FILL SFILL28760x55050 (
);

FILL FILL_0__7708_ (
);

DFFSR _9814_ (
    .Q(\datapath_1.regfile_1.regOut[23] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_1433_[0])
);

FILL FILL_1__8771_ (
);

FILL FILL_1__8351_ (
);

FILL FILL_4__14927_ (
);

FILL FILL_4__14507_ (
);

FILL FILL_2__15961_ (
);

FILL FILL_2__15541_ (
);

FILL FILL_2__15121_ (
);

FILL FILL_3__8697_ (
);

FILL FILL_3__8277_ (
);

FILL SFILL64120x29050 (
);

FILL SFILL3640x8050 (
);

FILL SFILL49240x82050 (
);

FILL FILL_1__14954_ (
);

FILL FILL_1__14534_ (
);

FILL FILL_1__14114_ (
);

FILL FILL_0__13947_ (
);

FILL SFILL89320x78050 (
);

INVX1 _13812_ (
    .A(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_4317_)
);

FILL FILL_0__13527_ (
);

FILL FILL_0__13107_ (
);

FILL FILL_5__9984_ (
);

FILL FILL_5__9144_ (
);

AOI22X1 _16284_ (
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [31]),
    .C(\datapath_1.regfile_1.regOut[22] [31]),
    .D(_5650_),
    .Y(_6733_)
);

FILL SFILL49640x51050 (
);

FILL FILL_1__9976_ (
);

FILL FILL_5__11854_ (
);

FILL FILL_1__9556_ (
);

FILL FILL_5__11434_ (
);

FILL FILL_1__9136_ (
);

FILL FILL_5__11014_ (
);

FILL SFILL28760x10050 (
);

FILL FILL_4__7981_ (
);

FILL FILL_2__16326_ (
);

FILL FILL_4__7561_ (
);

FILL SFILL89720x47050 (
);

FILL FILL_4__10427_ (
);

FILL FILL_2__11881_ (
);

FILL FILL_4__10007_ (
);

FILL FILL_2__11461_ (
);

FILL FILL_2__11041_ (
);

FILL FILL_6__7487_ (
);

FILL FILL_1__15739_ (
);

FILL FILL_1__15319_ (
);

FILL FILL_1__10874_ (
);

FILL FILL_1__10034_ (
);

FILL SFILL33960x73050 (
);

FILL FILL_0__7881_ (
);

FILL FILL_2__7479_ (
);

FILL FILL_0__7461_ (
);

FILL FILL_0__7041_ (
);

FILL FILL_2__7059_ (
);

FILL FILL_4__14680_ (
);

FILL FILL_4__14260_ (
);

FILL FILL_2__8840_ (
);

FILL FILL_5__12639_ (
);

FILL FILL_3__13673_ (
);

FILL FILL_5__12219_ (
);

FILL FILL_3__13253_ (
);

FILL FILL_2__8000_ (
);

NAND2X1 _6939_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_27_)
);

FILL SFILL18760x53050 (
);

FILL FILL_4__8766_ (
);

FILL FILL_4__8346_ (
);

FILL FILL_2__12246_ (
);

FILL FILL_0__13280_ (
);

FILL SFILL58840x49050 (
);

FILL SFILL54120x27050 (
);

FILL FILL_1__11659_ (
);

FILL FILL_1__11239_ (
);

FILL FILL_5__16052_ (
);

INVX2 _10937_ (
    .A(\control_1.op [2]),
    .Y(_2071_)
);

FILL FILL_0__8246_ (
);

NAND2X1 _10517_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1843_)
);

FILL SFILL79320x76050 (
);

FILL FILL_4__15885_ (
);

FILL FILL_1__12600_ (
);

FILL FILL_4__15465_ (
);

FILL FILL_4__15045_ (
);

FILL FILL_4__10180_ (
);

FILL FILL_3__14878_ (
);

FILL FILL_2__9625_ (
);

FILL FILL_3__14458_ (
);

FILL FILL_3__14038_ (
);

FILL FILL_1__15492_ (
);

FILL FILL_1__15072_ (
);

FILL FILL_5__7630_ (
);

FILL FILL_5__7210_ (
);

FILL FILL_0__14485_ (
);

INVX1 _14770_ (
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_5255_)
);

FILL FILL_0__14065_ (
);

INVX1 _14350_ (
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_4844_)
);

FILL FILL_1__7622_ (
);

FILL FILL_1__7202_ (
);

FILL FILL_2__14812_ (
);

FILL FILL_3__7968_ (
);

FILL FILL_3__7548_ (
);

FILL FILL_5__12392_ (
);

FILL FILL_1__13805_ (
);

FILL SFILL33960x9050 (
);

FILL SFILL79320x31050 (
);

FILL SFILL18680x15050 (
);

FILL FILL_4__11385_ (
);

FILL FILL_1__16277_ (
);

FILL FILL_5__8835_ (
);

FILL FILL_3__10798_ (
);

FILL FILL_3__10378_ (
);

FILL FILL111960x44050 (
);

NOR2X1 _15975_ (
    .A(_6431_),
    .B(_6429_),
    .Y(_6432_)
);

FILL FILL_6__11712_ (
);

NOR2X1 _15555_ (
    .A(_6019_),
    .B(_6022_),
    .Y(_6023_)
);

NOR2X1 _15135_ (
    .A(_5612_),
    .B(_5610_),
    .Y(_5613_)
);

NAND2X1 _10690_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1938_)
);

NAND2X1 _10270_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1719_)
);

FILL FILL_5__10705_ (
);

FILL FILL_1__8827_ (
);

FILL SFILL79240x38050 (
);

FILL FILL_0__16211_ (
);

FILL FILL_5__13597_ (
);

FILL FILL_2__10312_ (
);

DFFSR _7897_ (
    .Q(\datapath_1.regfile_1.regOut[8] [3]),
    .CLK(clk_bF$buf1),
    .R(rst_bF$buf104),
    .S(vdd),
    .D(_458_[3])
);

INVX1 _7477_ (
    .A(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_304_)
);

INVX1 _7057_ (
    .A(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_85_)
);

FILL FILL_1__12197_ (
);

FILL FILL_4__13951_ (
);

FILL FILL_4__13531_ (
);

FILL FILL_4__13111_ (
);

OAI21X1 _11895_ (
    .A(_2970_),
    .B(IorD_bF$buf6),
    .C(_2971_),
    .Y(_1_[2])
);

OAI21X1 _11475_ (
    .A(_2569_),
    .B(_2436_),
    .C(_2589_),
    .Y(_2590_)
);

NAND2X1 _11055_ (
    .A(_2170_),
    .B(_2173_),
    .Y(_2174_)
);

FILL FILL_3__12524_ (
);

FILL FILL_3__12104_ (
);

FILL FILL_4__7617_ (
);

FILL FILL_2__11937_ (
);

FILL FILL_0__12971_ (
);

FILL FILL_2__11517_ (
);

FILL FILL_0__12131_ (
);

FILL FILL_5__15743_ (
);

FILL FILL_0__7937_ (
);

FILL FILL_5__15323_ (
);

INVX1 _9623_ (
    .A(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_1389_)
);

DFFSR _9203_ (
    .Q(\datapath_1.regfile_1.regOut[18] [29]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_1108_[29])
);

FILL FILL_1__8580_ (
);

FILL FILL_4__14736_ (
);

FILL FILL_4__14316_ (
);

FILL FILL_2__15770_ (
);

FILL SFILL109400x19050 (
);

FILL FILL_2__15350_ (
);

FILL FILL_3__8086_ (
);

FILL FILL_3__13729_ (
);

FILL FILL_3__13309_ (
);

FILL FILL_1__14763_ (
);

FILL FILL_1__14343_ (
);

FILL FILL_5__6901_ (
);

FILL SFILL69240x36050 (
);

FILL FILL_0__13756_ (
);

FILL FILL_0__13336_ (
);

AOI22X1 _13621_ (
    .A(\datapath_1.regfile_1.regOut[27] [3]),
    .B(_4129_),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_4130_)
);

DFFSR _13201_ (
    .Q(\datapath_1.mux_iord.din0 [26]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3685_[26])
);

FILL FILL_5__9793_ (
);

FILL FILL_5__9373_ (
);

NOR3X1 _16093_ (
    .A(_6543_),
    .B(_6544_),
    .C(_6546_),
    .Y(_6547_)
);

FILL SFILL59320x72050 (
);

FILL FILL_5__16108_ (
);

FILL FILL_1__9785_ (
);

FILL FILL_5__11663_ (
);

FILL FILL_5__11243_ (
);

FILL FILL_1__9365_ (
);

FILL SFILL99400x68050 (
);

FILL FILL_2__16135_ (
);

FILL FILL_4__7370_ (
);

FILL FILL_4__10656_ (
);

FILL FILL_2__11690_ (
);

FILL FILL_4__10236_ (
);

FILL FILL_2__11270_ (
);

FILL FILL_1__15968_ (
);

FILL FILL_6__7296_ (
);

FILL FILL_1__15548_ (
);

FILL FILL_1__15128_ (
);

FILL FILL_1__10683_ (
);

FILL FILL_1__10263_ (
);

INVX1 _14826_ (
    .A(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_5310_)
);

INVX1 _14406_ (
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_4898_)
);

FILL FILL_0__7690_ (
);

FILL FILL_2__7288_ (
);

FILL SFILL104360x61050 (
);

FILL FILL_0__15902_ (
);

FILL FILL_5__12868_ (
);

FILL FILL_5__12448_ (
);

FILL SFILL43240x80050 (
);

FILL FILL_5__12028_ (
);

FILL FILL_3__13482_ (
);

FILL SFILL69080x9050 (
);

FILL FILL_4__8995_ (
);

FILL FILL_4__8575_ (
);

FILL FILL_2__12895_ (
);

FILL FILL_2__12475_ (
);

FILL FILL_2__12055_ (
);

FILL SFILL99400x23050 (
);

FILL SFILL104280x68050 (
);

FILL FILL_1__11888_ (
);

FILL FILL_1__11468_ (
);

FILL FILL_1__11048_ (
);

FILL FILL_0__8895_ (
);

FILL FILL_3__6992_ (
);

FILL FILL_5__16281_ (
);

FILL FILL_0__8475_ (
);

FILL FILL_0__8055_ (
);

NAND2X1 _10746_ (
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1955_)
);

DFFSR _10326_ (
    .Q(\datapath_1.regfile_1.regOut[27] [0]),
    .CLK(clk_bF$buf92),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_1693_[0])
);

FILL FILL_6__9022_ (
);

FILL FILL_4__15694_ (
);

FILL FILL_4__15274_ (
);

FILL FILL_2__9854_ (
);

FILL FILL_0__11822_ (
);

FILL FILL_3__14687_ (
);

FILL FILL_2__9014_ (
);

FILL FILL_3__14267_ (
);

FILL FILL_0__11402_ (
);

FILL FILL_0__14294_ (
);

FILL SFILL89400x66050 (
);

FILL FILL_1__7851_ (
);

FILL FILL_1__7431_ (
);

FILL SFILL104280x23050 (
);

FILL FILL_2__14621_ (
);

FILL FILL_2__14201_ (
);

FILL FILL_3__7357_ (
);

FILL FILL_1__13614_ (
);

FILL FILL_4__16059_ (
);

FILL FILL_4__11194_ (
);

FILL FILL_0__12607_ (
);

FILL FILL_1__16086_ (
);

FILL FILL_1_BUFX2_insert225 (
);

FILL FILL_1_BUFX2_insert226 (
);

FILL FILL_5__8644_ (
);

FILL FILL_1_BUFX2_insert227 (
);

FILL FILL_3__10187_ (
);

FILL FILL_5__8224_ (
);

FILL FILL_6_BUFX2_insert781 (
);

FILL FILL_1_BUFX2_insert228 (
);

FILL FILL_1_BUFX2_insert229 (
);

FILL FILL_0__15499_ (
);

NOR2X1 _15784_ (
    .A(_6245_),
    .B(_6242_),
    .Y(_6246_)
);

INVX1 _15364_ (
    .A(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_5837_)
);

FILL FILL_0__15079_ (
);

FILL FILL_6_BUFX2_insert787 (
);

FILL FILL_3__16413_ (
);

FILL FILL_5__10934_ (
);

FILL SFILL89400x21050 (
);

FILL FILL_1__8636_ (
);

FILL FILL_5__10514_ (
);

FILL FILL_1__8216_ (
);

FILL SFILL94280x72050 (
);

FILL FILL_2__15826_ (
);

FILL FILL_2__15406_ (
);

FILL FILL_0__16020_ (
);

FILL FILL_2__10961_ (
);

FILL FILL_2__10541_ (
);

FILL FILL_2__10121_ (
);

FILL FILL_1__14819_ (
);

INVX1 _7286_ (
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_261_)
);

FILL FILL_4__12399_ (
);

FILL FILL_3__9923_ (
);

FILL FILL_3__9503_ (
);

FILL SFILL33960x68050 (
);

FILL FILL_0__6961_ (
);

FILL FILL_2__6979_ (
);

FILL FILL_5__9849_ (
);

FILL FILL_5__9429_ (
);

FILL FILL_5__9009_ (
);

FILL FILL_4__13760_ (
);

FILL FILL_4__13340_ (
);

OAI21X1 _16149_ (
    .A(_5232_),
    .B(_5535__bF$buf3),
    .C(_6601_),
    .Y(_6602_)
);

NOR2X1 _11284_ (
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2403_)
);

FILL FILL_5__11719_ (
);

FILL FILL_3__12753_ (
);

FILL FILL_2__7500_ (
);

FILL FILL_3__12333_ (
);

FILL FILL_4__7846_ (
);

FILL FILL_4__7426_ (
);

FILL FILL_2__11746_ (
);

FILL FILL_0__12780_ (
);

FILL FILL_2__11326_ (
);

FILL FILL_0__12360_ (
);

FILL FILL_1__10319_ (
);

FILL FILL_5__15972_ (
);

FILL FILL_5__15552_ (
);

FILL FILL_5__15132_ (
);

FILL FILL_0__7746_ (
);

FILL FILL_6__8713_ (
);

FILL FILL_0__7326_ (
);

INVX1 _9852_ (
    .A(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_1501_)
);

DFFSR _9432_ (
    .Q(\datapath_1.regfile_1.regOut[20] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_1238_[2])
);

OAI21X1 _9012_ (
    .A(_1082_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1083_),
    .Y(_1043_[20])
);

FILL SFILL33960x23050 (
);

FILL FILL_4__14965_ (
);

FILL FILL_4__14545_ (
);

FILL FILL_4__14125_ (
);

OAI21X1 _12489_ (
    .A(_3391_),
    .B(vdd),
    .C(_3392_),
    .Y(_3360_[16])
);

AOI22X1 _12069_ (
    .A(\datapath_1.ALUResult [20]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3098_)
);

FILL FILL_2__8705_ (
);

FILL FILL_3__13958_ (
);

FILL FILL_1__14992_ (
);

FILL FILL_3__13538_ (
);

FILL FILL_1__14572_ (
);

FILL FILL_3__13118_ (
);

FILL FILL_1__14152_ (
);

FILL SFILL84280x70050 (
);

FILL FILL_0__13985_ (
);

NOR2X1 _13850_ (
    .A(_4353_),
    .B(_3977__bF$buf1),
    .Y(_4354_)
);

FILL FILL_0__13565_ (
);

INVX8 _13430_ (
    .A(_3941_),
    .Y(_3942_)
);

FILL FILL_0__13145_ (
);

OAI21X1 _13010_ (
    .A(_3657_),
    .B(vdd),
    .C(_3658_),
    .Y(_3620_[19])
);

FILL FILL_5__16337_ (
);

FILL FILL_5__11892_ (
);

FILL FILL_1__9594_ (
);

FILL FILL_5__11472_ (
);

FILL FILL_5__11052_ (
);

FILL SFILL79320x26050 (
);

FILL FILL_2__16364_ (
);

FILL FILL_4__10885_ (
);

FILL FILL_4__10045_ (
);

FILL FILL_1__15777_ (
);

FILL FILL_1__15357_ (
);

FILL FILL_1__10492_ (
);

INVX1 _14635_ (
    .A(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_5123_)
);

NAND3X1 _14215_ (
    .A(_4710_),
    .B(_4711_),
    .C(_4709_),
    .Y(_4712_)
);

FILL FILL_2__7097_ (
);

FILL FILL_6__13684_ (
);

FILL FILL_0__15711_ (
);

FILL FILL_5__12257_ (
);

FILL FILL_3__13291_ (
);

INVX1 _6977_ (
    .A(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_52_)
);

FILL FILL_4__8384_ (
);

FILL FILL_2__12284_ (
);

FILL SFILL114440x51050 (
);

FILL FILL_1__11697_ (
);

FILL FILL_1__11277_ (
);

FILL FILL_4__12611_ (
);

FILL FILL_5__16090_ (
);

INVX1 _10975_ (
    .A(\control_1.reg_state.dout [1]),
    .Y(_2101_)
);

INVX1 _10555_ (
    .A(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_1868_)
);

INVX1 _10135_ (
    .A(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_1649_)
);

FILL FILL_3__11604_ (
);

FILL FILL_4__15083_ (
);

FILL FILL_2__9663_ (
);

FILL FILL_3__14496_ (
);

FILL FILL_2__9243_ (
);

FILL FILL_0__11631_ (
);

FILL FILL_0__11211_ (
);

FILL FILL_3__14076_ (
);

FILL FILL_4__9169_ (
);

FILL FILL_2__13489_ (
);

FILL FILL_5__14823_ (
);

FILL FILL_5__14403_ (
);

INVX1 _8703_ (
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_918_)
);

FILL FILL_1__7240_ (
);

FILL FILL_4__13816_ (
);

FILL FILL_2__14850_ (
);

FILL FILL_2__14430_ (
);

FILL FILL_3__7586_ (
);

FILL FILL_2__14010_ (
);

FILL FILL_0__9489_ (
);

FILL FILL_3__7166_ (
);

FILL FILL_1__13843_ (
);

FILL FILL_1__13423_ (
);

FILL FILL_4__16288_ (
);

FILL FILL_1__13003_ (
);

FILL FILL_0__12836_ (
);

INVX1 _12701_ (
    .A(\aluControl_1.inst [2]),
    .Y(_3493_)
);

FILL FILL_0__12416_ (
);

FILL FILL_5__8873_ (
);

FILL FILL_5__8453_ (
);

NOR2X1 _15593_ (
    .A(_6056_),
    .B(_6059_),
    .Y(_6060_)
);

INVX8 _15173_ (
    .A(_5552__bF$buf2),
    .Y(_5650_)
);

FILL FILL_5__15608_ (
);

FILL FILL_3__16222_ (
);

OAI21X1 _9908_ (
    .A(_1537_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1538_),
    .Y(_1498_[20])
);

FILL FILL_1__8865_ (
);

FILL FILL_5__10743_ (
);

FILL FILL_5__10323_ (
);

FILL FILL_1__8445_ (
);

FILL FILL_2__15635_ (
);

FILL FILL_2__15215_ (
);

FILL FILL_4__6870_ (
);

FILL SFILL19160x78050 (
);

FILL FILL_2__10770_ (
);

FILL FILL_1__14628_ (
);

OAI21X1 _7095_ (
    .A(_109_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .C(_110_),
    .Y(_68_[21])
);

FILL FILL_1__14208_ (
);

FILL FILL_3__9732_ (
);

NOR2X1 _13906_ (
    .A(_4408_),
    .B(_4405_),
    .Y(_4409_)
);

FILL SFILL104360x56050 (
);

FILL FILL_5__9658_ (
);

FILL FILL_5__9238_ (
);

FILL FILL_6__12955_ (
);

INVX1 _16378_ (
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_6806_)
);

FILL FILL_5__11948_ (
);

INVX1 _11093_ (
    .A(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2212_)
);

FILL FILL_3__12982_ (
);

FILL FILL_5__11528_ (
);

FILL FILL_5__11108_ (
);

FILL FILL_3__12142_ (
);

FILL FILL_4__7235_ (
);

FILL FILL_2__11975_ (
);

FILL FILL_2__11555_ (
);

FILL SFILL99400x18050 (
);

FILL FILL_2__11135_ (
);

FILL FILL_1__10968_ (
);

FILL FILL_1__10548_ (
);

FILL FILL_1__10128_ (
);

FILL FILL_5__15781_ (
);

FILL FILL_0__7975_ (
);

FILL FILL_5__15361_ (
);

FILL FILL_0__7555_ (
);

FILL FILL112440x62050 (
);

OAI21X1 _9661_ (
    .A(_1413_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1414_),
    .Y(_1368_[23])
);

FILL FILL_5_CLKBUF1_insert1074 (
);

FILL FILL_6__8102_ (
);

OAI21X1 _9241_ (
    .A(_1194_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1195_),
    .Y(_1173_[11])
);

FILL FILL_5_CLKBUF1_insert1075 (
);

FILL FILL_5_CLKBUF1_insert1076 (
);

FILL FILL_5_CLKBUF1_insert1077 (
);

FILL FILL_5_CLKBUF1_insert1078 (
);

FILL FILL_4__14774_ (
);

FILL SFILL104360x11050 (
);

FILL FILL_4__14354_ (
);

FILL FILL_5_CLKBUF1_insert1079 (
);

NAND3X1 _12298_ (
    .A(_3260_),
    .B(_3261_),
    .C(_3262_),
    .Y(\datapath_1.alu_1.ALUInB [20])
);

FILL FILL_0__10902_ (
);

FILL FILL_3__13767_ (
);

FILL FILL_2__8514_ (
);

FILL FILL_3__13347_ (
);

FILL FILL_1__14381_ (
);

FILL FILL_0__13794_ (
);

FILL FILL_0__13374_ (
);

FILL FILL_1__6931_ (
);

FILL FILL_4__9801_ (
);

FILL FILL_2__13701_ (
);

FILL FILL_3__6857_ (
);

FILL FILL_5__16146_ (
);

FILL FILL_5__11281_ (
);

FILL FILL_4__15979_ (
);

FILL FILL_4__15559_ (
);

FILL FILL_4__15139_ (
);

FILL FILL_2__16173_ (
);

FILL FILL_4__10694_ (
);

FILL FILL_4__10274_ (
);

FILL FILL_2__9719_ (
);

FILL FILL_1__15586_ (
);

FILL FILL_1__15166_ (
);

FILL FILL_5__7724_ (
);

FILL FILL_5__7304_ (
);

FILL FILL_0__14999_ (
);

INVX1 _14864_ (
    .A(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_5347_)
);

FILL FILL_0__14579_ (
);

FILL FILL_0__14159_ (
);

OAI22X1 _14444_ (
    .A(_4935_),
    .B(_3941_),
    .C(_3966__bF$buf1),
    .D(_4934_),
    .Y(_4936_)
);

AOI21X1 _14024_ (
    .A(_4524_),
    .B(_4499_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [11])
);

FILL FILL_3__15913_ (
);

FILL SFILL89400x16050 (
);

FILL FILL_1__7716_ (
);

FILL FILL_2__14906_ (
);

FILL FILL_0__15940_ (
);

FILL FILL_0__15520_ (
);

FILL FILL_0__15100_ (
);

FILL FILL_5__12486_ (
);

FILL FILL_5__12066_ (
);

FILL SFILL49240x27050 (
);

FILL FILL_4__8193_ (
);

FILL FILL_4__11899_ (
);

FILL FILL_4__11479_ (
);

FILL FILL_4__11059_ (
);

FILL FILL_2__12093_ (
);

FILL FILL_5__8509_ (
);

FILL FILL_1__11086_ (
);

NAND2X1 _15649_ (
    .A(_6111_),
    .B(_6114_),
    .Y(_6115_)
);

FILL FILL_4__12840_ (
);

NAND3X1 _15229_ (
    .A(_5699_),
    .B(_5701_),
    .C(_5704_),
    .Y(_5705_)
);

FILL FILL_4__12420_ (
);

FILL FILL_4__12000_ (
);

INVX1 _10784_ (
    .A(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_1980_)
);

FILL FILL_0__10499_ (
);

FILL FILL_0__8093_ (
);

INVX1 _10364_ (
    .A(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_1761_)
);

FILL SFILL79400x59050 (
);

FILL FILL_3__11833_ (
);

FILL FILL_6__14278_ (
);

FILL FILL_3__11413_ (
);

FILL FILL_4__6926_ (
);

FILL FILL_0__16305_ (
);

FILL SFILL94280x22050 (
);

FILL FILL_2__9892_ (
);

FILL FILL_2__10826_ (
);

FILL FILL_2__9472_ (
);

FILL FILL_2__10406_ (
);

FILL FILL_0__11860_ (
);

FILL FILL_0__11440_ (
);

FILL FILL_0__11020_ (
);

FILL FILL_4__9398_ (
);

FILL FILL_2__13298_ (
);

FILL FILL_5__14632_ (
);

FILL FILL_5__14212_ (
);

DFFSR _8932_ (
    .Q(\datapath_1.regfile_1.regOut[16] [14]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf59),
    .S(vdd),
    .D(_978_[14])
);

OAI21X1 _8512_ (
    .A(_830_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .C(_831_),
    .Y(_783_[24])
);

FILL SFILL33960x18050 (
);

FILL FILL_4__13625_ (
);

AOI22X1 _11989_ (
    .A(\datapath_1.ALUResult [0]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3038_)
);

FILL FILL_0__9298_ (
);

OAI21X1 _11569_ (
    .A(_2676_),
    .B(_2520_),
    .C(_2275_),
    .Y(_2677_)
);

OAI21X1 _11149_ (
    .A(_2251_),
    .B(_2252_),
    .C(_2267_),
    .Y(_2268_)
);

FILL FILL_3_BUFX2_insert40 (
);

FILL FILL_3__12618_ (
);

FILL FILL_1__13652_ (
);

FILL FILL_3_BUFX2_insert41 (
);

FILL FILL_1__13232_ (
);

FILL FILL_3_BUFX2_insert42 (
);

FILL FILL_4__16097_ (
);

FILL FILL_3_BUFX2_insert43 (
);

FILL FILL_3_BUFX2_insert44 (
);

FILL FILL_3_BUFX2_insert45 (
);

FILL SFILL84280x65050 (
);

FILL FILL_3_BUFX2_insert46 (
);

FILL FILL_1_BUFX2_insert600 (
);

FILL FILL_3_BUFX2_insert47 (
);

FILL FILL_1_BUFX2_insert601 (
);

FILL FILL_0__12645_ (
);

FILL FILL_3_BUFX2_insert48 (
);

DFFSR _12930_ (
    .Q(\datapath_1.a [11]),
    .CLK(clk_bF$buf26),
    .R(rst_bF$buf7),
    .S(vdd),
    .D(_3555_[11])
);

FILL FILL_1_BUFX2_insert602 (
);

FILL FILL_1_BUFX2_insert603 (
);

OAI21X1 _12510_ (
    .A(_3405_),
    .B(vdd),
    .C(_3406_),
    .Y(_3360_[23])
);

FILL FILL_3_BUFX2_insert49 (
);

FILL FILL_0__12225_ (
);

FILL FILL_1_BUFX2_insert604 (
);

FILL FILL_1_BUFX2_insert605 (
);

FILL FILL_1_BUFX2_insert606 (
);

FILL FILL_1_BUFX2_insert607 (
);

FILL FILL_5__8262_ (
);

FILL FILL_1_BUFX2_insert608 (
);

FILL FILL_1_BUFX2_insert609 (
);

FILL FILL_5__15837_ (
);

FILL FILL_5__15417_ (
);

FILL FILL_3__16451_ (
);

FILL FILL_3__16031_ (
);

DFFSR _9717_ (
    .Q(\datapath_1.regfile_1.regOut[22] [31]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_1368_[31])
);

FILL FILL_5__10972_ (
);

FILL FILL_5__10552_ (
);

FILL FILL_1__8254_ (
);

FILL FILL_5__10132_ (
);

FILL FILL_2__15864_ (
);

FILL FILL_2__15444_ (
);

FILL SFILL29320x61050 (
);

FILL FILL_2__15024_ (
);

FILL FILL_1__14857_ (
);

FILL FILL_1__14437_ (
);

FILL FILL_1__14017_ (
);

FILL FILL_3__9541_ (
);

FILL FILL_3__9121_ (
);

INVX1 _13715_ (
    .A(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_4222_)
);

FILL SFILL84280x20050 (
);

FILL FILL_5__9887_ (
);

FILL FILL_5__9467_ (
);

FILL SFILL13640x83050 (
);

INVX1 _16187_ (
    .A(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_6639_)
);

FILL FILL_1__9879_ (
);

FILL FILL_5__11757_ (
);

FILL FILL_5__11337_ (
);

FILL FILL_1__9039_ (
);

FILL FILL_3__12371_ (
);

FILL SFILL53720x79050 (
);

FILL SFILL84600x32050 (
);

FILL FILL_2__16229_ (
);

FILL FILL_4__7884_ (
);

FILL FILL_4__7464_ (
);

FILL FILL_4__7044_ (
);

FILL FILL_2__11784_ (
);

FILL FILL_2__11364_ (
);

FILL FILL_1__10777_ (
);

FILL FILL_5__15590_ (
);

FILL FILL_5__15170_ (
);

FILL SFILL74280x63050 (
);

OAI21X1 _9890_ (
    .A(_1525_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1526_),
    .Y(_1498_[14])
);

FILL FILL_0__7364_ (
);

OAI21X1 _9470_ (
    .A(_1306_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .C(_1307_),
    .Y(_1303_[2])
);

DFFSR _9050_ (
    .Q(\datapath_1.regfile_1.regOut[17] [4]),
    .CLK(clk_bF$buf25),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_1043_[4])
);

FILL FILL_4__14583_ (
);

FILL FILL_4__14163_ (
);

FILL FILL_2__8743_ (
);

FILL FILL_3__13996_ (
);

FILL FILL_2__8323_ (
);

FILL FILL_3__13576_ (
);

FILL FILL_3__13156_ (
);

FILL FILL_1__14190_ (
);

FILL FILL_4__8249_ (
);

FILL FILL_2__12989_ (
);

FILL FILL_2__12569_ (
);

FILL FILL_2__12149_ (
);

FILL FILL_5__13903_ (
);

FILL FILL_4_BUFX2_insert110 (
);

FILL FILL_4__9610_ (
);

FILL FILL_2__13930_ (
);

FILL FILL_5__16375_ (
);

FILL FILL_2__13510_ (
);

FILL FILL_0__8989_ (
);

FILL SFILL74200x61050 (
);

FILL FILL_0__8569_ (
);

FILL FILL_0__8149_ (
);

FILL FILL_6__9116_ (
);

FILL FILL_5__11090_ (
);

FILL FILL_4__15788_ (
);

FILL FILL_4__15368_ (
);

FILL FILL_1__12503_ (
);

FILL FILL_0__9930_ (
);

FILL SFILL19240x66050 (
);

FILL FILL_0__9510_ (
);

FILL FILL_0__11916_ (
);

FILL FILL_2__9528_ (
);

FILL FILL_2__9108_ (
);

FILL FILL_1__15395_ (
);

FILL FILL_5__7953_ (
);

FILL FILL_5__7113_ (
);

FILL FILL_0__14388_ (
);

INVX1 _14673_ (
    .A(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_5160_)
);

NAND3X1 _14253_ (
    .A(_4747_),
    .B(_4748_),
    .C(_4746_),
    .Y(_4749_)
);

FILL FILL_3__15722_ (
);

FILL FILL_3__15302_ (
);

FILL FILL_1__7945_ (
);

FILL FILL_1__7105_ (
);

FILL FILL_2__14715_ (
);

FILL FILL_5__12295_ (
);

FILL FILL112120x81050 (
);

FILL FILL_1__13708_ (
);

FILL FILL_4__11288_ (
);

FILL FILL_5__8738_ (
);

FILL FILL_5__8318_ (
);

INVX1 _15878_ (
    .A(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_6338_)
);

FILL FILL_6__11615_ (
);

NOR2X1 _15458_ (
    .A(_4467_),
    .B(_5534__bF$buf1),
    .Y(_5928_)
);

NAND3X1 _15038_ (
    .A(_5459__bF$buf3),
    .B(_5477_),
    .C(_5468_),
    .Y(_5518_)
);

DFFSR _10593_ (
    .Q(\datapath_1.regfile_1.regOut[29] [11]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf107),
    .S(vdd),
    .D(_1823_[11])
);

OAI21X1 _10173_ (
    .A(_1673_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .C(_1674_),
    .Y(_1628_[23])
);

FILL FILL_3__11642_ (
);

FILL SFILL95080x21050 (
);

FILL FILL_3__11222_ (
);

FILL FILL_0__16114_ (
);

FILL FILL_2__10635_ (
);

FILL FILL_2__9281_ (
);

FILL FILL_5__14861_ (
);

FILL FILL_5__14441_ (
);

FILL FILL112440x57050 (
);

FILL FILL_5__14021_ (
);

OAI21X1 _8741_ (
    .A(_942_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_943_),
    .Y(_913_[15])
);

OAI21X1 _8321_ (
    .A(_723_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .C(_724_),
    .Y(_718_[3])
);

FILL FILL_4__13854_ (
);

FILL FILL_4__13434_ (
);

FILL FILL_4__13014_ (
);

OAI21X1 _11798_ (
    .A(_2889_),
    .B(_2890_),
    .C(_2886_),
    .Y(_2891_)
);

NOR2X1 _11378_ (
    .A(_2140_),
    .B(_2145_),
    .Y(_2495_)
);

FILL SFILL33720x75050 (
);

FILL FILL_3__12847_ (
);

FILL FILL_1__13881_ (
);

FILL FILL_3__12427_ (
);

FILL FILL_1__13461_ (
);

FILL FILL_3__12007_ (
);

FILL FILL_1__13041_ (
);

FILL FILL_0__12874_ (
);

FILL FILL_0__12454_ (
);

FILL FILL_0__12034_ (
);

FILL FILL_5__8491_ (
);

FILL FILL_5__8071_ (
);

FILL FILL_5__15646_ (
);

FILL FILL_5__15226_ (
);

DFFSR _9946_ (
    .Q(\datapath_1.regfile_1.regOut[24] [4]),
    .CLK(clk_bF$buf66),
    .R(rst_bF$buf84),
    .S(vdd),
    .D(_1498_[4])
);

FILL FILL_3__16260_ (
);

NAND2X1 _9526_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1345_)
);

FILL FILL_5__10781_ (
);

NAND2X1 _9106_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1126_)
);

FILL FILL_1__8483_ (
);

FILL FILL_5__10361_ (
);

FILL FILL_1__8063_ (
);

FILL FILL112440x12050 (
);

FILL FILL_4__14639_ (
);

FILL FILL_2__15673_ (
);

FILL FILL_4__14219_ (
);

FILL FILL_2__15253_ (
);

FILL FILL_1__14666_ (
);

FILL FILL_1__14246_ (
);

FILL SFILL33720x30050 (
);

FILL FILL_0_BUFX2_insert260 (
);

FILL FILL_0_BUFX2_insert261 (
);

FILL FILL_0_BUFX2_insert262 (
);

FILL FILL_3__9770_ (
);

FILL FILL_0_BUFX2_insert263 (
);

FILL FILL_0__13659_ (
);

FILL FILL_0_BUFX2_insert264 (
);

FILL FILL_3__9350_ (
);

INVX1 _13944_ (
    .A(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_4446_)
);

FILL FILL_0__13239_ (
);

FILL FILL_0_BUFX2_insert265 (
);

INVX1 _13524_ (
    .A(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_4035_)
);

NAND2X1 _13104_ (
    .A(PCEn_bF$buf6),
    .B(\datapath_1.mux_pcsrc.dout [8]),
    .Y(_3701_)
);

FILL FILL_0_BUFX2_insert266 (
);

FILL FILL_0_BUFX2_insert267 (
);

FILL FILL_0_BUFX2_insert268 (
);

FILL FILL_5__9276_ (
);

FILL FILL_0_BUFX2_insert269 (
);

FILL SFILL2680x82050 (
);

FILL FILL_6__12573_ (
);

FILL FILL_0__14600_ (
);

FILL FILL_5__11986_ (
);

FILL FILL_5__11566_ (
);

FILL FILL_1__9268_ (
);

FILL FILL_5__11146_ (
);

FILL FILL_3__12180_ (
);

FILL FILL_4__7693_ (
);

FILL FILL_2__16038_ (
);

FILL FILL_4__10979_ (
);

FILL FILL_4__10559_ (
);

FILL FILL_2__11593_ (
);

FILL FILL_4__10139_ (
);

FILL FILL_2__11173_ (
);

FILL SFILL23720x73050 (
);

FILL FILL_1__10166_ (
);

FILL SFILL37960x45050 (
);

FILL FILL_4__11920_ (
);

NOR2X1 _14729_ (
    .A(_5211_),
    .B(_5214_),
    .Y(_5215_)
);

AOI21X1 _14309_ (
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .B(_4090_),
    .C(_4803_),
    .Y(_4804_)
);

FILL FILL_4__11500_ (
);

FILL FILL_0__7593_ (
);

FILL FILL_0__7173_ (
);

FILL FILL_3__10913_ (
);

FILL FILL_4__14392_ (
);

FILL FILL_0__15805_ (
);

FILL SFILL94280x17050 (
);

FILL FILL_2__8972_ (
);

FILL FILL_0__10940_ (
);

FILL FILL_3__13385_ (
);

FILL FILL_0__10520_ (
);

FILL FILL_2__8132_ (
);

FILL FILL_4__8898_ (
);

FILL FILL_4__8478_ (
);

FILL FILL_4__8058_ (
);

FILL FILL_2__12378_ (
);

FILL FILL_5__13712_ (
);

FILL SFILL8680x79050 (
);

FILL FILL_4__12705_ (
);

FILL SFILL39320x13050 (
);

FILL FILL_5__16184_ (
);

FILL FILL_3__6895_ (
);

FILL FILL_0__8378_ (
);

OAI21X1 _10649_ (
    .A(_1909_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .C(_1910_),
    .Y(_1888_[11])
);

DFFSR _10229_ (
    .Q(\datapath_1.regfile_1.regOut[26] [31]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_1628_[31])
);

FILL FILL_1__12732_ (
);

FILL FILL_4__15597_ (
);

FILL FILL_4__15177_ (
);

FILL FILL_1__12312_ (
);

FILL FILL_2__9757_ (
);

FILL FILL_2__9337_ (
);

FILL FILL_0__11725_ (
);

FILL FILL_0__11305_ (
);

FILL FILL_5__7762_ (
);

FILL FILL_5__7342_ (
);

FILL FILL_0__14197_ (
);

AOI22X1 _14482_ (
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_4973_)
);

NOR2X1 _14062_ (
    .A(_4558_),
    .B(_4561_),
    .Y(_4562_)
);

FILL FILL_5__14917_ (
);

FILL FILL_3__15951_ (
);

FILL SFILL8600x77050 (
);

FILL FILL_3__15531_ (
);

FILL FILL_3__15111_ (
);

FILL FILL_1__7754_ (
);

FILL FILL_1__7334_ (
);

FILL SFILL8680x34050 (
);

FILL FILL_2__14944_ (
);

FILL SFILL13720x71050 (
);

FILL SFILL29320x56050 (
);

FILL FILL_2__14524_ (
);

FILL FILL_2__14104_ (
);

FILL SFILL109560x51050 (
);

FILL FILL_1__13937_ (
);

FILL FILL_1__13517_ (
);

FILL SFILL84200x58050 (
);

FILL FILL_4__11097_ (
);

FILL FILL_3__8621_ (
);

FILL SFILL99480x3050 (
);

FILL FILL_3__8201_ (
);

FILL SFILL84280x15050 (
);

FILL FILL_5__8967_ (
);

FILL FILL_5__8127_ (
);

OAI22X1 _15687_ (
    .A(_5463__bF$buf0),
    .B(_4704_),
    .C(_4703_),
    .D(_5504__bF$buf4),
    .Y(_6152_)
);

AOI22X1 _15267_ (
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_5742_)
);

FILL SFILL69000x38050 (
);

FILL FILL_3__16316_ (
);

FILL FILL_1__8959_ (
);

FILL FILL_5__10837_ (
);

FILL FILL_3__11871_ (
);

FILL FILL_5__10417_ (
);

FILL FILL_1__8119_ (
);

FILL FILL_3__11451_ (
);

FILL SFILL8600x32050 (
);

FILL FILL_3__11031_ (
);

FILL FILL_2__15729_ (
);

FILL FILL_2__15309_ (
);

FILL FILL_4__6964_ (
);

FILL FILL_0__16343_ (
);

FILL FILL_2__10444_ (
);

FILL FILL_2__9090_ (
);

FILL FILL_2__10024_ (
);

FILL FILL_1__9900_ (
);

NAND2X1 _7189_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_153_)
);

FILL FILL_3__9406_ (
);

FILL SFILL84200x13050 (
);

FILL FILL_5__14670_ (
);

FILL FILL_5__14250_ (
);

FILL FILL_0__6864_ (
);

OAI21X1 _8970_ (
    .A(_1054_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .C(_1055_),
    .Y(_1043_[6])
);

DFFSR _8550_ (
    .Q(\datapath_1.regfile_1.regOut[13] [16]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_783_[16])
);

NAND2X1 _8130_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_638_)
);

FILL FILL_6__12629_ (
);

FILL FILL_4__13663_ (
);

FILL FILL_4__13243_ (
);

FILL SFILL13640x33050 (
);

INVX1 _11187_ (
    .A(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2306_)
);

FILL FILL_2__7823_ (
);

FILL FILL_3__12656_ (
);

FILL FILL_3__12236_ (
);

FILL FILL_1__13690_ (
);

FILL SFILL109480x13050 (
);

FILL FILL_1__13270_ (
);

FILL FILL_4__7749_ (
);

FILL FILL_4__7329_ (
);

FILL FILL_2__11649_ (
);

FILL SFILL38840x82050 (
);

FILL FILL_2__11229_ (
);

FILL FILL_0__12263_ (
);

FILL FILL_5__15875_ (
);

FILL FILL_5__15455_ (
);

FILL FILL_5__15035_ (
);

FILL FILL_0__7229_ (
);

NAND2X1 _9755_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1457_)
);

NAND2X1 _9335_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .Y(_1302_)
);

FILL FILL_5__10170_ (
);

FILL SFILL74280x13050 (
);

FILL FILL_4__14868_ (
);

FILL FILL_4__14448_ (
);

FILL FILL_4__14028_ (
);

FILL FILL_2__15482_ (
);

FILL FILL_2__15062_ (
);

FILL FILL_2__8608_ (
);

FILL FILL_1__14895_ (
);

FILL FILL_1__14475_ (
);

FILL SFILL99480x62050 (
);

FILL FILL_1__14055_ (
);

FILL FILL_0__13888_ (
);

INVX1 _13753_ (
    .A(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_4259_)
);

FILL FILL_0__13468_ (
);

NOR2X1 _13333_ (
    .A(_3798_),
    .B(_3857_),
    .Y(\datapath_1.regfile_1.regEn [19])
);

FILL FILL_3__14802_ (
);

FILL FILL_5__9085_ (
);

FILL FILL_6__12382_ (
);

FILL SFILL65000x4050 (
);

FILL FILL_5__11795_ (
);

FILL FILL112120x76050 (
);

FILL FILL_1__9497_ (
);

FILL FILL_5__11375_ (
);

FILL SFILL74200x11050 (
);

FILL FILL_2__16267_ (
);

FILL FILL_4__10788_ (
);

FILL FILL_4__7082_ (
);

FILL FILL_4__10368_ (
);

FILL FILL_4_BUFX2_insert90 (
);

FILL FILL_4_BUFX2_insert91 (
);

FILL FILL_4_BUFX2_insert92 (
);

FILL FILL_4_BUFX2_insert93 (
);

FILL FILL_4_BUFX2_insert94 (
);

FILL FILL_5__7818_ (
);

FILL FILL_4_BUFX2_insert95 (
);

FILL FILL_4_BUFX2_insert96 (
);

FILL FILL_1__10395_ (
);

FILL FILL_4_BUFX2_insert97 (
);

FILL FILL_4_BUFX2_insert98 (
);

FILL FILL_4_BUFX2_insert99 (
);

INVX1 _14958_ (
    .A(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_5439_)
);

AOI22X1 _14538_ (
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .B(_3891__bF$buf0),
    .C(_3998__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_5028_)
);

OAI22X1 _14118_ (
    .A(_4615_),
    .B(_3925_),
    .C(_3983__bF$buf2),
    .D(_4616_),
    .Y(_4617_)
);

FILL SFILL43720x27050 (
);

FILL SFILL28840x80050 (
);

FILL FILL_1__16201_ (
);

FILL FILL_6__13587_ (
);

FILL FILL_3__10302_ (
);

FILL FILL_0__15614_ (
);

FILL FILL_2__8781_ (
);

FILL FILL_2__8361_ (
);

FILL SFILL64200x54050 (
);

FILL FILL112120x31050 (
);

FILL FILL_2__12187_ (
);

FILL FILL_5__13941_ (
);

FILL FILL_5__13521_ (
);

FILL FILL_5__13101_ (
);

OAI21X1 _7821_ (
    .A(_471_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .C(_472_),
    .Y(_458_[7])
);

DFFSR _7401_ (
    .Q(\datapath_1.regfile_1.regOut[4] [19]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf82),
    .S(vdd),
    .D(_198_[19])
);

FILL FILL_4__12514_ (
);

FILL FILL_6__9994_ (
);

NAND2X1 _10878_ (
    .A(ALUOp[1]),
    .B(_2025_),
    .Y(_2026_)
);

FILL FILL_0__8187_ (
);

DFFSR _10458_ (
    .Q(\datapath_1.regfile_1.regOut[28] [4]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_1758_[4])
);

NAND2X1 _10038_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1605_)
);

FILL FILL_3__11927_ (
);

FILL FILL_1__12961_ (
);

FILL FILL_3__11507_ (
);

FILL SFILL113960x65050 (
);

FILL FILL112040x38050 (
);

FILL FILL_1__12121_ (
);

FILL FILL_2__9986_ (
);

FILL FILL_0__11954_ (
);

FILL FILL_2__9146_ (
);

FILL FILL_3__14399_ (
);

FILL FILL_0__11534_ (
);

FILL FILL_0__11114_ (
);

FILL FILL_5__7991_ (
);

FILL FILL_5__7571_ (
);

INVX1 _14291_ (
    .A(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_4786_)
);

FILL FILL_5__14726_ (
);

FILL FILL_3__15760_ (
);

FILL FILL_5__14306_ (
);

FILL FILL_3__15340_ (
);

NAND2X1 _8606_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_874_)
);

FILL FILL_1__7983_ (
);

FILL FILL_1__7563_ (
);

FILL FILL_4__13719_ (
);

FILL FILL_2__14753_ (
);

FILL FILL_2__14333_ (
);

FILL FILL_3__7489_ (
);

FILL FILL_3__7069_ (
);

FILL FILL_1__13746_ (
);

FILL FILL_1__13326_ (
);

FILL SFILL33720x25050 (
);

FILL FILL_3__8850_ (
);

FILL FILL_0__12739_ (
);

NAND2X1 _12604_ (
    .A(vdd),
    .B(memoryOutData[12]),
    .Y(_3449_)
);

FILL FILL_3__8010_ (
);

FILL FILL_0__12319_ (
);

FILL FILL_5__8776_ (
);

FILL FILL_5__8356_ (
);

NOR2X1 _15496_ (
    .A(_5951_),
    .B(_5965_),
    .Y(_5966_)
);

NOR3X1 _15076_ (
    .A(_5522_),
    .B(_5555_),
    .C(_5538_),
    .Y(_5556_)
);

FILL FILL_3__16125_ (
);

FILL FILL_1__8768_ (
);

FILL FILL_5__10646_ (
);

FILL FILL_1__8348_ (
);

FILL FILL_3__11680_ (
);

FILL FILL_3__11260_ (
);

FILL FILL_2__15958_ (
);

FILL FILL_2__15538_ (
);

FILL FILL_2__15118_ (
);

FILL FILL_0__16152_ (
);

FILL FILL_2__10673_ (
);

FILL FILL_2__10253_ (
);

FILL SFILL23720x68050 (
);

FILL FILL_3__9635_ (
);

FILL FILL_3_BUFX2_insert510 (
);

FILL FILL_3__9215_ (
);

FILL FILL_3_BUFX2_insert511 (
);

INVX1 _13809_ (
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_4314_)
);

FILL FILL_3_BUFX2_insert512 (
);

FILL FILL_3_BUFX2_insert513 (
);

FILL FILL_3_BUFX2_insert514 (
);

FILL FILL_3_BUFX2_insert515 (
);

FILL FILL_3_BUFX2_insert516 (
);

FILL FILL_3_BUFX2_insert517 (
);

FILL FILL_3_BUFX2_insert518 (
);

FILL FILL_3_BUFX2_insert519 (
);

FILL FILL_6__12438_ (
);

FILL FILL_4__13892_ (
);

FILL FILL_4__13472_ (
);

FILL FILL_2__7632_ (
);

FILL FILL_3__12885_ (
);

FILL FILL_3__12465_ (
);

FILL FILL_2__7212_ (
);

FILL FILL_3__12045_ (
);

FILL FILL_4__7978_ (
);

FILL FILL_4__7558_ (
);

FILL FILL_2__11878_ (
);

FILL FILL_2__11458_ (
);

FILL FILL_0__12492_ (
);

FILL FILL_2__11038_ (
);

FILL FILL_0__12072_ (
);

FILL SFILL74120x2050 (
);

FILL SFILL23720x23050 (
);

FILL FILL_5__15684_ (
);

FILL FILL_0__7878_ (
);

FILL FILL_5__15264_ (
);

NAND2X1 _9984_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1569_)
);

FILL FILL_0__7458_ (
);

DFFSR _9564_ (
    .Q(\datapath_1.regfile_1.regOut[21] [6]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf30),
    .S(vdd),
    .D(_1303_[6])
);

FILL FILL_0__7038_ (
);

INVX1 _9144_ (
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_1151_)
);

FILL FILL_1__11812_ (
);

FILL FILL_4__14677_ (
);

FILL FILL_4__14257_ (
);

FILL SFILL48920x72050 (
);

FILL FILL_2__15291_ (
);

FILL SFILL69880x70050 (
);

FILL FILL_2__8837_ (
);

FILL SFILL109160x77050 (
);

FILL FILL_0__10805_ (
);

FILL FILL_1__14284_ (
);

FILL FILL_5__6842_ (
);

FILL FILL_0_BUFX2_insert640 (
);

FILL FILL_0_BUFX2_insert641 (
);

FILL FILL_0_BUFX2_insert642 (
);

FILL FILL_0_BUFX2_insert643 (
);

FILL FILL_0_BUFX2_insert644 (
);

OAI22X1 _13982_ (
    .A(_4481_),
    .B(_3930__bF$buf1),
    .C(_3977__bF$buf3),
    .D(_4482_),
    .Y(_4483_)
);

FILL FILL_0__13697_ (
);

FILL FILL_0__13277_ (
);

FILL FILL_0_BUFX2_insert645 (
);

INVX1 _13562_ (
    .A(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_4072_)
);

INVX1 _13142_ (
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3726_)
);

FILL FILL_0_BUFX2_insert646 (
);

FILL FILL_0_BUFX2_insert647 (
);

FILL FILL_3__14611_ (
);

FILL FILL_0_BUFX2_insert648 (
);

FILL FILL_0_BUFX2_insert649 (
);

FILL SFILL48840x79050 (
);

FILL SFILL13720x66050 (
);

FILL FILL_2__13604_ (
);

FILL FILL_5__16049_ (
);

FILL SFILL109560x46050 (
);

FILL FILL_5__11184_ (
);

FILL FILL_2__16076_ (
);

FILL FILL_4__10177_ (
);

FILL FILL_0__9604_ (
);

FILL FILL_3__7701_ (
);

FILL FILL_1__15489_ (
);

FILL FILL_1__15069_ (
);

FILL FILL_5__7627_ (
);

FILL FILL_5__7207_ (
);

FILL FILL_4__16403_ (
);

INVX1 _14767_ (
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_5252_)
);

INVX1 _14347_ (
    .A(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_4841_)
);

FILL FILL_3__15816_ (
);

FILL FILL_1__16010_ (
);

FILL FILL_3__10951_ (
);

FILL FILL_1__7619_ (
);

FILL SFILL8600x27050 (
);

FILL FILL_3__10531_ (
);

FILL FILL_3__10111_ (
);

FILL FILL_2__14809_ (
);

FILL FILL_0__15843_ (
);

FILL FILL_0__15423_ (
);

FILL FILL_0__15003_ (
);

FILL SFILL13720x21050 (
);

FILL FILL_2__8590_ (
);

FILL FILL_5__12389_ (
);

FILL FILL_4__8096_ (
);

FILL FILL_3__8906_ (
);

FILL SFILL38920x70050 (
);

FILL FILL_5__13750_ (
);

FILL FILL_5__13330_ (
);

NAND2X1 _7630_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_386_)
);

FILL SFILL48440x20050 (
);

NAND2X1 _7210_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_167_)
);

FILL FILL_4__12743_ (
);

FILL FILL_4__12323_ (
);

FILL SFILL13640x28050 (
);

NAND2X1 _10687_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1936_)
);

NAND2X1 _10267_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1717_)
);

FILL FILL_2__6903_ (
);

FILL FILL_3__11736_ (
);

FILL FILL_1__12770_ (
);

FILL FILL_3__11316_ (
);

FILL FILL_1__12350_ (
);

FILL FILL_0__16208_ (
);

FILL FILL_2__9795_ (
);

FILL FILL_2__10309_ (
);

FILL FILL_0__11763_ (
);

FILL FILL_2__9375_ (
);

FILL FILL_0__11343_ (
);

FILL FILL_5__7380_ (
);

FILL FILL_6__15122_ (
);

FILL FILL_5__14955_ (
);

FILL FILL_5__14535_ (
);

FILL FILL_5__14115_ (
);

NAND2X1 _8835_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_986_)
);

DFFSR _8415_ (
    .Q(\datapath_1.regfile_1.regOut[12] [9]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf66),
    .S(vdd),
    .D(_718_[9])
);

FILL FILL_1__7372_ (
);

FILL FILL_4__13948_ (
);

FILL FILL_2__14982_ (
);

FILL FILL_4__13528_ (
);

FILL FILL_2__14562_ (
);

FILL FILL_4__13108_ (
);

FILL FILL_2__14142_ (
);

FILL FILL_3__7298_ (
);

FILL SFILL44120x1050 (
);

FILL FILL112200x64050 (
);

FILL FILL_1__13975_ (
);

FILL SFILL99480x57050 (
);

FILL FILL_1__13555_ (
);

FILL FILL_1__13135_ (
);

FILL SFILL44040x6050 (
);

FILL FILL_0__12968_ (
);

NAND2X1 _12833_ (
    .A(vdd),
    .B(\datapath_1.rd1 [3]),
    .Y(_3561_)
);

NAND2X1 _12413_ (
    .A(MemToReg_bF$buf2),
    .B(\datapath_1.Data [23]),
    .Y(_3341_)
);

FILL FILL_0__12128_ (
);

FILL FILL_5__8585_ (
);

FILL FILL_6__11042_ (
);

FILL FILL_3__16354_ (
);

FILL FILL_1__8997_ (
);

FILL FILL_5__10875_ (
);

FILL FILL_1__8577_ (
);

FILL FILL_5__10035_ (
);

FILL FILL_2__15767_ (
);

FILL FILL_2__15347_ (
);

FILL FILL_0__16381_ (
);

FILL FILL_2__10062_ (
);

FILL SFILL99480x12050 (
);

FILL FILL_3__9864_ (
);

NOR2X1 _13618_ (
    .A(_4126_),
    .B(_4123_),
    .Y(_4127_)
);

FILL FILL_3__9024_ (
);

FILL SFILL28840x75050 (
);

FILL FILL_1__15701_ (
);

FILL FILL_4__13281_ (
);

FILL SFILL33800x58050 (
);

FILL FILL_2__7861_ (
);

FILL FILL_2__7441_ (
);

FILL FILL_3__12274_ (
);

FILL FILL112120x26050 (
);

FILL FILL_4__7367_ (
);

FILL FILL_2__11687_ (
);

FILL FILL_2__11267_ (
);

FILL FILL_5__12601_ (
);

BUFX2 _6901_ (
    .A(_2_[31]),
    .Y(memoryWriteData[31])
);

FILL FILL_5__15493_ (
);

FILL FILL_5__15073_ (
);

FILL FILL_0__7687_ (
);

INVX1 _9793_ (
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_1482_)
);

INVX1 _9373_ (
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_1263_)
);

FILL FILL_4__14486_ (
);

FILL FILL_1__11621_ (
);

FILL SFILL28840x30050 (
);

FILL FILL_4__14066_ (
);

FILL FILL_1__11201_ (
);

FILL FILL_2__8646_ (
);

FILL FILL_3__13899_ (
);

FILL FILL_2__8226_ (
);

FILL FILL_0__10614_ (
);

FILL FILL_3__13479_ (
);

FILL FILL_1__14093_ (
);

FILL SFILL89880x24050 (
);

NAND2X1 _13791_ (
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .B(_4102_),
    .Y(_4296_)
);

NOR2X1 _13371_ (
    .A(\datapath_1.PCJump [18]),
    .B(_3878_),
    .Y(_3883_)
);

FILL FILL_0__13086_ (
);

FILL FILL_5__13806_ (
);

FILL FILL_3__14840_ (
);

FILL FILL_3__14420_ (
);

FILL FILL_3__14000_ (
);

FILL FILL_4__9933_ (
);

FILL FILL_4__9513_ (
);

FILL FILL_2__13833_ (
);

FILL FILL_3__6989_ (
);

FILL FILL_2__13413_ (
);

FILL FILL_5__16278_ (
);

FILL FILL_1__12826_ (
);

FILL FILL_1__12406_ (
);

FILL SFILL18840x73050 (
);

FILL FILL_3__7930_ (
);

FILL FILL_0__9413_ (
);

FILL FILL_0__11819_ (
);

FILL FILL_1__15298_ (
);

FILL FILL_5__7856_ (
);

FILL FILL_5__7436_ (
);

FILL FILL_4__16212_ (
);

NOR2X1 _14996_ (
    .A(\datapath_1.PCJump [23]),
    .B(_5475_),
    .Y(_5476_)
);

INVX1 _14576_ (
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_5065_)
);

FILL SFILL13800x3050 (
);

INVX1 _14156_ (
    .A(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_4654_)
);

FILL FILL_3__15625_ (
);

FILL FILL_3__15205_ (
);

FILL SFILL13720x8050 (
);

FILL FILL_1__7848_ (
);

FILL FILL_1__7428_ (
);

FILL FILL_3__10760_ (
);

FILL FILL_2__14618_ (
);

FILL FILL_0__15652_ (
);

FILL FILL_0__15232_ (
);

FILL FILL_5__12198_ (
);

FILL FILL_3__8715_ (
);

FILL FILL_4__12972_ (
);

FILL FILL_6__11518_ (
);

FILL FILL_4__12132_ (
);

NAND2X1 _10496_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1829_)
);

DFFSR _10076_ (
    .Q(\datapath_1.regfile_1.regOut[25] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_1563_[6])
);

FILL FILL_3__11965_ (
);

FILL FILL_3__11545_ (
);

FILL FILL_3__11125_ (
);

FILL FILL_0__16017_ (
);

NOR2X1 _16302_ (
    .A(_6748_),
    .B(_6750_),
    .Y(_6751_)
);

FILL FILL_2__10958_ (
);

FILL FILL_0__11992_ (
);

FILL FILL_2__10538_ (
);

FILL FILL_0__11572_ (
);

FILL FILL_2__10118_ (
);

FILL FILL_0__11152_ (
);

FILL SFILL23720x18050 (
);

FILL FILL_5__14764_ (
);

FILL FILL_0__6958_ (
);

FILL FILL_5__14344_ (
);

FILL SFILL103960x13050 (
);

INVX1 _8644_ (
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_899_)
);

FILL SFILL69080x82050 (
);

INVX1 _8224_ (
    .A(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_680_)
);

FILL FILL_1__7181_ (
);

FILL FILL_4__13757_ (
);

FILL SFILL48920x67050 (
);

FILL FILL_4__13337_ (
);

FILL FILL_2__14791_ (
);

FILL FILL_2__14371_ (
);

FILL FILL_1__13784_ (
);

FILL FILL_1__13364_ (
);

FILL FILL_0__12777_ (
);

INVX1 _12642_ (
    .A(\datapath_1.Data [25]),
    .Y(_3474_)
);

FILL FILL_0__12357_ (
);

NAND3X1 _12222_ (
    .A(_3203_),
    .B(_3204_),
    .C(_3205_),
    .Y(\datapath_1.alu_1.ALUInB [1])
);

FILL FILL_5__8394_ (
);

FILL SFILL109240x20050 (
);

FILL FILL_6__11691_ (
);

FILL FILL_5__15969_ (
);

FILL FILL_5__15549_ (
);

FILL FILL_5__15129_ (
);

FILL FILL_3__16163_ (
);

INVX1 _9849_ (
    .A(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_1499_)
);

OAI21X1 _9429_ (
    .A(_1299_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1300_),
    .Y(_1238_[31])
);

FILL FILL_5__10684_ (
);

OAI21X1 _9009_ (
    .A(_1080_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .C(_1081_),
    .Y(_1043_[19])
);

FILL FILL_5__10264_ (
);

FILL FILL_1__8386_ (
);

FILL FILL_2__15996_ (
);

FILL FILL_2__15576_ (
);

FILL FILL_2__15156_ (
);

FILL FILL_0__16190_ (
);

FILL SFILL48920x22050 (
);

FILL FILL_2__10291_ (
);

FILL FILL_1__14989_ (
);

FILL FILL_1__14569_ (
);

FILL FILL_1__14149_ (
);

FILL FILL_4__15903_ (
);

FILL FILL_3__9673_ (
);

NOR2X1 _13847_ (
    .A(_4347_),
    .B(_4350_),
    .Y(_4351_)
);

FILL FILL_3__9253_ (
);

NAND2X1 _13427_ (
    .A(_3938_),
    .B(_3927_),
    .Y(_3939_)
);

OAI21X1 _13007_ (
    .A(_3655_),
    .B(vdd),
    .C(_3656_),
    .Y(_3620_[18])
);

FILL FILL_5__9599_ (
);

FILL FILL_1__15930_ (
);

FILL FILL_1__15510_ (
);

FILL FILL_4__13090_ (
);

FILL FILL_0__14923_ (
);

FILL FILL_0__14503_ (
);

FILL SFILL48840x29050 (
);

FILL SFILL13720x16050 (
);

FILL FILL_5__11889_ (
);

FILL FILL_2__7670_ (
);

FILL FILL_5__11469_ (
);

FILL FILL_2__7250_ (
);

FILL FILL_5__11049_ (
);

FILL FILL_3__12083_ (
);

FILL FILL_4__7596_ (
);

FILL FILL_4__7176_ (
);

FILL FILL_2__11496_ (
);

FILL SFILL38920x65050 (
);

FILL FILL_2__11076_ (
);

FILL FILL_5__12830_ (
);

FILL FILL_5__12410_ (
);

FILL FILL_1__10489_ (
);

FILL FILL_1__10069_ (
);

FILL FILL_4__11823_ (
);

FILL FILL_4__11403_ (
);

FILL FILL_0__7496_ (
);

FILL FILL_6__8883_ (
);

FILL FILL_0__7076_ (
);

DFFSR _9182_ (
    .Q(\datapath_1.regfile_1.regOut[18] [8]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf44),
    .S(vdd),
    .D(_1108_[8])
);

FILL FILL_3__10816_ (
);

FILL FILL_1__11850_ (
);

FILL FILL_4__14295_ (
);

FILL FILL_1__11430_ (
);

FILL FILL_1__11010_ (
);

FILL FILL_0__15708_ (
);

FILL FILL_2__8875_ (
);

FILL FILL_2__8455_ (
);

FILL FILL_0__10423_ (
);

FILL FILL_3__13288_ (
);

FILL FILL_0__10003_ (
);

FILL FILL_5__6880_ (
);

FILL SFILL3560x64050 (
);

DFFSR _13180_ (
    .Q(\datapath_1.mux_iord.din0 [5]),
    .CLK(clk_bF$buf71),
    .R(rst_bF$buf62),
    .S(vdd),
    .D(_3685_[5])
);

FILL FILL_5__13615_ (
);

DFFSR _7915_ (
    .Q(\datapath_1.regfile_1.regOut[8] [21]),
    .CLK(clk_bF$buf29),
    .R(rst_bF$buf2),
    .S(vdd),
    .D(_458_[21])
);

FILL SFILL38920x20050 (
);

FILL SFILL104440x81050 (
);

FILL FILL_1__6872_ (
);

FILL FILL_4__9742_ (
);

FILL FILL_4__12608_ (
);

FILL FILL_2__13642_ (
);

FILL FILL_2__13222_ (
);

FILL FILL_5__16087_ (
);

FILL FILL_6__9668_ (
);

FILL FILL112200x59050 (
);

FILL FILL_1__12635_ (
);

FILL FILL_1__12215_ (
);

FILL FILL_0__9642_ (
);

OAI21X1 _11913_ (
    .A(_2982_),
    .B(IorD_bF$buf0),
    .C(_2983_),
    .Y(_1_[8])
);

FILL FILL_0__9222_ (
);

FILL FILL_0__11628_ (
);

FILL FILL_0__11208_ (
);

FILL FILL_5__7245_ (
);

FILL FILL_4__16021_ (
);

INVX1 _14385_ (
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_4878_)
);

FILL FILL_3__15854_ (
);

FILL FILL_3__15434_ (
);

FILL FILL_3__15014_ (
);

FILL SFILL28920x63050 (
);

FILL SFILL3080x57050 (
);

FILL FILL_1__7237_ (
);

FILL FILL_2__14847_ (
);

FILL FILL_6_BUFX2_insert403 (
);

FILL FILL_0__15881_ (
);

FILL FILL_2__14427_ (
);

FILL FILL_2__14007_ (
);

FILL FILL_0__15461_ (
);

FILL FILL_0__15041_ (
);

FILL FILL_6_BUFX2_insert408 (
);

FILL FILL112200x14050 (
);

FILL FILL_3__8524_ (
);

FILL FILL_3__8104_ (
);

FILL SFILL3480x26050 (
);

FILL FILL_4__12781_ (
);

FILL FILL_4__12361_ (
);

FILL FILL_3__16219_ (
);

FILL FILL_2__6941_ (
);

FILL FILL_3__11774_ (
);

FILL FILL_5__9811_ (
);

FILL FILL_3__11354_ (
);

FILL FILL_4__6867_ (
);

FILL FILL_0__16246_ (
);

NAND3X1 _16111_ (
    .A(_6557_),
    .B(_6564_),
    .C(_6559_),
    .Y(_6565_)
);

FILL FILL_2__10767_ (
);

FILL FILL_0__11381_ (
);

FILL FILL_1__9803_ (
);

FILL FILL_3__9729_ (
);

FILL FILL_5__14993_ (
);

FILL FILL_5__14573_ (
);

FILL FILL_5__14153_ (
);

INVX1 _8873_ (
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_1011_)
);

INVX1 _8453_ (
    .A(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_792_)
);

DFFSR _8033_ (
    .Q(\datapath_1.regfile_1.regOut[9] [11]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_523_[11])
);

FILL FILL_4__13986_ (
);

FILL FILL_1__10701_ (
);

FILL FILL_4__13566_ (
);

FILL FILL_4__13146_ (
);

FILL FILL_2__14180_ (
);

FILL FILL_2__7726_ (
);

FILL FILL_3__12979_ (
);

FILL FILL_2__7306_ (
);

FILL FILL_1__13593_ (
);

FILL FILL_3__12139_ (
);

FILL FILL_1__13173_ (
);

FILL FILL_0__12586_ (
);

INVX1 _12871_ (
    .A(\datapath_1.a [16]),
    .Y(_3586_)
);

INVX1 _12451_ (
    .A(ALUOut[4]),
    .Y(_3367_)
);

FILL FILL_0__12166_ (
);

NAND3X1 _12031_ (
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[11]),
    .C(_3032__bF$buf3),
    .Y(_3069_)
);

FILL FILL_3__13920_ (
);

FILL FILL_6__16365_ (
);

FILL FILL_3__13500_ (
);

FILL FILL_5_BUFX2_insert420 (
);

FILL FILL_5_BUFX2_insert421 (
);

FILL FILL_5__15778_ (
);

FILL FILL_2__12913_ (
);

FILL FILL_5__15358_ (
);

FILL FILL_5_BUFX2_insert422 (
);

FILL FILL_5_BUFX2_insert423 (
);

FILL FILL_3__16392_ (
);

FILL FILL_5_BUFX2_insert424 (
);

OAI21X1 _9658_ (
    .A(_1411_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1412_),
    .Y(_1368_[22])
);

FILL FILL_5_BUFX2_insert425 (
);

OAI21X1 _9238_ (
    .A(_1192_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .C(_1193_),
    .Y(_1173_[10])
);

FILL FILL_5_BUFX2_insert426 (
);

FILL FILL_5__10493_ (
);

FILL FILL_1__8195_ (
);

FILL FILL_5_BUFX2_insert427 (
);

FILL FILL_1__11906_ (
);

FILL FILL_5_BUFX2_insert428 (
);

FILL FILL_5_BUFX2_insert429 (
);

FILL FILL_2__15385_ (
);

FILL FILL_0__8913_ (
);

FILL FILL_1__14798_ (
);

FILL FILL_1__14378_ (
);

FILL FILL_5__6936_ (
);

FILL FILL_4__15712_ (
);

FILL FILL_3__9482_ (
);

INVX1 _13656_ (
    .A(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_4164_)
);

OAI21X1 _13236_ (
    .A(_3773_),
    .B(_3776_),
    .C(_3778_),
    .Y(_3779_)
);

FILL FILL_3__14705_ (
);

FILL FILL_1__6928_ (
);

FILL FILL_6__12285_ (
);

FILL FILL_0__14732_ (
);

FILL FILL_0__14312_ (
);

FILL FILL_5__11698_ (
);

FILL FILL_5__11278_ (
);

FILL FILL_2_BUFX2_insert550 (
);

FILL FILL_1__10298_ (
);

FILL FILL_2_BUFX2_insert551 (
);

FILL FILL_2_BUFX2_insert552 (
);

FILL FILL_2_BUFX2_insert553 (
);

FILL FILL_2_BUFX2_insert554 (
);

FILL FILL_4__11632_ (
);

FILL FILL_4__11212_ (
);

FILL FILL_2_BUFX2_insert555 (
);

FILL FILL_2_BUFX2_insert556 (
);

FILL FILL_2_BUFX2_insert557 (
);

FILL FILL_2_BUFX2_insert558 (
);

FILL FILL_2_BUFX2_insert559 (
);

FILL FILL_1__16104_ (
);

FILL FILL_3__10625_ (
);

FILL FILL_0__15937_ (
);

FILL FILL_0__15517_ (
);

OAI22X1 _15802_ (
    .A(_5472__bF$buf2),
    .B(_4835_),
    .C(_4832_),
    .D(_5526__bF$buf4),
    .Y(_6264_)
);

FILL FILL_0__10652_ (
);

FILL FILL_2__8264_ (
);

FILL FILL_3__13097_ (
);

FILL FILL_0__10232_ (
);

FILL FILL_6__14851_ (
);

FILL FILL_6__14431_ (
);

FILL FILL_5__13844_ (
);

FILL FILL_5__13424_ (
);

FILL FILL_5__13004_ (
);

INVX1 _7724_ (
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_428_)
);

INVX1 _7304_ (
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_209_)
);

FILL FILL_4__9551_ (
);

FILL FILL_4__12837_ (
);

FILL FILL_4__9131_ (
);

FILL FILL_2__13871_ (
);

FILL FILL_4__12417_ (
);

FILL FILL_2__13451_ (
);

FILL FILL_2__13031_ (
);

FILL FILL_1__12864_ (
);

FILL FILL_1__12444_ (
);

FILL FILL_1__12024_ (
);

FILL FILL_0__9871_ (
);

FILL FILL_2__9889_ (
);

FILL FILL_0__11857_ (
);

FILL FILL_2__9469_ (
);

FILL FILL_0__9031_ (
);

FILL FILL_0__11437_ (
);

AOI22X1 _11722_ (
    .A(_2191_),
    .B(_2481__bF$buf3),
    .C(_2341__bF$buf1),
    .D(_2192_),
    .Y(_2820_)
);

FILL SFILL114520x71050 (
);

FILL FILL_0__11017_ (
);

NAND2X1 _11302_ (
    .A(_2420_),
    .B(_2417_),
    .Y(_2421_)
);

FILL FILL_5__7474_ (
);

FILL FILL_5__7054_ (
);

FILL FILL_4__16250_ (
);

NAND3X1 _14194_ (
    .A(_4682_),
    .B(_4690_),
    .C(_4683_),
    .Y(_4691_)
);

FILL FILL_5__14629_ (
);

FILL FILL_3__15663_ (
);

FILL FILL_5__14209_ (
);

DFFSR _8929_ (
    .Q(\datapath_1.regfile_1.regOut[16] [11]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_978_[11])
);

FILL FILL_3__15243_ (
);

OAI21X1 _8509_ (
    .A(_828_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .C(_829_),
    .Y(_783_[23])
);

FILL FILL_1__7886_ (
);

FILL FILL_1__7466_ (
);

FILL FILL_1__7046_ (
);

FILL SFILL69080x32050 (
);

FILL FILL_2__14656_ (
);

FILL FILL_0__15690_ (
);

FILL FILL_2__14236_ (
);

FILL FILL_0__15270_ (
);

FILL FILL_1__13649_ (
);

FILL FILL_1__13229_ (
);

FILL FILL_1_BUFX2_insert570 (
);

FILL FILL_1_BUFX2_insert571 (
);

FILL FILL_3__8753_ (
);

FILL FILL_3__8333_ (
);

FILL FILL_1_BUFX2_insert572 (
);

DFFSR _12927_ (
    .Q(\datapath_1.a [8]),
    .CLK(clk_bF$buf102),
    .R(rst_bF$buf38),
    .S(vdd),
    .D(_3555_[8])
);

FILL FILL_1_BUFX2_insert573 (
);

OAI21X1 _12507_ (
    .A(_3403_),
    .B(vdd),
    .C(_3404_),
    .Y(_3360_[22])
);

FILL FILL_1_BUFX2_insert574 (
);

FILL FILL_1_BUFX2_insert575 (
);

FILL FILL_1_BUFX2_insert576 (
);

FILL FILL_1_BUFX2_insert577 (
);

FILL FILL_5__8259_ (
);

FILL FILL_1_BUFX2_insert578 (
);

FILL FILL_1_BUFX2_insert579 (
);

FILL FILL_4__12590_ (
);

NAND3X1 _15399_ (
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5871_)
);

FILL FILL_4__12170_ (
);

FILL FILL_3__16028_ (
);

FILL FILL_5__10969_ (
);

FILL FILL_5__10549_ (
);

FILL FILL_5__9620_ (
);

FILL FILL_5__10129_ (
);

FILL FILL_3__11583_ (
);

FILL SFILL38120x77050 (
);

FILL FILL_3__11163_ (
);

FILL SFILL59080x75050 (
);

NAND2X1 _16340_ (
    .A(gnd),
    .B(gnd),
    .Y(_6781_)
);

FILL FILL_0__16055_ (
);

FILL FILL_2__10996_ (
);

FILL FILL_2__10576_ (
);

FILL FILL_2__10156_ (
);

FILL FILL_0__11190_ (
);

FILL FILL_5__11910_ (
);

FILL FILL_1__9612_ (
);

FILL FILL_3__9538_ (
);

FILL FILL_4__10903_ (
);

FILL FILL_3__9118_ (
);

FILL SFILL3640x52050 (
);

FILL FILL_0__6996_ (
);

FILL FILL_5__14382_ (
);

FILL FILL_6__7963_ (
);

DFFSR _8682_ (
    .Q(\datapath_1.regfile_1.regOut[14] [20]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_848_[20])
);

OAI21X1 _8262_ (
    .A(_704_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .C(_705_),
    .Y(_653_[26])
);

FILL FILL_1__10930_ (
);

FILL FILL_4__13795_ (
);

FILL FILL_1__10510_ (
);

FILL FILL_4__13375_ (
);

FILL FILL_2__7955_ (
);

FILL FILL_3__12788_ (
);

BUFX2 BUFX2_insert240 (
    .A(_5545_),
    .Y(_5545__bF$buf2)
);

FILL FILL_3__12368_ (
);

FILL FILL_2__7115_ (
);

BUFX2 BUFX2_insert241 (
    .A(_5545_),
    .Y(_5545__bF$buf1)
);

BUFX2 BUFX2_insert242 (
    .A(_5545_),
    .Y(_5545__bF$buf0)
);

FILL SFILL59000x73050 (
);

BUFX2 BUFX2_insert243 (
    .A(_3972_),
    .Y(_3972__bF$buf3)
);

BUFX2 BUFX2_insert244 (
    .A(_3972_),
    .Y(_3972__bF$buf2)
);

BUFX2 BUFX2_insert245 (
    .A(_3972_),
    .Y(_3972__bF$buf1)
);

BUFX2 BUFX2_insert246 (
    .A(_3972_),
    .Y(_3972__bF$buf0)
);

FILL SFILL38120x32050 (
);

BUFX2 BUFX2_insert247 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf7)
);

BUFX2 BUFX2_insert248 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf6)
);

FILL SFILL59080x30050 (
);

DFFSR _12680_ (
    .Q(\datapath_1.Data [17]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3425_[17])
);

FILL FILL_0__12395_ (
);

BUFX2 BUFX2_insert249 (
    .A(RegWrite),
    .Y(RegWrite_bF$buf5)
);

NAND3X1 _12260_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [13]),
    .C(_3198__bF$buf3),
    .Y(_3234_)
);

FILL SFILL104440x76050 (
);

FILL FILL_4__8822_ (
);

FILL FILL_4__8402_ (
);

FILL FILL_2__12722_ (
);

FILL FILL_5__15587_ (
);

FILL FILL_2__12302_ (
);

FILL FILL_5__15167_ (
);

FILL FILL_6__8748_ (
);

OAI21X1 _9887_ (
    .A(_1523_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .C(_1524_),
    .Y(_1498_[13])
);

OAI21X1 _9467_ (
    .A(_1304_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .C(_1305_),
    .Y(_1303_[1])
);

DFFSR _9047_ (
    .Q(\datapath_1.regfile_1.regOut[17] [1]),
    .CLK(clk_bF$buf69),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_1043_[1])
);

FILL FILL_1__11715_ (
);

FILL FILL_2__15194_ (
);

FILL FILL_0__8722_ (
);

FILL FILL_0__10708_ (
);

FILL FILL_1__14187_ (
);

FILL FILL_6__14907_ (
);

FILL FILL_4__15941_ (
);

FILL FILL_4__15521_ (
);

FILL FILL_4__15101_ (
);

FILL SFILL83960x10050 (
);

NAND3X1 _13885_ (
    .A(_4387_),
    .B(_4388_),
    .C(_4384_),
    .Y(_4389_)
);

FILL FILL_3__9291_ (
);

FILL SFILL49080x73050 (
);

NAND3X1 _13465_ (
    .A(_3898_),
    .B(_3888_),
    .C(_3879_),
    .Y(_3977_)
);

NAND2X1 _13045_ (
    .A(vdd),
    .B(\datapath_1.rd2 [31]),
    .Y(_3682_)
);

FILL FILL_3__14934_ (
);

FILL FILL_3__14514_ (
);

FILL SFILL3560x14050 (
);

FILL FILL_4__9607_ (
);

FILL FILL_2__13927_ (
);

FILL SFILL104440x31050 (
);

FILL FILL_0__14961_ (
);

FILL FILL_2__13507_ (
);

FILL FILL_0__14541_ (
);

FILL FILL_0__14121_ (
);

FILL FILL_5__11087_ (
);

FILL FILL_2__16399_ (
);

FILL SFILL28520x44050 (
);

FILL FILL_0__9927_ (
);

FILL FILL_0__9507_ (
);

FILL FILL_3__7604_ (
);

FILL FILL_4__16306_ (
);

FILL SFILL18600x80050 (
);

FILL FILL_6__10827_ (
);

FILL FILL_4__11861_ (
);

FILL FILL_4__11441_ (
);

FILL FILL_4__11021_ (
);

FILL FILL_3__15719_ (
);

FILL FILL_1__16333_ (
);

FILL FILL_3__10434_ (
);

FILL FILL_3__10014_ (
);

FILL SFILL28920x13050 (
);

FILL FILL_0__15746_ (
);

FILL FILL_0__15326_ (
);

OAI22X1 _15611_ (
    .A(_5504__bF$buf3),
    .B(_4664_),
    .C(_5527__bF$buf0),
    .D(_4638_),
    .Y(_6077_)
);

FILL FILL_0__10881_ (
);

FILL FILL_2__8493_ (
);

FILL FILL_2__8073_ (
);

FILL FILL_0__10041_ (
);

FILL SFILL115240x7050 (
);

FILL FILL_5__13653_ (
);

FILL FILL_5__13233_ (
);

INVX1 _7953_ (
    .A(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_540_)
);

DFFSR _7533_ (
    .Q(\datapath_1.regfile_1.regOut[5] [23]),
    .CLK(clk_bF$buf80),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_263_[23])
);

OAI21X1 _7113_ (
    .A(_121_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_122_),
    .Y(_68_[27])
);

FILL FILL_4__9780_ (
);

FILL FILL_4__9360_ (
);

FILL FILL_4__12646_ (
);

FILL FILL_2__13680_ (
);

FILL FILL_4__12226_ (
);

FILL FILL_2__13260_ (
);

FILL FILL_6__9286_ (
);

FILL FILL_3__11639_ (
);

FILL FILL_3__11219_ (
);

FILL FILL_1__12253_ (
);

FILL FILL_0__9680_ (
);

FILL SFILL79160x67050 (
);

FILL FILL_2__9278_ (
);

NAND2X1 _11951_ (
    .A(IorD_bF$buf5),
    .B(ALUOut[21]),
    .Y(_3009_)
);

FILL FILL_0__9260_ (
);

FILL FILL_0__11666_ (
);

FILL FILL_0__11246_ (
);

AOI21X1 _11531_ (
    .A(_2433_),
    .B(_2620_),
    .C(_2641_),
    .Y(_2642_)
);

NOR2X1 _11111_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2230_)
);

FILL FILL_6__15025_ (
);

FILL FILL_6__10160_ (
);

FILL FILL_5__14858_ (
);

FILL FILL_3__15892_ (
);

FILL FILL_5__14438_ (
);

FILL FILL_5__14018_ (
);

FILL FILL_3__15472_ (
);

OAI21X1 _8738_ (
    .A(_940_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_941_),
    .Y(_913_[14])
);

FILL FILL_3__15052_ (
);

OAI21X1 _8318_ (
    .A(_721_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .C(_722_),
    .Y(_718_[2])
);

FILL FILL_1__7695_ (
);

FILL FILL_2__14885_ (
);

FILL FILL_2__14465_ (
);

FILL FILL_2__14045_ (
);

FILL SFILL94360x42050 (
);

FILL FILL_1__13878_ (
);

FILL FILL_1__13458_ (
);

FILL FILL_1__13038_ (
);

FILL FILL_3__8982_ (
);

FILL FILL_3__8142_ (
);

OAI21X1 _12736_ (
    .A(_3515_),
    .B(IRWrite_bF$buf3),
    .C(_3516_),
    .Y(_3490_[13])
);

NAND3X1 _12316_ (
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf4),
    .Y(_3276_)
);

FILL FILL_5__8488_ (
);

FILL SFILL79160x22050 (
);

FILL FILL_5__8068_ (
);

FILL FILL_0__13812_ (
);

FILL FILL_3__16257_ (
);

FILL FILL_5__10778_ (
);

FILL FILL_5__10358_ (
);

FILL FILL_3__11392_ (
);

FILL FILL_0__16284_ (
);

FILL SFILL18840x18050 (
);

FILL FILL_2__10385_ (
);

FILL FILL_1__9421_ (
);

FILL FILL_1__9001_ (
);

FILL FILL_3__9767_ (
);

FILL FILL_3__9347_ (
);

FILL FILL_5__14191_ (
);

OAI21X1 _8491_ (
    .A(_816_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_817_),
    .Y(_783_[17])
);

FILL FILL_1__15604_ (
);

OAI21X1 _8071_ (
    .A(_597_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_598_),
    .Y(_588_[5])
);

FILL FILL_2__7764_ (
);

FILL FILL_3__12597_ (
);

FILL FILL_2__7344_ (
);

FILL FILL_3__12177_ (
);

FILL FILL_5__12504_ (
);

FILL SFILL84360x40050 (
);

FILL FILL_4__8631_ (
);

FILL FILL_5_BUFX2_insert800 (
);

FILL FILL_4__11917_ (
);

FILL FILL_4__8211_ (
);

FILL FILL_5_BUFX2_insert801 (
);

FILL FILL_2__12951_ (
);

FILL FILL_5__15396_ (
);

FILL FILL_2__12531_ (
);

FILL FILL_5_BUFX2_insert802 (
);

FILL FILL_2__12111_ (
);

FILL FILL_5_BUFX2_insert803 (
);

FILL FILL_5_BUFX2_insert804 (
);

DFFSR _9696_ (
    .Q(\datapath_1.regfile_1.regOut[22] [10]),
    .CLK(clk_bF$buf27),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1368_[10])
);

NAND2X1 _9276_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1219_)
);

FILL FILL_5_BUFX2_insert805 (
);

FILL FILL_5_BUFX2_insert806 (
);

FILL FILL_5_BUFX2_insert807 (
);

FILL FILL_1__11944_ (
);

FILL FILL_5_BUFX2_insert808 (
);

FILL FILL_5_BUFX2_insert809 (
);

FILL FILL_4__14389_ (
);

FILL FILL_1__11524_ (
);

FILL FILL_1__11104_ (
);

FILL FILL_2__8969_ (
);

FILL FILL_0__8951_ (
);

FILL FILL_0__10937_ (
);

FILL FILL_0__8531_ (
);

FILL SFILL114520x66050 (
);

FILL FILL_0__8111_ (
);

INVX1 _10802_ (
    .A(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_1992_)
);

FILL FILL_0__10517_ (
);

FILL FILL_2__8129_ (
);

FILL FILL_5__6974_ (
);

FILL FILL_4__15750_ (
);

FILL FILL_4__15330_ (
);

INVX1 _13694_ (
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_4201_)
);

NAND3X1 _13274_ (
    .A(RegWrite_bF$buf0),
    .B(_3814_),
    .C(_3808_),
    .Y(_3815_)
);

FILL FILL_2__9910_ (
);

FILL FILL_5__13709_ (
);

FILL FILL_3__14743_ (
);

FILL FILL_3__14323_ (
);

FILL FILL_1__6966_ (
);

FILL FILL_4__9416_ (
);

FILL SFILL69080x27050 (
);

FILL FILL_2__13736_ (
);

FILL FILL_2__13316_ (
);

FILL FILL_0__14770_ (
);

FILL FILL_0__14350_ (
);

FILL FILL_1__12729_ (
);

FILL FILL_1__12309_ (
);

FILL FILL_0__9736_ (
);

FILL FILL_3__7833_ (
);

FILL FILL_5__7759_ (
);

FILL FILL_5__7339_ (
);

FILL FILL_2_BUFX2_insert930 (
);

FILL FILL_4__16115_ (
);

FILL FILL_2_BUFX2_insert931 (
);

FILL FILL_2_BUFX2_insert932 (
);

FILL FILL_6__10636_ (
);

FILL FILL_2_BUFX2_insert933 (
);

INVX1 _14899_ (
    .A(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_5381_)
);

OAI22X1 _14479_ (
    .A(_4969_),
    .B(_3931__bF$buf2),
    .C(_3983__bF$buf4),
    .D(_4968_),
    .Y(_4970_)
);

FILL FILL_2_BUFX2_insert934 (
);

FILL FILL_4__11670_ (
);

FILL FILL_2_BUFX2_insert935 (
);

INVX1 _14059_ (
    .A(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_4559_)
);

FILL FILL_4__11250_ (
);

FILL FILL_2_BUFX2_insert936 (
);

FILL FILL_3__15948_ (
);

FILL SFILL3720x40050 (
);

FILL FILL_3__15528_ (
);

FILL FILL_2_BUFX2_insert937 (
);

FILL FILL_2_BUFX2_insert938 (
);

FILL FILL_3__15108_ (
);

FILL FILL_2_BUFX2_insert939 (
);

FILL FILL_1__16142_ (
);

FILL FILL_3__10663_ (
);

FILL FILL_5__8700_ (
);

FILL FILL_3__10243_ (
);

FILL FILL_0__15975_ (
);

FILL FILL_0__15555_ (
);

NAND2X1 _15840_ (
    .A(_6294_),
    .B(_6300_),
    .Y(_6301_)
);

NOR2X1 _15420_ (
    .A(_5890_),
    .B(_5549__bF$buf0),
    .Y(_5891_)
);

FILL FILL_0__15135_ (
);

NAND3X1 _15000_ (
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5462_),
    .C(_5476_),
    .Y(_5480_)
);

FILL FILL_0__10690_ (
);

FILL FILL_0__10270_ (
);

FILL FILL_3__8618_ (
);

FILL SFILL3640x47050 (
);

FILL FILL_5__13882_ (
);

FILL FILL_5__13462_ (
);

FILL FILL_5__13042_ (
);

OAI21X1 _7762_ (
    .A(_452_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_453_),
    .Y(_393_[30])
);

OAI21X1 _7342_ (
    .A(_233_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_234_),
    .Y(_198_[18])
);

FILL SFILL104520x64050 (
);

FILL SFILL43880x54050 (
);

FILL FILL_4__12875_ (
);

FILL FILL_4__12455_ (
);

FILL FILL_4__12035_ (
);

FILL FILL_6__9095_ (
);

OAI21X1 _10399_ (
    .A(_1783_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .C(_1784_),
    .Y(_1758_[13])
);

FILL FILL_5__9905_ (
);

FILL FILL_3__11868_ (
);

FILL FILL_3__11448_ (
);

FILL SFILL59000x68050 (
);

FILL FILL_1__12482_ (
);

FILL FILL_3__11028_ (
);

FILL FILL_1__12062_ (
);

AOI22X1 _16205_ (
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [29]),
    .C(\datapath_1.regfile_1.regOut[11] [29]),
    .D(_5496_),
    .Y(_6656_)
);

FILL SFILL59080x25050 (
);

FILL FILL_0__11895_ (
);

FILL FILL_2__9087_ (
);

OAI21X1 _11760_ (
    .A(_2138_),
    .B(_2139_),
    .C(_2851_),
    .Y(_2855_)
);

FILL FILL_0__11475_ (
);

AOI21X1 _11340_ (
    .A(_2110_),
    .B(_2457_),
    .C(_2458_),
    .Y(_2459_)
);

FILL FILL_0__11055_ (
);

FILL FILL_6__15674_ (
);

FILL FILL_5__7092_ (
);

FILL FILL_2__11802_ (
);

FILL FILL_5__14667_ (
);

FILL FILL_5__14247_ (
);

FILL FILL_3__15281_ (
);

OAI21X1 _8967_ (
    .A(_1052_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .C(_1053_),
    .Y(_1043_[5])
);

DFFSR _8547_ (
    .Q(\datapath_1.regfile_1.regOut[13] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf70),
    .S(vdd),
    .D(_783_[13])
);

NAND2X1 _8127_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_636_)
);

FILL FILL_1__7084_ (
);

FILL FILL_2__14694_ (
);

FILL FILL_2__14274_ (
);

FILL FILL_0__7802_ (
);

FILL FILL_1__13687_ (
);

FILL FILL_1__13267_ (
);

FILL FILL_4__14601_ (
);

FILL FILL_1_BUFX2_insert950 (
);

FILL SFILL59000x23050 (
);

FILL FILL_1_BUFX2_insert951 (
);

OAI21X1 _12965_ (
    .A(_3627_),
    .B(vdd),
    .C(_3628_),
    .Y(_3620_[4])
);

FILL FILL_1_BUFX2_insert952 (
);

FILL FILL_3__8371_ (
);

DFFSR _12545_ (
    .Q(ALUOut[10]),
    .CLK(clk_bF$buf22),
    .R(rst_bF$buf28),
    .S(vdd),
    .D(_3360_[10])
);

FILL FILL_1_BUFX2_insert953 (
);

FILL FILL_1_BUFX2_insert954 (
);

NAND2X1 _12125_ (
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [3]),
    .Y(_3137_)
);

FILL FILL_1_BUFX2_insert955 (
);

FILL FILL_1_BUFX2_insert956 (
);

FILL FILL_1_BUFX2_insert957 (
);

FILL FILL_1_BUFX2_insert958 (
);

FILL FILL_1_BUFX2_insert959 (
);

FILL FILL_6__11594_ (
);

FILL SFILL104440x26050 (
);

FILL FILL_0__13621_ (
);

FILL FILL_3__16066_ (
);

FILL FILL_5__10167_ (
);

FILL FILL_2__15899_ (
);

FILL FILL_2__15479_ (
);

FILL FILL_2__15059_ (
);

FILL FILL_0__16093_ (
);

FILL SFILL33880x52050 (
);

FILL FILL_2__10194_ (
);

FILL FILL_1__9650_ (
);

FILL FILL_1__9230_ (
);

FILL FILL_4__15806_ (
);

FILL FILL_3__9996_ (
);

FILL SFILL49000x66050 (
);

FILL FILL_2__16000_ (
);

FILL FILL_4__10941_ (
);

FILL FILL_3__9156_ (
);

FILL FILL_4__10521_ (
);

FILL SFILL28120x25050 (
);

FILL FILL_1__15833_ (
);

FILL SFILL49080x23050 (
);

FILL FILL_1__15413_ (
);

FILL SFILL94440x75050 (
);

FILL FILL_0__14826_ (
);

FILL FILL_0__14406_ (
);

FILL SFILL89160x19050 (
);

FILL FILL_2__7993_ (
);

BUFX2 BUFX2_insert620 (
    .A(_3942_),
    .Y(_3942__bF$buf1)
);

FILL FILL_2__7573_ (
);

BUFX2 BUFX2_insert621 (
    .A(_3942_),
    .Y(_3942__bF$buf0)
);

BUFX2 BUFX2_insert622 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf4 )
);

BUFX2 BUFX2_insert623 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf3 )
);

BUFX2 BUFX2_insert624 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf2 )
);

FILL FILL_4__7499_ (
);

BUFX2 BUFX2_insert625 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf1 )
);

FILL FILL_4__7079_ (
);

BUFX2 BUFX2_insert626 (
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf0 )
);

BUFX2 BUFX2_insert627 (
    .A(_3977_),
    .Y(_3977__bF$buf4)
);

BUFX2 BUFX2_insert628 (
    .A(_3977_),
    .Y(_3977__bF$buf3)
);

FILL FILL_2__11399_ (
);

BUFX2 BUFX2_insert629 (
    .A(_3977_),
    .Y(_3977__bF$buf2)
);

FILL FILL_5__12733_ (
);

FILL FILL_5__12313_ (
);

FILL FILL_4__8860_ (
);

FILL FILL_4__8440_ (
);

FILL FILL_4__8020_ (
);

FILL FILL_4__11726_ (
);

FILL FILL_2__12760_ (
);

FILL FILL_4__11306_ (
);

FILL FILL_2__12340_ (
);

FILL SFILL49000x21050 (
);

FILL FILL_6__8366_ (
);

NAND2X1 _9085_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1112_)
);

FILL FILL_1__11753_ (
);

FILL FILL_4__14198_ (
);

FILL FILL_1__11333_ (
);

FILL FILL_0__8760_ (
);

FILL FILL_2__8778_ (
);

FILL FILL_2__8358_ (
);

FILL FILL_0__10746_ (
);

FILL FILL_0__8340_ (
);

DFFSR _10611_ (
    .Q(\datapath_1.regfile_1.regOut[29] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf78),
    .S(vdd),
    .D(_1823_[29])
);

NAND2X1 _13083_ (
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [1]),
    .Y(_3687_)
);

FILL FILL_5__13938_ (
);

FILL FILL_3__14972_ (
);

FILL FILL_5__13518_ (
);

FILL FILL_3__14552_ (
);

OAI21X1 _7818_ (
    .A(_469_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_470_),
    .Y(_458_[6])
);

FILL FILL_3__14132_ (
);

FILL FILL_4_BUFX2_insert460 (
);

FILL FILL_4_BUFX2_insert461 (
);

FILL FILL_4__9645_ (
);

FILL FILL_4__9225_ (
);

FILL FILL_4_BUFX2_insert462 (
);

FILL FILL_4_BUFX2_insert463 (
);

FILL FILL_2__13965_ (
);

FILL FILL111800x66050 (
);

FILL FILL_4_BUFX2_insert464 (
);

FILL FILL_2__13545_ (
);

FILL FILL_2__13125_ (
);

FILL FILL_4_BUFX2_insert465 (
);

FILL FILL_4_BUFX2_insert466 (
);

FILL SFILL39000x64050 (
);

FILL SFILL94360x37050 (
);

FILL FILL_4_BUFX2_insert467 (
);

FILL FILL_4_BUFX2_insert468 (
);

FILL FILL_4_BUFX2_insert469 (
);

FILL FILL_1__12958_ (
);

FILL FILL_1__12118_ (
);

FILL FILL_0__9545_ (
);

FILL FILL_3__7222_ (
);

FILL FILL_0__9125_ (
);

AOI21X1 _11816_ (
    .A(_2133_),
    .B(_2359_),
    .C(_2351_),
    .Y(_2907_)
);

FILL FILL_5__7988_ (
);

FILL FILL_5__7568_ (
);

FILL FILL_4__16344_ (
);

NOR2X1 _14288_ (
    .A(_4770_),
    .B(_4782_),
    .Y(_4783_)
);

FILL FILL_3__15757_ (
);

FILL FILL_3__15337_ (
);

FILL FILL_1__16371_ (
);

FILL FILL_3__10892_ (
);

FILL FILL_3__10052_ (
);

FILL FILL_0__15784_ (
);

FILL FILL_0__15364_ (
);

FILL SFILL79240x2050 (
);

FILL FILL111800x21050 (
);

FILL SFILL79160x7050 (
);

FILL FILL_1__8501_ (
);

FILL SFILL29080x64050 (
);

FILL SFILL53880x3050 (
);

FILL FILL_3__8847_ (
);

FILL FILL_3__8007_ (
);

FILL FILL_5__13691_ (
);

FILL FILL_5__13271_ (
);

OAI21X1 _7991_ (
    .A(_564_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .C(_565_),
    .Y(_523_[21])
);

OAI21X1 _7571_ (
    .A(_345_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_346_),
    .Y(_328_[9])
);

DFFSR _7151_ (
    .Q(\datapath_1.regfile_1.regOut[2] [25]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_68_[25])
);

FILL FILL_4__12264_ (
);

FILL SFILL8760x54050 (
);

FILL FILL_2__6844_ (
);

FILL FILL_3__11677_ (
);

FILL FILL_3__11257_ (
);

FILL FILL_1__12291_ (
);

FILL FILL_0__16149_ (
);

DFFSR _16434_ (
    .Q(\datapath_1.regfile_1.regOut[0] [17]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf81),
    .S(vdd),
    .D(_6769_[17])
);

AOI22X1 _16014_ (
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_6470_)
);

FILL FILL_0__11284_ (
);

FILL SFILL114600x54050 (
);

FILL SFILL53960x44050 (
);

FILL FILL_3_BUFX2_insert480 (
);

FILL FILL_4__7711_ (
);

FILL FILL_3_BUFX2_insert481 (
);

FILL FILL_3_BUFX2_insert482 (
);

FILL FILL_5__14896_ (
);

FILL FILL_5__14476_ (
);

FILL FILL_3_BUFX2_insert483 (
);

FILL FILL_2__11611_ (
);

FILL FILL_5__14056_ (
);

FILL FILL_3_BUFX2_insert484 (
);

FILL FILL_3__15090_ (
);

FILL FILL_6__7637_ (
);

NAND2X1 _8776_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_967_)
);

FILL FILL_3_BUFX2_insert485 (
);

NAND2X1 _8356_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_748_)
);

FILL FILL_3_BUFX2_insert486 (
);

FILL FILL_3_BUFX2_insert487 (
);

FILL FILL_3_BUFX2_insert488 (
);

FILL FILL_3_BUFX2_insert489 (
);

FILL FILL_4__13889_ (
);

FILL FILL_4__13469_ (
);

FILL FILL_2__14083_ (
);

FILL FILL_0__7611_ (
);

FILL FILL_2__7629_ (
);

FILL FILL_2__7209_ (
);

FILL FILL_1__13496_ (
);

FILL FILL_4__14830_ (
);

FILL FILL_4__14410_ (
);

NAND2X1 _12774_ (
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[26]),
    .Y(_3542_)
);

FILL FILL_0__12489_ (
);

OAI21X1 _12354_ (
    .A(_3300_),
    .B(MemToReg_bF$buf2),
    .C(_3301_),
    .Y(\datapath_1.mux_wd3.dout [3])
);

FILL FILL_0__12069_ (
);

FILL FILL_3__13823_ (
);

FILL FILL_3__13403_ (
);

FILL FILL_6__16268_ (
);

FILL FILL_4__8916_ (
);

FILL FILL_0__13850_ (
);

FILL FILL_0__13430_ (
);

FILL FILL_3__16295_ (
);

FILL FILL_0__13010_ (
);

FILL FILL_5__10396_ (
);

FILL FILL_1__8098_ (
);

FILL SFILL34680x51050 (
);

FILL FILL_1__11809_ (
);

FILL FILL_2__15288_ (
);

FILL FILL_3__6913_ (
);

FILL FILL_5__16202_ (
);

FILL FILL_5__6839_ (
);

FILL SFILL114520x16050 (
);

FILL FILL_4__15615_ (
);

AOI21X1 _13979_ (
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .B(_4115_),
    .C(_4479_),
    .Y(_4480_)
);

FILL FILL_3__9385_ (
);

NAND2X1 _13559_ (
    .A(_4061_),
    .B(_4068_),
    .Y(_4069_)
);

FILL FILL_4__10750_ (
);

INVX1 _13139_ (
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3724_)
);

FILL SFILL3720x35050 (
);

FILL FILL_3__14608_ (
);

FILL FILL_1__15642_ (
);

FILL FILL_1__15222_ (
);

FILL SFILL43960x42050 (
);

FILL FILL_6__12188_ (
);

FILL FILL_0__14635_ (
);

OAI22X1 _14920_ (
    .A(_5400_),
    .B(_3893__bF$buf3),
    .C(_3944__bF$buf1),
    .D(_5401_),
    .Y(_5402_)
);

AOI21X1 _14500_ (
    .A(_4990_),
    .B(_4964_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [21])
);

FILL FILL_0__14215_ (
);

FILL FILL_5__12962_ (
);

FILL FILL_5__12122_ (
);

BUFX2 _6842_ (
    .A(_1_[4]),
    .Y(memoryAddress[4])
);

FILL SFILL104520x59050 (
);

FILL SFILL48920x4050 (
);

FILL FILL_4__11955_ (
);

FILL FILL_4__11535_ (
);

FILL FILL_4__11115_ (
);

FILL FILL_1__16007_ (
);

FILL FILL_3__10948_ (
);

FILL FILL_3__10528_ (
);

FILL FILL_1__11982_ (
);

FILL FILL_1__11562_ (
);

FILL FILL_3__10108_ (
);

FILL FILL_1__11142_ (
);

NAND3X1 _15705_ (
    .A(_6167_),
    .B(_6168_),
    .C(_6166_),
    .Y(_6169_)
);

FILL FILL112280x53050 (
);

FILL FILL_2__8587_ (
);

FILL FILL_0__10975_ (
);

FILL FILL_0__10555_ (
);

DFFSR _10840_ (
    .Q(\datapath_1.regfile_1.regOut[31] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_1953_[2])
);

FILL FILL_0__10135_ (
);

OAI21X1 _10420_ (
    .A(_1797_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .C(_1798_),
    .Y(_1758_[20])
);

OAI21X1 _10000_ (
    .A(_1578_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .C(_1579_),
    .Y(_1563_[8])
);

FILL FILL_6__14334_ (
);

FILL FILL_5__13747_ (
);

FILL FILL_5__13327_ (
);

FILL FILL_3__14781_ (
);

FILL FILL_3__14361_ (
);

NAND2X1 _7627_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_384_)
);

NAND2X1 _7207_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_165_)
);

FILL FILL_4__9874_ (
);

FILL FILL_4__9034_ (
);

FILL FILL_2__13774_ (
);

FILL SFILL104520x14050 (
);

FILL FILL_2__13354_ (
);

FILL FILL_1__12767_ (
);

FILL FILL_1__12347_ (
);

FILL SFILL59000x18050 (
);

FILL FILL_3__7871_ (
);

FILL FILL_0__9774_ (
);

FILL FILL_0__9354_ (
);

FILL FILL_3__7451_ (
);

FILL SFILL108840x22050 (
);

FILL FILL_3__7031_ (
);

NOR2X1 _11625_ (
    .A(_2419_),
    .B(_2729_),
    .Y(_2730_)
);

INVX2 _11205_ (
    .A(_2323_),
    .Y(_2324_)
);

FILL FILL_5__7377_ (
);

FILL FILL_4__16153_ (
);

FILL FILL_6__10254_ (
);

AOI22X1 _14097_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [13]),
    .C(\datapath_1.regfile_1.regOut[6] [13]),
    .D(_4001__bF$buf1),
    .Y(_4596_)
);

FILL FILL_3__15986_ (
);

FILL FILL_0__12701_ (
);

FILL FILL_3__15566_ (
);

FILL FILL_3__15146_ (
);

FILL FILL_1__16180_ (
);

FILL FILL_1__7369_ (
);

FILL FILL_3__10281_ (
);

FILL FILL_2__14979_ (
);

FILL FILL_2__14559_ (
);

FILL FILL_2__14139_ (
);

FILL FILL_0__15593_ (
);

FILL SFILL33880x47050 (
);

FILL FILL_0__15173_ (
);

FILL FILL_1__8730_ (
);

FILL FILL_1__8310_ (
);

FILL FILL_2__15920_ (
);

FILL FILL_2__15500_ (
);

FILL FILL_3__8656_ (
);

FILL FILL_3__8236_ (
);

FILL FILL_5__13080_ (
);

FILL SFILL49080x18050 (
);

FILL FILL_1__14913_ (
);

NAND2X1 _7380_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_260_)
);

FILL FILL_4__12493_ (
);

FILL FILL_4__12073_ (
);

FILL FILL_0__13906_ (
);

FILL FILL_5__9523_ (
);

FILL FILL_3__11486_ (
);

FILL FILL_5__9103_ (
);

FILL FILL_3__11066_ (
);

FILL FILL_0__16378_ (
);

NOR3X1 _16243_ (
    .A(_6693_),
    .B(_6672_),
    .C(_6682_),
    .Y(_6694_)
);

FILL FILL_2__10899_ (
);

FILL FILL_2__10059_ (
);

FILL FILL_0__11093_ (
);

FILL FILL_1__9935_ (
);

FILL FILL_5__11813_ (
);

FILL FILL_1__9515_ (
);

FILL FILL_4__7940_ (
);

FILL FILL_4__7100_ (
);

FILL FILL_4__10806_ (
);

FILL FILL_2__11840_ (
);

FILL SFILL18600x25050 (
);

FILL FILL_0__6899_ (
);

FILL FILL_5__14285_ (
);

FILL FILL_2__11420_ (
);

FILL SFILL49000x16050 (
);

FILL FILL_2__11000_ (
);

NAND2X1 _8585_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_860_)
);

FILL FILL_6__7446_ (
);

DFFSR _8165_ (
    .Q(\datapath_1.regfile_1.regOut[10] [15]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_588_[15])
);

FILL FILL_1__10833_ (
);

FILL FILL_4__13698_ (
);

FILL FILL_4__13278_ (
);

FILL FILL_1__10413_ (
);

FILL SFILL94440x25050 (
);

FILL FILL_0__7840_ (
);

FILL FILL_2__7858_ (
);

FILL FILL_2__7438_ (
);

FILL FILL_0__7420_ (
);

FILL SFILL18840x8050 (
);

NAND2X1 _12583_ (
    .A(vdd),
    .B(memoryOutData[5]),
    .Y(_3435_)
);

FILL FILL_0__12298_ (
);

FILL SFILL84520x61050 (
);

INVX1 _12163_ (
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_3162_)
);

FILL SFILL23880x45050 (
);

FILL FILL_3__13632_ (
);

FILL FILL_3__13212_ (
);

FILL FILL_4__8725_ (
);

FILL FILL_2__12625_ (
);

FILL FILL_2__12205_ (
);

FILL SFILL39000x59050 (
);

FILL FILL_1__11618_ (
);

FILL FILL_2__15097_ (
);

FILL FILL_5__16011_ (
);

FILL FILL_0__8625_ (
);

FILL FILL_0__8205_ (
);

FILL SFILL48680x80050 (
);

FILL FILL_4__15844_ (
);

FILL FILL_4__15424_ (
);

FILL FILL_4__15004_ (
);

NOR2X1 _13788_ (
    .A(_4293_),
    .B(_4278_),
    .Y(_4294_)
);

AND2X2 _13368_ (
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3880_)
);

FILL FILL_3__14837_ (
);

FILL FILL_3__14417_ (
);

FILL FILL_1__15871_ (
);

FILL FILL_1__15451_ (
);

FILL FILL_1__15031_ (
);

FILL FILL_0__14864_ (
);

FILL FILL_0__14444_ (
);

FILL FILL_0__14024_ (
);

FILL FILL_2__7191_ (
);

CLKBUF1 CLKBUF1_insert160 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf64)
);

CLKBUF1 CLKBUF1_insert161 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf63)
);

CLKBUF1 CLKBUF1_insert162 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf62)
);

CLKBUF1 CLKBUF1_insert163 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf61)
);

FILL FILL_3__7927_ (
);

CLKBUF1 CLKBUF1_insert164 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf60)
);

FILL FILL_3__7507_ (
);

CLKBUF1 CLKBUF1_insert165 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf59)
);

FILL FILL_5__12771_ (
);

CLKBUF1 CLKBUF1_insert166 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf58)
);

FILL FILL_5__12351_ (
);

CLKBUF1 CLKBUF1_insert167 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert168 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf56)
);

FILL SFILL84440x23050 (
);

CLKBUF1 CLKBUF1_insert169 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf55)
);

FILL FILL_4__16209_ (
);

FILL FILL_4__11764_ (
);

FILL SFILL8760x49050 (
);

FILL FILL_4__11344_ (
);

FILL FILL_1__16236_ (
);

FILL FILL_3__10757_ (
);

FILL FILL_1__11791_ (
);

FILL FILL_1__11371_ (
);

FILL FILL_0__15649_ (
);

AOI22X1 _15934_ (
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .B(_5494_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_6392_)
);

FILL FILL_0__15229_ (
);

OAI21X1 _15514_ (
    .A(_5524__bF$buf1),
    .B(_4482_),
    .C(_5982_),
    .Y(_5983_)
);

FILL FILL_2__8396_ (
);

FILL FILL_0__10784_ (
);

FILL FILL_0__10364_ (
);

FILL SFILL53960x39050 (
);

FILL FILL_5__13976_ (
);

FILL FILL_5__13556_ (
);

FILL FILL_3__14590_ (
);

FILL FILL_5__13136_ (
);

FILL FILL_3__14170_ (
);

NAND2X1 _7856_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_496_)
);

NAND2X1 _7436_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_277_)
);

DFFSR _7016_ (
    .Q(\datapath_1.regfile_1.regOut[1] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_3_[18])
);

FILL FILL_4_BUFX2_insert840 (
);

FILL FILL_4__9683_ (
);

FILL FILL_4_BUFX2_insert841 (
);

FILL FILL_4_BUFX2_insert842 (
);

FILL FILL_4__9263_ (
);

FILL FILL_4__12969_ (
);

FILL FILL_4_BUFX2_insert843 (
);

FILL FILL_4__12129_ (
);

FILL FILL_4_BUFX2_insert844 (
);

FILL FILL_2__13583_ (
);

FILL FILL_2__13163_ (
);

FILL FILL_4_BUFX2_insert845 (
);

FILL FILL_4_BUFX2_insert846 (
);

FILL FILL_4_BUFX2_insert847 (
);

FILL FILL_4_BUFX2_insert848 (
);

FILL FILL_4_BUFX2_insert849 (
);

FILL FILL_1__12996_ (
);

FILL FILL_1__12576_ (
);

FILL FILL_1__12156_ (
);

FILL FILL_4__13910_ (
);

FILL FILL_3__7680_ (
);

FILL FILL_0__11989_ (
);

FILL FILL_0__9163_ (
);

NOR2X1 _11854_ (
    .A(\datapath_1.ALUResult [9]),
    .B(_2940_),
    .Y(_2941_)
);

FILL FILL_0__11569_ (
);

FILL FILL_0__11149_ (
);

NAND2X1 _11434_ (
    .A(_2220_),
    .B(_2225_),
    .Y(_2550_)
);

OR2X2 _11014_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2133_)
);

FILL FILL_3__12903_ (
);

FILL FILL_4__16382_ (
);

FILL FILL_5__7186_ (
);

FILL FILL_3__15795_ (
);

FILL FILL_3__15375_ (
);

FILL FILL_0__12510_ (
);

FILL FILL_1__7598_ (
);

FILL FILL_1__7178_ (
);

FILL FILL_2__14788_ (
);

FILL FILL_2__14368_ (
);

FILL FILL_5__15702_ (
);

FILL FILL_3__8885_ (
);

FILL FILL_3__8465_ (
);

INVX1 _12639_ (
    .A(\datapath_1.Data [24]),
    .Y(_3472_)
);

NAND3X1 _12219_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3203_)
);

FILL FILL_1__14722_ (
);

FILL FILL_1__14302_ (
);

FILL FILL_0__13715_ (
);

FILL FILL_2__6882_ (
);

FILL FILL_5__9752_ (
);

FILL FILL_3__11295_ (
);

FILL FILL_0__16187_ (
);

NOR2X1 _16052_ (
    .A(_6506_),
    .B(_5549__bF$buf0),
    .Y(_6507_)
);

FILL SFILL78680x36050 (
);

FILL FILL112360x41050 (
);

FILL FILL_2__10288_ (
);

FILL FILL_1__9744_ (
);

FILL FILL_5__11622_ (
);

FILL FILL_5__11202_ (
);

FILL FILL_3_BUFX2_insert860 (
);

FILL FILL_3_BUFX2_insert861 (
);

FILL FILL_3_BUFX2_insert862 (
);

FILL FILL_4__10615_ (
);

FILL FILL_3_BUFX2_insert863 (
);

FILL SFILL64040x50050 (
);

FILL FILL_3_BUFX2_insert864 (
);

FILL FILL_5__14094_ (
);

FILL FILL_1__15927_ (
);

FILL FILL_3_BUFX2_insert865 (
);

INVX1 _8394_ (
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_773_)
);

FILL FILL_1__15507_ (
);

FILL FILL_3_BUFX2_insert866 (
);

FILL FILL_3_BUFX2_insert867 (
);

FILL FILL_3_BUFX2_insert868 (
);

FILL FILL_3_BUFX2_insert869 (
);

FILL FILL_1__10642_ (
);

FILL FILL_4__13087_ (
);

FILL FILL112280x48050 (
);

FILL FILL_2__7247_ (
);

NAND2X1 _12392_ (
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [16]),
    .Y(_3327_)
);

FILL FILL_5__12827_ (
);

FILL FILL_5__12407_ (
);

FILL FILL_3__13861_ (
);

FILL FILL_3__13441_ (
);

FILL FILL_3__13021_ (
);

FILL FILL_4__8954_ (
);

FILL FILL_4__8114_ (
);

FILL FILL_2__12854_ (
);

FILL FILL_2__12434_ (
);

FILL FILL_5__15299_ (
);

FILL FILL_2__12014_ (
);

INVX1 _9599_ (
    .A(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_1373_)
);

DFFSR _9179_ (
    .Q(\datapath_1.regfile_1.regOut[18] [5]),
    .CLK(clk_bF$buf77),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1108_[5])
);

FILL FILL_1__11847_ (
);

FILL FILL_1__11427_ (
);

FILL FILL_1__11007_ (
);

FILL FILL_3__6951_ (
);

FILL FILL_5__16240_ (
);

FILL FILL_0__8854_ (
);

FILL FILL_0__8014_ (
);

NAND2X1 _10705_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1948_)
);

FILL FILL_5__6877_ (
);

FILL FILL_0_BUFX2_insert990 (
);

FILL FILL_0_BUFX2_insert991 (
);

FILL FILL_4__15653_ (
);

FILL FILL_0_BUFX2_insert992 (
);

FILL FILL_4__15233_ (
);

FILL FILL_0_BUFX2_insert993 (
);

FILL FILL_0_BUFX2_insert994 (
);

INVX1 _13597_ (
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_4106_)
);

FILL FILL_0_BUFX2_insert995 (
);

DFFSR _13177_ (
    .Q(\datapath_1.mux_iord.din0 [2]),
    .CLK(clk_bF$buf40),
    .R(rst_bF$buf79),
    .S(vdd),
    .D(_3685_[2])
);

FILL FILL_0_BUFX2_insert996 (
);

FILL FILL_0_BUFX2_insert997 (
);

FILL FILL_2__9813_ (
);

FILL FILL_3__14646_ (
);

FILL FILL_0_BUFX2_insert998 (
);

FILL FILL_1__15680_ (
);

FILL FILL_3__14226_ (
);

FILL FILL_0_BUFX2_insert999 (
);

FILL FILL_1__15260_ (
);

FILL FILL_1__6869_ (
);

FILL FILL_4__9739_ (
);

FILL FILL_2__13639_ (
);

FILL FILL_2__13219_ (
);

FILL FILL_0__14673_ (
);

FILL FILL_0__14253_ (
);

FILL FILL_1__7810_ (
);

FILL FILL_0__9639_ (
);

FILL FILL_3__7736_ (
);

FILL FILL_0__9219_ (
);

FILL FILL_3__7316_ (
);

FILL FILL_5__12580_ (
);

FILL FILL_5__12160_ (
);

BUFX2 _6880_ (
    .A(_2_[10]),
    .Y(memoryWriteData[10])
);

FILL FILL_4__16018_ (
);

FILL FILL_4__11993_ (
);

FILL FILL_4__11573_ (
);

FILL FILL_6__10119_ (
);

FILL FILL_4__11153_ (
);

FILL FILL_1__16045_ (
);

FILL FILL_5__8603_ (
);

FILL FILL_3__10566_ (
);

FILL FILL_3__10146_ (
);

FILL FILL_6_BUFX2_insert372 (
);

FILL FILL_1__11180_ (
);

FILL SFILL33080x14050 (
);

FILL FILL_0__15878_ (
);

AOI22X1 _15743_ (
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_6206_)
);

FILL FILL_0__15458_ (
);

NOR2X1 _15323_ (
    .A(_5795_),
    .B(_5796_),
    .Y(_5797_)
);

FILL FILL_0__15038_ (
);

FILL FILL_6_BUFX2_insert377 (
);

FILL FILL_0__10173_ (
);

FILL FILL_2__10920_ (
);

FILL FILL_5__13785_ (
);

FILL FILL_5__13365_ (
);

FILL FILL_2__10500_ (
);

DFFSR _7665_ (
    .Q(\datapath_1.regfile_1.regOut[6] [27]),
    .CLK(clk_bF$buf57),
    .R(rst_bF$buf109),
    .S(vdd),
    .D(_328_[27])
);

INVX1 _7245_ (
    .A(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_190_)
);

FILL FILL_4__9492_ (
);

FILL FILL_4__12778_ (
);

FILL FILL_4__12358_ (
);

FILL FILL_2__13392_ (
);

FILL FILL_0__6920_ (
);

FILL FILL_2__6938_ (
);

FILL FILL_5__9808_ (
);

FILL FILL_1__12385_ (
);

INVX1 _16108_ (
    .A(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_6562_)
);

FILL FILL_0__9392_ (
);

FILL FILL_0__11798_ (
);

FILL FILL_0__11378_ (
);

OAI21X1 _11663_ (
    .A(_2764_),
    .B(_2186_),
    .C(_2209_),
    .Y(_2765_)
);

INVX1 _11243_ (
    .A(_2361_),
    .Y(_2362_)
);

FILL FILL_6__15997_ (
);

FILL FILL_3__12712_ (
);

FILL FILL_6__15577_ (
);

FILL FILL_4__16191_ (
);

FILL FILL_4__7805_ (
);

FILL FILL_2__11705_ (
);

FILL FILL_3__15184_ (
);

FILL FILL_2__14597_ (
);

FILL FILL_2__14177_ (
);

FILL FILL_5__15931_ (
);

FILL FILL_5__15511_ (
);

FILL FILL_0__7705_ (
);

INVX1 _9811_ (
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_1494_)
);

FILL FILL_4__14924_ (
);

FILL FILL_4__14504_ (
);

FILL FILL_3__8694_ (
);

INVX1 _12868_ (
    .A(\datapath_1.a [15]),
    .Y(_3584_)
);

FILL FILL_3__8274_ (
);

INVX1 _12448_ (
    .A(ALUOut[3]),
    .Y(_3365_)
);

NAND3X1 _12028_ (
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [10]),
    .C(_3034__bF$buf3),
    .Y(_3067_)
);

FILL FILL_3__13917_ (
);

FILL FILL_1__14951_ (
);

FILL FILL_1__14531_ (
);

FILL FILL_1__14111_ (
);

FILL FILL_6__11497_ (
);

FILL FILL_5_BUFX2_insert390 (
);

FILL FILL_5_BUFX2_insert391 (
);

FILL SFILL8840x37050 (
);

FILL FILL_5_BUFX2_insert392 (
);

FILL FILL_0__13944_ (
);

FILL FILL_3__16389_ (
);

FILL FILL_5_BUFX2_insert393 (
);

FILL FILL_0__13524_ (
);

FILL FILL_0__13104_ (
);

FILL FILL_5_BUFX2_insert394 (
);

FILL FILL_5_BUFX2_insert395 (
);

FILL FILL_5_BUFX2_insert396 (
);

FILL FILL_5__9981_ (
);

FILL FILL_5_BUFX2_insert397 (
);

FILL FILL_5__9141_ (
);

FILL FILL_5_BUFX2_insert398 (
);

FILL FILL_5_BUFX2_insert399 (
);

NAND3X1 _16281_ (
    .A(_6723_),
    .B(_6730_),
    .C(_6718_),
    .Y(_6731_)
);

FILL FILL_5__11851_ (
);

FILL FILL_1__9553_ (
);

FILL FILL_5__11431_ (
);

FILL FILL_1__9133_ (
);

FILL FILL_5__11011_ (
);

FILL FILL_4__15709_ (
);

FILL FILL_2__16323_ (
);

FILL FILL_3__9899_ (
);

FILL SFILL109320x40050 (
);

FILL FILL_3__9479_ (
);

FILL FILL_4__10424_ (
);

FILL FILL_4__10004_ (
);

FILL FILL_1__15736_ (
);

FILL FILL_1__15316_ (
);

FILL FILL_6__7064_ (
);

FILL FILL_1__10871_ (
);

FILL FILL_1__10451_ (
);

FILL FILL_1__10031_ (
);

FILL FILL_0__14729_ (
);

FILL FILL_0__14309_ (
);

FILL FILL_2__7476_ (
);

FILL FILL_2__7056_ (
);

FILL FILL_6__13643_ (
);

FILL SFILL74120x40050 (
);

FILL FILL_5__12636_ (
);

FILL FILL_3__13670_ (
);

FILL FILL_5__12216_ (
);

FILL FILL_3__13250_ (
);

NAND2X1 _6936_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_25_)
);

FILL FILL_4__8763_ (
);

FILL FILL_4__8343_ (
);

FILL FILL_4__11629_ (
);

FILL FILL_4__11209_ (
);

FILL FILL_2__12243_ (
);

FILL FILL_1__11656_ (
);

FILL FILL_1__11236_ (
);

NAND3X1 _10934_ (
    .A(\control_1.op [2]),
    .B(_2066_),
    .C(_2067_),
    .Y(_2068_)
);

FILL FILL_0__10649_ (
);

FILL FILL_0__8243_ (
);

NAND2X1 _10514_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1841_)
);

FILL FILL_4__15882_ (
);

FILL FILL_4__15462_ (
);

FILL FILL_4__15042_ (
);

FILL SFILL34360x20050 (
);

FILL FILL_3__14875_ (
);

FILL FILL_2__9622_ (
);

FILL FILL_3__14455_ (
);

FILL FILL_3_CLKBUF1_insert1080 (
);

FILL FILL_3_CLKBUF1_insert1081 (
);

FILL FILL_3__14035_ (
);

FILL FILL_3_CLKBUF1_insert1082 (
);

FILL FILL_3_CLKBUF1_insert1083 (
);

FILL FILL_4__9548_ (
);

FILL FILL_4__9128_ (
);

FILL FILL_2__13868_ (
);

FILL FILL_2__13448_ (
);

FILL FILL_0__14482_ (
);

FILL FILL_2__13028_ (
);

FILL FILL_0__14062_ (
);

FILL FILL_0__9868_ (
);

FILL FILL_3__7965_ (
);

FILL FILL_3__7545_ (
);

FILL FILL_0__9028_ (
);

FILL FILL_3__7125_ (
);

NOR2X1 _11719_ (
    .A(_2509_),
    .B(_2801_),
    .Y(_2817_)
);

FILL FILL_1__13802_ (
);

FILL FILL_4__16247_ (
);

FILL FILL_4__11382_ (
);

FILL FILL_1__16274_ (
);

FILL FILL_5__8832_ (
);

FILL FILL_3__10795_ (
);

FILL FILL_3__10375_ (
);

OAI22X1 _15972_ (
    .A(_6428_),
    .B(_5545__bF$buf0),
    .C(_5527__bF$buf1),
    .D(_5055_),
    .Y(_6429_)
);

FILL FILL_0__15687_ (
);

INVX1 _15552_ (
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_6020_)
);

FILL FILL_0__15267_ (
);

OAI22X1 _15132_ (
    .A(_5478__bF$buf2),
    .B(_5609_),
    .C(_5552__bF$buf3),
    .D(_4065_),
    .Y(_5610_)
);

FILL FILL112360x36050 (
);

FILL FILL_5__10702_ (
);

FILL FILL_1__8824_ (
);

FILL FILL_1__8404_ (
);

FILL SFILL64040x45050 (
);

FILL FILL_5__13594_ (
);

FILL FILL_5__13174_ (
);

DFFSR _7894_ (
    .Q(\datapath_1.regfile_1.regOut[8] [0]),
    .CLK(clk_bF$buf91),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_458_[0])
);

INVX1 _7474_ (
    .A(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_302_)
);

INVX1 _7054_ (
    .A(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_83_)
);

FILL FILL_4__12587_ (
);

FILL FILL_4__12167_ (
);

FILL SFILL54120x81050 (
);

FILL FILL_5__9617_ (
);

FILL FILL_1__12194_ (
);

NAND2X1 _16337_ (
    .A(gnd),
    .B(gnd),
    .Y(_6779_)
);

OAI21X1 _11892_ (
    .A(_2968_),
    .B(IorD_bF$buf1),
    .C(_2969_),
    .Y(_1_[1])
);

FILL FILL_0__11187_ (
);

OAI21X1 _11472_ (
    .A(_2586_),
    .B(_2447_),
    .C(_2288_),
    .Y(_2587_)
);

FILL FILL_5__11907_ (
);

XOR2X1 _11052_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2171_)
);

FILL FILL_1__9609_ (
);

FILL FILL_3__12521_ (
);

FILL FILL_3__12101_ (
);

FILL FILL_4__7614_ (
);

FILL FILL_2__11934_ (
);

FILL FILL_5__14799_ (
);

FILL FILL_5__14379_ (
);

FILL FILL_2__11514_ (
);

DFFSR _8679_ (
    .Q(\datapath_1.regfile_1.regOut[14] [17]),
    .CLK(clk_bF$buf31),
    .R(rst_bF$buf25),
    .S(vdd),
    .D(_848_[17])
);

OAI21X1 _8259_ (
    .A(_702_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_703_),
    .Y(_653_[25])
);

FILL FILL_1__10927_ (
);

FILL FILL_1__10507_ (
);

FILL FILL_5__15740_ (
);

FILL FILL_5__15320_ (
);

FILL FILL_0__7934_ (
);

INVX1 _9620_ (
    .A(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_1387_)
);

FILL FILL_1__13399_ (
);

DFFSR _9200_ (
    .Q(\datapath_1.regfile_1.regOut[18] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1108_[26])
);

FILL FILL_4__14733_ (
);

FILL FILL_4__14313_ (
);

FILL SFILL54440x57050 (
);

DFFSR _12677_ (
    .Q(\datapath_1.Data [14]),
    .CLK(clk_bF$buf12),
    .R(rst_bF$buf86),
    .S(vdd),
    .D(_3425_[14])
);

FILL FILL_3__8083_ (
);

AOI22X1 _12257_ (
    .A(_2_[10]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [10]),
    .Y(_3232_)
);

FILL FILL_3__13726_ (
);

FILL FILL_3__13306_ (
);

FILL FILL_1__14760_ (
);

FILL FILL_1__14340_ (
);

FILL FILL_2__12719_ (
);

FILL FILL_0__13753_ (
);

FILL FILL_0__13333_ (
);

FILL FILL_3__16198_ (
);

FILL FILL_5__9790_ (
);

FILL FILL_5__10299_ (
);

FILL SFILL54040x43050 (
);

FILL FILL_5__9370_ (
);

NOR2X1 _16090_ (
    .A(_5181_),
    .B(_5535__bF$buf4),
    .Y(_6544_)
);

FILL FILL_0__8719_ (
);

FILL FILL_5__16105_ (
);

FILL FILL_1__9782_ (
);

FILL FILL_5__11660_ (
);

FILL FILL_5__11240_ (
);

FILL FILL_1__9362_ (
);

FILL FILL_4__15938_ (
);

FILL FILL_4__15518_ (
);

FILL FILL_2__16132_ (
);

FILL FILL_3__9288_ (
);

FILL FILL_4__10653_ (
);

FILL FILL_4__10233_ (
);

FILL FILL_1__15965_ (
);

FILL FILL_1__15545_ (
);

FILL FILL_1__15125_ (
);

FILL FILL_1__10680_ (
);

FILL FILL_1__10260_ (
);

FILL FILL_0__14958_ (
);

AOI22X1 _14823_ (
    .A(\datapath_1.regfile_1.regOut[28] [28]),
    .B(_3894_),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_5307_)
);

FILL FILL_0__14538_ (
);

AOI22X1 _14403_ (
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .B(_4154_),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_4895_)
);

FILL FILL_0__14118_ (
);

FILL FILL_6__13032_ (
);

FILL FILL_5__12865_ (
);

FILL FILL_5__12445_ (
);

FILL FILL_5__12025_ (
);

FILL FILL_4__8992_ (
);

FILL FILL_4__8572_ (
);

FILL FILL_4__11858_ (
);

FILL FILL_2__12892_ (
);

FILL FILL_4__11438_ (
);

FILL FILL_2__12472_ (
);

FILL FILL_4__11018_ (
);

FILL FILL_2__12052_ (
);

FILL FILL_1__11885_ (
);

FILL FILL_1__11465_ (
);

FILL FILL_1__11045_ (
);

NAND2X1 _15608_ (
    .A(_6069_),
    .B(_6074_),
    .Y(_6075_)
);

FILL FILL_0__8892_ (
);

FILL FILL_0__8472_ (
);

FILL FILL_0__10878_ (
);

NAND2X1 _10743_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .Y(_2017_)
);

FILL FILL_0__10038_ (
);

INVX1 _10323_ (
    .A(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_1754_)
);

FILL SFILL109400x73050 (
);

FILL FILL_4__15691_ (
);

FILL FILL_6__14237_ (
);

FILL FILL_4__15271_ (
);

FILL SFILL44040x41050 (
);

FILL FILL_2__9851_ (
);

FILL FILL_3__14684_ (
);

FILL FILL_3__14264_ (
);

FILL FILL_2__9011_ (
);

FILL FILL_4__9777_ (
);

FILL FILL112200x1050 (
);

FILL FILL_4__9357_ (
);

FILL FILL_2__13677_ (
);

FILL FILL_2__13257_ (
);

FILL FILL_0__14291_ (
);

FILL FILL112120x6050 (
);

FILL FILL_0__9677_ (
);

NAND2X1 _11948_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[20]),
    .Y(_3007_)
);

FILL FILL_3__7354_ (
);

FILL FILL_0__9257_ (
);

NAND3X1 _11528_ (
    .A(_2462__bF$buf1),
    .B(_2633_),
    .C(_2638_),
    .Y(_2639_)
);

INVX1 _11108_ (
    .A(\datapath_1.alu_1.ALUInA [21]),
    .Y(_2227_)
);

FILL SFILL8520x11050 (
);

FILL FILL_1__13611_ (
);

FILL FILL_4__16056_ (
);

FILL FILL_4__11191_ (
);

FILL FILL_3__15889_ (
);

FILL FILL_0__12604_ (
);

FILL FILL_3__15469_ (
);

FILL FILL_3__15049_ (
);

FILL FILL_1__16083_ (
);

FILL FILL_5__8641_ (
);

FILL FILL_6_BUFX2_insert751 (
);

FILL FILL_3__10184_ (
);

FILL FILL_5__8221_ (
);

INVX1 _15781_ (
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_6243_)
);

FILL FILL_0__15496_ (
);

NAND3X1 _15361_ (
    .A(_5829_),
    .B(_5830_),
    .C(_5833_),
    .Y(_5834_)
);

FILL FILL_0__15076_ (
);

FILL FILL_6_BUFX2_insert756 (
);

FILL FILL_3__16410_ (
);

FILL FILL_5__10931_ (
);

FILL FILL_5__10511_ (
);

FILL FILL_1__8633_ (
);

FILL FILL_1__8213_ (
);

FILL FILL_2__15823_ (
);

FILL FILL_2__15403_ (
);

FILL FILL_3__8979_ (
);

FILL FILL_3__8139_ (
);

FILL FILL_1__14816_ (
);

DFFSR _7283_ (
    .Q(\datapath_1.regfile_1.regOut[3] [29]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_133_[29])
);

FILL FILL_4__12396_ (
);

FILL FILL_3__9920_ (
);

FILL SFILL69160x52050 (
);

FILL FILL_0__13809_ (
);

FILL FILL_3__9500_ (
);

FILL FILL_2__6976_ (
);

FILL FILL_5__9846_ (
);

FILL FILL_5__9426_ (
);

FILL FILL_3__11389_ (
);

FILL FILL_5__9006_ (
);

FILL SFILL74120x35050 (
);

OAI22X1 _16146_ (
    .A(_6597_),
    .B(_5544__bF$buf0),
    .C(_5499__bF$buf3),
    .D(_6598_),
    .Y(_6599_)
);

FILL SFILL13480x19050 (
);

AOI21X1 _11281_ (
    .A(_2399_),
    .B(_2184_),
    .C(_2397_),
    .Y(_2400_)
);

FILL FILL_5__11716_ (
);

FILL FILL_3__12750_ (
);

FILL FILL_1__9418_ (
);

FILL FILL_3__12330_ (
);

FILL FILL_4__7843_ (
);

FILL FILL_4__7423_ (
);

FILL FILL_4__10709_ (
);

FILL FILL_2__11743_ (
);

FILL FILL_5__14188_ (
);

FILL FILL_2__11323_ (
);

OAI21X1 _8488_ (
    .A(_814_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .C(_815_),
    .Y(_783_[16])
);

OAI21X1 _8068_ (
    .A(_595_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .C(_596_),
    .Y(_588_[4])
);

FILL FILL_1__10316_ (
);

FILL FILL_0__7743_ (
);

FILL FILL_0__7323_ (
);

FILL FILL_4__14962_ (
);

FILL FILL_4__14542_ (
);

FILL SFILL64120x78050 (
);

FILL FILL_4__14122_ (
);

OAI21X1 _12486_ (
    .A(_3389_),
    .B(vdd),
    .C(_3390_),
    .Y(_3360_[15])
);

NAND3X1 _12066_ (
    .A(_3093_),
    .B(_3094_),
    .C(_3095_),
    .Y(\datapath_1.mux_pcsrc.dout [19])
);

FILL FILL_3__13955_ (
);

FILL FILL_2__8702_ (
);

FILL FILL_3__13535_ (
);

FILL FILL_3__13115_ (
);

FILL FILL_4__8628_ (
);

FILL FILL_4__8208_ (
);

FILL FILL_5_BUFX2_insert770 (
);

FILL FILL_5_BUFX2_insert771 (
);

FILL FILL_2__12528_ (
);

FILL FILL_0__13982_ (
);

FILL FILL_5_BUFX2_insert772 (
);

FILL FILL_5_BUFX2_insert773 (
);

FILL FILL_2__12108_ (
);

FILL FILL_0__13562_ (
);

FILL FILL_5_BUFX2_insert774 (
);

FILL FILL_0__13142_ (
);

FILL FILL_5_BUFX2_insert775 (
);

FILL FILL_5_BUFX2_insert776 (
);

FILL FILL_5_BUFX2_insert777 (
);

FILL FILL_5_BUFX2_insert778 (
);

FILL FILL_5_BUFX2_insert779 (
);

FILL FILL_5__16334_ (
);

FILL FILL_0__8528_ (
);

FILL FILL_0__8108_ (
);

FILL SFILL59160x50050 (
);

FILL FILL_1__9591_ (
);

FILL FILL_1__9171_ (
);

FILL FILL_4__15747_ (
);

FILL FILL_4__15327_ (
);

FILL FILL_2__16361_ (
);

FILL FILL_3__9097_ (
);

FILL FILL_4__10882_ (
);

FILL FILL_4__10042_ (
);

FILL FILL_2__9907_ (
);

FILL SFILL64120x33050 (
);

FILL FILL_1__15774_ (
);

FILL SFILL84920x7050 (
);

FILL FILL_1__15354_ (
);

FILL FILL_0__14767_ (
);

INVX1 _14632_ (
    .A(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_5120_)
);

FILL FILL_0__14347_ (
);

FILL SFILL89320x82050 (
);

NOR2X1 _14212_ (
    .A(_4705_),
    .B(_4708_),
    .Y(_4709_)
);

FILL FILL_2__7094_ (
);

FILL SFILL14040x80050 (
);

FILL FILL_5__12254_ (
);

FILL SFILL113880x44050 (
);

INVX1 _6974_ (
    .A(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_50_)
);

FILL FILL_4__8381_ (
);

FILL FILL_4__11667_ (
);

FILL FILL_4__11247_ (
);

FILL FILL_2__12281_ (
);

FILL FILL_1__16139_ (
);

FILL FILL_1__11694_ (
);

FILL FILL_1__11274_ (
);

INVX1 _15837_ (
    .A(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_6298_)
);

INVX1 _15417_ (
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_5888_)
);

FILL FILL_0__10687_ (
);

INVX1 _10972_ (
    .A(\control_1.reg_state.dout [0]),
    .Y(_2099_)
);

INVX1 _10552_ (
    .A(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_1866_)
);

FILL FILL_0__10267_ (
);

INVX1 _10132_ (
    .A(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_1647_)
);

FILL FILL_6__14886_ (
);

FILL FILL_3__11601_ (
);

FILL FILL_4__15080_ (
);

FILL FILL_5__13879_ (
);

FILL FILL_2__9660_ (
);

FILL FILL_5__13459_ (
);

FILL FILL_3__14493_ (
);

FILL FILL_5__13039_ (
);

FILL FILL_2__9240_ (
);

OAI21X1 _7759_ (
    .A(_450_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_451_),
    .Y(_393_[29])
);

FILL FILL_3__14073_ (
);

OAI21X1 _7339_ (
    .A(_231_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_232_),
    .Y(_198_[17])
);

FILL FILL_4__9166_ (
);

FILL FILL_2__13486_ (
);

FILL FILL_5__14820_ (
);

FILL FILL_5__14400_ (
);

FILL FILL_1__12899_ (
);

INVX1 _8700_ (
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_916_)
);

FILL FILL_1__12479_ (
);

FILL FILL_1__12059_ (
);

FILL FILL_4__13813_ (
);

FILL FILL_0__9486_ (
);

FILL FILL_3__7583_ (
);

AND2X2 _11757_ (
    .A(_2851_),
    .B(_2558_),
    .Y(_2852_)
);

FILL FILL_3__7163_ (
);

AOI21X1 _11337_ (
    .A(_2453_),
    .B(_2450_),
    .C(_2455_),
    .Y(_2456_)
);

FILL SFILL18680x64050 (
);

FILL FILL_1__13840_ (
);

FILL FILL_1__13420_ (
);

FILL FILL_4__16285_ (
);

FILL FILL_5__7089_ (
);

FILL FILL_1__13000_ (
);

FILL FILL_3__15698_ (
);

FILL FILL_0__12833_ (
);

FILL FILL_0__12413_ (
);

FILL FILL_3__15278_ (
);

FILL FILL_5__8870_ (
);

FILL FILL_5__8450_ (
);

INVX1 _15590_ (
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_6057_)
);

OAI22X1 _15170_ (
    .A(_5466__bF$buf0),
    .B(_4105_),
    .C(_4141_),
    .D(_5526__bF$buf2),
    .Y(_5647_)
);

FILL FILL_5__15605_ (
);

OAI21X1 _9905_ (
    .A(_1535_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1536_),
    .Y(_1498_[19])
);

FILL FILL_1__8862_ (
);

FILL FILL_1__8442_ (
);

FILL FILL_5__10320_ (
);

FILL FILL_2__15632_ (
);

FILL FILL_2__15212_ (
);

FILL FILL_3__8788_ (
);

FILL FILL_3__8368_ (
);

FILL FILL_1__14625_ (
);

FILL FILL_1__14205_ (
);

OAI21X1 _7092_ (
    .A(_107_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_108_),
    .Y(_68_[20])
);

FILL FILL_0__13618_ (
);

INVX1 _13903_ (
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_4406_)
);

FILL FILL_5__9655_ (
);

FILL FILL_3__11198_ (
);

FILL FILL_5__9235_ (
);

INVX1 _16375_ (
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_6804_)
);

FILL FILL_5__11945_ (
);

AOI21X1 _11090_ (
    .A(_2208_),
    .B(_2181_),
    .C(_2207_),
    .Y(_2209_)
);

FILL FILL_1__9647_ (
);

FILL FILL_5__11525_ (
);

FILL FILL_1__9227_ (
);

FILL FILL_5__11105_ (
);

FILL SFILL79240x42050 (
);

FILL FILL_4__10938_ (
);

FILL FILL_4__7232_ (
);

FILL FILL_2__11972_ (
);

FILL FILL_4__10518_ (
);

FILL FILL_2__11552_ (
);

FILL FILL_2__11132_ (
);

DFFSR _8297_ (
    .Q(\datapath_1.regfile_1.regOut[11] [19]),
    .CLK(clk_bF$buf90),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_653_[19])
);

FILL FILL_1__10965_ (
);

FILL FILL_1__10545_ (
);

FILL FILL_1__10125_ (
);

FILL FILL_0__7972_ (
);

FILL FILL_0__7552_ (
);

BUFX2 BUFX2_insert590 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf17)
);

BUFX2 BUFX2_insert591 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf16)
);

BUFX2 BUFX2_insert592 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf15)
);

BUFX2 BUFX2_insert593 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf14)
);

BUFX2 BUFX2_insert594 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf13)
);

BUFX2 BUFX2_insert595 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf12)
);

FILL FILL_4__14771_ (
);

FILL SFILL44040x36050 (
);

BUFX2 BUFX2_insert596 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf11)
);

FILL FILL_4__14351_ (
);

BUFX2 BUFX2_insert597 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf10)
);

FILL SFILL94360x2050 (
);

BUFX2 BUFX2_insert598 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf9)
);

BUFX2 BUFX2_insert599 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf8)
);

NAND3X1 _12295_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3260_)
);

FILL SFILL54040x9050 (
);

FILL FILL_2__8511_ (
);

FILL FILL_3__13764_ (
);

FILL FILL_3__13344_ (
);

FILL FILL_4__8857_ (
);

FILL FILL_4__8017_ (
);

FILL FILL_2__12757_ (
);

FILL FILL_0__13791_ (
);

FILL FILL_2__12337_ (
);

FILL FILL_0__13371_ (
);

FILL FILL111880x10050 (
);

FILL FILL_0__8757_ (
);

FILL FILL_3__6854_ (
);

FILL FILL_5__16143_ (
);

FILL FILL_0__8337_ (
);

DFFSR _10608_ (
    .Q(\datapath_1.regfile_1.regOut[29] [26]),
    .CLK(clk_bF$buf55),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_1823_[26])
);

FILL SFILL104520x5050 (
);

FILL FILL_4__15976_ (
);

FILL FILL_4__15556_ (
);

FILL SFILL34040x79050 (
);

FILL FILL_4__15136_ (
);

FILL FILL_2__16170_ (
);

FILL SFILL109400x23050 (
);

FILL FILL_4__10691_ (
);

FILL FILL_4__10271_ (
);

FILL FILL_3__14969_ (
);

FILL FILL_3__14549_ (
);

FILL FILL_3__14129_ (
);

FILL FILL_1__15583_ (
);

FILL FILL_1__15163_ (
);

FILL FILL_5__7721_ (
);

FILL FILL_5__7301_ (
);

FILL FILL_0__14996_ (
);

INVX1 _14861_ (
    .A(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_5344_)
);

FILL FILL_0__14576_ (
);

FILL SFILL69240x40050 (
);

FILL FILL_0__14156_ (
);

OAI22X1 _14441_ (
    .A(_4931_),
    .B(_3893__bF$buf3),
    .C(_3959_),
    .D(_4932_),
    .Y(_4933_)
);

AOI22X1 _14021_ (
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[18] [11]),
    .C(\datapath_1.regfile_1.regOut[31] [11]),
    .D(_3995__bF$buf1),
    .Y(_4522_)
);

FILL FILL_3__15910_ (
);

FILL FILL_1__7713_ (
);

FILL FILL_6__13490_ (
);

FILL FILL_2__14903_ (
);

FILL SFILL114680x43050 (
);

FILL FILL_3__7219_ (
);

FILL FILL_5__12483_ (
);

FILL FILL_5__12063_ (
);

FILL FILL_4__11896_ (
);

FILL FILL_4__8190_ (
);

FILL SFILL38760x56050 (
);

FILL FILL_4__11476_ (
);

FILL SFILL69160x47050 (
);

FILL FILL_4__11056_ (
);

FILL FILL_2__12090_ (
);

FILL FILL_1__16368_ (
);

FILL FILL_3__10889_ (
);

FILL FILL_5__8506_ (
);

FILL FILL_3__10049_ (
);

FILL FILL_1__11083_ (
);

OAI22X1 _15646_ (
    .A(_5478__bF$buf1),
    .B(_4649_),
    .C(_4663_),
    .D(_5534__bF$buf0),
    .Y(_6112_)
);

OAI22X1 _15226_ (
    .A(_5526__bF$buf0),
    .B(_4158_),
    .C(_4150_),
    .D(_5527__bF$buf0),
    .Y(_5702_)
);

FILL FILL_0__8090_ (
);

FILL FILL_0__10496_ (
);

INVX1 _10781_ (
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_1978_)
);

INVX1 _10361_ (
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .Y(_1759_)
);

FILL FILL_3__11830_ (
);

FILL FILL_3__11410_ (
);

FILL FILL_4__6923_ (
);

FILL FILL_0__16302_ (
);

FILL FILL_2__10823_ (
);

FILL FILL_5__13688_ (
);

FILL FILL_5__13268_ (
);

FILL FILL_2__10403_ (
);

OAI21X1 _7988_ (
    .A(_562_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .C(_563_),
    .Y(_523_[20])
);

OAI21X1 _7568_ (
    .A(_343_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .C(_344_),
    .Y(_328_[8])
);

DFFSR _7148_ (
    .Q(\datapath_1.regfile_1.regOut[2] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf34),
    .S(vdd),
    .D(_68_[22])
);

FILL FILL_4__9395_ (
);

FILL FILL_2__13295_ (
);

FILL SFILL104280x72050 (
);

FILL FILL_1__12288_ (
);

FILL FILL_4__13622_ (
);

FILL FILL_0__9295_ (
);

NAND3X1 _11986_ (
    .A(PCSource_1_bF$buf3),
    .B(gnd),
    .C(_3034__bF$buf2),
    .Y(_3035_)
);

AOI21X1 _11566_ (
    .A(_2674_),
    .B(_2672_),
    .C(_2667_),
    .Y(_2675_)
);

NOR2X1 _11146_ (
    .A(_2263_),
    .B(_2264_),
    .Y(_2265_)
);

FILL FILL_3__12615_ (
);

FILL FILL_3_BUFX2_insert10 (
);

FILL FILL_3_BUFX2_insert11 (
);

FILL FILL_4__16094_ (
);

FILL FILL_3_BUFX2_insert12 (
);

FILL FILL_3_BUFX2_insert13 (
);

FILL FILL_4__7708_ (
);

FILL FILL_3_BUFX2_insert14 (
);

FILL FILL_3_BUFX2_insert15 (
);

FILL FILL_3_BUFX2_insert16 (
);

FILL FILL_3_BUFX2_insert17 (
);

FILL FILL_2__11608_ (
);

FILL SFILL99320x34050 (
);

FILL FILL_0__12642_ (
);

FILL FILL_3_BUFX2_insert18 (
);

FILL FILL_3_BUFX2_insert19 (
);

FILL FILL_0__12222_ (
);

FILL FILL_3__15087_ (
);

FILL SFILL23800x6050 (
);

FILL SFILL63960x9050 (
);

FILL FILL_5__15834_ (
);

FILL SFILL89400x70050 (
);

FILL FILL_5__15414_ (
);

FILL SFILL28760x54050 (
);

FILL FILL_0__7608_ (
);

FILL SFILL59160x45050 (
);

DFFSR _9714_ (
    .Q(\datapath_1.regfile_1.regOut[22] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1368_[28])
);

FILL FILL_1__8251_ (
);

FILL FILL_4__14827_ (
);

FILL SFILL3720x2050 (
);

FILL FILL_4__14407_ (
);

FILL FILL_2__15861_ (
);

FILL FILL_2__15441_ (
);

FILL FILL_2__15021_ (
);

FILL FILL_3__8597_ (
);

FILL SFILL64120x28050 (
);

FILL SFILL3640x7050 (
);

FILL FILL_1__14854_ (
);

FILL FILL_1__14434_ (
);

FILL FILL_1__14014_ (
);

FILL FILL_0__13847_ (
);

FILL FILL_0__13427_ (
);

NOR2X1 _13712_ (
    .A(_4218_),
    .B(_4215_),
    .Y(_4219_)
);

FILL FILL_0__13007_ (
);

FILL FILL_5__9884_ (
);

FILL FILL_5__9464_ (
);

FILL FILL_5__9044_ (
);

FILL FILL_6__12341_ (
);

NOR2X1 _16184_ (
    .A(_6635_),
    .B(_6633_),
    .Y(_6636_)
);

FILL FILL_5__11754_ (
);

FILL FILL_1__9876_ (
);

FILL SFILL113880x39050 (
);

FILL FILL_5__11334_ (
);

FILL FILL_1__9036_ (
);

FILL FILL_2__16226_ (
);

FILL FILL_4__7881_ (
);

FILL FILL_4__7461_ (
);

FILL FILL_4__7041_ (
);

FILL FILL_4__10747_ (
);

FILL FILL_2__11781_ (
);

FILL FILL_2__11361_ (
);

FILL FILL_1__15639_ (
);

FILL FILL_1__15219_ (
);

FILL FILL_1__10774_ (
);

NAND3X1 _14917_ (
    .A(_5390_),
    .B(_5391_),
    .C(_5398_),
    .Y(_5399_)
);

FILL SFILL33960x72050 (
);

FILL FILL_2__7799_ (
);

FILL FILL_2__7379_ (
);

FILL FILL_0__7361_ (
);

FILL SFILL89320x32050 (
);

FILL FILL_6__13966_ (
);

FILL FILL_6__13546_ (
);

FILL FILL_4__14580_ (
);

FILL FILL_4__14160_ (
);

FILL FILL_5__12959_ (
);

FILL FILL_2__8740_ (
);

FILL FILL_3__13993_ (
);

FILL FILL_2__8320_ (
);

FILL FILL_5__12119_ (
);

FILL FILL_3__13573_ (
);

FILL FILL_3__13153_ (
);

BUFX2 _6839_ (
    .A(_1_[1]),
    .Y(memoryAddress[1])
);

FILL FILL_4__8246_ (
);

FILL FILL_2__12986_ (
);

FILL FILL_2__12146_ (
);

FILL FILL_5__13900_ (
);

FILL SFILL89240x39050 (
);

FILL FILL_1__11979_ (
);

FILL FILL_1__11559_ (
);

FILL FILL_1__11139_ (
);

FILL FILL_0__8986_ (
);

FILL FILL_5__16372_ (
);

FILL FILL_0__8566_ (
);

OAI21X1 _10837_ (
    .A(_2014_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_2015_),
    .Y(_1953_[31])
);

FILL FILL_0__8146_ (
);

OAI21X1 _10417_ (
    .A(_1795_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .C(_1796_),
    .Y(_1758_[19])
);

FILL SFILL79320x75050 (
);

FILL SFILL18680x59050 (
);

FILL FILL_4__15785_ (
);

FILL FILL_4__15365_ (
);

FILL FILL_1__12500_ (
);

FILL FILL_2__9525_ (
);

FILL FILL_0__11913_ (
);

FILL FILL_3__14778_ (
);

FILL FILL_3__14358_ (
);

FILL FILL_2__9105_ (
);

FILL FILL_1__15392_ (
);

FILL FILL_5__7950_ (
);

FILL FILL_5__7110_ (
);

FILL FILL_0__14385_ (
);

INVX1 _14670_ (
    .A(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_5157_)
);

NOR2X1 _14250_ (
    .A(_4745_),
    .B(_4742_),
    .Y(_4746_)
);

FILL FILL_1__7942_ (
);

FILL FILL_1__7102_ (
);

FILL FILL_2__14712_ (
);

FILL FILL_3__7868_ (
);

FILL FILL_3__7448_ (
);

FILL FILL_5__12292_ (
);

FILL SFILL23960x70050 (
);

FILL FILL_1__13705_ (
);

FILL SFILL79320x30050 (
);

FILL SFILL18680x14050 (
);

FILL SFILL59000x1050 (
);

FILL FILL_4__11285_ (
);

FILL FILL_1__16177_ (
);

FILL FILL_3__10698_ (
);

FILL FILL_5__8735_ (
);

FILL FILL_3__10278_ (
);

FILL FILL_5__8315_ (
);

OAI22X1 _15875_ (
    .A(_6334_),
    .B(_5545__bF$buf2),
    .C(_5466__bF$buf4),
    .D(_4934_),
    .Y(_6335_)
);

NOR2X1 _15455_ (
    .A(_5911_),
    .B(_5925_),
    .Y(_5926_)
);

OAI21X1 _15035_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5514_),
    .C(_5512_),
    .Y(_5515_)
);

DFFSR _10590_ (
    .Q(\datapath_1.regfile_1.regOut[29] [8]),
    .CLK(clk_bF$buf8),
    .R(rst_bF$buf48),
    .S(vdd),
    .D(_1823_[8])
);

OAI21X1 _10170_ (
    .A(_1671_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1672_),
    .Y(_1628_[22])
);

FILL FILL_1__8727_ (
);

FILL SFILL79240x37050 (
);

FILL FILL_2__15917_ (
);

FILL FILL_0__16111_ (
);

FILL FILL_2__10632_ (
);

FILL FILL_5__13497_ (
);

DFFSR _7797_ (
    .Q(\datapath_1.regfile_1.regOut[7] [31]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_393_[31])
);

NAND2X1 _7377_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_258_)
);

FILL SFILL69320x73050 (
);

FILL SFILL39560x10050 (
);

FILL FILL_3_BUFX2_insert100 (
);

FILL FILL_3_BUFX2_insert101 (
);

FILL FILL_3_BUFX2_insert102 (
);

FILL FILL_3_BUFX2_insert103 (
);

FILL FILL_3_BUFX2_insert104 (
);

FILL FILL_3_BUFX2_insert105 (
);

FILL FILL_3_BUFX2_insert106 (
);

FILL FILL_3_BUFX2_insert107 (
);

FILL FILL_1__12097_ (
);

FILL FILL_3_BUFX2_insert108 (
);

FILL FILL_4__13851_ (
);

FILL FILL_3_BUFX2_insert109 (
);

FILL FILL_4__13431_ (
);

FILL FILL_4__13011_ (
);

AOI21X1 _11795_ (
    .A(_2887_),
    .B(_2363_),
    .C(_2143_),
    .Y(_2888_)
);

OAI22X1 _11375_ (
    .A(_2490_),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .C(_2491_),
    .D(_2357_),
    .Y(_2492_)
);

FILL FILL_3__12844_ (
);

FILL FILL_3__12424_ (
);

FILL FILL_3__12004_ (
);

FILL FILL_4__7937_ (
);

FILL FILL_2__11837_ (
);

FILL FILL_0__12871_ (
);

FILL FILL_2__11417_ (
);

FILL FILL_0__12451_ (
);

FILL FILL_0__12031_ (
);

FILL FILL_5__15643_ (
);

FILL FILL_5__15223_ (
);

FILL FILL_0__7837_ (
);

FILL FILL_0__7417_ (
);

DFFSR _9943_ (
    .Q(\datapath_1.regfile_1.regOut[24] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf95),
    .S(vdd),
    .D(_1498_[1])
);

NAND2X1 _9523_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1343_)
);

NAND2X1 _9103_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1124_)
);

FILL FILL_1__8480_ (
);

FILL FILL_1__8060_ (
);

FILL FILL_4__14636_ (
);

FILL FILL_2__15670_ (
);

FILL FILL_4__14216_ (
);

FILL SFILL109400x18050 (
);

FILL FILL_2__15250_ (
);

FILL FILL_3__13629_ (
);

FILL FILL_3__13209_ (
);

FILL FILL_1__14663_ (
);

FILL FILL_1__14243_ (
);

FILL FILL_0_BUFX2_insert230 (
);

FILL FILL_0_BUFX2_insert231 (
);

FILL FILL_0_BUFX2_insert232 (
);

FILL FILL_0_BUFX2_insert233 (
);

FILL FILL_0__13656_ (
);

NOR2X1 _13941_ (
    .A(_4442_),
    .B(_4439_),
    .Y(_4443_)
);

FILL FILL_0_BUFX2_insert234 (
);

FILL FILL_0__13236_ (
);

INVX1 _13521_ (
    .A(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_4032_)
);

FILL FILL_0_BUFX2_insert235 (
);

NAND2X1 _13101_ (
    .A(PCEn_bF$buf4),
    .B(\datapath_1.mux_pcsrc.dout [7]),
    .Y(_3699_)
);

FILL FILL_0_BUFX2_insert236 (
);

FILL FILL_0_BUFX2_insert237 (
);

FILL FILL_0_BUFX2_insert238 (
);

FILL FILL_5__9273_ (
);

FILL FILL_0_BUFX2_insert239 (
);

FILL FILL_5__16008_ (
);

FILL FILL_5__11983_ (
);

FILL FILL_1__9685_ (
);

FILL FILL_5__11563_ (
);

FILL FILL_1__9265_ (
);

FILL FILL_5__11143_ (
);

FILL SFILL99400x67050 (
);

FILL FILL_4__7690_ (
);

FILL FILL_2__16035_ (
);

FILL FILL_4__10976_ (
);

FILL FILL_4__10556_ (
);

FILL FILL_4__10136_ (
);

FILL FILL_2__11590_ (
);

FILL FILL_2__11170_ (
);

FILL FILL_1__15868_ (
);

FILL FILL_1__15448_ (
);

FILL FILL_1__15028_ (
);

FILL FILL_1__10163_ (
);

INVX1 _14726_ (
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_5212_)
);

AOI22X1 _14306_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [17]),
    .C(\datapath_1.regfile_1.regOut[2] [17]),
    .D(_3998__bF$buf0),
    .Y(_4801_)
);

FILL FILL_0__7590_ (
);

BUFX2 BUFX2_insert970 (
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf0 )
);

FILL FILL_0__7170_ (
);

BUFX2 BUFX2_insert971 (
    .A(PCEn),
    .Y(PCEn_bF$buf7)
);

FILL FILL_2__7188_ (
);

BUFX2 BUFX2_insert972 (
    .A(PCEn),
    .Y(PCEn_bF$buf6)
);

BUFX2 BUFX2_insert973 (
    .A(PCEn),
    .Y(PCEn_bF$buf5)
);

FILL FILL_3__10910_ (
);

BUFX2 BUFX2_insert974 (
    .A(PCEn),
    .Y(PCEn_bF$buf4)
);

BUFX2 BUFX2_insert975 (
    .A(PCEn),
    .Y(PCEn_bF$buf3)
);

BUFX2 BUFX2_insert976 (
    .A(PCEn),
    .Y(PCEn_bF$buf2)
);

BUFX2 BUFX2_insert977 (
    .A(PCEn),
    .Y(PCEn_bF$buf1)
);

BUFX2 BUFX2_insert978 (
    .A(PCEn),
    .Y(PCEn_bF$buf0)
);

FILL FILL_0__15802_ (
);

BUFX2 BUFX2_insert979 (
    .A(_3967_),
    .Y(_3967__bF$buf3)
);

FILL SFILL69160x3050 (
);

FILL FILL_5__12768_ (
);

FILL FILL_5__12348_ (
);

FILL FILL_3__13382_ (
);

FILL SFILL69080x8050 (
);

FILL FILL_4__8895_ (
);

FILL FILL_4__8475_ (
);

FILL FILL_4__8055_ (
);

FILL FILL_2__12375_ (
);

FILL SFILL99400x22050 (
);

FILL FILL_1__11788_ (
);

FILL FILL_1__11368_ (
);

FILL FILL_4__12702_ (
);

FILL FILL_5__16181_ (
);

FILL FILL_3__6892_ (
);

FILL FILL_0__8375_ (
);

FILL FILL_6__9762_ (
);

OAI21X1 _10646_ (
    .A(_1907_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1908_),
    .Y(_1888_[10])
);

DFFSR _10226_ (
    .Q(\datapath_1.regfile_1.regOut[26] [28]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf9),
    .S(vdd),
    .D(_1628_[28])
);

FILL FILL_4__15594_ (
);

FILL FILL_4__15174_ (
);

FILL SFILL99320x29050 (
);

FILL FILL_2__9754_ (
);

FILL FILL_3__14587_ (
);

FILL FILL_2__9334_ (
);

FILL FILL_0__11722_ (
);

FILL FILL_3__14167_ (
);

FILL FILL_0__11302_ (
);

FILL FILL_0__14194_ (
);

FILL SFILL73800x80050 (
);

FILL FILL_5__14914_ (
);

FILL SFILL28760x49050 (
);

FILL FILL_1__7751_ (
);

FILL FILL_1__7331_ (
);

FILL SFILL104280x22050 (
);

FILL FILL_4__13907_ (
);

FILL FILL_2__14941_ (
);

FILL FILL_2__14521_ (
);

FILL FILL_2__14101_ (
);

FILL FILL_3__7677_ (
);

FILL FILL_1__13934_ (
);

FILL FILL_4__16379_ (
);

FILL FILL_1__13514_ (
);

FILL FILL_4__11094_ (
);

FILL FILL_0__12507_ (
);

FILL FILL_5__8964_ (
);

FILL FILL_5__8124_ (
);

NOR2X1 _15684_ (
    .A(_6148_),
    .B(_6146_),
    .Y(_6149_)
);

FILL FILL_0__15399_ (
);

FILL FILL_6__11001_ (
);

NOR2X1 _15264_ (
    .A(_5738_),
    .B(_5737_),
    .Y(_5739_)
);

FILL FILL_3__16313_ (
);

FILL FILL_5__10834_ (
);

FILL FILL_1__8956_ (
);

FILL FILL_5__10414_ (
);

FILL FILL_1__8116_ (
);

FILL SFILL94280x71050 (
);

FILL FILL_2__15726_ (
);

FILL FILL_2__15306_ (
);

FILL FILL_4__6961_ (
);

FILL FILL_0__16340_ (
);

FILL FILL_2__10441_ (
);

FILL FILL_2__10021_ (
);

FILL FILL_1__14719_ (
);

NAND2X1 _7186_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_151_)
);

FILL FILL_4__12299_ (
);

FILL FILL_3__9403_ (
);

FILL FILL_0__6861_ (
);

FILL FILL_2__6879_ (
);

FILL FILL_5__9749_ (
);

FILL SFILL89320x27050 (
);

FILL FILL_4__13660_ (
);

FILL FILL_4__13240_ (
);

INVX1 _16049_ (
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_6504_)
);

NOR2X1 _11184_ (
    .A(_2302_),
    .B(_2293_),
    .Y(_2303_)
);

FILL FILL_2__7820_ (
);

FILL FILL_5__11619_ (
);

FILL FILL_3__12653_ (
);

FILL SFILL18760x47050 (
);

FILL FILL_3__12233_ (
);

FILL FILL_4__7746_ (
);

FILL FILL_4__7326_ (
);

FILL FILL_2__11646_ (
);

FILL FILL_2__11226_ (
);

FILL FILL_0__12260_ (
);

FILL FILL_1__10639_ (
);

FILL FILL_5__15872_ (
);

FILL FILL_5__15452_ (
);

FILL FILL_5__15032_ (
);

NAND2X1 _9752_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1455_)
);

FILL FILL_0__7226_ (
);

DFFSR _9332_ (
    .Q(\datapath_1.regfile_1.regOut[19] [30]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_1173_[30])
);

FILL FILL_4__14865_ (
);

FILL FILL_4__14445_ (
);

FILL FILL_4__14025_ (
);

NAND2X1 _12389_ (
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [15]),
    .Y(_3325_)
);

FILL FILL_3__13858_ (
);

FILL FILL_2__8605_ (
);

FILL FILL_3__13438_ (
);

FILL FILL_1__14892_ (
);

FILL FILL_1__14472_ (
);

FILL FILL_3__13018_ (
);

FILL FILL_1__14052_ (
);

FILL FILL_0__13885_ (
);

NAND3X1 _13750_ (
    .A(_4247_),
    .B(_4248_),
    .C(_4255_),
    .Y(_4256_)
);

FILL FILL_0__13465_ (
);

INVX2 _13330_ (
    .A(_3798_),
    .Y(_3856_)
);

FILL FILL_0__13045_ (
);

FILL SFILL79720x39050 (
);

FILL FILL_5__9082_ (
);

FILL FILL_5__16237_ (
);

FILL FILL_3__6948_ (
);

FILL FILL_5__11792_ (
);

FILL FILL_5__11372_ (
);

FILL FILL_1__9494_ (
);

FILL SFILL79320x25050 (
);

FILL FILL_2__16264_ (
);

FILL FILL_4__10785_ (
);

FILL FILL_4__10365_ (
);

FILL FILL_4_BUFX2_insert60 (
);

FILL FILL_4_BUFX2_insert61 (
);

FILL FILL_1__15677_ (
);

FILL FILL_4_BUFX2_insert62 (
);

FILL FILL_1__15257_ (
);

FILL FILL_4_BUFX2_insert63 (
);

FILL FILL_4_BUFX2_insert64 (
);

FILL FILL_4_BUFX2_insert65 (
);

FILL FILL_5__7815_ (
);

FILL FILL111960x38050 (
);

FILL FILL_4_BUFX2_insert66 (
);

FILL FILL_1__10392_ (
);

FILL FILL_4_BUFX2_insert67 (
);

FILL FILL_4_BUFX2_insert68 (
);

FILL FILL_4_BUFX2_insert69 (
);

AOI21X1 _14955_ (
    .A(\datapath_1.regfile_1.regOut[14] [31]),
    .B(_4154_),
    .C(_5435_),
    .Y(_5436_)
);

OAI22X1 _14535_ (
    .A(_5024_),
    .B(_3941_),
    .C(_3949_),
    .D(_5023_),
    .Y(_5025_)
);

OAI22X1 _14115_ (
    .A(_4612_),
    .B(_3955__bF$buf2),
    .C(_3954__bF$buf2),
    .D(_4613_),
    .Y(_4614_)
);

FILL FILL_1__7807_ (
);

FILL FILL_0__15611_ (
);

FILL FILL_5__12997_ (
);

FILL FILL_5__12577_ (
);

FILL FILL_5__12157_ (
);

BUFX2 _6877_ (
    .A(_2_[7]),
    .Y(memoryWriteData[7])
);

FILL FILL_2__12184_ (
);

FILL SFILL114440x50050 (
);

FILL FILL_1__11597_ (
);

FILL FILL_1__11177_ (
);

FILL FILL_4__12511_ (
);

FILL FILL_0__8184_ (
);

INVX1 _10875_ (
    .A(_2022_),
    .Y(_2023_)
);

FILL FILL_6__9151_ (
);

DFFSR _10455_ (
    .Q(\datapath_1.regfile_1.regOut[28] [1]),
    .CLK(clk_bF$buf35),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_1758_[1])
);

NAND2X1 _10035_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1603_)
);

FILL FILL_3__11924_ (
);

FILL FILL_6__14789_ (
);

FILL FILL_3__11504_ (
);

FILL FILL_2__9983_ (
);

FILL FILL_2__10917_ (
);

FILL FILL_0__11951_ (
);

FILL FILL_2__9143_ (
);

FILL FILL_3__14396_ (
);

FILL FILL_0__11531_ (
);

FILL FILL_0__11111_ (
);

FILL FILL_4__9489_ (
);

FILL FILL_2__13389_ (
);

FILL FILL_5__14723_ (
);

FILL FILL_5__14303_ (
);

FILL FILL_0__6917_ (
);

NAND2X1 _8603_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_872_)
);

FILL FILL_1__7980_ (
);

FILL FILL_1__7560_ (
);

FILL FILL_4__13716_ (
);

FILL SFILL93800x34050 (
);

FILL FILL_2__14750_ (
);

FILL FILL_2__14330_ (
);

FILL FILL_3__7486_ (
);

FILL FILL_0__9389_ (
);

FILL FILL_3__7066_ (
);

FILL FILL_3__12709_ (
);

FILL FILL_1__13743_ (
);

FILL FILL_1__13323_ (
);

FILL FILL_4__16188_ (
);

FILL FILL_6__10289_ (
);

FILL FILL_0__12736_ (
);

NAND2X1 _12601_ (
    .A(vdd),
    .B(memoryOutData[11]),
    .Y(_3447_)
);

FILL FILL_0__12316_ (
);

FILL SFILL114360x12050 (
);

FILL FILL_5__8773_ (
);

FILL FILL_5__8353_ (
);

OAI22X1 _15493_ (
    .A(_5463__bF$buf2),
    .B(_5962_),
    .C(_5961_),
    .D(_5504__bF$buf2),
    .Y(_5963_)
);

FILL FILL_5__15928_ (
);

OAI21X1 _15073_ (
    .A(_5552__bF$buf2),
    .B(_3952_),
    .C(_5551_),
    .Y(_5553_)
);

FILL FILL_5__15508_ (
);

FILL FILL_3__16122_ (
);

INVX1 _9808_ (
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_1492_)
);

FILL FILL_1__8765_ (
);

FILL FILL_5__10643_ (
);

FILL FILL_1__8345_ (
);

FILL FILL_2__15955_ (
);

FILL FILL_2__15535_ (
);

FILL FILL_2__15115_ (
);

FILL FILL_2__10670_ (
);

FILL FILL_2__10250_ (
);

FILL FILL_1__14948_ (
);

FILL FILL_1__14528_ (
);

FILL FILL_1__14108_ (
);

FILL SFILL59720x35050 (
);

FILL FILL_3__9632_ (
);

AOI22X1 _13806_ (
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .B(_3894_),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_4311_)
);

FILL FILL_3__9212_ (
);

FILL FILL_5__9978_ (
);

FILL SFILL104360x55050 (
);

FILL FILL_5__9138_ (
);

INVX1 _16278_ (
    .A(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_6728_)
);

FILL FILL_5__11848_ (
);

FILL FILL_3__12882_ (
);

FILL FILL_5__11428_ (
);

FILL FILL_3__12462_ (
);

FILL FILL_5__11008_ (
);

FILL FILL_3__12042_ (
);

FILL SFILL108680x63050 (
);

FILL FILL_4__7975_ (
);

FILL FILL_4__7555_ (
);

FILL FILL_2__11875_ (
);

FILL FILL_2__11455_ (
);

FILL SFILL99400x17050 (
);

FILL FILL_2__11035_ (
);

FILL FILL_1__10448_ (
);

FILL FILL_1__10028_ (
);

FILL FILL_5__15681_ (
);

FILL FILL_5__15261_ (
);

FILL FILL_0__7875_ (
);

FILL FILL_6__8842_ (
);

NAND2X1 _9981_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1567_)
);

FILL FILL_0__7455_ (
);

FILL SFILL59240x28050 (
);

FILL FILL112440x61050 (
);

DFFSR _9561_ (
    .Q(\datapath_1.regfile_1.regOut[21] [3]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_1303_[3])
);

FILL FILL_0__7035_ (
);

INVX1 _9141_ (
    .A(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_1149_)
);

FILL FILL_4__14674_ (
);

FILL SFILL104360x10050 (
);

FILL FILL_4__14254_ (
);

OAI21X1 _12198_ (
    .A(_3184_),
    .B(ALUSrcA_bF$buf5),
    .C(_3185_),
    .Y(\datapath_1.alu_1.ALUInA [27])
);

FILL FILL_2__8834_ (
);

FILL FILL_3__13667_ (
);

FILL FILL_0__10802_ (
);

FILL FILL_3__13247_ (
);

FILL FILL_1__14281_ (
);

FILL FILL_0_BUFX2_insert610 (
);

FILL FILL_0_BUFX2_insert611 (
);

FILL FILL_0_BUFX2_insert612 (
);

FILL FILL_0_BUFX2_insert613 (
);

FILL FILL_0_BUFX2_insert614 (
);

FILL FILL_0__13694_ (
);

FILL FILL_0__13274_ (
);

FILL FILL_0_BUFX2_insert615 (
);

FILL FILL_0_BUFX2_insert616 (
);

FILL FILL_0_BUFX2_insert617 (
);

FILL FILL_0_BUFX2_insert618 (
);

FILL FILL_0_BUFX2_insert619 (
);

FILL FILL_2__13601_ (
);

FILL FILL_5__16046_ (
);

FILL FILL_6__9627_ (
);

FILL FILL_5__11181_ (
);

FILL FILL_4__15879_ (
);

FILL FILL_4__15459_ (
);

FILL FILL_4__15039_ (
);

FILL FILL_2__16073_ (
);

FILL FILL_4__10174_ (
);

FILL FILL_0__9601_ (
);

FILL FILL_2__9619_ (
);

FILL FILL_1__15486_ (
);

FILL FILL_1__15066_ (
);

FILL FILL_5__7624_ (
);

FILL FILL_5__7204_ (
);

FILL FILL_4__16400_ (
);

FILL FILL_0__14899_ (
);

FILL FILL_0__14479_ (
);

NAND3X1 _14764_ (
    .A(_5247_),
    .B(_5248_),
    .C(_5246_),
    .Y(_5249_)
);

FILL FILL_0__14059_ (
);

AOI22X1 _14344_ (
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .B(_4102_),
    .C(_3998__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_4838_)
);

FILL FILL_3__15813_ (
);

FILL SFILL89400x15050 (
);

FILL FILL_1__7616_ (
);

FILL SFILL94280x66050 (
);

FILL FILL_6__13393_ (
);

FILL FILL_2__14806_ (
);

FILL FILL_0__15840_ (
);

FILL FILL_0__15420_ (
);

FILL FILL_0__15000_ (
);

FILL FILL_5__12386_ (
);

FILL FILL_4__11799_ (
);

FILL FILL_4__8093_ (
);

FILL FILL_4__11379_ (
);

FILL FILL_3__8903_ (
);

FILL FILL_5__8829_ (
);

AOI22X1 _15969_ (
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .B(_5606_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_6426_)
);

FILL FILL_4__12740_ (
);

NOR2X1 _15549_ (
    .A(_6016_),
    .B(_6010_),
    .Y(_6017_)
);

FILL FILL_4__12320_ (
);

AOI22X1 _15129_ (
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .B(_5606_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_5607_)
);

NAND2X1 _10684_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1934_)
);

FILL FILL_0__10399_ (
);

NAND2X1 _10264_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1715_)
);

FILL FILL_2__6900_ (
);

FILL FILL_3__11733_ (
);

FILL FILL_3__11313_ (
);

FILL FILL_0__16205_ (
);

FILL FILL_2__9792_ (
);

FILL FILL_2__9372_ (
);

FILL FILL_0__11760_ (
);

FILL FILL_2__10306_ (
);

FILL FILL_0__11340_ (
);

FILL FILL_4__9298_ (
);

FILL FILL_5__14952_ (
);

FILL FILL_5__14532_ (
);

FILL FILL_5__14112_ (
);

NAND2X1 _8832_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_984_)
);

FILL SFILL8680x83050 (
);

DFFSR _8412_ (
    .Q(\datapath_1.regfile_1.regOut[12] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_718_[6])
);

FILL SFILL33960x17050 (
);

FILL FILL_4__13945_ (
);

FILL FILL_4__13525_ (
);

FILL FILL_4__13105_ (
);

FILL FILL_3__7295_ (
);

OAI21X1 _11889_ (
    .A(_3030_),
    .B(IorD_bF$buf2),
    .C(_3031_),
    .Y(_1_[0])
);

OAI21X1 _11469_ (
    .A(_2344__bF$buf0),
    .B(_2291_),
    .C(_2347__bF$buf0),
    .Y(_2584_)
);

XOR2X1 _11049_ (
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2168_)
);

FILL FILL_3__12518_ (
);

FILL FILL_1__13972_ (
);

FILL FILL_1__13552_ (
);

FILL FILL_1__13132_ (
);

FILL SFILL84280x64050 (
);

FILL FILL_0__12965_ (
);

NAND2X1 _12830_ (
    .A(vdd),
    .B(\datapath_1.rd1 [2]),
    .Y(_3559_)
);

NAND2X1 _12410_ (
    .A(MemToReg_bF$buf2),
    .B(\datapath_1.Data [22]),
    .Y(_3339_)
);

FILL FILL_0__12125_ (
);

FILL FILL_6__16324_ (
);

FILL FILL_5__8582_ (
);

FILL FILL_5__15737_ (
);

FILL FILL_5__15317_ (
);

FILL FILL_3__16351_ (
);

FILL SFILL8600x81050 (
);

INVX1 _9617_ (
    .A(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_1385_)
);

FILL FILL_1__8994_ (
);

FILL FILL_5__10872_ (
);

FILL FILL_5__10452_ (
);

FILL FILL_1__8574_ (
);

FILL FILL_5__10032_ (
);

FILL FILL_2__15764_ (
);

FILL FILL_2__15344_ (
);

FILL FILL_1__14757_ (
);

FILL FILL_1__14337_ (
);

FILL SFILL69400x56050 (
);

FILL SFILL84200x62050 (
);

FILL SFILL23560x46050 (
);

FILL FILL_3__9861_ (
);

INVX1 _13615_ (
    .A(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_4124_)
);

FILL FILL_3__9021_ (
);

FILL FILL_5__9787_ (
);

FILL FILL_5__9367_ (
);

FILL FILL_6__12244_ (
);

FILL SFILL13640x82050 (
);

AOI21X1 _16087_ (
    .A(_6541_),
    .B(_6522_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [25])
);

FILL SFILL23160x32050 (
);

FILL FILL_1__9779_ (
);

FILL FILL_5__11657_ (
);

FILL FILL_1__9359_ (
);

FILL FILL_5__11237_ (
);

FILL FILL_3__12271_ (
);

FILL FILL_2__16129_ (
);

FILL FILL_4__7364_ (
);

FILL FILL_2__11684_ (
);

FILL SFILL114440x45050 (
);

FILL FILL_2__11264_ (
);

FILL FILL_1__10677_ (
);

FILL FILL_1__10257_ (
);

FILL FILL_5__15490_ (
);

FILL FILL_0__7684_ (
);

FILL FILL_5__15070_ (
);

FILL SFILL74280x62050 (
);

INVX1 _9790_ (
    .A(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_1480_)
);

INVX1 _9370_ (
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_1261_)
);

FILL FILL_6__13449_ (
);

FILL FILL_4__14483_ (
);

FILL FILL_4__14063_ (
);

FILL SFILL114840x14050 (
);

FILL FILL_3__13896_ (
);

FILL FILL_2__8643_ (
);

FILL FILL_3__13476_ (
);

FILL FILL_2__8223_ (
);

FILL FILL_1__14090_ (
);

FILL FILL_6__14810_ (
);

FILL FILL_4__8989_ (
);

FILL FILL_4__8569_ (
);

FILL FILL_4__8149_ (
);

FILL FILL_2__12889_ (
);

FILL FILL_2__12469_ (
);

FILL FILL_2__12049_ (
);

FILL FILL_0__13083_ (
);

FILL FILL_5__13803_ (
);

FILL FILL_4__9930_ (
);

FILL FILL_4__9510_ (
);

FILL FILL_2__13830_ (
);

FILL FILL_3__6986_ (
);

FILL FILL_2__13410_ (
);

FILL FILL_0__8889_ (
);

FILL FILL_5__16275_ (
);

FILL SFILL74200x60050 (
);

FILL FILL_0__8469_ (
);

FILL SFILL13560x44050 (
);

FILL FILL_4__15688_ (
);

FILL FILL_1__12823_ (
);

FILL FILL_1__12403_ (
);

FILL FILL_4__15268_ (
);

FILL FILL_2__9848_ (
);

FILL FILL_2__9428_ (
);

FILL FILL_0__11816_ (
);

FILL FILL_0__9410_ (
);

FILL FILL_2__9008_ (
);

FILL FILL_1__15295_ (
);

FILL FILL_5__7853_ (
);

FILL FILL_5__7433_ (
);

OAI22X1 _14993_ (
    .A(_3897_),
    .B(_5469__bF$buf1),
    .C(_5472__bF$buf3),
    .D(_3953_),
    .Y(_5473_)
);

INVX1 _14573_ (
    .A(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_5062_)
);

FILL FILL_6__10310_ (
);

FILL FILL_0__14288_ (
);

NOR2X1 _14153_ (
    .A(_4650_),
    .B(_4647_),
    .Y(_4651_)
);

FILL FILL_3__15622_ (
);

FILL FILL_3__15202_ (
);

FILL FILL_1__7845_ (
);

FILL FILL_1__7425_ (
);

FILL FILL_2__14615_ (
);

FILL FILL_5__12195_ (
);

FILL FILL_1__13608_ (
);

FILL FILL_4__11188_ (
);

FILL FILL_3__8712_ (
);

FILL FILL_5__8638_ (
);

FILL FILL_5__8218_ (
);

NAND2X1 _15778_ (
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .B(_5490_),
    .Y(_6240_)
);

INVX1 _15358_ (
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_5831_)
);

FILL FILL_3__16407_ (
);

NAND2X1 _10493_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1827_)
);

DFFSR _10073_ (
    .Q(\datapath_1.regfile_1.regOut[25] [3]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf58),
    .S(vdd),
    .D(_1563_[3])
);

FILL FILL_5__10928_ (
);

FILL FILL_5__10508_ (
);

FILL FILL_3__11962_ (
);

FILL FILL_3__11542_ (
);

FILL FILL_3__11122_ (
);

FILL FILL_0__16014_ (
);

FILL FILL_2__10955_ (
);

FILL FILL_2__10535_ (
);

FILL FILL_2__10115_ (
);

FILL FILL_3__9917_ (
);

FILL FILL_5__14761_ (
);

FILL FILL_5__14341_ (
);

FILL FILL_0__6955_ (
);

FILL FILL112440x56050 (
);

FILL FILL_6__7502_ (
);

INVX1 _8641_ (
    .A(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_897_)
);

INVX1 _8221_ (
    .A(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_678_)
);

FILL FILL_4__13754_ (
);

FILL FILL_4__13334_ (
);

NAND3X1 _11698_ (
    .A(_2794_),
    .B(_2795_),
    .C(_2797_),
    .Y(_2798_)
);

NOR2X1 _11278_ (
    .A(_2396_),
    .B(_2206_),
    .Y(_2397_)
);

FILL SFILL49320x59050 (
);

FILL FILL_3__12747_ (
);

FILL FILL_1__13781_ (
);

FILL FILL_3__12327_ (
);

FILL FILL_1__13361_ (
);

FILL FILL112040x42050 (
);

FILL FILL_0__12774_ (
);

FILL FILL_0__12354_ (
);

FILL FILL_5__8391_ (
);

FILL FILL_5__15966_ (
);

FILL FILL_5__15546_ (
);

FILL FILL_5__15126_ (
);

FILL FILL_6__8707_ (
);

INVX1 _9846_ (
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_1561_)
);

FILL FILL_3__16160_ (
);

OAI21X1 _9426_ (
    .A(_1297_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .C(_1298_),
    .Y(_1238_[30])
);

FILL FILL_5__10681_ (
);

OAI21X1 _9006_ (
    .A(_1078_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .C(_1079_),
    .Y(_1043_[18])
);

FILL FILL_1__8383_ (
);

FILL FILL_5__10261_ (
);

FILL FILL_4__14959_ (
);

FILL FILL112440x11050 (
);

FILL FILL_2__15993_ (
);

FILL FILL_4__14539_ (
);

FILL FILL_2__15573_ (
);

FILL FILL_4__14119_ (
);

FILL FILL_2__15153_ (
);

FILL FILL_1__14986_ (
);

FILL FILL_1__14566_ (
);

FILL FILL_1__14146_ (
);

FILL FILL_4__15900_ (
);

FILL FILL_0__13979_ (
);

FILL FILL_3__9670_ (
);

INVX1 _13844_ (
    .A(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_4348_)
);

FILL FILL_3__9250_ (
);

FILL FILL_0__13559_ (
);

NAND3X1 _13424_ (
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3892_),
    .C(_3904_),
    .Y(_3936_)
);

FILL FILL_0__13139_ (
);

OAI21X1 _13004_ (
    .A(_3653_),
    .B(vdd),
    .C(_3654_),
    .Y(_3620_[17])
);

FILL FILL_5__9596_ (
);

FILL SFILL73800x25050 (
);

FILL FILL_0__14920_ (
);

FILL FILL_0__14500_ (
);

FILL FILL_5__11886_ (
);

FILL FILL_5__11466_ (
);

FILL FILL_1__9168_ (
);

FILL FILL_5__11046_ (
);

FILL FILL_3__12080_ (
);

FILL FILL_2__16358_ (
);

FILL FILL_4__7593_ (
);

FILL FILL_4__10879_ (
);

FILL FILL_4__7173_ (
);

FILL FILL_4__10039_ (
);

FILL FILL_2__11493_ (
);

FILL FILL_2__11073_ (
);

FILL FILL_6__7099_ (
);

FILL FILL_1__10486_ (
);

FILL FILL_1__10066_ (
);

AOI21X1 _14629_ (
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .B(_4246_),
    .C(_5116_),
    .Y(_5117_)
);

FILL FILL_4__11820_ (
);

INVX1 _14209_ (
    .A(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_4706_)
);

FILL FILL_4__11400_ (
);

FILL FILL_0__7493_ (
);

FILL FILL_0__7073_ (
);

FILL FILL_3__10813_ (
);

FILL FILL_4__14292_ (
);

FILL FILL_0__15705_ (
);

FILL FILL_2__8872_ (
);

FILL FILL_2__8452_ (
);

FILL FILL_3__13285_ (
);

FILL FILL_0__10420_ (
);

FILL FILL_0__10000_ (
);

FILL FILL_4__8378_ (
);

FILL FILL_2__12698_ (
);

FILL FILL_2__12278_ (
);

FILL FILL_5__13612_ (
);

FILL SFILL8680x78050 (
);

DFFSR _7912_ (
    .Q(\datapath_1.regfile_1.regOut[8] [18]),
    .CLK(clk_bF$buf5),
    .R(rst_bF$buf83),
    .S(vdd),
    .D(_458_[18])
);

FILL FILL_4__12605_ (
);

FILL FILL_5__16084_ (
);

FILL FILL_0__8698_ (
);

OAI22X1 _10969_ (
    .A(_2065_),
    .B(_2068_),
    .C(_2092_),
    .D(_2043_),
    .Y(_2044_)
);

INVX1 _10549_ (
    .A(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_1864_)
);

FILL FILL_6__9245_ (
);

INVX1 _10129_ (
    .A(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_1645_)
);

FILL FILL_1__12632_ (
);

FILL FILL_4__15497_ (
);

FILL FILL_4__15077_ (
);

FILL FILL_1__12212_ (
);

FILL SFILL94200x14050 (
);

FILL SFILL84280x59050 (
);

FILL FILL_2__9657_ (
);

OAI21X1 _11910_ (
    .A(_2980_),
    .B(IorD_bF$buf5),
    .C(_2981_),
    .Y(_1_[7])
);

FILL FILL_2__9237_ (
);

FILL FILL_0__11625_ (
);

FILL FILL_0__11205_ (
);

FILL FILL_5__7242_ (
);

INVX1 _14382_ (
    .A(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_4875_)
);

FILL FILL_0__14097_ (
);

FILL FILL_5__14817_ (
);

FILL FILL_3__15851_ (
);

FILL SFILL8600x76050 (
);

FILL FILL_3__15431_ (
);

FILL FILL_3__15011_ (
);

FILL SFILL59640x5050 (
);

FILL FILL_1__7234_ (
);

FILL SFILL8680x33050 (
);

FILL FILL_2__14844_ (
);

FILL SFILL13720x70050 (
);

FILL FILL_2__14424_ (
);

FILL FILL_2__14004_ (
);

FILL SFILL109560x50050 (
);

FILL FILL_1__13837_ (
);

FILL FILL_1__13417_ (
);

FILL SFILL84200x57050 (
);

FILL FILL_3__8521_ (
);

FILL SFILL99480x2050 (
);

FILL FILL_3__8101_ (
);

FILL SFILL84280x14050 (
);

FILL FILL_5__8867_ (
);

FILL FILL_5__8447_ (
);

FILL SFILL13640x77050 (
);

NOR3X1 _15587_ (
    .A(_5515__bF$buf2),
    .B(_4598_),
    .C(_5521__bF$buf1),
    .Y(_6054_)
);

AOI21X1 _15167_ (
    .A(_5622_),
    .B(_5644_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [2])
);

FILL SFILL109480x57050 (
);

FILL FILL_3__16216_ (
);

FILL FILL_1__8859_ (
);

FILL FILL_5__10317_ (
);

FILL FILL_1__8439_ (
);

FILL FILL_3__11771_ (
);

FILL FILL_1__8019_ (
);

FILL FILL_3__11351_ (
);

FILL FILL_2__15629_ (
);

FILL FILL_4__6864_ (
);

FILL FILL_2__15209_ (
);

FILL FILL_0__16243_ (
);

FILL FILL_2__10764_ (
);

OAI21X1 _7089_ (
    .A(_105_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_106_),
    .Y(_68_[19])
);

FILL FILL_1__9800_ (
);

FILL FILL_3__9726_ (
);

FILL FILL_5__14990_ (
);

FILL SFILL84200x12050 (
);

FILL FILL_5__14570_ (
);

FILL SFILL74280x57050 (
);

FILL FILL_5__14150_ (
);

INVX1 _8870_ (
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_1009_)
);

INVX1 _8450_ (
    .A(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_790_)
);

DFFSR _8030_ (
    .Q(\datapath_1.regfile_1.regOut[9] [8]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_523_[8])
);

FILL FILL_4__13983_ (
);

FILL FILL_4__13563_ (
);

FILL FILL_4__13143_ (
);

FILL SFILL13640x32050 (
);

FILL SFILL29240x17050 (
);

INVX2 _11087_ (
    .A(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2206_)
);

FILL FILL_3__12976_ (
);

FILL FILL_2__7723_ (
);

FILL FILL_2__7303_ (
);

FILL FILL_1__13590_ (
);

FILL FILL_3__12136_ (
);

FILL FILL_1__13170_ (
);

FILL FILL_4__7229_ (
);

FILL FILL_2__11969_ (
);

FILL FILL_2__11549_ (
);

FILL SFILL38840x81050 (
);

FILL FILL_0__12583_ (
);

FILL FILL_2__11129_ (
);

FILL FILL_0__12163_ (
);

FILL SFILL78920x77050 (
);

FILL FILL_2__12910_ (
);

FILL FILL_5__15775_ (
);

FILL SFILL74200x55050 (
);

FILL FILL_5__15355_ (
);

FILL FILL_0__7969_ (
);

FILL FILL_0__7549_ (
);

OAI21X1 _9655_ (
    .A(_1409_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1410_),
    .Y(_1368_[21])
);

FILL FILL_6__8516_ (
);

OAI21X1 _9235_ (
    .A(_1190_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1191_),
    .Y(_1173_[9])
);

FILL FILL_5__10490_ (
);

FILL FILL_1__8192_ (
);

FILL SFILL74280x12050 (
);

FILL FILL_1__11903_ (
);

FILL FILL_4__14768_ (
);

FILL FILL_4__14348_ (
);

FILL FILL_2__15382_ (
);

FILL FILL_0__8910_ (
);

FILL FILL_2__8508_ (
);

FILL FILL_1__14795_ (
);

FILL FILL_1__14375_ (
);

FILL FILL_5__6933_ (
);

FILL FILL_0__13788_ (
);

INVX1 _13653_ (
    .A(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_4161_)
);

FILL FILL_0__13368_ (
);

FILL SFILL3480x80050 (
);

INVX2 _13233_ (
    .A(_3770_),
    .Y(_3776_)
);

FILL FILL_3__14702_ (
);

FILL FILL_1__6925_ (
);

FILL FILL_5__11695_ (
);

FILL FILL112120x75050 (
);

FILL FILL_1__9397_ (
);

FILL FILL_5__11275_ (
);

FILL SFILL74200x10050 (
);

FILL FILL_2__16167_ (
);

FILL FILL_4__10688_ (
);

FILL FILL_4__10268_ (
);

FILL FILL_5__7718_ (
);

FILL FILL_2_BUFX2_insert520 (
);

FILL FILL_1__10295_ (
);

FILL FILL_2_BUFX2_insert521 (
);

FILL FILL_2_BUFX2_insert522 (
);

NAND3X1 _14858_ (
    .A(_5330_),
    .B(_5333_),
    .C(_5340_),
    .Y(_5341_)
);

FILL FILL_2_BUFX2_insert523 (
);

FILL FILL_2_BUFX2_insert524 (
);

NAND2X1 _14438_ (
    .A(_4929_),
    .B(_4922_),
    .Y(_4930_)
);

OAI22X1 _14018_ (
    .A(_3982__bF$buf1),
    .B(_4518_),
    .C(_3966__bF$buf0),
    .D(_4517_),
    .Y(_4519_)
);

FILL FILL_2_BUFX2_insert525 (
);

FILL FILL_3__15907_ (
);

FILL FILL_2_BUFX2_insert526 (
);

FILL FILL_2_BUFX2_insert527 (
);

FILL SFILL43720x26050 (
);

FILL FILL_2_BUFX2_insert528 (
);

FILL FILL_2_BUFX2_insert529 (
);

FILL FILL_1__16101_ (
);

FILL FILL_3__10622_ (
);

FILL FILL_0_CLKBUF1_insert220 (
);

FILL FILL_0_CLKBUF1_insert221 (
);

FILL FILL_0__15934_ (
);

FILL FILL_0_CLKBUF1_insert222 (
);

FILL FILL_0_CLKBUF1_insert223 (
);

FILL FILL_0__15514_ (
);

FILL FILL_0_CLKBUF1_insert224 (
);

FILL SFILL33800x62050 (
);

FILL FILL_2__8261_ (
);

FILL FILL_3__13094_ (
);

FILL FILL112120x30050 (
);

FILL FILL_4__8187_ (
);

FILL FILL_2__12087_ (
);

FILL FILL_5__13841_ (
);

FILL FILL_5__13421_ (
);

FILL FILL_5__13001_ (
);

INVX1 _7721_ (
    .A(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_426_)
);

INVX1 _7301_ (
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .Y(_207_)
);

FILL FILL_4__12834_ (
);

FILL FILL_4__12414_ (
);

FILL FILL_0__8087_ (
);

INVX1 _10778_ (
    .A(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_1976_)
);

INVX1 _10358_ (
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_1821_)
);

FILL FILL_3__11827_ (
);

FILL FILL_1__12861_ (
);

FILL FILL_3__11407_ (
);

FILL FILL_1__12441_ (
);

FILL FILL112040x37050 (
);

FILL FILL_1__12021_ (
);

FILL FILL_2__9886_ (
);

FILL FILL_0__11854_ (
);

FILL FILL_2__9466_ (
);

FILL FILL_3__14299_ (
);

FILL FILL_0__11434_ (
);

FILL FILL_0__11014_ (
);

FILL FILL_6__15633_ (
);

FILL FILL_5__7891_ (
);

FILL FILL_5__7471_ (
);

FILL FILL_5__7051_ (
);

INVX1 _14191_ (
    .A(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_4688_)
);

FILL FILL_5__14626_ (
);

FILL FILL_3__15660_ (
);

FILL FILL_5__14206_ (
);

DFFSR _8926_ (
    .Q(\datapath_1.regfile_1.regOut[16] [8]),
    .CLK(clk_bF$buf56),
    .R(rst_bF$buf92),
    .S(vdd),
    .D(_978_[8])
);

FILL FILL_3__15240_ (
);

OAI21X1 _8506_ (
    .A(_826_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_827_),
    .Y(_783_[22])
);

FILL FILL_1__7883_ (
);

FILL FILL_1__7463_ (
);

FILL FILL_1__7043_ (
);

FILL FILL_4__13619_ (
);

FILL FILL_2__14653_ (
);

FILL FILL_2__14233_ (
);

FILL FILL_1__13646_ (
);

FILL FILL_1__13226_ (
);

FILL FILL_1_BUFX2_insert540 (
);

FILL FILL_3__8750_ (
);

FILL FILL_1_BUFX2_insert541 (
);

FILL FILL_0__12639_ (
);

FILL FILL_3__8330_ (
);

FILL FILL_1_BUFX2_insert542 (
);

DFFSR _12924_ (
    .Q(\datapath_1.a [5]),
    .CLK(clk_bF$buf24),
    .R(rst_bF$buf105),
    .S(vdd),
    .D(_3555_[5])
);

OAI21X1 _12504_ (
    .A(_3401_),
    .B(vdd),
    .C(_3402_),
    .Y(_3360_[21])
);

FILL FILL_1_BUFX2_insert543 (
);

FILL FILL_0__12219_ (
);

FILL FILL_1_BUFX2_insert544 (
);

FILL FILL_1_BUFX2_insert545 (
);

FILL FILL_1_BUFX2_insert546 (
);

FILL FILL_5__8256_ (
);

FILL FILL_1_BUFX2_insert547 (
);

FILL FILL_1_BUFX2_insert548 (
);

FILL FILL_1_BUFX2_insert549 (
);

FILL FILL_6__11973_ (
);

FILL FILL_6__11553_ (
);

OAI22X1 _15396_ (
    .A(_5466__bF$buf0),
    .B(_4359_),
    .C(_4348_),
    .D(_5483__bF$buf3),
    .Y(_5868_)
);

FILL FILL_3__16025_ (
);

FILL FILL_5__10966_ (
);

FILL FILL_5__10546_ (
);

FILL FILL_5__10126_ (
);

FILL FILL_1__8248_ (
);

FILL FILL_3__11580_ (
);

FILL FILL_3__11160_ (
);

FILL FILL_2__15858_ (
);

FILL FILL_2__15438_ (
);

FILL FILL_2__15018_ (
);

FILL FILL_0__16052_ (
);

FILL FILL_2__10993_ (
);

FILL FILL_2__10573_ (
);

FILL FILL_2__10153_ (
);

FILL FILL_3__9535_ (
);

FILL FILL_4__10900_ (
);

FILL FILL_3__9115_ (
);

INVX1 _13709_ (
    .A(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_4216_)
);

FILL FILL_0__6993_ (
);

FILL FILL_6__7120_ (
);

FILL FILL_6__12758_ (
);

FILL FILL_4__13792_ (
);

FILL FILL_4__13372_ (
);

FILL FILL_2__7952_ (
);

FILL FILL_3__12785_ (
);

FILL FILL_3__12365_ (
);

FILL FILL_2__7112_ (
);

FILL FILL_4__7878_ (
);

FILL FILL_4__7458_ (
);

FILL FILL_4__7038_ (
);

FILL FILL_2__11778_ (
);

FILL FILL_2__11358_ (
);

FILL FILL_0__12392_ (
);

FILL FILL_6__16171_ (
);

FILL SFILL74120x1050 (
);

FILL SFILL23720x22050 (
);

FILL FILL_5__15584_ (
);

FILL FILL_5__15164_ (
);

FILL FILL_0__7358_ (
);

OAI21X1 _9884_ (
    .A(_1521_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .C(_1522_),
    .Y(_1498_[12])
);

OAI21X1 _9464_ (
    .A(_1366_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1367_),
    .Y(_1303_[0])
);

FILL FILL_6__8325_ (
);

NAND2X1 _9044_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1105_)
);

FILL FILL_4__14997_ (
);

FILL FILL_4__14577_ (
);

FILL FILL_1__11712_ (
);

FILL FILL_4__14157_ (
);

FILL FILL_2__15191_ (
);

FILL FILL_2__8737_ (
);

FILL FILL_0__10705_ (
);

FILL FILL_2__8317_ (
);

FILL FILL_1__14184_ (
);

FILL SFILL23640x29050 (
);

FILL FILL_0__13597_ (
);

NOR2X1 _13882_ (
    .A(_4385_),
    .B(_3971__bF$buf4),
    .Y(_4386_)
);

NOR2X1 _13462_ (
    .A(_3968_),
    .B(_3973_),
    .Y(_3974_)
);

NAND2X1 _13042_ (
    .A(vdd),
    .B(\datapath_1.rd2 [30]),
    .Y(_3680_)
);

FILL FILL_3__14931_ (
);

FILL FILL_3__14511_ (
);

FILL FILL_4__9604_ (
);

FILL FILL_2__13924_ (
);

FILL SFILL44120x56050 (
);

FILL FILL_5__16369_ (
);

FILL FILL_2__13504_ (
);

FILL SFILL109560x45050 (
);

FILL FILL_5__11084_ (
);

FILL FILL_1__12917_ (
);

FILL FILL_2__16396_ (
);

FILL FILL_4__10497_ (
);

FILL FILL_0__9924_ (
);

FILL FILL_0__9504_ (
);

FILL FILL_3__7601_ (
);

FILL FILL_1__15389_ (
);

FILL FILL_5__7947_ (
);

FILL SFILL109160x31050 (
);

FILL FILL_4__16303_ (
);

FILL FILL_5__7107_ (
);

NAND3X1 _14667_ (
    .A(_5145_),
    .B(_5146_),
    .C(_5153_),
    .Y(_5154_)
);

INVX1 _14247_ (
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_4743_)
);

FILL FILL_3__15716_ (
);

FILL FILL_1__16330_ (
);

FILL FILL_1__7939_ (
);

FILL FILL_3__10431_ (
);

FILL FILL_3__10011_ (
);

FILL FILL_2__14709_ (
);

FILL FILL_0__15743_ (
);

FILL FILL_0__15323_ (
);

FILL SFILL13720x20050 (
);

FILL FILL_5__12289_ (
);

FILL FILL_2__8490_ (
);

FILL FILL_2__8070_ (
);

FILL FILL_5__13650_ (
);

FILL FILL_5__13230_ (
);

INVX1 _7950_ (
    .A(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_538_)
);

DFFSR _7530_ (
    .Q(\datapath_1.regfile_1.regOut[5] [20]),
    .CLK(clk_bF$buf53),
    .R(rst_bF$buf80),
    .S(vdd),
    .D(_263_[20])
);

OAI21X1 _7110_ (
    .A(_119_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .C(_120_),
    .Y(_68_[26])
);

FILL FILL_4__12643_ (
);

FILL FILL_4__12223_ (
);

FILL SFILL13640x27050 (
);

DFFSR _10587_ (
    .Q(\datapath_1.regfile_1.regOut[29] [5]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf18),
    .S(vdd),
    .D(_1823_[5])
);

OAI21X1 _10167_ (
    .A(_1669_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .C(_1670_),
    .Y(_1628_[21])
);

FILL FILL_3__11636_ (
);

FILL FILL_3__11216_ (
);

FILL FILL_1__12250_ (
);

FILL FILL_0__16108_ (
);

FILL FILL_2__10629_ (
);

FILL FILL_2__9275_ (
);

FILL FILL_0__11663_ (
);

FILL FILL_0__11243_ (
);

FILL FILL_5__14855_ (
);

FILL FILL_5__14435_ (
);

FILL FILL_5__14015_ (
);

OAI21X1 _8735_ (
    .A(_938_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .C(_939_),
    .Y(_913_[13])
);

OAI21X1 _8315_ (
    .A(_719_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .C(_720_),
    .Y(_718_[1])
);

FILL FILL_1__7692_ (
);

FILL FILL_4__13848_ (
);

FILL FILL_4__13428_ (
);

FILL FILL_2__14882_ (
);

FILL FILL_2__14462_ (
);

FILL FILL_4__13008_ (
);

FILL FILL_2__14042_ (
);

FILL FILL_3__7198_ (
);

FILL FILL112200x63050 (
);

FILL FILL_1__13875_ (
);

FILL SFILL83880x71050 (
);

FILL SFILL99480x56050 (
);

FILL FILL_1__13455_ (
);

FILL FILL_1__13035_ (
);

FILL SFILL44040x5050 (
);

FILL FILL_0__12868_ (
);

OAI21X1 _12733_ (
    .A(_3513_),
    .B(IRWrite_bF$buf6),
    .C(_3514_),
    .Y(_3490_[12])
);

FILL FILL_0__12448_ (
);

FILL FILL_0__12028_ (
);

AOI22X1 _12313_ (
    .A(_2_[24]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3274_)
);

FILL FILL_6__16227_ (
);

FILL FILL_5__8485_ (
);

FILL FILL_5__8065_ (
);

FILL FILL_3__16254_ (
);

FILL SFILL43800x14050 (
);

FILL FILL_5__10775_ (
);

FILL FILL_1__8897_ (
);

FILL FILL_1__8477_ (
);

FILL FILL_1__8057_ (
);

FILL SFILL68200x80050 (
);

FILL FILL_2__15667_ (
);

FILL FILL_2__15247_ (
);

FILL FILL_0__16281_ (
);

FILL FILL_2__10382_ (
);

FILL SFILL99480x11050 (
);

FILL FILL_3__9764_ (
);

FILL FILL_3__9344_ (
);

INVX1 _13938_ (
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_4440_)
);

NOR2X1 _13518_ (
    .A(_4025_),
    .B(_4028_),
    .Y(_4029_)
);

FILL SFILL28840x74050 (
);

FILL FILL_1__15601_ (
);

FILL FILL_6__12147_ (
);

FILL FILL_2__7761_ (
);

FILL SFILL64200x48050 (
);

FILL FILL_3__12594_ (
);

FILL FILL_2__7341_ (
);

FILL FILL_3__12174_ (
);

FILL FILL112120x25050 (
);

FILL FILL_4__7687_ (
);

FILL FILL_2__11587_ (
);

FILL FILL_2__11167_ (
);

FILL FILL_5__12501_ (
);

FILL FILL_4__11914_ (
);

FILL FILL_5__15393_ (
);

FILL FILL_0__7587_ (
);

FILL FILL_0__7167_ (
);

DFFSR _9693_ (
    .Q(\datapath_1.regfile_1.regOut[22] [7]),
    .CLK(clk_bF$buf19),
    .R(rst_bF$buf101),
    .S(vdd),
    .D(_1368_[7])
);

NAND2X1 _9273_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1217_)
);

FILL FILL_3__10907_ (
);

FILL FILL_1__11941_ (
);

FILL FILL_4__14386_ (
);

FILL FILL_1__11521_ (
);

FILL FILL_1__11101_ (
);

FILL FILL_2__8966_ (
);

FILL FILL_3__13799_ (
);

FILL FILL_0__10934_ (
);

FILL FILL_2__8126_ (
);

FILL FILL_3__13379_ (
);

FILL FILL_0__10514_ (
);

FILL FILL_5__6971_ (
);

FILL FILL_6__14713_ (
);

FILL SFILL33800x12050 (
);

INVX1 _13691_ (
    .A(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_4198_)
);

INVX2 _13271_ (
    .A(_3764_),
    .Y(_3812_)
);

FILL FILL_5__13706_ (
);

FILL FILL_3__14740_ (
);

FILL FILL_3__14320_ (
);

FILL FILL_1__6963_ (
);

FILL FILL_4__9413_ (
);

FILL FILL_2__13733_ (
);

FILL FILL_2__13313_ (
);

FILL FILL_5__16178_ (
);

FILL FILL_3__6889_ (
);

FILL FILL_1__12726_ (
);

FILL FILL_1__12306_ (
);

FILL SFILL18840x72050 (
);

FILL FILL_0__9733_ (
);

FILL FILL_3__7830_ (
);

FILL FILL_0__11719_ (
);

FILL FILL_1__15198_ (
);

FILL FILL_5__7756_ (
);

FILL FILL_5__7336_ (
);

FILL FILL_2_BUFX2_insert900 (
);

FILL FILL_4__16112_ (
);

FILL FILL_2_BUFX2_insert901 (
);

FILL FILL_2_BUFX2_insert902 (
);

FILL FILL_2_BUFX2_insert903 (
);

INVX1 _14896_ (
    .A(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_5378_)
);

FILL FILL_2_BUFX2_insert904 (
);

OAI22X1 _14476_ (
    .A(_4965_),
    .B(_3890_),
    .C(_3960_),
    .D(_4966_),
    .Y(_4967_)
);

FILL FILL_2_BUFX2_insert905 (
);

INVX1 _14056_ (
    .A(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_4556_)
);

FILL FILL_2_BUFX2_insert906 (
);

FILL FILL_3__15945_ (
);

FILL FILL_2_BUFX2_insert907 (
);

FILL FILL_3__15525_ (
);

FILL FILL_2_BUFX2_insert908 (
);

FILL FILL_3__15105_ (
);

FILL FILL_2_BUFX2_insert909 (
);

FILL SFILL13720x7050 (
);

FILL FILL_1__7748_ (
);

FILL FILL_3__10660_ (
);

FILL FILL_1__7328_ (
);

FILL FILL_3__10240_ (
);

FILL FILL_2__14938_ (
);

FILL FILL_0__15972_ (
);

FILL FILL_2__14518_ (
);

FILL FILL_0__15552_ (
);

FILL FILL_0__15132_ (
);

FILL FILL_5__12098_ (
);

FILL FILL_3__8615_ (
);

FILL FILL_4__12872_ (
);

FILL SFILL58920x23050 (
);

FILL FILL_4__12452_ (
);

FILL FILL_4__12032_ (
);

OAI21X1 _10396_ (
    .A(_1781_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1782_),
    .Y(_1758_[12])
);

FILL FILL_3__11865_ (
);

FILL FILL_5__9902_ (
);

FILL FILL_3__11445_ (
);

FILL FILL_3__11025_ (
);

FILL FILL_4__6958_ (
);

FILL FILL_0__16337_ (
);

NOR3X1 _16202_ (
    .A(_6653_),
    .B(_6632_),
    .C(_6642_),
    .Y(_6654_)
);

FILL FILL_2__10438_ (
);

FILL FILL_0__11892_ (
);

FILL FILL_2__10018_ (
);

FILL FILL_2__9084_ (
);

FILL FILL_0__11472_ (
);

FILL FILL_0__11052_ (
);

FILL SFILL23720x17050 (
);

FILL FILL_5__14664_ (
);

FILL FILL_5__14244_ (
);

FILL FILL_0__6858_ (
);

OAI21X1 _8964_ (
    .A(_1050_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1051_),
    .Y(_1043_[4])
);

DFFSR _8544_ (
    .Q(\datapath_1.regfile_1.regOut[13] [10]),
    .CLK(clk_bF$buf87),
    .R(rst_bF$buf43),
    .S(vdd),
    .D(_783_[10])
);

NAND2X1 _8124_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_634_)
);

FILL FILL_1__7081_ (
);

FILL FILL_4__13657_ (
);

FILL SFILL48920x66050 (
);

FILL FILL_4__13237_ (
);

FILL FILL_2__14691_ (
);

FILL FILL_2__14271_ (
);

FILL FILL_2__7817_ (
);

FILL FILL_1__13684_ (
);

FILL FILL_1__13264_ (
);

FILL FILL_1_BUFX2_insert920 (
);

FILL FILL_1_BUFX2_insert921 (
);

OAI21X1 _12962_ (
    .A(_3625_),
    .B(vdd),
    .C(_3626_),
    .Y(_3620_[3])
);

FILL FILL_1_BUFX2_insert922 (
);

DFFSR _12542_ (
    .Q(ALUOut[7]),
    .CLK(clk_bF$buf39),
    .R(rst_bF$buf73),
    .S(vdd),
    .D(_3360_[7])
);

FILL FILL_1_BUFX2_insert923 (
);

FILL FILL_0__12257_ (
);

FILL FILL_1_BUFX2_insert924 (
);

NAND2X1 _12122_ (
    .A(ALUSrcA_bF$buf0),
    .B(\datapath_1.a [2]),
    .Y(_3135_)
);

FILL FILL_1_BUFX2_insert925 (
);

FILL FILL_1_BUFX2_insert926 (
);

FILL FILL_1_BUFX2_insert927 (
);

FILL FILL_1_BUFX2_insert928 (
);

FILL FILL_1_BUFX2_insert929 (
);

FILL FILL_5__15869_ (
);

FILL FILL_5__15449_ (
);

FILL FILL_5__15029_ (
);

FILL FILL_3__16063_ (
);

NAND2X1 _9749_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1453_)
);

DFFSR _9329_ (
    .Q(\datapath_1.regfile_1.regOut[19] [27]),
    .CLK(clk_bF$buf54),
    .R(rst_bF$buf21),
    .S(vdd),
    .D(_1173_[27])
);

FILL FILL_5__10164_ (
);

FILL FILL_2__15896_ (
);

FILL FILL_2__15476_ (
);

FILL FILL_2__15056_ (
);

FILL FILL_0__16090_ (
);

FILL SFILL48920x21050 (
);

FILL FILL_2__10191_ (
);

FILL FILL_1__14889_ (
);

FILL FILL_1__14469_ (
);

FILL FILL_1__14049_ (
);

FILL FILL_4__15803_ (
);

FILL FILL_3__9993_ (
);

INVX1 _13747_ (
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_4253_)
);

FILL FILL_3__9153_ (
);

AND2X2 _13327_ (
    .A(_3784_),
    .B(RegWrite_bF$buf0),
    .Y(\datapath_1.regfile_1.regEn [16])
);

FILL FILL_5__9499_ (
);

FILL FILL_1__15830_ (
);

FILL FILL_1__15410_ (
);

FILL FILL_5__9079_ (
);

FILL FILL_0__14823_ (
);

FILL FILL_0__14403_ (
);

FILL SFILL13720x15050 (
);

FILL FILL_2__7990_ (
);

FILL FILL_5__11789_ (
);

FILL FILL_5__11369_ (
);

FILL FILL_2__7570_ (
);

FILL FILL_4__7496_ (
);

FILL FILL_4__7076_ (
);

FILL FILL_2__11396_ (
);

FILL SFILL38920x64050 (
);

FILL FILL_5__12730_ (
);

FILL FILL_5__12310_ (
);

FILL FILL_1__10389_ (
);

FILL FILL_4__11723_ (
);

FILL FILL_4__11303_ (
);

NAND2X1 _9082_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1110_)
);

FILL FILL_1__11750_ (
);

FILL FILL_4__14195_ (
);

FILL FILL_1__11330_ (
);

FILL FILL_0__15608_ (
);

FILL FILL_2__8775_ (
);

FILL FILL_2__8355_ (
);

FILL FILL_0__10743_ (
);

FILL FILL_0__10323_ (
);

FILL SFILL3560x63050 (
);

NAND2X1 _13080_ (
    .A(\datapath_1.mux_pcsrc.dout [0]),
    .B(PCEn_bF$buf4),
    .Y(_3749_)
);

FILL FILL_5__13935_ (
);

FILL FILL_5__13515_ (
);

OAI21X1 _7815_ (
    .A(_467_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_468_),
    .Y(_458_[5])
);

FILL FILL_4_BUFX2_insert430 (
);

FILL FILL_4_BUFX2_insert431 (
);

FILL FILL_4__9642_ (
);

FILL FILL_4__9222_ (
);

FILL FILL_4_BUFX2_insert432 (
);

FILL FILL_4_BUFX2_insert433 (
);

FILL FILL_4__12508_ (
);

FILL FILL_2__13962_ (
);

FILL FILL_4_BUFX2_insert434 (
);

FILL FILL_2__13542_ (
);

FILL FILL_2__13122_ (
);

FILL FILL_4_BUFX2_insert435 (
);

FILL FILL_4_BUFX2_insert436 (
);

FILL FILL_4_BUFX2_insert437 (
);

FILL FILL_4_BUFX2_insert438 (
);

FILL FILL112200x58050 (
);

FILL FILL_4_BUFX2_insert439 (
);

FILL FILL_1__12955_ (
);

FILL FILL_1__12115_ (
);

FILL FILL_0__11948_ (
);

FILL FILL_0__9542_ (
);

FILL FILL_0__9122_ (
);

OAI22X1 _11813_ (
    .A(_2124_),
    .B(_2344__bF$buf3),
    .C(_2480_),
    .D(_2123_),
    .Y(_2904_)
);

FILL FILL_0__11528_ (
);

FILL FILL_0__11108_ (
);

FILL SFILL38840x26050 (
);

FILL FILL_5__7985_ (
);

FILL FILL_5__7565_ (
);

FILL FILL_4__16341_ (
);

NOR2X1 _14285_ (
    .A(_4779_),
    .B(_3955__bF$buf2),
    .Y(_4780_)
);

FILL FILL_3__15754_ (
);

FILL FILL_3__15334_ (
);

FILL FILL_1__7977_ (
);

FILL FILL_1__7557_ (
);

FILL FILL_2__14747_ (
);

FILL SFILL89160x73050 (
);

FILL FILL_0__15781_ (
);

FILL FILL_2__14327_ (
);

FILL FILL_0__15361_ (
);

FILL FILL112200x13050 (
);

FILL FILL_3__8844_ (
);

FILL FILL_3__8004_ (
);

FILL SFILL28840x69050 (
);

FILL SFILL68600x44050 (
);

FILL FILL_4__12261_ (
);

FILL FILL_3__16119_ (
);

FILL FILL_2__6841_ (
);

FILL FILL_3__11674_ (
);

FILL FILL_3__11254_ (
);

DFFSR _16431_ (
    .Q(\datapath_1.regfile_1.regOut[0] [14]),
    .CLK(clk_bF$buf48),
    .R(rst_bF$buf85),
    .S(vdd),
    .D(_6769_[14])
);

FILL FILL_0__16146_ (
);

AOI22X1 _16011_ (
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [24]),
    .C(\datapath_1.regfile_1.regOut[10] [24]),
    .D(_6314_),
    .Y(_6467_)
);

FILL FILL_2__10667_ (
);

FILL FILL_2__10247_ (
);

FILL FILL_0__11281_ (
);

FILL FILL_6__15480_ (
);

FILL FILL_6__15060_ (
);

FILL SFILL115000x46050 (
);

FILL FILL_3_BUFX2_insert450 (
);

FILL FILL_3__9629_ (
);

FILL FILL_3_BUFX2_insert451 (
);

FILL FILL_3__9209_ (
);

FILL FILL_5__14893_ (
);

FILL FILL_3_BUFX2_insert452 (
);

FILL FILL_3_BUFX2_insert453 (
);

FILL FILL_5__14473_ (
);

FILL FILL_3_BUFX2_insert454 (
);

FILL FILL_5__14053_ (
);

NAND2X1 _8773_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_965_)
);

FILL FILL_3_BUFX2_insert455 (
);

NAND2X1 _8353_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_746_)
);

FILL FILL_3_BUFX2_insert456 (
);

FILL FILL_3_BUFX2_insert457 (
);

FILL FILL_3_BUFX2_insert458 (
);

FILL FILL_4__13886_ (
);

FILL FILL_3_BUFX2_insert459 (
);

FILL FILL_4__13466_ (
);

FILL FILL_4__13046_ (
);

FILL FILL_2__14080_ (
);

FILL FILL_2__7626_ (
);

FILL FILL_3__12879_ (
);

FILL FILL_3__12459_ (
);

FILL FILL_2__7206_ (
);

FILL FILL_3__12039_ (
);

FILL FILL_1__13493_ (
);

NAND2X1 _12771_ (
    .A(IRWrite_bF$buf3),
    .B(memoryOutData[25]),
    .Y(_3540_)
);

FILL FILL_0__12486_ (
);

OAI21X1 _12351_ (
    .A(_3298_),
    .B(MemToReg_bF$buf0),
    .C(_3299_),
    .Y(\datapath_1.mux_wd3.dout [2])
);

FILL FILL_0__12066_ (
);

FILL FILL_3__13820_ (
);

FILL FILL_3__13400_ (
);

FILL FILL_4__8913_ (
);

FILL FILL_5__15678_ (
);

FILL FILL_5__15258_ (
);

FILL FILL_3__16292_ (
);

NAND2X1 _9978_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1565_)
);

DFFSR _9558_ (
    .Q(\datapath_1.regfile_1.regOut[21] [0]),
    .CLK(clk_bF$buf49),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_1303_[0])
);

INVX1 _9138_ (
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_1147_)
);

FILL FILL_5__10393_ (
);

FILL FILL_1__8095_ (
);

FILL FILL_1__11806_ (
);

FILL SFILL18840x67050 (
);

FILL FILL_2__15285_ (
);

FILL FILL_3__6910_ (
);

FILL FILL_1__14698_ (
);

FILL FILL_1__14278_ (
);

FILL FILL_5__6836_ (
);

FILL FILL_0_BUFX2_insert580 (
);

FILL FILL_0_BUFX2_insert581 (
);

FILL FILL_4__15612_ (
);

FILL FILL_0_BUFX2_insert582 (
);

FILL FILL_0_BUFX2_insert583 (
);

FILL FILL_3__9382_ (
);

AOI22X1 _13976_ (
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .B(_3891__bF$buf0),
    .C(_3998__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_4477_)
);

FILL FILL_0_BUFX2_insert584 (
);

FILL FILL_0_BUFX2_insert585 (
);

INVX1 _13556_ (
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_4066_)
);

INVX1 _13136_ (
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3722_)
);

FILL FILL_0_BUFX2_insert586 (
);

FILL FILL_0_BUFX2_insert587 (
);

FILL FILL_3__14605_ (
);

FILL FILL_0_BUFX2_insert588 (
);

FILL FILL_0_BUFX2_insert589 (
);

FILL FILL_0__14632_ (
);

FILL FILL_0__14212_ (
);

FILL FILL_5__11598_ (
);

FILL FILL_5__11178_ (
);

FILL SFILL18840x22050 (
);

FILL SFILL79080x33050 (
);

FILL FILL_4__11952_ (
);

FILL FILL_4__11532_ (
);

FILL FILL_4__11112_ (
);

FILL FILL_1__16004_ (
);

FILL FILL_3__10945_ (
);

FILL FILL_3__10525_ (
);

FILL FILL_3__10105_ (
);

FILL FILL_0__15837_ (
);

NOR3X1 _15702_ (
    .A(_6163_),
    .B(_6165_),
    .C(_6164_),
    .Y(_6166_)
);

FILL FILL_0__15417_ (
);

FILL FILL_2__8584_ (
);

FILL FILL_0__10972_ (
);

FILL FILL_0__10552_ (
);

FILL FILL_0__10132_ (
);

FILL FILL_5__13744_ (
);

FILL SFILL48600x40050 (
);

FILL FILL_5__13324_ (
);

NAND2X1 _7624_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_382_)
);

NAND2X1 _7204_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_163_)
);

FILL FILL_4__9871_ (
);

FILL FILL_4__12737_ (
);

FILL FILL_4__9031_ (
);

FILL FILL_2__13771_ (
);

FILL FILL_4__12317_ (
);

FILL FILL_2__13351_ (
);

FILL FILL_6__9797_ (
);

FILL FILL_1__12764_ (
);

FILL FILL_1__12344_ (
);

FILL FILL_2__9789_ (
);

FILL FILL_0__9771_ (
);

FILL FILL_2__9369_ (
);

FILL FILL_0__11757_ (
);

FILL FILL_0__9351_ (
);

FILL FILL_0__11337_ (
);

NOR2X1 _11622_ (
    .A(_2726_),
    .B(_2725_),
    .Y(_2727_)
);

FILL SFILL114520x70050 (
);

AND2X2 _11202_ (
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2321_)
);

FILL FILL_6__15956_ (
);

FILL FILL_6__15536_ (
);

FILL FILL_5__7374_ (
);

FILL SFILL109240x14050 (
);

FILL FILL_4__16150_ (
);

FILL FILL_5__14949_ (
);

AOI22X1 _14094_ (
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .B(_3885_),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_4593_)
);

FILL FILL_3__15983_ (
);

FILL FILL_5__14529_ (
);

FILL FILL_3__15563_ (
);

FILL FILL_5__14109_ (
);

FILL SFILL69000x74050 (
);

FILL FILL_3__15143_ (
);

NAND2X1 _8829_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_982_)
);

DFFSR _8409_ (
    .Q(\datapath_1.regfile_1.regOut[12] [3]),
    .CLK(clk_bF$buf28),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_718_[3])
);

FILL FILL_1__7366_ (
);

FILL FILL_2__14976_ (
);

FILL SFILL69080x31050 (
);

FILL FILL_2__14556_ (
);

FILL FILL_2__14136_ (
);

FILL FILL_0__15590_ (
);

FILL FILL_0__15170_ (
);

FILL SFILL48920x16050 (
);

FILL FILL_1__13969_ (
);

FILL FILL_1__13549_ (
);

FILL FILL_1__13129_ (
);

FILL FILL_3__8653_ (
);

FILL FILL_3__8233_ (
);

NAND2X1 _12827_ (
    .A(vdd),
    .B(\datapath_1.rd1 [1]),
    .Y(_3557_)
);

NAND2X1 _12407_ (
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [21]),
    .Y(_3337_)
);

FILL FILL_5__8999_ (
);

FILL FILL_5__8579_ (
);

FILL FILL_1__14910_ (
);

FILL FILL_6__11876_ (
);

FILL FILL_6__11456_ (
);

OAI22X1 _15299_ (
    .A(_5466__bF$buf0),
    .B(_4252_),
    .C(_4249_),
    .D(_5483__bF$buf3),
    .Y(_5773_)
);

FILL FILL_4__12490_ (
);

FILL FILL_4__12070_ (
);

FILL FILL_0__13903_ (
);

FILL FILL_3__16348_ (
);

FILL FILL_5__9940_ (
);

FILL FILL_5__10449_ (
);

FILL FILL_5__10029_ (
);

FILL FILL_5__9520_ (
);

FILL FILL_3__11483_ (
);

FILL FILL_5__9100_ (
);

FILL FILL_3__11063_ (
);

FILL FILL_4__6996_ (
);

FILL FILL_0__16375_ (
);

OAI22X1 _16240_ (
    .A(_5485__bF$buf3),
    .B(_6690_),
    .C(_5483__bF$buf4),
    .D(_5322_),
    .Y(_6691_)
);

FILL FILL_2__10896_ (
);

FILL SFILL38920x59050 (
);

FILL FILL_2__10056_ (
);

FILL FILL_0__11090_ (
);

FILL FILL_1__9932_ (
);

FILL FILL_5__11810_ (
);

FILL FILL_1__9512_ (
);

FILL FILL_3__9858_ (
);

FILL FILL_3__9018_ (
);

FILL FILL_4__10803_ (
);

FILL SFILL3640x51050 (
);

FILL FILL_0__6896_ (
);

FILL FILL_5__14282_ (
);

NAND2X1 _8582_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_858_)
);

DFFSR _8162_ (
    .Q(\datapath_1.regfile_1.regOut[10] [12]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_588_[12])
);

FILL FILL_1__10830_ (
);

FILL FILL_4__13695_ (
);

FILL FILL_4__13275_ (
);

FILL FILL_1__10410_ (
);

FILL FILL_2__7855_ (
);

FILL FILL_2__7435_ (
);

FILL FILL_3__12268_ (
);

FILL FILL_6__13602_ (
);

FILL SFILL3560x58050 (
);

NAND2X1 _12580_ (
    .A(vdd),
    .B(memoryOutData[4]),
    .Y(_3433_)
);

FILL FILL_0__12295_ (
);

INVX1 _12160_ (
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_3160_)
);

FILL SFILL104440x75050 (
);

FILL FILL_4__8722_ (
);

FILL FILL_2__12622_ (
);

FILL FILL_5__15487_ (
);

FILL FILL_2__12202_ (
);

FILL FILL_5__15067_ (
);

INVX1 _9787_ (
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_1478_)
);

INVX1 _9367_ (
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_1259_)
);

FILL SFILL7880x66050 (
);

FILL FILL_1__11615_ (
);

FILL FILL_2__15094_ (
);

FILL FILL_0__8622_ (
);

FILL FILL_0__8202_ (
);

FILL FILL_1__14087_ (
);

FILL FILL_4__15841_ (
);

FILL FILL_4__15421_ (
);

FILL FILL_4__15001_ (
);

OAI22X1 _13785_ (
    .A(_4290_),
    .B(_3890_),
    .C(_3967__bF$buf3),
    .D(_4289_),
    .Y(_4291_)
);

FILL SFILL49080x72050 (
);

NOR2X1 _13365_ (
    .A(_3797_),
    .B(_3873_),
    .Y(\datapath_1.regfile_1.regEn [31])
);

FILL FILL_3__14834_ (
);

FILL FILL_3__14414_ (
);

FILL SFILL28920x57050 (
);

FILL SFILL3560x13050 (
);

FILL FILL_4__9927_ (
);

FILL FILL_4__9507_ (
);

FILL FILL_2__13827_ (
);

FILL SFILL104440x30050 (
);

FILL FILL_0__14861_ (
);

FILL FILL_2__13407_ (
);

FILL FILL_0__14441_ (
);

FILL FILL_0__14021_ (
);

FILL FILL_2__16299_ (
);

CLKBUF1 CLKBUF1_insert130 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf94)
);

FILL SFILL28520x43050 (
);

CLKBUF1 CLKBUF1_insert131 (
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf93)
);

CLKBUF1 CLKBUF1_insert132 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf92)
);

CLKBUF1 CLKBUF1_insert133 (
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf91)
);

FILL FILL_0__9407_ (
);

CLKBUF1 CLKBUF1_insert134 (
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf90)
);

FILL FILL_3__7504_ (
);

CLKBUF1 CLKBUF1_insert135 (
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf89)
);

CLKBUF1 CLKBUF1_insert136 (
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf88)
);

CLKBUF1 CLKBUF1_insert137 (
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf87)
);

CLKBUF1 CLKBUF1_insert138 (
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf86)
);

CLKBUF1 CLKBUF1_insert139 (
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf85)
);

FILL FILL_4__16206_ (
);

FILL FILL_4__11761_ (
);

FILL FILL_4__11341_ (
);

FILL FILL_3__15619_ (
);

FILL FILL_1__16233_ (
);

FILL SFILL14200x78050 (
);

FILL FILL_3__10754_ (
);

FILL FILL_0__15646_ (
);

INVX1 _15931_ (
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_6389_)
);

FILL FILL_0__15226_ (
);

NOR2X1 _15511_ (
    .A(_5979_),
    .B(_5973_),
    .Y(_5980_)
);

FILL FILL_2__8393_ (
);

FILL FILL_0__10781_ (
);

FILL FILL_0__10361_ (
);

FILL FILL_6__14140_ (
);

FILL FILL_3__8709_ (
);

FILL FILL_5__13973_ (
);

FILL FILL_5__13553_ (
);

FILL FILL_5__13133_ (
);

NAND2X1 _7853_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_494_)
);

NAND2X1 _7433_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_275_)
);

DFFSR _7013_ (
    .Q(\datapath_1.regfile_1.regOut[1] [15]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_3_[15])
);

FILL FILL_4_BUFX2_insert810 (
);

FILL FILL_4_BUFX2_insert811 (
);

FILL FILL_4__9680_ (
);

FILL SFILL28840x19050 (
);

FILL FILL_4__9260_ (
);

FILL FILL_4__12966_ (
);

FILL FILL_4_BUFX2_insert812 (
);

FILL FILL_4_BUFX2_insert813 (
);

FILL FILL_4_BUFX2_insert814 (
);

FILL FILL_4__12126_ (
);

FILL FILL_2__13580_ (
);

FILL FILL_2__13160_ (
);

FILL FILL_4_BUFX2_insert815 (
);

FILL FILL_4_BUFX2_insert816 (
);

FILL FILL_4_BUFX2_insert817 (
);

FILL FILL_4_BUFX2_insert818 (
);

FILL FILL_3__11959_ (
);

FILL FILL_4_BUFX2_insert819 (
);

FILL FILL_1__12993_ (
);

FILL FILL_3__11539_ (
);

FILL FILL_1__12573_ (
);

FILL FILL_3__11119_ (
);

FILL FILL_1__12153_ (
);

FILL FILL_0__11986_ (
);

FILL FILL_2__9598_ (
);

FILL SFILL79160x66050 (
);

NAND2X1 _11851_ (
    .A(_2919_),
    .B(_2937_),
    .Y(_2938_)
);

FILL FILL_0__11566_ (
);

FILL FILL_0__9160_ (
);

AOI21X1 _11431_ (
    .A(_2546_),
    .B(_2545_),
    .C(_2383_),
    .Y(_2547_)
);

FILL FILL_0__11146_ (
);

OR2X2 _11011_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2130_)
);

FILL FILL_3__12900_ (
);

FILL FILL_5__7183_ (
);

FILL FILL_5__14758_ (
);

FILL FILL_5__14338_ (
);

FILL FILL_3__15792_ (
);

FILL FILL_3__15372_ (
);

INVX1 _8638_ (
    .A(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_895_)
);

INVX1 _8218_ (
    .A(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_676_)
);

FILL FILL_1__7595_ (
);

FILL FILL_1__7175_ (
);

FILL FILL_2__14785_ (
);

FILL FILL_2__14365_ (
);

FILL SFILL94360x41050 (
);

FILL FILL_1__13778_ (
);

FILL FILL_1__13358_ (
);

FILL FILL_3__8882_ (
);

FILL FILL_3__8462_ (
);

INVX1 _12636_ (
    .A(\datapath_1.Data [23]),
    .Y(_3470_)
);

AND2X2 _12216_ (
    .A(ALUSrcB_0_bF$buf2),
    .B(ALUSrcB_1_bF$buf2),
    .Y(_3201_)
);

FILL FILL_5__8388_ (
);

FILL SFILL79160x21050 (
);

FILL FILL_0__13712_ (
);

FILL FILL_3__16157_ (
);

FILL FILL_5__10678_ (
);

FILL FILL_5__10258_ (
);

FILL FILL_3__11292_ (
);

FILL FILL_0__16184_ (
);

FILL SFILL18840x17050 (
);

FILL FILL_2__10285_ (
);

FILL FILL_1__9741_ (
);

FILL FILL_3_BUFX2_insert830 (
);

FILL FILL_3__9667_ (
);

FILL FILL_3_BUFX2_insert831 (
);

FILL FILL_3__9247_ (
);

FILL FILL_3_BUFX2_insert832 (
);

FILL FILL_3_BUFX2_insert833 (
);

FILL FILL_3_BUFX2_insert834 (
);

FILL FILL_5__14091_ (
);

FILL FILL_3_BUFX2_insert835 (
);

FILL FILL_1__15924_ (
);

FILL FILL_3_BUFX2_insert836 (
);

FILL FILL_1__15504_ (
);

INVX1 _8391_ (
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_771_)
);

FILL FILL_3_BUFX2_insert837 (
);

FILL FILL_3_BUFX2_insert838 (
);

FILL FILL_3_BUFX2_insert839 (
);

FILL FILL_4__13084_ (
);

FILL SFILL99800x7050 (
);

FILL FILL_0__14917_ (
);

FILL FILL_2__7244_ (
);

FILL FILL_3__12497_ (
);

FILL FILL_3__12077_ (
);

FILL SFILL48600x35050 (
);

FILL FILL_5__12824_ (
);

FILL SFILL99400x6050 (
);

FILL FILL_5__12404_ (
);

FILL FILL_4__8951_ (
);

FILL FILL_4__8531_ (
);

FILL FILL_4__8111_ (
);

FILL FILL_4__11817_ (
);

FILL SFILL79160x50 (
);

FILL FILL_2__12851_ (
);

FILL FILL_2__12431_ (
);

FILL FILL_5__15296_ (
);

FILL FILL_2__12011_ (
);

INVX1 _9596_ (
    .A(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_1371_)
);

DFFSR _9176_ (
    .Q(\datapath_1.regfile_1.regOut[18] [2]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf57),
    .S(vdd),
    .D(_1108_[2])
);

FILL FILL_1__11844_ (
);

FILL FILL_4__14289_ (
);

FILL FILL_1__11424_ (
);

FILL FILL_1__11004_ (
);

FILL FILL_2__8869_ (
);

FILL FILL_0__8851_ (
);

FILL FILL_2__8449_ (
);

FILL FILL_0__10837_ (
);

NAND2X1 _10702_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1946_)
);

FILL FILL_0__8011_ (
);

FILL FILL_0__10417_ (
);

FILL FILL_5__6874_ (
);

FILL FILL_0_BUFX2_insert960 (
);

FILL FILL_4__15650_ (
);

FILL FILL_0_BUFX2_insert961 (
);

FILL FILL_0_BUFX2_insert962 (
);

FILL FILL_4__15230_ (
);

FILL FILL_0_BUFX2_insert963 (
);

FILL FILL_0_BUFX2_insert964 (
);

FILL FILL_0_BUFX2_insert965 (
);

AOI22X1 _13594_ (
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .B(_4102_),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_4103_)
);

FILL FILL_0_BUFX2_insert966 (
);

OAI21X1 _13174_ (
    .A(_3746_),
    .B(PCEn_bF$buf0),
    .C(_3747_),
    .Y(_3685_[31])
);

FILL FILL_5__13609_ (
);

FILL FILL_0_BUFX2_insert967 (
);

FILL FILL_2__9810_ (
);

FILL FILL_0_BUFX2_insert968 (
);

FILL FILL_3__14643_ (
);

FILL FILL_0_BUFX2_insert969 (
);

DFFSR _7909_ (
    .Q(\datapath_1.regfile_1.regOut[8] [15]),
    .CLK(clk_bF$buf44),
    .R(rst_bF$buf12),
    .S(vdd),
    .D(_458_[15])
);

FILL FILL_3__14223_ (
);

FILL FILL_1__6866_ (
);

FILL FILL_4__9736_ (
);

FILL FILL_2__13636_ (
);

FILL FILL_2__13216_ (
);

FILL FILL_0__14670_ (
);

FILL FILL_0__14250_ (
);

FILL SFILL110200x12050 (
);

FILL FILL_1__12629_ (
);

FILL FILL_1__12209_ (
);

FILL FILL_3__7733_ (
);

FILL FILL_0__9636_ (
);

FILL FILL_0__9216_ (
);

OAI21X1 _11907_ (
    .A(_2978_),
    .B(IorD_bF$buf0),
    .C(_2979_),
    .Y(_1_[6])
);

FILL FILL_3__7313_ (
);

FILL FILL_5__7239_ (
);

FILL SFILL114520x20050 (
);

FILL FILL_4__16015_ (
);

FILL FILL_6__10956_ (
);

FILL FILL_4__11990_ (
);

OAI22X1 _14799_ (
    .A(_3935__bF$buf4),
    .B(_5282_),
    .C(_5281_),
    .D(_3944__bF$buf2),
    .Y(_5283_)
);

NAND3X1 _14379_ (
    .A(_4868_),
    .B(_4871_),
    .C(_4867_),
    .Y(_4872_)
);

FILL FILL_4__11570_ (
);

FILL FILL_4__11150_ (
);

FILL FILL_3__15848_ (
);

FILL FILL_3__15428_ (
);

FILL FILL_3__15008_ (
);

FILL FILL_1__16042_ (
);

FILL FILL_3__10983_ (
);

FILL FILL_5__8600_ (
);

FILL FILL_3__10563_ (
);

FILL FILL_6_BUFX2_insert341 (
);

FILL FILL_3__10143_ (
);

FILL SFILL59080x69050 (
);

FILL FILL_0__15875_ (
);

NAND3X1 _15740_ (
    .A(_6202_),
    .B(_6201_),
    .C(_6200_),
    .Y(_6203_)
);

FILL FILL_0__15455_ (
);

INVX1 _15320_ (
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_5794_)
);

FILL FILL_0__15035_ (
);

FILL FILL_6_BUFX2_insert347 (
);

FILL FILL_0__10170_ (
);

FILL FILL_3__8518_ (
);

FILL SFILL3640x46050 (
);

FILL FILL_5__13782_ (
);

FILL FILL_5__13362_ (
);

DFFSR _7662_ (
    .Q(\datapath_1.regfile_1.regOut[6] [24]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf68),
    .S(vdd),
    .D(_328_[24])
);

INVX1 _7242_ (
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_188_)
);

FILL SFILL104520x63050 (
);

FILL SFILL43880x53050 (
);

FILL FILL_4__12775_ (
);

FILL FILL_4__12355_ (
);

INVX1 _10299_ (
    .A(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_1738_)
);

FILL FILL_2__6935_ (
);

FILL FILL_5__9805_ (
);

FILL FILL_3__11768_ (
);

FILL FILL_3__11348_ (
);

FILL SFILL59000x67050 (
);

FILL FILL_1__12382_ (
);

AOI21X1 _16105_ (
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .B(_5567_),
    .C(_6558_),
    .Y(_6559_)
);

FILL SFILL59080x24050 (
);

FILL FILL_0__11795_ (
);

FILL FILL_0__11375_ (
);

NAND3X1 _11660_ (
    .A(_2470__bF$buf0),
    .B(_2762_),
    .C(_2761_),
    .Y(_2763_)
);

OAI21X1 _11240_ (
    .A(_2357_),
    .B(_2358_),
    .C(_2129_),
    .Y(_2359_)
);

FILL FILL_4__7802_ (
);

FILL FILL_5__14987_ (
);

FILL FILL_5__14567_ (
);

FILL FILL_2__11702_ (
);

FILL FILL_5__14147_ (
);

FILL FILL_3__15181_ (
);

INVX1 _8867_ (
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_1007_)
);

INVX1 _8447_ (
    .A(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_788_)
);

DFFSR _8027_ (
    .Q(\datapath_1.regfile_1.regOut[9] [5]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_523_[5])
);

FILL FILL_2__14594_ (
);

FILL FILL_2__14174_ (
);

FILL FILL_0__7702_ (
);

FILL FILL_1__13587_ (
);

FILL FILL_1__13167_ (
);

FILL FILL_4__14921_ (
);

FILL FILL_4__14501_ (
);

FILL SFILL59000x22050 (
);

FILL SFILL49080x67050 (
);

FILL FILL_3__8271_ (
);

INVX1 _12865_ (
    .A(\datapath_1.a [14]),
    .Y(_3582_)
);

INVX1 _12445_ (
    .A(ALUOut[2]),
    .Y(_3363_)
);

AOI22X1 _12025_ (
    .A(\datapath_1.ALUResult [9]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3065_)
);

FILL FILL_3__13914_ (
);

FILL FILL_5__8197_ (
);

FILL SFILL73560x78050 (
);

FILL FILL_5_BUFX2_insert360 (
);

FILL FILL_2__12907_ (
);

FILL FILL_5_BUFX2_insert361 (
);

FILL FILL_0__13941_ (
);

FILL FILL_5_BUFX2_insert362 (
);

FILL FILL_3__16386_ (
);

FILL FILL_0__13521_ (
);

FILL FILL_5_BUFX2_insert363 (
);

FILL FILL_0__13101_ (
);

FILL FILL_5_BUFX2_insert364 (
);

FILL FILL_5_BUFX2_insert365 (
);

FILL FILL_5__10487_ (
);

FILL FILL_5_BUFX2_insert366 (
);

FILL FILL_5__10067_ (
);

FILL FILL_5_BUFX2_insert367 (
);

FILL FILL_1__8189_ (
);

FILL FILL_5_BUFX2_insert368 (
);

FILL FILL_5_BUFX2_insert369 (
);

FILL FILL_2__15799_ (
);

FILL FILL_2__15379_ (
);

FILL FILL_0__8907_ (
);

FILL FILL_1__9550_ (
);

FILL FILL_1__9130_ (
);

FILL FILL_4__15706_ (
);

FILL FILL_3__9896_ (
);

FILL FILL_2__16320_ (
);

FILL SFILL49000x65050 (
);

FILL FILL_3__9476_ (
);

FILL FILL_4__10421_ (
);

FILL FILL_4__10001_ (
);

FILL FILL_1__15733_ (
);

FILL SFILL49080x22050 (
);

FILL FILL_1__15313_ (
);

FILL FILL_0__14726_ (
);

FILL FILL_0__14306_ (
);

FILL FILL_2__7893_ (
);

FILL FILL_2__7473_ (
);

FILL FILL_2__7053_ (
);

FILL FILL_2__11299_ (
);

FILL FILL_5__12633_ (
);

FILL FILL_5__12213_ (
);

NAND2X1 _6933_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_23_)
);

FILL FILL_2_BUFX2_insert490 (
);

FILL FILL_2_BUFX2_insert491 (
);

FILL FILL_4__8760_ (
);

FILL FILL_2_BUFX2_insert492 (
);

FILL FILL_2_BUFX2_insert493 (
);

FILL FILL_4__8340_ (
);

FILL FILL_2_BUFX2_insert494 (
);

FILL FILL_4__11626_ (
);

FILL FILL_2__12660_ (
);

FILL FILL_2_BUFX2_insert495 (
);

FILL FILL_4__11206_ (
);

FILL FILL_2_BUFX2_insert496 (
);

FILL FILL_2__12240_ (
);

FILL FILL_0__7299_ (
);

FILL FILL_2_BUFX2_insert497 (
);

FILL FILL_2_BUFX2_insert498 (
);

FILL FILL_2_BUFX2_insert499 (
);

FILL FILL_3__10619_ (
);

FILL FILL_0_CLKBUF1_insert190 (
);

FILL FILL_1__11653_ (
);

FILL FILL_0_CLKBUF1_insert191 (
);

FILL FILL_1__11233_ (
);

FILL FILL_4__14098_ (
);

FILL FILL_0_CLKBUF1_insert192 (
);

FILL FILL_0_CLKBUF1_insert193 (
);

FILL FILL_0_CLKBUF1_insert194 (
);

FILL FILL_0_CLKBUF1_insert195 (
);

FILL FILL_0_CLKBUF1_insert196 (
);

FILL FILL_0__8660_ (
);

INVX1 _10931_ (
    .A(_2064_),
    .Y(_2065_)
);

FILL FILL_0__8240_ (
);

FILL FILL_0_CLKBUF1_insert197 (
);

FILL FILL_0__10646_ (
);

FILL FILL_2__8258_ (
);

NAND2X1 _10511_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1839_)
);

FILL FILL_0_CLKBUF1_insert198 (
);

FILL FILL_0_CLKBUF1_insert199 (
);

FILL FILL_5__13838_ (
);

FILL FILL_3__14872_ (
);

FILL FILL_5__13418_ (
);

FILL FILL_3__14452_ (
);

INVX1 _7718_ (
    .A(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_424_)
);

FILL FILL_3__14032_ (
);

FILL FILL_4__9545_ (
);

FILL FILL_4__9125_ (
);

FILL FILL_2__13865_ (
);

FILL FILL111800x65050 (
);

FILL FILL_2__13445_ (
);

FILL FILL_2__13025_ (
);

FILL SFILL39000x63050 (
);

FILL SFILL94360x36050 (
);

FILL FILL_1__12858_ (
);

FILL FILL_1__12438_ (
);

FILL FILL_1__12018_ (
);

FILL FILL_0_BUFX2_insert0 (
);

FILL FILL_0_BUFX2_insert1 (
);

FILL FILL_0_BUFX2_insert2 (
);

FILL FILL_0__9865_ (
);

FILL FILL_0_BUFX2_insert3 (
);

FILL FILL_3__7962_ (
);

FILL FILL_0_BUFX2_insert4 (
);

FILL FILL_3__7542_ (
);

FILL FILL_0_BUFX2_insert5 (
);

FILL FILL_3__7122_ (
);

FILL FILL_0__9025_ (
);

OAI21X1 _11716_ (
    .A(_2813_),
    .B(_2814_),
    .C(_2809_),
    .Y(_2815_)
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_5__7888_ (
);

FILL SFILL79160x16050 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_5__7468_ (
);

FILL FILL_4__16244_ (
);

FILL FILL_5__7048_ (
);

FILL FILL_6__10765_ (
);

INVX1 _14188_ (
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_4685_)
);

FILL FILL_3__15657_ (
);

FILL FILL_3__15237_ (
);

FILL FILL_1__16271_ (
);

FILL FILL_3__10792_ (
);

FILL FILL_3__10372_ (
);

FILL FILL_0__15684_ (
);

FILL FILL_0__15264_ (
);

FILL SFILL79240x1050 (
);

FILL FILL_1__8401_ (
);

FILL SFILL53880x2050 (
);

FILL FILL_3__8747_ (
);

FILL FILL_3__8327_ (
);

FILL FILL_5__13591_ (
);

FILL FILL_5__13171_ (
);

INVX1 _7891_ (
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_519_)
);

FILL SFILL53560x74050 (
);

INVX1 _7471_ (
    .A(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_300_)
);

INVX1 _7051_ (
    .A(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_81_)
);

FILL FILL_4__12584_ (
);

FILL FILL_4__12164_ (
);

FILL SFILL8760x53050 (
);

FILL FILL111720x27050 (
);

FILL FILL_3__11997_ (
);

FILL FILL_5__9614_ (
);

FILL FILL_3__11577_ (
);

FILL FILL_3__11157_ (
);

FILL FILL_1__12191_ (
);

NAND2X1 _16334_ (
    .A(gnd),
    .B(gnd),
    .Y(_6777_)
);

FILL FILL_0__16049_ (
);

FILL FILL_0__11184_ (
);

FILL FILL_5__11904_ (
);

FILL SFILL53960x43050 (
);

FILL FILL_1__9606_ (
);

FILL FILL_6__15383_ (
);

FILL FILL_4__7611_ (
);

FILL FILL_5__14796_ (
);

FILL FILL_2__11931_ (
);

FILL FILL_5__14376_ (
);

FILL FILL_2__11511_ (
);

DFFSR _8676_ (
    .Q(\datapath_1.regfile_1.regOut[14] [14]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_848_[14])
);

OAI21X1 _8256_ (
    .A(_700_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .C(_701_),
    .Y(_653_[24])
);

FILL FILL_1__10924_ (
);

FILL FILL_4__13789_ (
);

FILL FILL_4__13369_ (
);

FILL FILL_1__10504_ (
);

FILL FILL_2__7949_ (
);

FILL FILL_0__7931_ (
);

FILL FILL_2__7109_ (
);

FILL FILL_1__13396_ (
);

FILL FILL_4__14730_ (
);

FILL SFILL3720x79050 (
);

FILL FILL_4__14310_ (
);

FILL FILL_3__8080_ (
);

DFFSR _12674_ (
    .Q(\datapath_1.Data [11]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3425_[11])
);

FILL FILL_0__12389_ (
);

NAND3X1 _12254_ (
    .A(_3227_),
    .B(_3228_),
    .C(_3229_),
    .Y(\datapath_1.alu_1.ALUInB [9])
);

FILL FILL_3__13723_ (
);

FILL FILL_3__13303_ (
);

FILL FILL_2__12716_ (
);

FILL FILL_0__13750_ (
);

FILL FILL_0__13330_ (
);

FILL FILL_3__16195_ (
);

FILL FILL_5__10296_ (
);

FILL FILL_1__11709_ (
);

FILL FILL_2__15188_ (
);

FILL FILL_0__8716_ (
);

FILL FILL_5__16102_ (
);

FILL FILL_4__15935_ (
);

FILL FILL_4__15515_ (
);

OAI22X1 _13879_ (
    .A(_4382_),
    .B(_3916_),
    .C(_3881_),
    .D(_4381_),
    .Y(_4383_)
);

FILL FILL_3__9285_ (
);

NAND3X1 _13459_ (
    .A(_3898_),
    .B(_3919_),
    .C(_3879_),
    .Y(_3971_)
);

FILL FILL_4__10650_ (
);

NAND2X1 _13039_ (
    .A(vdd),
    .B(\datapath_1.rd2 [29]),
    .Y(_3678_)
);

FILL FILL_4__10230_ (
);

FILL SFILL3720x34050 (
);

FILL FILL_3__14928_ (
);

FILL FILL_3__14508_ (
);

FILL FILL_1__15962_ (
);

FILL FILL_1__15542_ (
);

FILL FILL_1__15122_ (
);

FILL SFILL43960x41050 (
);

FILL FILL_0__14955_ (
);

AOI22X1 _14820_ (
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [28]),
    .C(\datapath_1.regfile_1.regOut[6] [28]),
    .D(_4001__bF$buf2),
    .Y(_5304_)
);

FILL FILL_0__14535_ (
);

NAND3X1 _14400_ (
    .A(_4891_),
    .B(_4892_),
    .C(_4890_),
    .Y(_4893_)
);

FILL FILL_0__14115_ (
);

FILL FILL_5__12862_ (
);

FILL FILL_5__12442_ (
);

FILL FILL_5__12022_ (
);

FILL SFILL104520x58050 (
);

FILL SFILL48920x3050 (
);

FILL FILL_4__11855_ (
);

FILL FILL_4__11435_ (
);

FILL FILL_4__11015_ (
);

FILL FILL_6__8495_ (
);

FILL FILL_1__16327_ (
);

FILL FILL_3__10428_ (
);

FILL FILL_1__11882_ (
);

FILL FILL_3__10008_ (
);

FILL FILL_1__11462_ (
);

FILL FILL_1__11042_ (
);

INVX1 _15605_ (
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_6072_)
);

FILL SFILL59080x19050 (
);

FILL FILL112280x52050 (
);

FILL FILL_2__8487_ (
);

FILL FILL_0__10875_ (
);

FILL FILL_2__8067_ (
);

DFFSR _10740_ (
    .Q(\datapath_1.regfile_1.regOut[30] [30]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_1888_[30])
);

INVX1 _10320_ (
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_1752_)
);

FILL FILL_0__10035_ (
);

FILL FILL_5__13647_ (
);

FILL FILL_5__13227_ (
);

FILL FILL_3__14681_ (
);

INVX1 _7947_ (
    .A(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_536_)
);

FILL FILL_3__14261_ (
);

DFFSR _7527_ (
    .Q(\datapath_1.regfile_1.regOut[5] [17]),
    .CLK(clk_bF$buf95),
    .R(rst_bF$buf76),
    .S(vdd),
    .D(_263_[17])
);

OAI21X1 _7107_ (
    .A(_117_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .C(_118_),
    .Y(_68_[25])
);

FILL FILL_4__9774_ (
);

FILL FILL_4__9354_ (
);

FILL FILL_2__13674_ (
);

FILL FILL_2__13254_ (
);

FILL FILL_1__12247_ (
);

FILL SFILL59000x17050 (
);

FILL FILL_0__9674_ (
);

FILL FILL_3__7351_ (
);

FILL FILL_0__9254_ (
);

NAND2X1 _11945_ (
    .A(IorD_bF$buf6),
    .B(ALUOut[19]),
    .Y(_3005_)
);

OAI21X1 _11525_ (
    .A(_2635_),
    .B(_2524_),
    .C(_2237_),
    .Y(_2636_)
);

NOR2X1 _11105_ (
    .A(\datapath_1.alu_1.ALUInA [23]),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2224_)
);

FILL FILL_6__15859_ (
);

FILL FILL_5__7697_ (
);

FILL FILL_6__15439_ (
);

FILL FILL_4__16053_ (
);

FILL FILL_3__15886_ (
);

FILL FILL_0__12601_ (
);

FILL FILL_3__15466_ (
);

FILL FILL_3__15046_ (
);

FILL FILL_1__16080_ (
);

FILL FILL_1__7689_ (
);

FILL FILL_6_BUFX2_insert720 (
);

FILL FILL_3__10181_ (
);

FILL FILL_2__14879_ (
);

FILL FILL_2__14459_ (
);

FILL FILL_2__14039_ (
);

FILL FILL_0__15493_ (
);

FILL SFILL33880x46050 (
);

FILL FILL_0__15073_ (
);

FILL FILL_6_BUFX2_insert725 (
);

FILL FILL_1__8630_ (
);

FILL FILL_1__8210_ (
);

FILL FILL_2__15820_ (
);

FILL FILL_2__15400_ (
);

FILL FILL_3__8976_ (
);

FILL FILL_3__8136_ (
);

FILL FILL_6__6981_ (
);

FILL SFILL49080x17050 (
);

FILL FILL_1__14813_ (
);

DFFSR _7280_ (
    .Q(\datapath_1.regfile_1.regOut[3] [26]),
    .CLK(clk_bF$buf104),
    .R(rst_bF$buf11),
    .S(vdd),
    .D(_133_[26])
);

FILL FILL_6__11359_ (
);

FILL SFILL94440x69050 (
);

FILL FILL_4__12393_ (
);

FILL FILL_0__13806_ (
);

FILL FILL_2__6973_ (
);

FILL FILL_5__9423_ (
);

FILL FILL_3__11386_ (
);

FILL FILL_5__9003_ (
);

FILL FILL_4__6899_ (
);

FILL FILL_6__12300_ (
);

FILL FILL_0__16278_ (
);

OAI21X1 _16143_ (
    .A(_5524__bF$buf2),
    .B(_5228_),
    .C(_6595_),
    .Y(_6596_)
);

FILL FILL_2__10799_ (
);

FILL FILL_2__10379_ (
);

FILL FILL_5__11713_ (
);

FILL FILL_1__9415_ (
);

FILL FILL_4__7840_ (
);

FILL FILL_4__7420_ (
);

FILL FILL_4__10706_ (
);

FILL FILL_2__11740_ (
);

FILL FILL_5__14185_ (
);

FILL FILL_2__11320_ (
);

FILL SFILL49000x15050 (
);

OAI21X1 _8485_ (
    .A(_812_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .C(_813_),
    .Y(_783_[15])
);

OAI21X1 _8065_ (
    .A(_593_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .C(_594_),
    .Y(_588_[3])
);

FILL FILL_4__13598_ (
);

FILL FILL_1__10313_ (
);

FILL FILL_2__7758_ (
);

FILL FILL_0__7740_ (
);

FILL FILL_0__7320_ (
);

FILL FILL_2__7338_ (
);

FILL FILL_6__13925_ (
);

FILL SFILL18840x7050 (
);

FILL FILL_6__13505_ (
);

OAI21X1 _12483_ (
    .A(_3387_),
    .B(vdd),
    .C(_3388_),
    .Y(_3360_[14])
);

FILL FILL_0__12198_ (
);

NAND3X1 _12063_ (
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[19]),
    .C(_3032__bF$buf2),
    .Y(_3093_)
);

FILL FILL_5__12918_ (
);

FILL FILL_3__13952_ (
);

FILL FILL_3__13532_ (
);

FILL FILL_3__13112_ (
);

FILL FILL_4__8625_ (
);

FILL FILL_4__8205_ (
);

FILL FILL_5_BUFX2_insert740 (
);

FILL FILL_5_BUFX2_insert741 (
);

FILL FILL_2__12525_ (
);

FILL FILL_5_BUFX2_insert742 (
);

FILL FILL_2__12105_ (
);

FILL FILL_5_BUFX2_insert743 (
);

FILL FILL_5_BUFX2_insert744 (
);

FILL FILL_5_BUFX2_insert745 (
);

FILL FILL_5_BUFX2_insert746 (
);

FILL FILL_5_BUFX2_insert747 (
);

FILL FILL_1__11938_ (
);

FILL FILL_5_BUFX2_insert748 (
);

FILL FILL_5_BUFX2_insert749 (
);

FILL FILL_1__11518_ (
);

FILL FILL_5__16331_ (
);

FILL FILL_0__8525_ (
);

FILL FILL_0__8105_ (
);

FILL FILL_5__6968_ (
);

FILL FILL_4__15744_ (
);

FILL FILL_4__15324_ (
);

INVX1 _13688_ (
    .A(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_4195_)
);

FILL FILL_3__9094_ (
);

OR2X2 _13268_ (
    .A(_3796_),
    .B(_3809_),
    .Y(_3810_)
);

FILL SFILL23800x42050 (
);

FILL FILL_2__9904_ (
);

FILL FILL_3__14737_ (
);

FILL FILL_3__14317_ (
);

FILL FILL_1__15771_ (
);

FILL FILL_1__15351_ (
);

FILL FILL_0__14764_ (
);

FILL FILL_0__14344_ (
);

FILL FILL_2__7091_ (
);

FILL FILL_3__7827_ (
);

FILL FILL_5__12251_ (
);

INVX1 _6971_ (
    .A(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_48_)
);

FILL FILL_2_BUFX2_insert870 (
);

FILL FILL_2_BUFX2_insert871 (
);

FILL FILL_4__16109_ (
);

FILL FILL_2_BUFX2_insert872 (
);

FILL FILL_2_BUFX2_insert873 (
);

FILL FILL_2_BUFX2_insert874 (
);

FILL FILL_4__11664_ (
);

FILL SFILL8760x48050 (
);

FILL FILL_2_BUFX2_insert875 (
);

FILL FILL_4__11244_ (
);

FILL FILL_2_BUFX2_insert876 (
);

FILL FILL_2_BUFX2_insert877 (
);

FILL FILL_2_BUFX2_insert878 (
);

FILL FILL_2_BUFX2_insert879 (
);

FILL FILL_1__16136_ (
);

FILL FILL_3__10657_ (
);

FILL FILL_3__10237_ (
);

FILL FILL_1__11691_ (
);

FILL SFILL44280x33050 (
);

FILL FILL_1__11271_ (
);

FILL FILL_0__15969_ (
);

FILL FILL_0__15549_ (
);

INVX1 _15834_ (
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_6295_)
);

AOI21X1 _15414_ (
    .A(_5885_),
    .B(_5861_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [8])
);

FILL FILL_0__15129_ (
);

FILL FILL_0__10684_ (
);

FILL SFILL114600x48050 (
);

FILL FILL_0__10264_ (
);

FILL SFILL84360x29050 (
);

FILL FILL_5__13876_ (
);

FILL FILL_5__13456_ (
);

FILL FILL_3__14490_ (
);

FILL FILL_5__13036_ (
);

OAI21X1 _7756_ (
    .A(_448_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .C(_449_),
    .Y(_393_[28])
);

FILL FILL_3__14070_ (
);

OAI21X1 _7336_ (
    .A(_229_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_230_),
    .Y(_198_[16])
);

FILL FILL_4__9163_ (
);

FILL FILL_4__12869_ (
);

FILL FILL_4__12449_ (
);

FILL FILL_4__12029_ (
);

FILL FILL_2__13483_ (
);

FILL SFILL13800x40050 (
);

FILL FILL_1__12896_ (
);

FILL FILL_1__12476_ (
);

FILL FILL_1__12056_ (
);

FILL FILL_4__13810_ (
);

FILL SFILL74040x51050 (
);

FILL FILL_0__9483_ (
);

FILL FILL_0__11889_ (
);

FILL FILL_3__7580_ (
);

FILL FILL_3__7160_ (
);

INVX1 _11754_ (
    .A(_2849_),
    .Y(\datapath_1.ALUResult [8])
);

FILL FILL_0__11469_ (
);

NOR2X1 _11334_ (
    .A(_2324_),
    .B(_2452_),
    .Y(_2453_)
);

FILL FILL_0__11049_ (
);

FILL FILL_5__7086_ (
);

FILL FILL_4__16282_ (
);

FILL FILL_6__10383_ (
);

FILL FILL_3__15695_ (
);

FILL FILL_0__12830_ (
);

FILL FILL_0__12410_ (
);

FILL FILL_3__15275_ (
);

FILL FILL_1__7498_ (
);

FILL FILL_1__7078_ (
);

FILL FILL_2__14688_ (
);

FILL FILL_2__14268_ (
);

FILL FILL_5__15602_ (
);

OAI21X1 _9902_ (
    .A(_1533_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .C(_1534_),
    .Y(_1498_[18])
);

FILL FILL_1_BUFX2_insert890 (
);

FILL FILL_1_BUFX2_insert891 (
);

FILL FILL_3__8785_ (
);

FILL FILL_1_BUFX2_insert892 (
);

FILL FILL_3__8365_ (
);

OAI21X1 _12959_ (
    .A(_3623_),
    .B(vdd),
    .C(_3624_),
    .Y(_3620_[2])
);

FILL FILL_1_BUFX2_insert893 (
);

DFFSR _12539_ (
    .Q(ALUOut[4]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[4])
);

FILL SFILL3720x29050 (
);

FILL FILL_1_BUFX2_insert894 (
);

NAND2X1 _12119_ (
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [1]),
    .Y(_3133_)
);

FILL FILL_1_BUFX2_insert895 (
);

FILL FILL_1_BUFX2_insert896 (
);

FILL FILL_1__14622_ (
);

FILL FILL_1_BUFX2_insert897 (
);

FILL FILL_1__14202_ (
);

FILL FILL_1_BUFX2_insert898 (
);

FILL FILL_1_BUFX2_insert899 (
);

FILL SFILL43960x36050 (
);

FILL FILL_0__13615_ (
);

INVX1 _13900_ (
    .A(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_4403_)
);

FILL FILL_5__9652_ (
);

FILL FILL_5__9232_ (
);

FILL FILL_3__11195_ (
);

FILL FILL_0__16087_ (
);

INVX1 _16372_ (
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_6802_)
);

FILL SFILL78680x35050 (
);

FILL FILL_2__10188_ (
);

FILL FILL_5__11942_ (
);

FILL FILL_1__9644_ (
);

FILL FILL_5__11522_ (
);

FILL FILL_1__9224_ (
);

FILL FILL_5__11102_ (
);

FILL FILL_2__16414_ (
);

FILL FILL_4__10935_ (
);

FILL FILL_4__10515_ (
);

FILL FILL_1__15827_ (
);

FILL FILL_6__7575_ (
);

FILL FILL_1__15407_ (
);

DFFSR _8294_ (
    .Q(\datapath_1.regfile_1.regOut[11] [16]),
    .CLK(clk_bF$buf64),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_653_[16])
);

FILL FILL_1__10962_ (
);

FILL FILL_1__10542_ (
);

FILL FILL_1__10122_ (
);

FILL FILL112280x47050 (
);

FILL FILL_2__7987_ (
);

FILL FILL_2__7567_ (
);

BUFX2 BUFX2_insert560 (
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf47)
);

BUFX2 BUFX2_insert561 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf46)
);

BUFX2 BUFX2_insert562 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf45)
);

BUFX2 BUFX2_insert563 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf44)
);

BUFX2 BUFX2_insert564 (
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf43)
);

BUFX2 BUFX2_insert565 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf42)
);

BUFX2 BUFX2_insert566 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf41)
);

BUFX2 BUFX2_insert567 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf40)
);

BUFX2 BUFX2_insert568 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf39)
);

BUFX2 BUFX2_insert569 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf38)
);

NAND3X1 _12292_ (
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3198__bF$buf1),
    .Y(_3258_)
);

FILL FILL_5__12727_ (
);

FILL FILL_3__13761_ (
);

FILL FILL_5__12307_ (
);

FILL FILL_3__13341_ (
);

FILL FILL_4__8854_ (
);

FILL FILL_4__8014_ (
);

FILL FILL_2__12754_ (
);

FILL FILL_5__15199_ (
);

FILL FILL_2__12334_ (
);

NAND2X1 _9499_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1327_)
);

NAND2X1 _9079_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .Y(_1172_)
);

FILL FILL_1__11747_ (
);

FILL FILL_1__11327_ (
);

FILL FILL_3__6851_ (
);

FILL FILL_5__16140_ (
);

FILL FILL_0__8754_ (
);

FILL FILL_0__8334_ (
);

FILL FILL_6__9721_ (
);

DFFSR _10605_ (
    .Q(\datapath_1.regfile_1.regOut[29] [23]),
    .CLK(clk_bF$buf38),
    .R(rst_bF$buf32),
    .S(vdd),
    .D(_1823_[23])
);

FILL FILL_6__9301_ (
);

FILL FILL_0_BUFX2_insert80 (
);

FILL FILL_0_BUFX2_insert81 (
);

FILL FILL_4__15973_ (
);

FILL FILL_0_BUFX2_insert82 (
);

FILL FILL_0_BUFX2_insert83 (
);

FILL FILL_4__15553_ (
);

FILL FILL_0_BUFX2_insert84 (
);

FILL FILL_4__15133_ (
);

FILL FILL_0_BUFX2_insert85 (
);

FILL FILL_0_BUFX2_insert86 (
);

FILL FILL_0_BUFX2_insert87 (
);

INVX1 _13497_ (
    .A(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_4008_)
);

FILL FILL_0_BUFX2_insert88 (
);

DFFSR _13077_ (
    .Q(_2_[30]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3620_[30])
);

FILL FILL_0_BUFX2_insert89 (
);

FILL FILL_3__14966_ (
);

FILL FILL_3__14546_ (
);

FILL FILL_3__14126_ (
);

FILL FILL_1__15580_ (
);

FILL FILL_1__15160_ (
);

FILL FILL_4__9639_ (
);

FILL FILL_4__9219_ (
);

FILL FILL_2__13959_ (
);

FILL SFILL94520x57050 (
);

FILL FILL_0__14993_ (
);

FILL FILL_2__13539_ (
);

FILL FILL_0__14573_ (
);

FILL FILL_2__13119_ (
);

FILL FILL_0__14153_ (
);

FILL FILL_1__7710_ (
);

FILL FILL_2__14900_ (
);

FILL FILL_3__7636_ (
);

FILL FILL_0__9539_ (
);

FILL FILL_3__7216_ (
);

FILL FILL_0__9119_ (
);

FILL FILL_5__12480_ (
);

FILL FILL_5__12060_ (
);

FILL FILL_4__16338_ (
);

FILL FILL_4__11893_ (
);

FILL FILL_6__10439_ (
);

FILL FILL_4__11473_ (
);

FILL FILL_4__11053_ (
);

FILL FILL_1__16365_ (
);

FILL FILL_3__10886_ (
);

FILL FILL_5__8503_ (
);

FILL FILL_3__10046_ (
);

FILL FILL_1__11080_ (
);

FILL FILL_0__15778_ (
);

FILL FILL_0__15358_ (
);

INVX1 _15643_ (
    .A(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_6109_)
);

AOI22X1 _15223_ (
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_5699_)
);

FILL SFILL94520x12050 (
);

FILL FILL_0__10493_ (
);

FILL FILL_1__8915_ (
);

FILL FILL_6__14692_ (
);

FILL FILL_4__6920_ (
);

FILL FILL_5__13685_ (
);

FILL FILL_2__10820_ (
);

FILL FILL_5__13265_ (
);

FILL FILL_2__10400_ (
);

OAI21X1 _7985_ (
    .A(_560_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .C(_561_),
    .Y(_523_[19])
);

OAI21X1 _7565_ (
    .A(_341_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_342_),
    .Y(_328_[7])
);

DFFSR _7145_ (
    .Q(\datapath_1.regfile_1.regOut[2] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_68_[19])
);

FILL FILL_4__9392_ (
);

FILL FILL_4__12258_ (
);

FILL FILL_2__13292_ (
);

FILL SFILL94440x19050 (
);

FILL FILL_2__6838_ (
);

FILL FILL_1__12285_ (
);

DFFSR _16428_ (
    .Q(\datapath_1.regfile_1.regOut[0] [11]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf71),
    .S(vdd),
    .D(_6769_[11])
);

OAI22X1 _16008_ (
    .A(_5099_),
    .B(_5544__bF$buf2),
    .C(_5523_),
    .D(_5107_),
    .Y(_6464_)
);

INVX8 _11983_ (
    .A(PCSource_1_bF$buf0),
    .Y(_3032_)
);

FILL FILL_0__9292_ (
);

FILL FILL_0__11698_ (
);

NAND3X1 _11563_ (
    .A(_2231_),
    .B(_2668_),
    .C(_2671_),
    .Y(_2672_)
);

FILL FILL_0__11278_ (
);

NAND2X1 _11143_ (
    .A(_2226_),
    .B(_2237_),
    .Y(_2262_)
);

FILL FILL_3__12612_ (
);

FILL FILL_4__16091_ (
);

FILL FILL_4__7705_ (
);

FILL FILL_2__11605_ (
);

FILL FILL_3__15084_ (
);

FILL FILL_2__14497_ (
);

FILL FILL_2__14077_ (
);

FILL FILL_5__15831_ (
);

FILL FILL_5__15411_ (
);

FILL FILL_0__7605_ (
);

DFFSR _9711_ (
    .Q(\datapath_1.regfile_1.regOut[22] [25]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_1368_[25])
);

FILL FILL_4__14824_ (
);

FILL FILL_4__14404_ (
);

FILL FILL_3__8594_ (
);

NAND2X1 _12768_ (
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[24]),
    .Y(_3538_)
);

FILL SFILL23800x37050 (
);

OAI21X1 _12348_ (
    .A(_3296_),
    .B(MemToReg_bF$buf4),
    .C(_3297_),
    .Y(\datapath_1.mux_wd3.dout [1])
);

FILL FILL_3__13817_ (
);

FILL FILL_1__14851_ (
);

FILL FILL_1__14431_ (
);

FILL FILL_1__14011_ (
);

FILL FILL_0__13844_ (
);

FILL FILL_0__13424_ (
);

FILL FILL_3__16289_ (
);

FILL FILL_0__13004_ (
);

FILL FILL_5__9881_ (
);

FILL SFILL109720x53050 (
);

FILL FILL_5__9041_ (
);

OAI22X1 _16181_ (
    .A(_5310_),
    .B(_5501_),
    .C(_5524__bF$buf3),
    .D(_5292_),
    .Y(_6633_)
);

FILL FILL_3__6907_ (
);

FILL FILL_5__11751_ (
);

FILL FILL_1__9873_ (
);

FILL FILL_5__11331_ (
);

FILL FILL_1__9033_ (
);

FILL FILL_4__15609_ (
);

FILL FILL_2__16223_ (
);

FILL FILL_3__9799_ (
);

FILL FILL_3__9379_ (
);

FILL FILL_4__10744_ (
);

FILL FILL_4__10324_ (
);

FILL FILL_1__15636_ (
);

FILL FILL_1__15216_ (
);

FILL FILL_1__10771_ (
);

FILL FILL_0__14629_ (
);

INVX1 _14914_ (
    .A(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_5396_)
);

FILL FILL_0__14209_ (
);

FILL FILL_2__7376_ (
);

FILL FILL_5__12956_ (
);

FILL FILL_3__13990_ (
);

FILL FILL_5__12116_ (
);

FILL FILL_3__13570_ (
);

BUFX2 _6836_ (
    .A(gnd),
    .Y(MemRead)
);

FILL FILL_3__13150_ (
);

FILL FILL_4__11949_ (
);

FILL FILL_4__8243_ (
);

FILL FILL_2__12983_ (
);

FILL FILL_4__11529_ (
);

FILL FILL_4__11109_ (
);

FILL FILL_2__12143_ (
);

FILL FILL_6__8589_ (
);

FILL SFILL13800x35050 (
);

FILL FILL_1__11976_ (
);

FILL FILL_1__11556_ (
);

FILL FILL_1__11136_ (
);

FILL FILL_0__8983_ (
);

FILL FILL_0__10969_ (
);

FILL FILL_0__10549_ (
);

FILL FILL_0__8143_ (
);

OAI21X1 _10834_ (
    .A(_2012_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_2013_),
    .Y(_1953_[30])
);

OAI21X1 _10414_ (
    .A(_1793_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1794_),
    .Y(_1758_[18])
);

FILL FILL_0__10129_ (
);

FILL FILL_6__9110_ (
);

FILL FILL_6__14748_ (
);

FILL FILL_4__15782_ (
);

FILL FILL_4__15362_ (
);

FILL SFILL64120x82050 (
);

FILL FILL_0__11910_ (
);

FILL FILL_2__9522_ (
);

FILL FILL_3__14775_ (
);

FILL FILL_2__9102_ (
);

FILL FILL_3__14355_ (
);

FILL FILL_4__9868_ (
);

FILL FILL_4__9028_ (
);

FILL FILL_2__13768_ (
);

FILL FILL_2__13348_ (
);

FILL FILL_0__14382_ (
);

FILL FILL_0__9768_ (
);

FILL FILL_3__7865_ (
);

FILL FILL_0__9348_ (
);

FILL FILL_3__7445_ (
);

AOI21X1 _11619_ (
    .A(_2719_),
    .B(_2722_),
    .C(_2458_),
    .Y(_2724_)
);

FILL FILL_1__13702_ (
);

FILL FILL_4__16147_ (
);

FILL FILL_6__10248_ (
);

FILL FILL_4__11282_ (
);

FILL FILL_1__16174_ (
);

FILL FILL_5__8732_ (
);

FILL FILL_3__10695_ (
);

FILL FILL_3__10275_ (
);

FILL FILL_5__8312_ (
);

FILL FILL_2_BUFX2_insert0 (
);

FILL FILL_2_BUFX2_insert1 (
);

NAND3X1 _15872_ (
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf1),
    .Y(_6332_)
);

FILL FILL_0__15587_ (
);

FILL FILL_2_BUFX2_insert2 (
);

OAI22X1 _15452_ (
    .A(_5463__bF$buf2),
    .B(_5922_),
    .C(_5921_),
    .D(_5504__bF$buf2),
    .Y(_5923_)
);

FILL FILL_0__15167_ (
);

FILL SFILL104200x27050 (
);

NAND2X1 _15032_ (
    .A(_5459__bF$buf3),
    .B(_5511_),
    .Y(_5512_)
);

FILL FILL_2_BUFX2_insert3 (
);

FILL FILL112360x35050 (
);

FILL FILL_2_BUFX2_insert4 (
);

FILL FILL_2_BUFX2_insert5 (
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_1__8724_ (
);

FILL FILL_2_BUFX2_insert9 (
);

FILL FILL_2__15914_ (
);

FILL SFILL64040x44050 (
);

FILL FILL_5__13494_ (
);

DFFSR _7794_ (
    .Q(\datapath_1.regfile_1.regOut[7] [28]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_393_[28])
);

FILL FILL_1__14907_ (
);

NAND2X1 _7374_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_256_)
);

FILL FILL_4__12487_ (
);

FILL FILL_4__12067_ (
);

FILL SFILL54120x80050 (
);

FILL FILL_5__9937_ (
);

FILL FILL_5__9517_ (
);

FILL FILL_1__12094_ (
);

NAND3X1 _16237_ (
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf2),
    .Y(_6688_)
);

OAI21X1 _11792_ (
    .A(_2148_),
    .B(_2344__bF$buf3),
    .C(_2884_),
    .Y(_2885_)
);

INVX1 _11372_ (
    .A(_2127_),
    .Y(_2489_)
);

FILL FILL_0__11087_ (
);

FILL FILL_1__9929_ (
);

FILL FILL_5__11807_ (
);

FILL FILL_1__9509_ (
);

FILL FILL_3__12841_ (
);

FILL FILL_3__12421_ (
);

FILL FILL_6__15286_ (
);

FILL FILL_3__12001_ (
);

FILL FILL_4__7934_ (
);

FILL FILL_5__14699_ (
);

FILL FILL_2__11834_ (
);

FILL FILL_5__14279_ (
);

FILL FILL_2__11414_ (
);

NAND2X1 _8999_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1075_)
);

NAND2X1 _8579_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_856_)
);

DFFSR _8159_ (
    .Q(\datapath_1.regfile_1.regOut[10] [9]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_588_[9])
);

FILL FILL_1__10827_ (
);

FILL FILL_1__10407_ (
);

FILL FILL_5__15640_ (
);

FILL FILL_5__15220_ (
);

FILL FILL_0__7834_ (
);

FILL FILL_0__7414_ (
);

NAND2X1 _9940_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1560_)
);

NAND2X1 _9520_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1341_)
);

NAND2X1 _9100_ (
    .A(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1122_)
);

FILL FILL_1__13299_ (
);

FILL FILL_4__14633_ (
);

FILL FILL_4__14213_ (
);

NAND2X1 _12997_ (
    .A(vdd),
    .B(\datapath_1.rd2 [15]),
    .Y(_3650_)
);

NAND2X1 _12577_ (
    .A(vdd),
    .B(memoryOutData[3]),
    .Y(_3431_)
);

INVX1 _12157_ (
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_3158_)
);

FILL FILL_3__13626_ (
);

FILL FILL_1__14660_ (
);

FILL FILL_1__14240_ (
);

FILL FILL_4__8719_ (
);

FILL FILL_2__12619_ (
);

FILL FILL_0__13653_ (
);

FILL FILL_0__13233_ (
);

FILL FILL_3__16098_ (
);

FILL FILL_5__9270_ (
);

FILL FILL_5__16005_ (
);

FILL FILL_0__8619_ (
);

FILL FILL_5__11980_ (
);

FILL FILL_1__9682_ (
);

FILL FILL_5__11560_ (
);

FILL FILL_1__9262_ (
);

FILL FILL_5__11140_ (
);

FILL FILL_4__15838_ (
);

FILL FILL_4__15418_ (
);

FILL FILL_2__16032_ (
);

FILL FILL_4__10973_ (
);

FILL FILL_4__10553_ (
);

FILL FILL_4__10133_ (
);

FILL FILL_1__15865_ (
);

FILL FILL_6__7193_ (
);

FILL FILL_1__15445_ (
);

FILL FILL_1__15025_ (
);

FILL FILL_1__10580_ (
);

FILL FILL_1__10160_ (
);

FILL FILL_0__14858_ (
);

INVX1 _14723_ (
    .A(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_5209_)
);

FILL FILL_0__14438_ (
);

FILL FILL_0__14018_ (
);

INVX1 _14303_ (
    .A(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_4798_)
);

BUFX2 BUFX2_insert940 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf4 )
);

BUFX2 BUFX2_insert941 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf3 )
);

FILL FILL_2__7185_ (
);

BUFX2 BUFX2_insert942 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf2 )
);

BUFX2 BUFX2_insert943 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf1 )
);

BUFX2 BUFX2_insert944 (
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf0 )
);

FILL SFILL58280x57050 (
);

FILL FILL_6__13352_ (
);

BUFX2 BUFX2_insert945 (
    .A(_3036_),
    .Y(_3036__bF$buf4)
);

BUFX2 BUFX2_insert946 (
    .A(_3036_),
    .Y(_3036__bF$buf3)
);

BUFX2 BUFX2_insert947 (
    .A(_3036_),
    .Y(_3036__bF$buf2)
);

BUFX2 BUFX2_insert948 (
    .A(_3036_),
    .Y(_3036__bF$buf1)
);

BUFX2 BUFX2_insert949 (
    .A(_3036_),
    .Y(_3036__bF$buf0)
);

FILL FILL_5__12765_ (
);

FILL FILL_5__12345_ (
);

FILL FILL_4__8892_ (
);

FILL FILL_4__8472_ (
);

FILL FILL_4__11758_ (
);

FILL FILL_4__11338_ (
);

FILL FILL_2__12372_ (
);

FILL FILL_1__11785_ (
);

FILL FILL_1__11365_ (
);

NOR2X1 _15928_ (
    .A(_6376_),
    .B(_6386_),
    .Y(_6387_)
);

AOI22X1 _15508_ (
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [11]),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_5977_)
);

FILL SFILL8520x55050 (
);

FILL FILL_0__10778_ (
);

FILL FILL_0__8372_ (
);

FILL FILL_0__10358_ (
);

OAI21X1 _10643_ (
    .A(_1905_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .C(_1906_),
    .Y(_1888_[9])
);

DFFSR _10223_ (
    .Q(\datapath_1.regfile_1.regOut[26] [25]),
    .CLK(clk_bF$buf70),
    .R(rst_bF$buf90),
    .S(vdd),
    .D(_1628_[25])
);

FILL SFILL109400x72050 (
);

FILL FILL_4__15591_ (
);

FILL FILL_4__15171_ (
);

FILL SFILL44040x40050 (
);

FILL FILL_2__9751_ (
);

FILL FILL_3__14584_ (
);

FILL FILL_3__14164_ (
);

FILL FILL_4_BUFX2_insert780 (
);

FILL FILL_4__9677_ (
);

FILL FILL_4_BUFX2_insert781 (
);

FILL FILL_4_BUFX2_insert782 (
);

FILL FILL_4__9257_ (
);

FILL FILL_2__13997_ (
);

FILL FILL_4_BUFX2_insert783 (
);

FILL FILL_4_BUFX2_insert784 (
);

FILL FILL_2__13577_ (
);

FILL FILL_2__13157_ (
);

FILL FILL_4_BUFX2_insert785 (
);

FILL FILL_0__14191_ (
);

FILL FILL_4_BUFX2_insert786 (
);

FILL FILL112120x5050 (
);

FILL FILL_4_BUFX2_insert787 (
);

FILL FILL_5__14911_ (
);

FILL FILL_4_BUFX2_insert788 (
);

FILL FILL_4_BUFX2_insert789 (
);

FILL FILL_4__13904_ (
);

FILL FILL_0__9997_ (
);

FILL FILL_3__7674_ (
);

FILL FILL_0__9157_ (
);

AOI22X1 _11848_ (
    .A(_2481__bF$buf1),
    .B(_2542_),
    .C(_2341__bF$buf2),
    .D(_2935_),
    .Y(_2936_)
);

NOR3X1 _11428_ (
    .A(_2541_),
    .B(_2124_),
    .C(_2543_),
    .Y(_2544_)
);

NOR2X1 _11008_ (
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(_2126_),
    .Y(_2127_)
);

FILL FILL_1__13931_ (
);

FILL FILL_4__16376_ (
);

FILL FILL_1__13511_ (
);

FILL SFILL34040x83050 (
);

FILL FILL_6__10057_ (
);

FILL FILL_4__11091_ (
);

FILL FILL_3__15789_ (
);

FILL FILL_3__15369_ (
);

FILL FILL_0__12504_ (
);

FILL FILL_5__8961_ (
);

FILL SFILL74120x79050 (
);

FILL FILL_5__8121_ (
);

OAI22X1 _15681_ (
    .A(_4696_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf0),
    .D(_4695_),
    .Y(_6146_)
);

FILL FILL_0__15396_ (
);

AOI22X1 _15261_ (
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .B(_5567_),
    .C(_5565__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_5736_)
);

FILL FILL_3__16310_ (
);

FILL FILL_5__10831_ (
);

FILL FILL_1__8953_ (
);

FILL FILL_1__8533_ (
);

FILL FILL_5__10411_ (
);

FILL FILL_1__8113_ (
);

FILL FILL_2__15723_ (
);

FILL FILL_2__15303_ (
);

FILL FILL_3__8879_ (
);

FILL FILL_3__8459_ (
);

FILL FILL_1__14716_ (
);

NAND2X1 _7183_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_149_)
);

FILL FILL_4__12296_ (
);

FILL SFILL69160x51050 (
);

FILL FILL_3__9400_ (
);

FILL FILL_0__13709_ (
);

FILL FILL_2__6876_ (
);

FILL FILL_5__9746_ (
);

FILL FILL_3__11289_ (
);

FILL FILL_6__12203_ (
);

FILL SFILL74120x34050 (
);

AOI21X1 _16046_ (
    .A(_6477_),
    .B(_6501_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [24])
);

NOR2X1 _11181_ (
    .A(_2298_),
    .B(_2299_),
    .Y(_2300_)
);

FILL FILL_1__9738_ (
);

FILL FILL_5__11616_ (
);

FILL FILL_3__12650_ (
);

FILL FILL_3__12230_ (
);

FILL SFILL99320x83050 (
);

FILL FILL_4__7743_ (
);

FILL FILL_4__7323_ (
);

FILL FILL_2__11643_ (
);

FILL FILL_2__11223_ (
);

FILL FILL_5__14088_ (
);

INVX1 _8388_ (
    .A(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_769_)
);

FILL FILL_6__7249_ (
);

FILL FILL_1__10636_ (
);

FILL FILL_0__7223_ (
);

FILL FILL_4__14862_ (
);

FILL FILL_6__13408_ (
);

FILL FILL_4__14442_ (
);

FILL SFILL64120x77050 (
);

FILL FILL_4__14022_ (
);

FILL SFILL95000x30050 (
);

NAND2X1 _12386_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [14]),
    .Y(_3323_)
);

FILL FILL_3__13855_ (
);

FILL FILL_2__8602_ (
);

FILL FILL_3__13435_ (
);

FILL FILL_3__13015_ (
);

FILL FILL_4__8528_ (
);

FILL FILL_4__8108_ (
);

FILL FILL_2__12848_ (
);

FILL FILL_2__12428_ (
);

FILL FILL_0__13882_ (
);

FILL FILL_0__13462_ (
);

FILL FILL_2__12008_ (
);

FILL FILL_0__13042_ (
);

FILL SFILL74040x50 (
);

FILL FILL_0__8848_ (
);

FILL FILL_5__16234_ (
);

FILL FILL_3__6945_ (
);

FILL FILL_0__8008_ (
);

FILL FILL_1__9491_ (
);

FILL FILL_4__15647_ (
);

FILL FILL_4__15227_ (
);

FILL FILL_2__16261_ (
);

FILL FILL_4__10782_ (
);

FILL FILL_4__10362_ (
);

FILL FILL_2__9807_ (
);

FILL FILL_4_BUFX2_insert30 (
);

FILL SFILL64120x32050 (
);

FILL FILL_4_BUFX2_insert31 (
);

FILL FILL_1__15674_ (
);

FILL FILL_4_BUFX2_insert32 (
);

FILL FILL_1__15254_ (
);

FILL FILL_4_BUFX2_insert33 (
);

FILL FILL_4_BUFX2_insert34 (
);

FILL FILL_5__7812_ (
);

FILL FILL_4_BUFX2_insert35 (
);

FILL FILL_4_BUFX2_insert36 (
);

FILL FILL_4_BUFX2_insert37 (
);

FILL FILL_4_BUFX2_insert38 (
);

NOR2X1 _14952_ (
    .A(_5432_),
    .B(_5420_),
    .Y(_5433_)
);

FILL FILL_4_BUFX2_insert39 (
);

FILL FILL_0__14667_ (
);

FILL FILL_0__14247_ (
);

OAI22X1 _14532_ (
    .A(_5020_),
    .B(_3916_),
    .C(_3983__bF$buf4),
    .D(_5021_),
    .Y(_5022_)
);

FILL SFILL89320x81050 (
);

AOI21X1 _14112_ (
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .B(_4225_),
    .C(_4610_),
    .Y(_4611_)
);

FILL FILL_1__7804_ (
);

FILL FILL_6__13161_ (
);

FILL FILL_5__12994_ (
);

FILL FILL_5__12574_ (
);

FILL FILL_5__12154_ (
);

BUFX2 _6874_ (
    .A(_2_[4]),
    .Y(memoryWriteData[4])
);

FILL FILL_4__11987_ (
);

FILL FILL_4__11567_ (
);

FILL FILL_4__11147_ (
);

FILL FILL_2__12181_ (
);

FILL SFILL54120x75050 (
);

FILL FILL_1__16039_ (
);

FILL FILL_1__11594_ (
);

FILL FILL_1__11174_ (
);

NAND2X1 _15737_ (
    .A(\datapath_1.regfile_1.regOut[6] [17]),
    .B(_5565__bF$buf2),
    .Y(_6200_)
);

NOR2X1 _15317_ (
    .A(_5790_),
    .B(_5535__bF$buf2),
    .Y(_5791_)
);

INVX1 _10872_ (
    .A(\aluControl_1.inst [3]),
    .Y(_2020_)
);

FILL FILL_2__8199_ (
);

FILL FILL_0__10167_ (
);

NAND2X1 _10452_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1820_)
);

NAND2X1 _10032_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1601_)
);

BUFX2 BUFX2_insert90 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf3 )
);

FILL FILL_3__11921_ (
);

BUFX2 BUFX2_insert91 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf2 )
);

FILL FILL_3__11501_ (
);

BUFX2 BUFX2_insert92 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf1 )
);

BUFX2 BUFX2_insert93 (
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf0 )
);

BUFX2 BUFX2_insert94 (
    .A(_5548_),
    .Y(_5548__bF$buf4)
);

BUFX2 BUFX2_insert95 (
    .A(_5548_),
    .Y(_5548__bF$buf3)
);

BUFX2 BUFX2_insert96 (
    .A(_5548_),
    .Y(_5548__bF$buf2)
);

FILL FILL_2__10914_ (
);

FILL FILL_5__13779_ (
);

BUFX2 BUFX2_insert97 (
    .A(_5548_),
    .Y(_5548__bF$buf1)
);

FILL FILL_2__9980_ (
);

FILL FILL_5__13359_ (
);

BUFX2 BUFX2_insert98 (
    .A(_5548_),
    .Y(_5548__bF$buf0)
);

BUFX2 BUFX2_insert99 (
    .A(_5489_),
    .Y(_5489__bF$buf3)
);

FILL FILL_3__14393_ (
);

FILL FILL_2__9140_ (
);

DFFSR _7659_ (
    .Q(\datapath_1.regfile_1.regOut[6] [21]),
    .CLK(clk_bF$buf68),
    .R(rst_bF$buf49),
    .S(vdd),
    .D(_328_[21])
);

INVX1 _7239_ (
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_186_)
);

FILL FILL_4__9486_ (
);

FILL FILL_2__13386_ (
);

FILL FILL_5__14720_ (
);

FILL FILL_0__6914_ (
);

FILL FILL_5__14300_ (
);

FILL SFILL89240x43050 (
);

NAND2X1 _8600_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_870_)
);

FILL SFILL54120x30050 (
);

FILL FILL_1__12379_ (
);

FILL FILL_4__13713_ (
);

FILL FILL_3__7483_ (
);

FILL FILL_0__9386_ (
);

FILL FILL_3__7063_ (
);

NOR2X1 _11657_ (
    .A(_2178_),
    .B(_2759_),
    .Y(_2760_)
);

NOR2X1 _11237_ (
    .A(_2355_),
    .B(_2354_),
    .Y(_2356_)
);

FILL FILL_3__12706_ (
);

FILL FILL_1__13740_ (
);

FILL FILL_1__13320_ (
);

FILL FILL_4__16185_ (
);

FILL FILL_0__12733_ (
);

FILL FILL_3__15598_ (
);

FILL FILL_3__15178_ (
);

FILL FILL_0__12313_ (
);

FILL SFILL54040x37050 (
);

FILL FILL_5__8770_ (
);

FILL FILL_5__8350_ (
);

OAI22X1 _15490_ (
    .A(_5958_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf0),
    .D(_5959_),
    .Y(_5960_)
);

FILL FILL_5__15925_ (
);

OAI22X1 _15070_ (
    .A(_3929_),
    .B(_5548__bF$buf2),
    .C(_5549__bF$buf3),
    .D(_3969_),
    .Y(_5550_)
);

FILL FILL_5__15505_ (
);

INVX1 _9805_ (
    .A(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_1490_)
);

FILL FILL_5__10640_ (
);

FILL FILL_1__8762_ (
);

FILL FILL_1__8342_ (
);

FILL FILL_4__14918_ (
);

FILL FILL_2__15952_ (
);

FILL FILL_2__15532_ (
);

FILL FILL_2__15112_ (
);

FILL FILL_3__8268_ (
);

FILL FILL_1__14945_ (
);

FILL FILL_1__14525_ (
);

FILL FILL_1__14105_ (
);

FILL FILL_0__13938_ (
);

OAI22X1 _13803_ (
    .A(_3905__bF$buf2),
    .B(_4306_),
    .C(_3902__bF$buf0),
    .D(_4307_),
    .Y(_4308_)
);

FILL FILL_0__13518_ (
);

FILL FILL_5__9975_ (
);

FILL FILL_5__9555_ (
);

FILL FILL_5__9135_ (
);

FILL FILL_3__11098_ (
);

FILL FILL_6__12852_ (
);

INVX1 _16275_ (
    .A(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_6725_)
);

FILL FILL_5__11845_ (
);

FILL FILL_1__9547_ (
);

FILL FILL_5__11425_ (
);

FILL FILL_1__9127_ (
);

FILL FILL_5__11005_ (
);

FILL SFILL79240x41050 (
);

FILL FILL_4__7972_ (
);

FILL FILL_2__16317_ (
);

FILL FILL_4__7552_ (
);

FILL FILL_2__11872_ (
);

FILL FILL_4__10418_ (
);

FILL FILL_2__11452_ (
);

FILL FILL_2__11032_ (
);

INVX1 _8197_ (
    .A(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_662_)
);

FILL FILL_1__10445_ (
);

FILL FILL_1__10025_ (
);

FILL SFILL94680x7050 (
);

FILL FILL_0__7872_ (
);

FILL FILL_0__7452_ (
);

FILL FILL_0__7032_ (
);

FILL FILL_4__14671_ (
);

FILL SFILL44040x35050 (
);

FILL FILL_4__14251_ (
);

OAI21X1 _12195_ (
    .A(_3182_),
    .B(ALUSrcA_bF$buf5),
    .C(_3183_),
    .Y(\datapath_1.alu_1.ALUInA [26])
);

FILL SFILL54040x8050 (
);

FILL FILL_2__8831_ (
);

FILL FILL_3__13664_ (
);

FILL SFILL94280x6050 (
);

FILL FILL_3__13244_ (
);

FILL FILL_4__8757_ (
);

FILL FILL_4__8337_ (
);

FILL FILL_2__12657_ (
);

FILL FILL_2__12237_ (
);

FILL FILL_0__13691_ (
);

FILL FILL_0__13271_ (
);

FILL FILL_5__16043_ (
);

FILL FILL_0__8657_ (
);

OAI22X1 _10928_ (
    .A(_2054_),
    .B(\control_1.reg_state.dout [2]),
    .C(_2057_),
    .D(_2049_),
    .Y(ALUSrcB[1])
);

FILL FILL_0__8237_ (
);

NAND2X1 _10508_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1837_)
);

FILL FILL_4__15876_ (
);

FILL FILL_4__15456_ (
);

FILL FILL_4__15036_ (
);

FILL SFILL104440x9050 (
);

FILL FILL_2__16070_ (
);

FILL FILL_4__10171_ (
);

FILL FILL_2__9616_ (
);

FILL FILL_3__14869_ (
);

FILL FILL_3__14449_ (
);

FILL FILL_3__14029_ (
);

FILL FILL_1__15483_ (
);

FILL FILL_1__15063_ (
);

FILL FILL_5__7621_ (
);

FILL FILL_5__7201_ (
);

FILL SFILL104120x3050 (
);

FILL FILL_0__14896_ (
);

FILL FILL_0__14476_ (
);

NOR2X1 _14761_ (
    .A(_5242_),
    .B(_5245_),
    .Y(_5246_)
);

FILL FILL_0__14056_ (
);

INVX1 _14341_ (
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_4835_)
);

FILL FILL_3__15810_ (
);

FILL FILL_1__7613_ (
);

FILL FILL_2__14803_ (
);

FILL FILL_3__7959_ (
);

FILL FILL_3__7119_ (
);

FILL FILL_5__12383_ (
);

FILL SFILL99400x71050 (
);

FILL FILL_4__8090_ (
);

FILL FILL_4__11796_ (
);

FILL FILL_4__11376_ (
);

FILL SFILL69160x46050 (
);

FILL FILL_3__8900_ (
);

FILL FILL_1__16268_ (
);

FILL FILL_3__10789_ (
);

FILL FILL_5__8826_ (
);

FILL FILL_3__10369_ (
);

NAND2X1 _15966_ (
    .A(_6417_),
    .B(_6423_),
    .Y(_6424_)
);

AOI22X1 _15546_ (
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .B(_5577_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_6014_)
);

NOR3X1 _15126_ (
    .A(_5604_),
    .B(_5583_),
    .C(_5592_),
    .Y(_5605_)
);

FILL FILL_0__10396_ (
);

NAND2X1 _10681_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1932_)
);

NAND2X1 _10261_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1713_)
);

FILL FILL_6__14595_ (
);

FILL FILL_3__11730_ (
);

FILL FILL_6__14175_ (
);

FILL FILL_3__11310_ (
);

FILL SFILL99320x78050 (
);

FILL FILL_0__16202_ (
);

FILL FILL_5__13588_ (
);

FILL FILL_2__10303_ (
);

FILL FILL_5__13168_ (
);

INVX1 _7888_ (
    .A(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_517_)
);

INVX1 _7468_ (
    .A(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_298_)
);

INVX1 _7048_ (
    .A(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_79_)
);

FILL FILL_4__9295_ (
);

FILL FILL_1__12188_ (
);

FILL FILL_6__12908_ (
);

FILL FILL_4__13942_ (
);

FILL FILL_4__13522_ (
);

FILL FILL_4__13102_ (
);

OAI21X1 _11886_ (
    .A(_2966_),
    .B(RegDst),
    .C(_2967_),
    .Y(\datapath_1.a3 [4])
);

FILL FILL_3__7292_ (
);

NAND3X1 _11466_ (
    .A(_2462__bF$buf2),
    .B(_2576_),
    .C(_2580_),
    .Y(_2581_)
);

XOR2X1 _11046_ (
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2165_)
);

FILL FILL_3__12515_ (
);

FILL FILL_4__7608_ (
);

FILL FILL_2__11928_ (
);

FILL FILL_0__12962_ (
);

FILL FILL_2__11508_ (
);

FILL SFILL99320x33050 (
);

FILL FILL_0__12122_ (
);

FILL SFILL89320x7050 (
);

FILL SFILL23800x5050 (
);

FILL FILL_5__15734_ (
);

FILL FILL_5__15314_ (
);

FILL FILL_0__7928_ (
);

FILL SFILL28760x53050 (
);

FILL FILL_0__7508_ (
);

INVX1 _9614_ (
    .A(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_1383_)
);

FILL SFILL24040x31050 (
);

FILL FILL_1__8991_ (
);

FILL FILL_1__8571_ (
);

FILL FILL_4__14727_ (
);

FILL SFILL3720x1050 (
);

FILL FILL_4__14307_ (
);

FILL FILL_2__15761_ (
);

FILL FILL_2__15341_ (
);

FILL FILL_3__8497_ (
);

FILL FILL_3__8077_ (
);

FILL SFILL64120x27050 (
);

FILL SFILL3640x6050 (
);

FILL FILL_1__14754_ (
);

FILL FILL_1__14334_ (
);

FILL FILL_0__13747_ (
);

FILL SFILL89320x76050 (
);

INVX1 _13612_ (
    .A(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_4121_)
);

FILL FILL_0__13327_ (
);

FILL FILL_5__9784_ (
);

FILL FILL_5__9364_ (
);

FILL SFILL9400x42050 (
);

NOR2X1 _16084_ (
    .A(_6537_),
    .B(_6538_),
    .Y(_6539_)
);

FILL FILL_1__9776_ (
);

FILL FILL_5__11654_ (
);

FILL SFILL113880x38050 (
);

FILL FILL_1__9356_ (
);

FILL FILL_5__11234_ (
);

FILL FILL_2__16126_ (
);

FILL FILL_4__7361_ (
);

FILL FILL_4__10647_ (
);

FILL FILL_2__11681_ (
);

FILL FILL_2__11261_ (
);

FILL FILL_1__15959_ (
);

FILL FILL_1__15539_ (
);

FILL FILL_1__15119_ (
);

FILL FILL_2_BUFX2_insert110 (
);

FILL FILL_1__10674_ (
);

FILL FILL_1__10254_ (
);

INVX1 _14817_ (
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_5301_)
);

FILL SFILL33960x71050 (
);

FILL FILL_0__7681_ (
);

FILL FILL_2__7699_ (
);

FILL SFILL89320x31050 (
);

FILL FILL_4__14480_ (
);

FILL FILL_4__14060_ (
);

FILL FILL_5__12859_ (
);

FILL FILL_2__8640_ (
);

FILL FILL_5__12439_ (
);

FILL FILL_3__13893_ (
);

FILL FILL_5__12019_ (
);

FILL FILL_3__13473_ (
);

FILL FILL_2__8220_ (
);

FILL SFILL18760x51050 (
);

FILL SFILL49160x42050 (
);

FILL FILL_4__8986_ (
);

FILL FILL_4__8566_ (
);

FILL FILL_4__8146_ (
);

FILL FILL_2__12886_ (
);

FILL FILL_2__12466_ (
);

FILL FILL_2__12046_ (
);

FILL FILL_0__13080_ (
);

FILL FILL_5__13800_ (
);

FILL SFILL54120x25050 (
);

FILL FILL_1__11879_ (
);

FILL FILL_1__11459_ (
);

FILL FILL_1__11039_ (
);

FILL FILL_0__8886_ (
);

FILL FILL_5__16272_ (
);

FILL FILL_3__6983_ (
);

FILL FILL_0__8466_ (
);

DFFSR _10737_ (
    .Q(\datapath_1.regfile_1.regOut[30] [27]),
    .CLK(clk_bF$buf109),
    .R(rst_bF$buf67),
    .S(vdd),
    .D(_1888_[27])
);

INVX1 _10317_ (
    .A(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_1750_)
);

FILL SFILL79320x74050 (
);

FILL SFILL18680x58050 (
);

FILL FILL_4__15685_ (
);

FILL FILL_1__12400_ (
);

FILL FILL_4__15265_ (
);

FILL FILL_2__9425_ (
);

FILL FILL_0__11813_ (
);

FILL FILL_3__14678_ (
);

FILL FILL_3__14258_ (
);

FILL FILL_2__9005_ (
);

FILL FILL_1__15292_ (
);

FILL FILL_5__7850_ (
);

FILL SFILL114520x50 (
);

FILL FILL_5__7430_ (
);

INVX2 _14990_ (
    .A(\datapath_1.PCJump [25]),
    .Y(_5470_)
);

NOR2X1 _14570_ (
    .A(_5058_),
    .B(_5048_),
    .Y(_5059_)
);

FILL FILL_0__14285_ (
);

INVX1 _14150_ (
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_4648_)
);

FILL FILL_1__7842_ (
);

FILL FILL_1__7422_ (
);

FILL FILL_2__14612_ (
);

FILL FILL_3__7348_ (
);

FILL FILL_5__12192_ (
);

FILL SFILL39560x54050 (
);

FILL SFILL89800x50 (
);

FILL FILL_1__13605_ (
);

FILL SFILL33960x7050 (
);

FILL SFILL18680x13050 (
);

FILL FILL_4__11185_ (
);

FILL FILL_1__16077_ (
);

FILL FILL_5__8635_ (
);

FILL FILL_5__8215_ (
);

FILL FILL_3__10178_ (
);

FILL FILL111960x42050 (
);

FILL FILL_6__11932_ (
);

FILL FILL_6_BUFX2_insert694 (
);

OAI22X1 _15775_ (
    .A(_4810_),
    .B(_5539__bF$buf2),
    .C(_5552__bF$buf3),
    .D(_4828_),
    .Y(_6237_)
);

FILL FILL_6__11512_ (
);

NOR2X1 _15355_ (
    .A(_5827_),
    .B(_5821_),
    .Y(_5828_)
);

FILL SFILL99080x8050 (
);

FILL FILL_3__16404_ (
);

NAND2X1 _10490_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1825_)
);

FILL FILL_5__10925_ (
);

DFFSR _10070_ (
    .Q(\datapath_1.regfile_1.regOut[25] [0]),
    .CLK(clk_bF$buf62),
    .R(rst_bF$buf33),
    .S(vdd),
    .D(_1563_[0])
);

FILL FILL_5__10505_ (
);

FILL FILL_1__8627_ (
);

FILL FILL_1__8207_ (
);

FILL FILL_2__15817_ (
);

FILL FILL_0__16011_ (
);

FILL FILL_2__10952_ (
);

FILL FILL_2__10532_ (
);

FILL FILL_5__13397_ (
);

FILL FILL_2__10112_ (
);

INVX1 _7697_ (
    .A(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_410_)
);

DFFSR _7277_ (
    .Q(\datapath_1.regfile_1.regOut[3] [23]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf60),
    .S(vdd),
    .D(_133_[23])
);

FILL FILL111880x49050 (
);

FILL FILL_4_BUFX2_insert0 (
);

FILL FILL_4_BUFX2_insert1 (
);

FILL FILL_3__9914_ (
);

FILL SFILL109320x6050 (
);

FILL FILL_4_BUFX2_insert2 (
);

FILL FILL_4_BUFX2_insert3 (
);

FILL FILL_4_BUFX2_insert4 (
);

FILL FILL_0__6952_ (
);

FILL FILL_4_BUFX2_insert5 (
);

FILL FILL_4_BUFX2_insert6 (
);

FILL FILL_4_BUFX2_insert7 (
);

FILL FILL_4_BUFX2_insert8 (
);

FILL FILL_4_BUFX2_insert9 (
);

FILL FILL_6__12717_ (
);

FILL FILL_4__13751_ (
);

FILL FILL_4__13331_ (
);

AOI22X1 _11695_ (
    .A(_2184_),
    .B(_2481__bF$buf3),
    .C(_2478_),
    .D(_2165_),
    .Y(_2795_)
);

AOI21X1 _11275_ (
    .A(_2393_),
    .B(_2191_),
    .C(_2392_),
    .Y(_2394_)
);

FILL FILL_3__12744_ (
);

FILL SFILL108600x8050 (
);

FILL FILL_3__12324_ (
);

FILL FILL_4__7837_ (
);

FILL FILL_4__7417_ (
);

FILL FILL_2__11737_ (
);

FILL FILL_0__12771_ (
);

FILL FILL_2__11317_ (
);

FILL FILL_0__12351_ (
);

FILL FILL_6__16130_ (
);

FILL FILL_5__15963_ (
);

FILL FILL_5__15543_ (
);

FILL FILL_0__7737_ (
);

FILL FILL_5__15123_ (
);

DFFSR _9843_ (
    .Q(\datapath_1.regfile_1.regOut[23] [29]),
    .CLK(clk_bF$buf67),
    .R(rst_bF$buf75),
    .S(vdd),
    .D(_1433_[29])
);

FILL FILL_0__7317_ (
);

OAI21X1 _9423_ (
    .A(_1295_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .C(_1296_),
    .Y(_1238_[29])
);

OAI21X1 _9003_ (
    .A(_1076_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .C(_1077_),
    .Y(_1043_[17])
);

FILL FILL_1__8380_ (
);

FILL FILL_4__14956_ (
);

FILL FILL_2__15990_ (
);

FILL FILL_4__14536_ (
);

FILL FILL_2__15570_ (
);

FILL FILL_4__14116_ (
);

FILL SFILL109400x17050 (
);

FILL FILL_2__15150_ (
);

FILL FILL_3__13949_ (
);

FILL FILL_1__14983_ (
);

FILL FILL_3__13529_ (
);

FILL FILL_1__14563_ (
);

FILL FILL_3__13109_ (
);

FILL FILL_1__14143_ (
);

FILL FILL_0__13976_ (
);

FILL SFILL69240x34050 (
);

INVX1 _13841_ (
    .A(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_4345_)
);

FILL FILL_0__13556_ (
);

INVX1 _13421_ (
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_3933_)
);

FILL FILL_0__13136_ (
);

OAI21X1 _13001_ (
    .A(_3651_),
    .B(vdd),
    .C(_3652_),
    .Y(_3620_[16])
);

FILL FILL_5__9593_ (
);

FILL FILL_5__9173_ (
);

FILL SFILL93720x45050 (
);

FILL FILL_6__12050_ (
);

FILL FILL_5__16328_ (
);

FILL FILL_5__11883_ (
);

FILL FILL_5__11463_ (
);

FILL FILL_1__9165_ (
);

FILL FILL_5__11043_ (
);

FILL FILL_2__16355_ (
);

FILL SFILL99400x66050 (
);

FILL FILL_4__7590_ (
);

FILL FILL_4__7170_ (
);

FILL FILL_4__10876_ (
);

FILL FILL_2__11490_ (
);

FILL FILL_4__10036_ (
);

FILL FILL_2__11070_ (
);

FILL FILL_1__15768_ (
);

FILL FILL_1__15348_ (
);

FILL FILL_1__10063_ (
);

AOI22X1 _14626_ (
    .A(_3891__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [24]),
    .C(\datapath_1.regfile_1.regOut[8] [24]),
    .D(_4090_),
    .Y(_5114_)
);

INVX1 _14206_ (
    .A(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_4703_)
);

FILL FILL_0__7490_ (
);

FILL FILL_2__7088_ (
);

FILL FILL_0__7070_ (
);

FILL FILL_3__10810_ (
);

FILL FILL_6__13255_ (
);

FILL FILL_0__15702_ (
);

FILL SFILL69160x2050 (
);

FILL FILL_5__12248_ (
);

FILL FILL_3__13282_ (
);

INVX1 _6968_ (
    .A(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_46_)
);

FILL SFILL69080x7050 (
);

FILL FILL_4__8375_ (
);

FILL SFILL59640x46050 (
);

FILL FILL_2__12695_ (
);

FILL FILL_2__12275_ (
);

FILL SFILL99400x21050 (
);

FILL FILL_1__11688_ (
);

FILL FILL_1__11268_ (
);

FILL FILL_4__12602_ (
);

FILL FILL_0__8695_ (
);

FILL FILL_5__16081_ (
);

NOR2X1 _10966_ (
    .A(_2089_),
    .B(_2081_),
    .Y(_2097_)
);

FILL FILL_0__8275_ (
);

INVX1 _10546_ (
    .A(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_1862_)
);

INVX1 _10126_ (
    .A(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_1643_)
);

FILL FILL_4__15494_ (
);

FILL FILL_4__15074_ (
);

FILL SFILL99320x28050 (
);

FILL FILL_2__9654_ (
);

FILL FILL_3__14487_ (
);

FILL FILL_0__11622_ (
);

FILL FILL_2__9234_ (
);

FILL FILL_3__14067_ (
);

FILL FILL_0__11202_ (
);

FILL FILL_0__14094_ (
);

FILL SFILL89400x64050 (
);

FILL FILL_5__14814_ (
);

FILL SFILL59160x39050 (
);

FILL FILL_1__7231_ (
);

FILL FILL_4__13807_ (
);

FILL FILL_2__14841_ (
);

FILL FILL_3__7997_ (
);

FILL FILL_2__14421_ (
);

FILL FILL_2__14001_ (
);

FILL FILL_3__7577_ (
);

FILL FILL_1__13834_ (
);

FILL FILL_1__13414_ (
);

FILL FILL_4__16279_ (
);

FILL FILL_0__12827_ (
);

FILL FILL_0__12407_ (
);

FILL FILL_5__8864_ (
);

FILL FILL_5__8444_ (
);

FILL FILL_0__15299_ (
);

AOI22X1 _15584_ (
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .B(_5577_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_6051_)
);

NOR2X1 _15164_ (
    .A(_5640_),
    .B(_5641_),
    .Y(_5642_)
);

FILL FILL_3__16213_ (
);

FILL FILL_1__8856_ (
);

FILL FILL_5__10314_ (
);

FILL FILL_1__8016_ (
);

FILL SFILL94280x70050 (
);

FILL FILL_2__15626_ (
);

FILL FILL_2__15206_ (
);

FILL FILL_4__6861_ (
);

FILL FILL_0__16240_ (
);

FILL FILL_2__10761_ (
);

FILL FILL_1__14619_ (
);

OAI21X1 _7086_ (
    .A(_103_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_104_),
    .Y(_68_[18])
);

FILL FILL_4__12199_ (
);

FILL FILL_3__9723_ (
);

FILL FILL_5__9649_ (
);

FILL FILL_5__9229_ (
);

FILL FILL_4__13980_ (
);

INVX1 _16369_ (
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_6800_)
);

FILL FILL_6__12106_ (
);

FILL FILL_4__13560_ (
);

FILL FILL_4__13140_ (
);

FILL FILL_5__11939_ (
);

NOR2X1 _11084_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(_2202_),
    .Y(_2203_)
);

FILL FILL_2__7720_ (
);

FILL FILL_3__12973_ (
);

FILL FILL_5__11519_ (
);

FILL FILL_2__7300_ (
);

FILL SFILL18760x46050 (
);

FILL FILL_3__12133_ (
);

FILL FILL_4__7226_ (
);

FILL FILL_2__11966_ (
);

FILL FILL_2__11546_ (
);

FILL FILL_0__12580_ (
);

FILL FILL_2__11126_ (
);

FILL FILL_0__12160_ (
);

FILL FILL_1__10959_ (
);

FILL FILL_1__10539_ (
);

FILL FILL_1__10119_ (
);

FILL FILL_5__15772_ (
);

FILL FILL_5__15352_ (
);

FILL FILL_0__7966_ (
);

FILL SFILL38760x9050 (
);

FILL FILL_0__7546_ (
);

OAI21X1 _9652_ (
    .A(_1407_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .C(_1408_),
    .Y(_1368_[20])
);

FILL SFILL79320x69050 (
);

OAI21X1 _9232_ (
    .A(_1188_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .C(_1189_),
    .Y(_1173_[8])
);

FILL SFILL33960x21050 (
);

FILL FILL_1__11900_ (
);

FILL FILL_4__14765_ (
);

FILL FILL_4__14345_ (
);

AOI22X1 _12289_ (
    .A(_2_[18]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3256_)
);

FILL FILL_2__8505_ (
);

FILL FILL_3__13758_ (
);

FILL FILL_3__13338_ (
);

FILL FILL_1__14792_ (
);

FILL FILL_1__14372_ (
);

FILL FILL_5__6930_ (
);

FILL FILL_0__13785_ (
);

FILL FILL_0__13365_ (
);

INVX1 _13650_ (
    .A(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_4158_)
);

INVX2 _13230_ (
    .A(_3772_),
    .Y(_3773_)
);

FILL FILL_1__6922_ (
);

FILL FILL_3__6848_ (
);

FILL FILL_5__16137_ (
);

FILL FILL_5__11692_ (
);

FILL FILL_1__9394_ (
);

FILL FILL_5__11272_ (
);

FILL SFILL79320x24050 (
);

FILL FILL_2__16164_ (
);

FILL FILL_4__10685_ (
);

FILL FILL_4__10265_ (
);

FILL FILL_1__15997_ (
);

FILL FILL_1__15577_ (
);

FILL FILL_1__15157_ (
);

FILL FILL_5__7715_ (
);

FILL FILL111960x37050 (
);

FILL FILL_1__10292_ (
);

INVX1 _14855_ (
    .A(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_5338_)
);

INVX1 _14435_ (
    .A(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_4927_)
);

OAI22X1 _14015_ (
    .A(_4515_),
    .B(_3949_),
    .C(_3978_),
    .D(_4514_),
    .Y(_4516_)
);

FILL FILL_3__15904_ (
);

FILL FILL_1__7707_ (
);

FILL FILL_0__15931_ (
);

FILL FILL_0__15511_ (
);

FILL FILL_5__12897_ (
);

FILL FILL_5__12477_ (
);

FILL FILL_5__12057_ (
);

FILL FILL_3__13091_ (
);

FILL SFILL69320x67050 (
);

FILL FILL_4__8184_ (
);

FILL FILL_2__12084_ (
);

FILL FILL_1__11497_ (
);

FILL FILL_1__11077_ (
);

FILL FILL_4__12831_ (
);

FILL FILL_4__12411_ (
);

FILL FILL_6__9891_ (
);

INVX1 _10775_ (
    .A(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_1974_)
);

FILL FILL_0__8084_ (
);

DFFSR _10355_ (
    .Q(\datapath_1.regfile_1.regOut[27] [29]),
    .CLK(clk_bF$buf17),
    .R(rst_bF$buf13),
    .S(vdd),
    .D(_1693_[29])
);

FILL FILL_3__11824_ (
);

FILL FILL_3__11404_ (
);

FILL FILL_4__6917_ (
);

FILL FILL_2__9883_ (
);

FILL FILL_2__10817_ (
);

FILL FILL_2__9463_ (
);

FILL FILL_0__11851_ (
);

FILL FILL_3__14296_ (
);

FILL FILL_2__9043_ (
);

FILL FILL_0__11431_ (
);

FILL FILL_0__11011_ (
);

FILL FILL_4__9389_ (
);

FILL FILL_2__13289_ (
);

FILL FILL_5__14623_ (
);

FILL FILL_5__14203_ (
);

DFFSR _8923_ (
    .Q(\datapath_1.regfile_1.regOut[16] [5]),
    .CLK(clk_bF$buf3),
    .R(rst_bF$buf56),
    .S(vdd),
    .D(_978_[5])
);

OAI21X1 _8503_ (
    .A(_824_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_825_),
    .Y(_783_[21])
);

FILL FILL_1__7880_ (
);

FILL FILL_1__7460_ (
);

FILL FILL_1__7040_ (
);

FILL FILL_4__13616_ (
);

FILL FILL_2__14650_ (
);

FILL FILL_2__14230_ (
);

FILL FILL_0__9289_ (
);

FILL FILL_3__12609_ (
);

FILL FILL_1__13643_ (
);

FILL FILL_1__13223_ (
);

FILL FILL_4__16088_ (
);

FILL FILL_1_BUFX2_insert510 (
);

FILL FILL_1_BUFX2_insert511 (
);

FILL FILL_0__12636_ (
);

DFFSR _12921_ (
    .Q(\datapath_1.a [2]),
    .CLK(clk_bF$buf50),
    .R(rst_bF$buf47),
    .S(vdd),
    .D(_3555_[2])
);

FILL FILL_1_BUFX2_insert512 (
);

OAI21X1 _12501_ (
    .A(_3399_),
    .B(vdd),
    .C(_3400_),
    .Y(_3360_[20])
);

FILL FILL_0__12216_ (
);

FILL FILL_1_BUFX2_insert513 (
);

FILL FILL_1_BUFX2_insert514 (
);

FILL FILL_1_BUFX2_insert515 (
);

FILL SFILL114360x11050 (
);

FILL FILL_1_BUFX2_insert516 (
);

FILL FILL_5__8253_ (
);

FILL FILL_1_BUFX2_insert517 (
);

FILL FILL_1_BUFX2_insert518 (
);

FILL FILL_1_BUFX2_insert519 (
);

INVX1 _15393_ (
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_5865_)
);

FILL FILL_5__15828_ (
);

FILL FILL_5__15408_ (
);

FILL FILL_3__16022_ (
);

DFFSR _9708_ (
    .Q(\datapath_1.regfile_1.regOut[22] [22]),
    .CLK(clk_bF$buf97),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1368_[22])
);

FILL FILL_5__10963_ (
);

FILL FILL_5__10543_ (
);

FILL FILL_5__10123_ (
);

FILL FILL_1__8245_ (
);

FILL FILL_2__15855_ (
);

FILL FILL_2__15435_ (
);

FILL FILL_2__15015_ (
);

FILL FILL_2__10990_ (
);

FILL FILL_2__10570_ (
);

FILL FILL_2__10150_ (
);

FILL FILL_1__14848_ (
);

FILL FILL_1__14428_ (
);

FILL FILL_1__14008_ (
);

FILL FILL_3__9532_ (
);

FILL FILL_3__9112_ (
);

INVX1 _13706_ (
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_4213_)
);

FILL FILL_0__6990_ (
);

FILL FILL_5__9878_ (
);

FILL FILL_5__9038_ (
);

NAND3X1 _16178_ (
    .A(_6628_),
    .B(_6629_),
    .C(_6627_),
    .Y(_6630_)
);

FILL FILL_5__11748_ (
);

FILL FILL_3__12782_ (
);

FILL FILL_5__11328_ (
);

FILL FILL_3__12362_ (
);

FILL FILL_4__7875_ (
);

FILL FILL_4__7455_ (
);

FILL FILL_4__7035_ (
);

FILL FILL_2__11775_ (
);

FILL FILL_2__11355_ (
);

FILL SFILL99400x16050 (
);

FILL FILL_1__10768_ (
);

FILL FILL_5__15581_ (
);

FILL FILL_5__15161_ (
);

FILL FILL_0__7355_ (
);

OAI21X1 _9881_ (
    .A(_1519_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1520_),
    .Y(_1498_[11])
);

FILL FILL112440x60050 (
);

DFFSR _9461_ (
    .Q(\datapath_1.regfile_1.regOut[20] [31]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf50),
    .S(vdd),
    .D(_1238_[31])
);

NAND2X1 _9041_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1103_)
);

FILL FILL_4__14994_ (
);

FILL FILL_4__14574_ (
);

FILL FILL_4__14154_ (
);

NAND3X1 _12098_ (
    .A(_3117_),
    .B(_3118_),
    .C(_3119_),
    .Y(\datapath_1.mux_pcsrc.dout [27])
);

FILL FILL_3__13987_ (
);

FILL FILL_2__8734_ (
);

FILL FILL_0__10702_ (
);

FILL FILL_3__13567_ (
);

FILL FILL_2__8314_ (
);

FILL FILL_3__13147_ (
);

FILL FILL_1__14181_ (
);

FILL FILL_0__13594_ (
);

FILL SFILL89400x59050 (
);

FILL FILL_0__13174_ (
);

FILL FILL_4__9601_ (
);

FILL FILL_2__13921_ (
);

FILL FILL_5__16366_ (
);

FILL FILL_2__13501_ (
);

FILL FILL_5__11081_ (
);

FILL FILL_4__15779_ (
);

FILL FILL_1__12914_ (
);

FILL FILL_4__15359_ (
);

FILL FILL_2__16393_ (
);

FILL FILL_4__10494_ (
);

FILL FILL_2__9939_ (
);

FILL FILL_0__9921_ (
);

FILL FILL_0__11907_ (
);

FILL FILL_2__9519_ (
);

FILL FILL_0__9501_ (
);

FILL FILL_1__15386_ (
);

FILL FILL_5__7944_ (
);

FILL FILL_5__7104_ (
);

FILL FILL_4__16300_ (
);

FILL FILL_0__14799_ (
);

FILL FILL_0__14379_ (
);

INVX1 _14664_ (
    .A(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_5151_)
);

INVX1 _14244_ (
    .A(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_4740_)
);

FILL FILL_3__15713_ (
);

FILL SFILL89400x14050 (
);

FILL FILL_1__7936_ (
);

FILL FILL_2__14706_ (
);

FILL FILL_0__15740_ (
);

FILL FILL_0__15320_ (
);

FILL FILL_5__12286_ (
);

FILL SFILL33640x40050 (
);

FILL FILL_4__11699_ (
);

FILL FILL_4__11279_ (
);

FILL FILL_5__8729_ (
);

OAI21X1 _15869_ (
    .A(_5524__bF$buf1),
    .B(_4908_),
    .C(_6328_),
    .Y(_6329_)
);

FILL FILL_4__12640_ (
);

OAI22X1 _15449_ (
    .A(_5918_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf0),
    .D(_5919_),
    .Y(_5920_)
);

NAND2X1 _15029_ (
    .A(\datapath_1.PCJump [25]),
    .B(_5464_),
    .Y(_5509_)
);

FILL FILL_4__12220_ (
);

FILL FILL_0__10299_ (
);

DFFSR _10584_ (
    .Q(\datapath_1.regfile_1.regOut[29] [2]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1823_[2])
);

OAI21X1 _10164_ (
    .A(_1667_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1668_),
    .Y(_1628_[20])
);

FILL FILL_6__14498_ (
);

FILL FILL_3__11633_ (
);

FILL FILL_3__11213_ (
);

FILL FILL_6__14078_ (
);

FILL FILL_0__16105_ (
);

FILL SFILL94280x20050 (
);

FILL FILL_2__10626_ (
);

FILL FILL_2__9272_ (
);

FILL FILL_0__11660_ (
);

FILL FILL_0__11240_ (
);

FILL FILL_2__13098_ (
);

FILL FILL_5__14852_ (
);

FILL FILL_5__14432_ (
);

FILL FILL_5__14012_ (
);

OAI21X1 _8732_ (
    .A(_936_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .C(_937_),
    .Y(_913_[12])
);

FILL SFILL8680x82050 (
);

OAI21X1 _8312_ (
    .A(_781_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_782_),
    .Y(_718_[0])
);

FILL SFILL33960x16050 (
);

FILL FILL_4__13845_ (
);

FILL FILL_4__13425_ (
);

FILL FILL_4__13005_ (
);

FILL FILL_0__9098_ (
);

FILL FILL_3__7195_ (
);

NOR2X1 _11789_ (
    .A(_2148_),
    .B(_2881_),
    .Y(_2882_)
);

INVX1 _11369_ (
    .A(_2328_),
    .Y(_2486_)
);

FILL FILL_3__12838_ (
);

FILL FILL_1__13872_ (
);

FILL FILL_3__12418_ (
);

FILL FILL_1__13452_ (
);

FILL FILL_1__13032_ (
);

FILL FILL_0__12865_ (
);

OAI21X1 _12730_ (
    .A(_3511_),
    .B(IRWrite_bF$buf5),
    .C(_3512_),
    .Y(_3490_[11])
);

FILL FILL_0__12445_ (
);

FILL FILL_0__12025_ (
);

NAND3X1 _12310_ (
    .A(_3269_),
    .B(_3270_),
    .C(_3271_),
    .Y(\datapath_1.alu_1.ALUInB [23])
);

FILL FILL_5__8482_ (
);

FILL FILL_5__8062_ (
);

FILL FILL_5__15637_ (
);

FILL FILL_5__15217_ (
);

NAND2X1 _9937_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1558_)
);

FILL FILL_3__16251_ (
);

NAND2X1 _9517_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1339_)
);

FILL FILL_1__8894_ (
);

FILL FILL_5__10772_ (
);

FILL FILL_1__8474_ (
);

FILL FILL_1__8054_ (
);

FILL SFILL63720x34050 (
);

FILL FILL_2__15664_ (
);

FILL FILL_2__15244_ (
);

FILL FILL_1__14657_ (
);

FILL FILL_1__14237_ (
);

FILL SFILL53800x70050 (
);

FILL FILL_3__9761_ (
);

INVX1 _13935_ (
    .A(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_4437_)
);

FILL FILL_3__9341_ (
);

INVX1 _13515_ (
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_4026_)
);

FILL FILL_5__9267_ (
);

FILL SFILL13640x81050 (
);

FILL SFILL69000x41050 (
);

FILL SFILL109480x61050 (
);

FILL FILL_5__11977_ (
);

FILL FILL_1__9679_ (
);

FILL FILL_5__11557_ (
);

FILL FILL_3__12591_ (
);

FILL FILL_1__9259_ (
);

FILL FILL_5__11137_ (
);

FILL FILL_3__12171_ (
);

BUFX2 BUFX2_insert1090 (
    .A(rst),
    .Y(rst_hier0_bF$buf3)
);

FILL FILL_2__16449_ (
);

BUFX2 BUFX2_insert1091 (
    .A(rst),
    .Y(rst_hier0_bF$buf2)
);

FILL FILL_2__16029_ (
);

FILL FILL_4__7684_ (
);

BUFX2 BUFX2_insert1092 (
    .A(rst),
    .Y(rst_hier0_bF$buf1)
);

BUFX2 BUFX2_insert1093 (
    .A(rst),
    .Y(rst_hier0_bF$buf0)
);

FILL FILL_2__11584_ (
);

FILL FILL_2__11164_ (
);

FILL FILL_1__10997_ (
);

FILL FILL_1__10577_ (
);

FILL FILL_1__10157_ (
);

FILL FILL_4__11911_ (
);

FILL FILL_5__15390_ (
);

FILL FILL_6__8971_ (
);

FILL FILL_0__7584_ (
);

FILL SFILL74280x61050 (
);

DFFSR _9690_ (
    .Q(\datapath_1.regfile_1.regOut[22] [4]),
    .CLK(clk_bF$buf51),
    .R(rst_bF$buf39),
    .S(vdd),
    .D(_1368_[4])
);

FILL FILL_0__7164_ (
);

NAND2X1 _9270_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1215_)
);

FILL FILL_1_CLKBUF1_insert220 (
);

FILL FILL_3__10904_ (
);

FILL FILL_1_CLKBUF1_insert221 (
);

FILL FILL_1_CLKBUF1_insert222 (
);

FILL FILL_1_CLKBUF1_insert223 (
);

FILL FILL_4__14383_ (
);

FILL FILL_1_CLKBUF1_insert224 (
);

FILL FILL_2__8963_ (
);

FILL FILL_0__10931_ (
);

FILL FILL_3__13796_ (
);

FILL FILL_0__10511_ (
);

FILL FILL_2__8123_ (
);

FILL FILL_3__13376_ (
);

FILL FILL_4__8889_ (
);

FILL FILL_4__8469_ (
);

FILL FILL_2__12789_ (
);

FILL FILL_2__12369_ (
);

FILL FILL_5__13703_ (
);

FILL FILL_1__6960_ (
);

FILL FILL_4__9410_ (
);

FILL FILL_2__13730_ (
);

FILL FILL_2__13310_ (
);

FILL FILL_5__16175_ (
);

FILL FILL_3__6886_ (
);

FILL FILL_0__8789_ (
);

FILL FILL_6__9756_ (
);

FILL FILL_0__8369_ (
);

FILL SFILL13560x43050 (
);

FILL FILL_1__12723_ (
);

FILL FILL_4__15588_ (
);

FILL FILL_4__15168_ (
);

FILL FILL_1__12303_ (
);

FILL FILL_0__9730_ (
);

FILL FILL_2__9748_ (
);

FILL FILL_0__11716_ (
);

FILL FILL_1__15195_ (
);

FILL FILL_6__15915_ (
);

FILL FILL_5__7753_ (
);

FILL FILL_5__7333_ (
);

INVX1 _14893_ (
    .A(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_5375_)
);

NOR2X1 _14473_ (
    .A(_4963_),
    .B(_4951_),
    .Y(_4964_)
);

FILL FILL_0__14188_ (
);

INVX1 _14053_ (
    .A(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_4553_)
);

FILL FILL_5__14908_ (
);

FILL FILL_3__15942_ (
);

FILL FILL_3__15522_ (
);

FILL FILL_3__15102_ (
);

FILL FILL_1__7745_ (
);

FILL FILL_1__7325_ (
);

FILL FILL_2__14935_ (
);

FILL FILL_2__14515_ (
);

FILL FILL_5__12095_ (
);

FILL FILL_1__13928_ (
);

FILL FILL_1__13508_ (
);

FILL FILL_4__11088_ (
);

FILL FILL_3__8612_ (
);

FILL SFILL104360x49050 (
);

FILL FILL_5__8958_ (
);

FILL FILL_5__8118_ (
);

FILL FILL_6__11835_ (
);

AOI21X1 _15678_ (
    .A(\datapath_1.regfile_1.regOut[27] [15]),
    .B(_5570__bF$buf3),
    .C(_6142_),
    .Y(_6143_)
);

FILL FILL_6__11415_ (
);

NOR2X1 _15258_ (
    .A(_5717_),
    .B(_5733_),
    .Y(_5734_)
);

FILL FILL_3__16307_ (
);

OAI21X1 _10393_ (
    .A(_1779_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .C(_1780_),
    .Y(_1758_[11])
);

FILL FILL_5__10828_ (
);

FILL FILL_5__10408_ (
);

FILL FILL_3__11862_ (
);

FILL FILL_3__11442_ (
);

FILL FILL_3__11022_ (
);

FILL FILL_4__6955_ (
);

FILL FILL_0__16334_ (
);

FILL FILL_2__10435_ (
);

FILL FILL_2__9081_ (
);

FILL FILL_2__10015_ (
);

FILL FILL_5__14661_ (
);

FILL FILL_5__14241_ (
);

FILL FILL_0__6855_ (
);

FILL FILL112440x55050 (
);

OAI21X1 _8961_ (
    .A(_1048_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1049_),
    .Y(_1043_[3])
);

DFFSR _8541_ (
    .Q(\datapath_1.regfile_1.regOut[13] [7]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_783_[7])
);

NAND2X1 _8121_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_632_)
);

FILL FILL_4__13654_ (
);

FILL FILL_4__13234_ (
);

OAI21X1 _11598_ (
    .A(_2704_),
    .B(_2241_),
    .C(_2264_),
    .Y(_2705_)
);

INVX2 _11178_ (
    .A(_2296_),
    .Y(_2297_)
);

FILL FILL_2__7814_ (
);

FILL FILL_3__12647_ (
);

FILL FILL_1__13681_ (
);

FILL FILL_3__12227_ (
);

FILL FILL_1__13261_ (
);

FILL SFILL89640x5050 (
);

FILL FILL_6_BUFX2_insert4 (
);

FILL FILL_0__12254_ (
);

FILL FILL_6_BUFX2_insert9 (
);

FILL FILL_5__15866_ (
);

FILL FILL_5__15446_ (
);

FILL FILL_5__15026_ (
);

NAND2X1 _9746_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1451_)
);

FILL FILL_3__16060_ (
);

DFFSR _9326_ (
    .Q(\datapath_1.regfile_1.regOut[19] [24]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf26),
    .S(vdd),
    .D(_1173_[24])
);

FILL FILL_5__10581_ (
);

FILL FILL_5__10161_ (
);

FILL FILL_4__14859_ (
);

FILL FILL112440x10050 (
);

FILL FILL_2__15893_ (
);

FILL FILL_4__14439_ (
);

FILL FILL_4__14019_ (
);

FILL FILL_2__15473_ (
);

FILL FILL_2__15053_ (
);

FILL FILL_1__14886_ (
);

FILL FILL_1__14466_ (
);

FILL FILL_1__14046_ (
);

FILL FILL_4__15800_ (
);

FILL FILL_3__9990_ (
);

FILL FILL_0__13879_ (
);

FILL FILL_3__9150_ (
);

INVX1 _13744_ (
    .A(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_4250_)
);

FILL FILL_0__13459_ (
);

NOR2X1 _13324_ (
    .A(_3781_),
    .B(_3853_),
    .Y(\datapath_1.regfile_1.regEn [14])
);

FILL FILL_0__13039_ (
);

FILL FILL_5__9496_ (
);

FILL FILL_0__14820_ (
);

FILL FILL_0__14400_ (
);

FILL FILL_5__11786_ (
);

FILL FILL_1__9488_ (
);

FILL FILL_5__11366_ (
);

FILL FILL_2__16258_ (
);

FILL FILL_4__7493_ (
);

FILL FILL_4__7073_ (
);

FILL FILL_4__10779_ (
);

FILL FILL_4__10359_ (
);

FILL FILL_2__11393_ (
);

FILL FILL_5__7809_ (
);

FILL FILL_1__10386_ (
);

OAI22X1 _14949_ (
    .A(_5428_),
    .B(_3930__bF$buf0),
    .C(_3971__bF$buf2),
    .D(_5429_),
    .Y(_5430_)
);

AOI22X1 _14529_ (
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .B(_3894_),
    .C(_4090_),
    .D(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_5019_)
);

FILL FILL_4__11720_ (
);

FILL FILL_4__11300_ (
);

AOI21X1 _14109_ (
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .B(_4115_),
    .C(_4607_),
    .Y(_4608_)
);

FILL FILL_4__14192_ (
);

FILL FILL_0__15605_ (
);

FILL SFILL94280x15050 (
);

FILL FILL_2__8772_ (
);

FILL FILL_2__8352_ (
);

FILL FILL_0__10320_ (
);

FILL FILL_4__8698_ (
);

FILL FILL_2__12598_ (
);

FILL FILL_2__12178_ (
);

FILL FILL_5__13932_ (
);

FILL FILL_5__13512_ (
);

FILL SFILL8680x77050 (
);

OAI21X1 _7812_ (
    .A(_465_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_466_),
    .Y(_458_[4])
);

FILL FILL_4_BUFX2_insert400 (
);

FILL FILL_4_BUFX2_insert401 (
);

FILL FILL_4_BUFX2_insert402 (
);

FILL FILL_4__12505_ (
);

FILL FILL_4_BUFX2_insert403 (
);

FILL FILL_4_BUFX2_insert404 (
);

FILL FILL_4_BUFX2_insert405 (
);

FILL FILL_0__8598_ (
);

FILL FILL_4_BUFX2_insert406 (
);

DFFSR _10869_ (
    .Q(\datapath_1.regfile_1.regOut[31] [31]),
    .CLK(clk_bF$buf86),
    .R(rst_bF$buf27),
    .S(vdd),
    .D(_1953_[31])
);

FILL FILL_4_BUFX2_insert407 (
);

NAND2X1 _10449_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1818_)
);

FILL FILL_4_BUFX2_insert408 (
);

NAND2X1 _10029_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1599_)
);

FILL FILL_4_BUFX2_insert409 (
);

FILL FILL_3__11918_ (
);

FILL FILL_1__12952_ (
);

FILL FILL_4__15397_ (
);

FILL FILL_1__12532_ (
);

FILL FILL_1__12112_ (
);

FILL SFILL84280x58050 (
);

FILL FILL_2__9977_ (
);

FILL FILL_0__11945_ (
);

FILL FILL_2__9557_ (
);

FILL FILL_2__9137_ (
);

OAI21X1 _11810_ (
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(_2120_),
    .C(_2900_),
    .Y(_2901_)
);

FILL FILL_0__11525_ (
);

FILL FILL_0__11105_ (
);

FILL FILL_5__7982_ (
);

FILL FILL_5__7562_ (
);

NOR2X1 _14282_ (
    .A(_4773_),
    .B(_4776_),
    .Y(_4777_)
);

FILL FILL_5__14717_ (
);

FILL FILL_3__15751_ (
);

FILL FILL_3__15331_ (
);

FILL FILL_1__7974_ (
);

FILL FILL_1__7554_ (
);

FILL SFILL8680x32050 (
);

FILL FILL_2__14744_ (
);

FILL FILL_2__14324_ (
);

FILL FILL_1__13737_ (
);

FILL FILL_1__13317_ (
);

FILL FILL_3__8841_ (
);

FILL FILL_3__8001_ (
);

FILL SFILL84280x13050 (
);

FILL FILL_5__8767_ (
);

FILL FILL_5__8347_ (
);

NOR2X1 _15487_ (
    .A(_5956_),
    .B(_5955_),
    .Y(_5957_)
);

NOR3X1 _15067_ (
    .A(_5546_),
    .B(_5540_),
    .C(_5542_),
    .Y(_5547_)
);

FILL SFILL109480x56050 (
);

FILL FILL_3__16116_ (
);

FILL FILL_5__10637_ (
);

FILL FILL_1__8759_ (
);

FILL FILL_1__8339_ (
);

FILL FILL_3__11671_ (
);

FILL FILL_3__11251_ (
);

FILL SFILL8600x30050 (
);

FILL FILL_2__15949_ (
);

FILL FILL_2__15529_ (
);

FILL FILL_2__15109_ (
);

FILL FILL_0__16143_ (
);

FILL FILL_2__10664_ (
);

FILL FILL_2__10244_ (
);

FILL FILL_3__9626_ (
);

FILL FILL_3_BUFX2_insert420 (
);

FILL SFILL109560x9050 (
);

FILL FILL_3_BUFX2_insert421 (
);

FILL FILL_3__9206_ (
);

FILL FILL_3_BUFX2_insert422 (
);

FILL FILL_5__14890_ (
);

FILL SFILL84200x11050 (
);

FILL FILL_5__14470_ (
);

FILL FILL_3_BUFX2_insert423 (
);

FILL FILL_3_BUFX2_insert424 (
);

FILL FILL_5__14050_ (
);

FILL FILL_3_BUFX2_insert425 (
);

NAND2X1 _8770_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_963_)
);

FILL FILL_3_BUFX2_insert426 (
);

NAND2X1 _8350_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_744_)
);

FILL FILL_3_BUFX2_insert427 (
);

FILL FILL_3_BUFX2_insert428 (
);

FILL FILL_4__13883_ (
);

FILL FILL_3_BUFX2_insert429 (
);

FILL FILL_4__13463_ (
);

FILL FILL_6__12009_ (
);

FILL FILL_4__13043_ (
);

FILL SFILL13640x31050 (
);

FILL FILL_3__12876_ (
);

FILL FILL_2__7623_ (
);

FILL FILL_2__7203_ (
);

FILL FILL_3__12456_ (
);

FILL FILL_1__13490_ (
);

FILL FILL_3__12036_ (
);

FILL SFILL109480x11050 (
);

FILL FILL_4__7969_ (
);

FILL FILL_4__7549_ (
);

FILL FILL_2__11869_ (
);

FILL FILL_2__11449_ (
);

FILL SFILL38840x80050 (
);

FILL FILL_0__12483_ (
);

FILL FILL_2__11029_ (
);

FILL FILL_0__12063_ (
);

FILL FILL_4__8910_ (
);

FILL FILL_5__15675_ (
);

FILL FILL_0__7869_ (
);

FILL FILL_5__15255_ (
);

NAND2X1 _9975_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .Y(_1627_)
);

FILL FILL_0__7449_ (
);

INVX1 _9555_ (
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_1364_)
);

INVX1 _9135_ (
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_1145_)
);

FILL FILL_5__10390_ (
);

FILL FILL_1__8092_ (
);

FILL SFILL74280x11050 (
);

FILL FILL_1__11803_ (
);

FILL FILL_4__14668_ (
);

FILL FILL_4__14248_ (
);

FILL FILL_2__15282_ (
);

FILL FILL_2__8828_ (
);

FILL FILL_1__14695_ (
);

FILL FILL_1__14275_ (
);

FILL SFILL99480x60050 (
);

FILL FILL_0_BUFX2_insert550 (
);

FILL FILL_0_BUFX2_insert551 (
);

FILL FILL_0_BUFX2_insert552 (
);

FILL FILL_0_BUFX2_insert553 (
);

FILL FILL_0_BUFX2_insert554 (
);

NAND3X1 _13973_ (
    .A(_4473_),
    .B(_4474_),
    .C(_4472_),
    .Y(_4475_)
);

FILL FILL_0__13688_ (
);

FILL FILL_0__13268_ (
);

INVX1 _13553_ (
    .A(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_4063_)
);

FILL FILL_0_BUFX2_insert555 (
);

FILL FILL_0_BUFX2_insert556 (
);

INVX1 _13133_ (
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3720_)
);

FILL FILL_0_BUFX2_insert557 (
);

FILL FILL_0_BUFX2_insert558 (
);

FILL FILL_3__14602_ (
);

FILL FILL_0_BUFX2_insert559 (
);

FILL FILL_5__11595_ (
);

FILL FILL_5__11175_ (
);

FILL FILL_1__9297_ (
);

FILL FILL_2__16067_ (
);

FILL FILL_4__10168_ (
);

FILL FILL_5__7618_ (
);

FILL FILL_1__10195_ (
);

FILL FILL_6__10915_ (
);

INVX1 _14758_ (
    .A(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_5243_)
);

INVX1 _14338_ (
    .A(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_4832_)
);

FILL FILL_3__15807_ (
);

FILL FILL_1__16001_ (
);

FILL FILL_3__10942_ (
);

FILL FILL_3__10522_ (
);

FILL FILL_3__10102_ (
);

FILL FILL_0__15834_ (
);

FILL FILL_0__15414_ (
);

FILL FILL_2__8581_ (
);

FILL SFILL33800x61050 (
);

FILL SFILL64200x52050 (
);

FILL FILL_4__8087_ (
);

FILL FILL_5__13741_ (
);

FILL FILL_5__13321_ (
);

NAND2X1 _7621_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_380_)
);

NAND2X1 _7201_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_161_)
);

FILL FILL_4__12734_ (
);

FILL FILL_4__12314_ (
);

NAND2X1 _10678_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1930_)
);

FILL FILL_6__9374_ (
);

NAND2X1 _10258_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1711_)
);

FILL FILL_3__11727_ (
);

FILL FILL_1__12761_ (
);

FILL FILL_3__11307_ (
);

FILL FILL_1__12341_ (
);

FILL FILL112040x36050 (
);

FILL FILL_2__9786_ (
);

FILL FILL_0__11754_ (
);

FILL FILL_2__9366_ (
);

FILL FILL_3__14199_ (
);

FILL FILL_0__11334_ (
);

FILL FILL_5__7371_ (
);

FILL FILL_5__14946_ (
);

OAI22X1 _14091_ (
    .A(_4589_),
    .B(_3949_),
    .C(_3881_),
    .D(_4588_),
    .Y(_4590_)
);

FILL FILL_3__15980_ (
);

FILL FILL_5__14526_ (
);

FILL FILL_3__15560_ (
);

FILL FILL_5__14106_ (
);

FILL FILL_3__15140_ (
);

NAND2X1 _8826_ (
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_980_)
);

DFFSR _8406_ (
    .Q(\datapath_1.regfile_1.regOut[12] [0]),
    .CLK(clk_bF$buf4),
    .R(rst_bF$buf63),
    .S(vdd),
    .D(_718_[0])
);

FILL FILL_1__7363_ (
);

FILL FILL_4__13939_ (
);

FILL FILL_2__14973_ (
);

FILL FILL_4__13519_ (
);

FILL FILL_2__14553_ (
);

FILL FILL_2__14133_ (
);

FILL FILL_3__7289_ (
);

FILL FILL_1__13966_ (
);

FILL FILL_1__13546_ (
);

FILL FILL_1__13126_ (
);

FILL FILL_3__8650_ (
);

FILL FILL_0__12959_ (
);

FILL FILL_3__8230_ (
);

NAND2X1 _12824_ (
    .A(\datapath_1.rd1 [0]),
    .B(vdd),
    .Y(_3619_)
);

NAND2X1 _12404_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [20]),
    .Y(_3335_)
);

FILL FILL_0__12119_ (
);

FILL FILL_5__8996_ (
);

FILL FILL_5__8576_ (
);

AOI21X1 _15296_ (
    .A(_5749_),
    .B(_5770_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [5])
);

FILL FILL_0__13900_ (
);

FILL FILL_3__16345_ (
);

FILL FILL_1__8988_ (
);

FILL FILL_5__10446_ (
);

FILL FILL_1__8568_ (
);

FILL FILL_1__8148_ (
);

FILL FILL_5__10026_ (
);

FILL FILL_3__11480_ (
);

FILL FILL_3__11060_ (
);

FILL FILL_2__15758_ (
);

FILL FILL_2__15338_ (
);

FILL FILL_4__6993_ (
);

FILL FILL_0__16372_ (
);

FILL FILL_2__10893_ (
);

FILL FILL_2__10053_ (
);

FILL SFILL23720x66050 (
);

FILL FILL_3__9855_ (
);

FILL FILL_3__9015_ (
);

AOI21X1 _13609_ (
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .B(_4115_),
    .C(_4117_),
    .Y(_4118_)
);

FILL FILL_4__10800_ (
);

FILL FILL_0__6893_ (
);

FILL FILL_4__13692_ (
);

FILL FILL_4__13272_ (
);

FILL FILL_2__7852_ (
);

FILL FILL_2__7432_ (
);

FILL FILL_3__12265_ (
);

FILL FILL_4__7358_ (
);

FILL FILL_2__11678_ (
);

FILL FILL_2__11258_ (
);

FILL FILL_0__12292_ (
);

FILL SFILL23720x21050 (
);

FILL FILL_5__15484_ (
);

FILL FILL_5__15064_ (
);

FILL FILL_0__7678_ (
);

FILL FILL_6__8645_ (
);

INVX1 _9784_ (
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_1476_)
);

FILL SFILL103480x54050 (
);

INVX1 _9364_ (
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_1257_)
);

FILL FILL_4__14897_ (
);

FILL FILL_4__14477_ (
);

FILL FILL_1__11612_ (
);

FILL FILL_4__14057_ (
);

FILL FILL_2__15091_ (
);

FILL FILL_2__8637_ (
);

FILL FILL_2__8217_ (
);

FILL FILL_1__14084_ (
);

FILL SFILL109960x58050 (
);

OAI22X1 _13782_ (
    .A(_4286_),
    .B(_3955__bF$buf1),
    .C(_3954__bF$buf1),
    .D(_4287_),
    .Y(_4288_)
);

FILL FILL_0__13497_ (
);

NOR2X1 _13362_ (
    .A(_3798_),
    .B(_3756_),
    .Y(\datapath_1.regfile_1.regEn [29])
);

FILL FILL_3__14831_ (
);

FILL FILL_3__14411_ (
);

FILL FILL_4__9924_ (
);

FILL FILL_4__9504_ (
);

FILL SFILL8680x27050 (
);

FILL FILL_2__13824_ (
);

FILL FILL_2__13404_ (
);

FILL FILL_5__16269_ (
);

FILL FILL_2__16296_ (
);

FILL FILL_4__10397_ (
);

FILL FILL_3__7501_ (
);

FILL FILL_0__9404_ (
);

FILL FILL_1__15289_ (
);

FILL FILL_5__7847_ (
);

FILL FILL_5__7427_ (
);

FILL FILL_4__16203_ (
);

OAI22X1 _14987_ (
    .A(_5463__bF$buf0),
    .B(_3975_),
    .C(_5466__bF$buf2),
    .D(_3965_),
    .Y(_5467_)
);

OAI22X1 _14567_ (
    .A(_3902__bF$buf0),
    .B(_5054_),
    .C(_5055_),
    .D(_3935__bF$buf4),
    .Y(_5056_)
);

INVX1 _14147_ (
    .A(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_4645_)
);

FILL FILL_3__15616_ (
);

FILL FILL_1__16230_ (
);

FILL FILL_1__7839_ (
);

FILL FILL_3__10751_ (
);

FILL FILL_1__7419_ (
);

FILL SFILL8600x25050 (
);

FILL FILL_2__14609_ (
);

FILL FILL_0__15643_ (
);

FILL FILL_0__15223_ (
);

FILL SFILL48840x32050 (
);

FILL FILL_5__12189_ (
);

FILL FILL_2__8390_ (
);

FILL FILL_3__8706_ (
);

FILL FILL_5__13970_ (
);

FILL FILL_5__13550_ (
);

FILL FILL_5__13130_ (
);

NAND2X1 _7850_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_492_)
);

NAND2X1 _7430_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_273_)
);

DFFSR _7010_ (
    .Q(\datapath_1.regfile_1.regOut[1] [12]),
    .CLK(clk_bF$buf103),
    .R(rst_bF$buf16),
    .S(vdd),
    .D(_3_[12])
);

FILL FILL_4__12963_ (
);

FILL FILL_4__12123_ (
);

FILL SFILL13640x26050 (
);

NAND2X1 _10487_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .Y(_1887_)
);

INVX1 _10067_ (
    .A(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_1624_)
);

FILL FILL_3__11956_ (
);

FILL FILL_1__12990_ (
);

FILL FILL_3__11536_ (
);

FILL FILL_1__12570_ (
);

FILL FILL_3__11116_ (
);

FILL FILL_1__12150_ (
);

FILL FILL_0__16008_ (
);

FILL FILL_2__10949_ (
);

FILL FILL_0__11983_ (
);

FILL FILL_2__10529_ (
);

FILL FILL_2__9595_ (
);

FILL FILL_0__11563_ (
);

FILL FILL_2__10109_ (
);

FILL FILL_0__11143_ (
);

FILL FILL_6__15342_ (
);

FILL FILL_5__7180_ (
);

FILL SFILL74200x49050 (
);

FILL FILL_5__14755_ (
);

FILL FILL_0__6949_ (
);

FILL FILL_5__14335_ (
);

INVX1 _8635_ (
    .A(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_893_)
);

INVX1 _8215_ (
    .A(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_674_)
);

FILL FILL_1__7592_ (
);

FILL FILL_1__7172_ (
);

FILL FILL_4__13748_ (
);

FILL FILL_4__13328_ (
);

FILL FILL_2__14782_ (
);

FILL FILL_2__14362_ (
);

FILL FILL_3__7098_ (
);

FILL FILL112200x62050 (
);

FILL FILL_1__13775_ (
);

FILL SFILL99480x55050 (
);

FILL FILL_1__13355_ (
);

FILL FILL_0__12768_ (
);

INVX1 _12633_ (
    .A(\datapath_1.Data [22]),
    .Y(_3468_)
);

FILL FILL_0__12348_ (
);

INVX8 _12213_ (
    .A(ALUSrcB_0_bF$buf2),
    .Y(_3198_)
);

FILL SFILL38840x30050 (
);

FILL FILL_5__8385_ (
);

FILL FILL_6__11262_ (
);

FILL FILL_3__16154_ (
);

FILL FILL112120x69050 (
);

FILL FILL_5__10675_ (
);

FILL FILL_5__10255_ (
);

FILL FILL_1__8377_ (
);

FILL FILL_2__15987_ (
);

FILL FILL_2__15567_ (
);

FILL FILL_2__15147_ (
);

FILL FILL_0__16181_ (
);

FILL FILL_2__10282_ (
);

FILL SFILL99480x10050 (
);

FILL FILL_3__9664_ (
);

FILL FILL_3_BUFX2_insert800 (
);

NAND3X1 _13838_ (
    .A(_4332_),
    .B(_4335_),
    .C(_4342_),
    .Y(_4343_)
);

FILL FILL_3__9244_ (
);

FILL FILL_3_BUFX2_insert801 (
);

NAND2X1 _13418_ (
    .A(_3904_),
    .B(_3889_),
    .Y(_3930_)
);

FILL FILL_3_BUFX2_insert802 (
);

FILL FILL_3_BUFX2_insert803 (
);

FILL FILL_3_BUFX2_insert804 (
);

FILL FILL_1__15921_ (
);

FILL FILL_3_BUFX2_insert805 (
);

FILL SFILL28840x73050 (
);

FILL FILL_1__15501_ (
);

FILL FILL_3_BUFX2_insert806 (
);

FILL FILL_3_BUFX2_insert807 (
);

FILL FILL_6__12887_ (
);

FILL FILL_3_BUFX2_insert808 (
);

FILL FILL_3_BUFX2_insert809 (
);

FILL FILL_4__13081_ (
);

FILL FILL_0__14914_ (
);

FILL SFILL68920x69050 (
);

FILL SFILL33800x56050 (
);

FILL SFILL64200x47050 (
);

FILL FILL_3__12494_ (
);

FILL FILL_2__7241_ (
);

FILL SFILL9160x50050 (
);

FILL FILL_3__12074_ (
);

FILL FILL_4__7587_ (
);

FILL FILL_4__7167_ (
);

FILL FILL_2__11487_ (
);

FILL FILL_2__11067_ (
);

FILL FILL_5__12401_ (
);

FILL FILL_4__11814_ (
);

FILL FILL_5__15293_ (
);

FILL FILL_0__7487_ (
);

FILL FILL_0__7067_ (
);

INVX1 _9593_ (
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_1369_)
);

FILL FILL_6__8454_ (
);

OAI21X1 _9173_ (
    .A(_1169_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .C(_1170_),
    .Y(_1108_[31])
);

FILL FILL_3__10807_ (
);

FILL FILL_1__11841_ (
);

FILL FILL_4__14286_ (
);

FILL FILL_1__11421_ (
);

FILL FILL_1__11001_ (
);

FILL FILL_2__8866_ (
);

FILL FILL_0__10834_ (
);

FILL FILL_2__8446_ (
);

FILL FILL_3__13699_ (
);

FILL FILL_3__13279_ (
);

FILL FILL_0__10414_ (
);

FILL FILL_0_BUFX2_insert930 (
);

FILL FILL_5__6871_ (
);

FILL SFILL33800x11050 (
);

FILL FILL_0_BUFX2_insert931 (
);

FILL FILL_0_BUFX2_insert932 (
);

FILL FILL_0_BUFX2_insert933 (
);

FILL FILL_0_BUFX2_insert934 (
);

NOR2X1 _13591_ (
    .A(_4096_),
    .B(_4099_),
    .Y(_4100_)
);

FILL FILL_0_BUFX2_insert935 (
);

FILL FILL_0_BUFX2_insert936 (
);

OAI21X1 _13171_ (
    .A(_3744_),
    .B(PCEn_bF$buf0),
    .C(_3745_),
    .Y(_3685_[30])
);

FILL FILL_5__13606_ (
);

FILL FILL_0_BUFX2_insert937 (
);

FILL FILL_3__14640_ (
);

FILL FILL_0_BUFX2_insert938 (
);

FILL FILL_3__14220_ (
);

DFFSR _7906_ (
    .Q(\datapath_1.regfile_1.regOut[8] [12]),
    .CLK(clk_bF$buf101),
    .R(rst_bF$buf102),
    .S(vdd),
    .D(_458_[12])
);

FILL FILL_0_BUFX2_insert939 (
);

FILL FILL_1__6863_ (
);

FILL FILL_4__9733_ (
);

FILL FILL_2__13633_ (
);

FILL SFILL103640x80050 (
);

FILL FILL_2__13213_ (
);

FILL FILL_5__16078_ (
);

FILL FILL_1__12626_ (
);

FILL FILL_1__12206_ (
);

FILL SFILL18840x71050 (
);

FILL FILL_0__9633_ (
);

FILL FILL_3__7730_ (
);

FILL FILL_3__7310_ (
);

OAI21X1 _11904_ (
    .A(_2976_),
    .B(IorD_bF$buf3),
    .C(_2977_),
    .Y(_1_[5])
);

FILL FILL_0__9213_ (
);

FILL FILL_0__11619_ (
);

FILL FILL_1__15098_ (
);

FILL FILL_6__15818_ (
);

FILL FILL_5__7236_ (
);

FILL FILL_4__16012_ (
);

OAI22X1 _14796_ (
    .A(_5279_),
    .B(_3936__bF$buf3),
    .C(_3905__bF$buf1),
    .D(_5278_),
    .Y(_5280_)
);

INVX1 _14376_ (
    .A(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_4869_)
);

FILL SFILL13800x1050 (
);

FILL FILL_3__15845_ (
);

FILL FILL_3__15425_ (
);

FILL FILL_3__15005_ (
);

FILL SFILL13720x6050 (
);

FILL FILL_3__10980_ (
);

FILL FILL_1__7228_ (
);

FILL FILL_3__10560_ (
);

FILL FILL_3__10140_ (
);

FILL FILL_6_BUFX2_insert311 (
);

FILL FILL_2__14838_ (
);

FILL FILL_2__14418_ (
);

FILL FILL_0__15872_ (
);

FILL FILL_0__15452_ (
);

FILL FILL_0__15032_ (
);

FILL FILL_6_BUFX2_insert316 (
);

FILL FILL_3__8515_ (
);

FILL FILL_6__6940_ (
);

FILL FILL_4__12772_ (
);

FILL FILL_6__11318_ (
);

FILL FILL_4__12352_ (
);

INVX1 _10296_ (
    .A(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_1736_)
);

FILL SFILL103560x42050 (
);

FILL FILL_2__6932_ (
);

FILL FILL_5__9802_ (
);

FILL FILL_3__11765_ (
);

FILL FILL_3__11345_ (
);

FILL FILL_4__6858_ (
);

FILL FILL_0__16237_ (
);

NOR2X1 _16102_ (
    .A(_6555_),
    .B(_6549_),
    .Y(_6556_)
);

FILL FILL_2__10758_ (
);

FILL FILL_0__11792_ (
);

FILL FILL_0__11372_ (
);

FILL SFILL23720x16050 (
);

FILL FILL_5__14984_ (
);

FILL FILL_5__14564_ (
);

FILL FILL_5__14144_ (
);

INVX1 _8864_ (
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_1005_)
);

FILL FILL_6__7725_ (
);

INVX1 _8444_ (
    .A(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_786_)
);

DFFSR _8024_ (
    .Q(\datapath_1.regfile_1.regOut[9] [2]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_523_[2])
);

FILL FILL_4__13977_ (
);

FILL FILL_4__13557_ (
);

FILL SFILL48920x65050 (
);

FILL FILL_2__14591_ (
);

FILL FILL_4__13137_ (
);

FILL FILL_2__14171_ (
);

FILL FILL_2__7717_ (
);

FILL FILL_1__13584_ (
);

FILL FILL_1__13164_ (
);

FILL FILL_0__12997_ (
);

FILL FILL_0__12577_ (
);

INVX1 _12862_ (
    .A(\datapath_1.a [13]),
    .Y(_3580_)
);

FILL FILL_0__12157_ (
);

INVX1 _12442_ (
    .A(ALUOut[1]),
    .Y(_3361_)
);

NAND3X1 _12022_ (
    .A(_3060_),
    .B(_3061_),
    .C(_3062_),
    .Y(\datapath_1.mux_pcsrc.dout [8])
);

FILL FILL_3__13911_ (
);

FILL FILL_5__8194_ (
);

FILL FILL_5_BUFX2_insert330 (
);

FILL FILL_2__12904_ (
);

FILL FILL_5__15769_ (
);

FILL FILL_5_BUFX2_insert331 (
);

FILL FILL_5__15349_ (
);

FILL FILL_5_BUFX2_insert332 (
);

FILL FILL_3__16383_ (
);

FILL FILL_5_BUFX2_insert333 (
);

FILL SFILL109560x39050 (
);

FILL FILL_5_BUFX2_insert334 (
);

OAI21X1 _9649_ (
    .A(_1405_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1406_),
    .Y(_1368_[19])
);

OAI21X1 _9229_ (
    .A(_1186_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .C(_1187_),
    .Y(_1173_[7])
);

FILL FILL_5_BUFX2_insert335 (
);

FILL FILL_5_BUFX2_insert336 (
);

FILL FILL_5_BUFX2_insert337 (
);

FILL FILL_1__8186_ (
);

FILL FILL_5__10064_ (
);

FILL FILL_5_BUFX2_insert338 (
);

FILL FILL_5_BUFX2_insert339 (
);

FILL FILL_2__15796_ (
);

FILL FILL_2__15376_ (
);

FILL FILL_0__8904_ (
);

FILL FILL_1__14789_ (
);

FILL FILL_1__14369_ (
);

FILL FILL_5__6927_ (
);

FILL FILL_4__15703_ (
);

FILL FILL_3__9893_ (
);

FILL FILL_3__9473_ (
);

AOI22X1 _13647_ (
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .B(_4005__bF$buf2),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_4155_)
);

NOR2X1 _13227_ (
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_3770_)
);

FILL FILL_5__9399_ (
);

FILL FILL_1__15730_ (
);

FILL FILL_1__15310_ (
);

FILL FILL_1__6919_ (
);

FILL FILL_0__14723_ (
);

FILL FILL_0__14303_ (
);

FILL SFILL13720x14050 (
);

FILL FILL_2__7890_ (
);

FILL FILL_5__11689_ (
);

FILL FILL_2__7470_ (
);

FILL FILL_5__11269_ (
);

FILL FILL_2__7050_ (
);

FILL FILL_2__11296_ (
);

FILL SFILL38920x63050 (
);

FILL FILL_5__12630_ (
);

FILL FILL_5__12210_ (
);

NAND2X1 _6930_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_21_)
);

FILL FILL_2_BUFX2_insert460 (
);

FILL FILL_2_BUFX2_insert461 (
);

FILL FILL_1__10289_ (
);

FILL FILL_2_BUFX2_insert462 (
);

FILL FILL_2_BUFX2_insert463 (
);

FILL FILL_2_BUFX2_insert464 (
);

FILL FILL_4__11623_ (
);

FILL FILL_4__11203_ (
);

FILL FILL_2_BUFX2_insert465 (
);

FILL FILL_2_BUFX2_insert466 (
);

FILL FILL_0__7296_ (
);

FILL FILL_2_BUFX2_insert467 (
);

FILL FILL_2_BUFX2_insert468 (
);

FILL FILL_2_BUFX2_insert469 (
);

FILL FILL_3__10616_ (
);

FILL FILL_0_CLKBUF1_insert160 (
);

FILL FILL_1__11650_ (
);

FILL FILL_1__11230_ (
);

FILL FILL_4__14095_ (
);

FILL FILL_0_CLKBUF1_insert161 (
);

FILL FILL_0__15928_ (
);

FILL FILL_0_CLKBUF1_insert162 (
);

FILL FILL_0__15508_ (
);

FILL FILL_0_CLKBUF1_insert163 (
);

FILL FILL_0_CLKBUF1_insert164 (
);

FILL FILL_0_CLKBUF1_insert165 (
);

FILL FILL_0_CLKBUF1_insert166 (
);

FILL FILL_2__8255_ (
);

FILL FILL_0__10643_ (
);

FILL FILL_0_CLKBUF1_insert167 (
);

FILL FILL_0_CLKBUF1_insert168 (
);

FILL FILL_3__13088_ (
);

FILL FILL_0_CLKBUF1_insert169 (
);

FILL FILL_5__13835_ (
);

FILL FILL_5__13415_ (
);

INVX1 _7715_ (
    .A(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_422_)
);

FILL FILL_4__9542_ (
);

FILL FILL_4__9122_ (
);

FILL FILL_4__12828_ (
);

FILL FILL_4__12408_ (
);

FILL FILL_2__13862_ (
);

FILL FILL_2__13442_ (
);

FILL FILL_2__13022_ (
);

FILL SFILL7880x70050 (
);

FILL FILL112200x57050 (
);

FILL FILL_1__12855_ (
);

FILL FILL_1__12435_ (
);

FILL FILL_1__12015_ (
);

FILL FILL_0__9862_ (
);

FILL FILL_0__11848_ (
);

FILL FILL_0__11428_ (
);

AOI21X1 _11713_ (
    .A(_2810_),
    .B(_2811_),
    .C(_2191_),
    .Y(_2812_)
);

FILL FILL_0__9022_ (
);

FILL FILL_0__11008_ (
);

FILL SFILL38840x25050 (
);

FILL FILL_5__7885_ (
);

FILL FILL_5__7465_ (
);

FILL FILL_4__16241_ (
);

FILL FILL_5__7045_ (
);

AOI21X1 _14185_ (
    .A(\datapath_1.regfile_1.regOut[6] [15]),
    .B(_4001__bF$buf2),
    .C(_4681_),
    .Y(_4682_)
);

FILL FILL_3__15654_ (
);

FILL FILL_3__15234_ (
);

FILL FILL_1__7877_ (
);

FILL FILL_1__7457_ (
);

FILL FILL_1__7037_ (
);

FILL FILL_2__14647_ (
);

FILL FILL_0__15681_ (
);

FILL FILL_2__14227_ (
);

FILL FILL_0__15261_ (
);

FILL SFILL89960x55050 (
);

FILL SFILL113640x77050 (
);

FILL FILL112200x12050 (
);

FILL FILL_1_BUFX2_insert480 (
);

FILL FILL_3__8744_ (
);

FILL FILL_1_BUFX2_insert481 (
);

FILL FILL_3__8324_ (
);

FILL FILL_1_BUFX2_insert482 (
);

OAI21X1 _12918_ (
    .A(_3616_),
    .B(vdd),
    .C(_3617_),
    .Y(_3555_[31])
);

FILL FILL_1_BUFX2_insert483 (
);

FILL FILL_1_BUFX2_insert484 (
);

FILL FILL_1_BUFX2_insert485 (
);

FILL SFILL28840x68050 (
);

FILL FILL_1_BUFX2_insert486 (
);

FILL SFILL3480x24050 (
);

FILL FILL_1_BUFX2_insert487 (
);

FILL FILL_1_BUFX2_insert488 (
);

FILL FILL_1_BUFX2_insert489 (
);

FILL FILL_4__12581_ (
);

FILL FILL_4__12161_ (
);

FILL FILL_3__16019_ (
);

FILL FILL_3__11994_ (
);

FILL FILL_5__9611_ (
);

FILL FILL_3__11574_ (
);

FILL FILL_3__11154_ (
);

FILL FILL112120x19050 (
);

NAND2X1 _16331_ (
    .A(gnd),
    .B(gnd),
    .Y(_6775_)
);

FILL FILL_0__16046_ (
);

FILL FILL_2__10567_ (
);

FILL FILL_2__10147_ (
);

FILL FILL_0__11181_ (
);

FILL FILL_5__11901_ (
);

FILL FILL_1__9603_ (
);

FILL SFILL89480x48050 (
);

FILL SFILL89960x10050 (
);

FILL FILL_3__9529_ (
);

FILL FILL_3__9109_ (
);

FILL FILL_5__14793_ (
);

FILL FILL_0__6987_ (
);

FILL FILL_5__14373_ (
);

DFFSR _8673_ (
    .Q(\datapath_1.regfile_1.regOut[14] [11]),
    .CLK(clk_bF$buf10),
    .R(rst_bF$buf61),
    .S(vdd),
    .D(_848_[11])
);

OAI21X1 _8253_ (
    .A(_698_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .C(_699_),
    .Y(_653_[23])
);

FILL FILL_1__10921_ (
);

FILL FILL_4__13786_ (
);

FILL SFILL28840x23050 (
);

FILL FILL_4__13366_ (
);

FILL FILL_1__10501_ (
);

FILL FILL_2__7946_ (
);

FILL FILL_3__12779_ (
);

FILL FILL_3__12359_ (
);

FILL FILL_2__7106_ (
);

FILL FILL_1__13393_ (
);

DFFSR _12671_ (
    .Q(\datapath_1.Data [8]),
    .CLK(clk_bF$buf37),
    .R(rst_bF$buf35),
    .S(vdd),
    .D(_3425_[8])
);

FILL FILL_0__12386_ (
);

NAND3X1 _12251_ (
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3227_)
);

FILL FILL_3__13720_ (
);

FILL FILL_3__13300_ (
);

FILL FILL_6__16165_ (
);

FILL FILL_5__15998_ (
);

FILL FILL_2__12713_ (
);

FILL FILL_5__15578_ (
);

FILL FILL_5__15158_ (
);

FILL FILL_3__16192_ (
);

OAI21X1 _9878_ (
    .A(_1517_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .C(_1518_),
    .Y(_1498_[10])
);

DFFSR _9458_ (
    .Q(\datapath_1.regfile_1.regOut[20] [28]),
    .CLK(clk_bF$buf46),
    .R(rst_bF$buf23),
    .S(vdd),
    .D(_1238_[28])
);

NAND2X1 _9038_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1101_)
);

FILL FILL_5__10293_ (
);

FILL FILL_1__11706_ (
);

FILL FILL_2__15185_ (
);

FILL FILL_0__8713_ (
);

FILL FILL_1__14598_ (
);

FILL FILL_1__14178_ (
);

FILL FILL_4__15932_ (
);

FILL FILL_4__15512_ (
);

OAI22X1 _13876_ (
    .A(_4379_),
    .B(_3972__bF$buf0),
    .C(_3920_),
    .D(_4378_),
    .Y(_4380_)
);

FILL FILL_3__9282_ (
);

OAI22X1 _13456_ (
    .A(_3967__bF$buf2),
    .B(_3964_),
    .C(_3966__bF$buf3),
    .D(_3965_),
    .Y(_3968_)
);

NAND2X1 _13036_ (
    .A(vdd),
    .B(\datapath_1.rd2 [28]),
    .Y(_3676_)
);

FILL FILL_6_BUFX2_insert1088 (
);

FILL FILL_3__14925_ (
);

FILL FILL_3__14505_ (
);

FILL FILL_6__12085_ (
);

FILL FILL_2__13918_ (
);

FILL FILL_0__14952_ (
);

FILL FILL_0__14532_ (
);

FILL SFILL63880x61050 (
);

FILL FILL_0__14112_ (
);

FILL FILL_5__11498_ (
);

FILL FILL_5__11078_ (
);

FILL FILL_0__9918_ (
);

FILL SFILL18840x21050 (
);

FILL SFILL58920x17050 (
);

FILL FILL_4__11852_ (
);

FILL FILL_4__11432_ (
);

FILL FILL_4__11012_ (
);

FILL FILL_6__8072_ (
);

FILL FILL_1__16324_ (
);

FILL FILL_3__10425_ (
);

FILL FILL_3__10005_ (
);

FILL FILL_0__15737_ (
);

FILL FILL_0__15317_ (
);

NOR2X1 _15602_ (
    .A(_6068_),
    .B(_6066_),
    .Y(_6069_)
);

FILL FILL_2__8484_ (
);

FILL FILL_0__10872_ (
);

FILL FILL_2__8064_ (
);

FILL FILL_0__10452_ (
);

FILL FILL_0__10032_ (
);

FILL FILL_6__14651_ (
);

FILL FILL_5__13644_ (
);

FILL FILL_5__13224_ (
);

INVX1 _7944_ (
    .A(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_534_)
);

FILL SFILL69080x75050 (
);

DFFSR _7524_ (
    .Q(\datapath_1.regfile_1.regOut[5] [14]),
    .CLK(clk_bF$buf13),
    .R(rst_bF$buf74),
    .S(vdd),
    .D(_263_[14])
);

OAI21X1 _7104_ (
    .A(_115_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .C(_116_),
    .Y(_68_[24])
);

FILL FILL_4__9771_ (
);

FILL FILL_4__9351_ (
);

FILL FILL_4__12637_ (
);

FILL FILL_2__13671_ (
);

FILL FILL_4__12217_ (
);

FILL FILL_2__13251_ (
);

FILL FILL_1__12244_ (
);

FILL FILL_0__9671_ (
);

FILL FILL_2__9269_ (
);

FILL FILL_0__9251_ (
);

NAND2X1 _11942_ (
    .A(IorD_bF$buf7),
    .B(ALUOut[18]),
    .Y(_3003_)
);

FILL FILL_0__11657_ (
);

FILL FILL_0__11237_ (
);

NAND3X1 _11522_ (
    .A(_2225_),
    .B(_2628_),
    .C(_2632_),
    .Y(_2633_)
);

INVX1 _11102_ (
    .A(\datapath_1.alu_1.ALUInA [23]),
    .Y(_2221_)
);

FILL FILL_5__7694_ (
);

FILL FILL_4__16050_ (
);

FILL FILL_6__10991_ (
);

FILL FILL_5__14849_ (
);

FILL FILL_3__15883_ (
);

FILL FILL_5__14429_ (
);

FILL FILL_5__14009_ (
);

FILL FILL_3__15463_ (
);

OAI21X1 _8729_ (
    .A(_934_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .C(_935_),
    .Y(_913_[11])
);

FILL FILL_3__15043_ (
);

DFFSR _8309_ (
    .Q(\datapath_1.regfile_1.regOut[11] [31]),
    .CLK(clk_bF$buf47),
    .R(rst_bF$buf53),
    .S(vdd),
    .D(_653_[31])
);

FILL FILL_1__7686_ (
);

FILL FILL_2__14876_ (
);

FILL SFILL69080x30050 (
);

FILL FILL_2__14456_ (
);

FILL FILL_2__14036_ (
);

FILL FILL_0__15490_ (
);

FILL FILL_0__15070_ (
);

FILL SFILL48920x15050 (
);

FILL FILL_1__13869_ (
);

FILL FILL_1__13449_ (
);

FILL FILL_1__13029_ (
);

FILL FILL_3__8973_ (
);

OAI21X1 _12727_ (
    .A(_3509_),
    .B(IRWrite_bF$buf1),
    .C(_3510_),
    .Y(_3490_[10])
);

FILL FILL_3__8133_ (
);

NAND3X1 _12307_ (
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3269_)
);

FILL FILL_5__8899_ (
);

FILL FILL_1__14810_ (
);

FILL FILL_5__8479_ (
);

FILL FILL_5__8059_ (
);

INVX1 _15199_ (
    .A(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_5676_)
);

FILL FILL_4__12390_ (
);

FILL FILL_0__13803_ (
);

FILL FILL_3__16248_ (
);

FILL FILL_2__6970_ (
);

FILL FILL_5__10769_ (
);

FILL FILL_5__9420_ (
);

FILL FILL_3__11383_ (
);

FILL FILL_5__9000_ (
);

FILL SFILL59080x73050 (
);

FILL FILL_4__6896_ (
);

FILL FILL_0__16275_ (
);

NOR2X1 _16140_ (
    .A(_6584_),
    .B(_6592_),
    .Y(_6593_)
);

FILL FILL_2__10796_ (
);

FILL FILL_2__10376_ (
);

FILL FILL_5__11710_ (
);

FILL FILL_1__9412_ (
);

FILL FILL_3__9758_ (
);

FILL FILL_3__9338_ (
);

FILL FILL_4__10703_ (
);

FILL SFILL3640x50050 (
);

FILL FILL_5__14182_ (
);

OAI21X1 _8482_ (
    .A(_810_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .C(_811_),
    .Y(_783_[14])
);

FILL FILL_6__7343_ (
);

OAI21X1 _8062_ (
    .A(_591_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_592_),
    .Y(_588_[2])
);

FILL FILL_4__13595_ (
);

FILL FILL_1__10310_ (
);

FILL FILL_2__7755_ (
);

FILL FILL_3__12588_ (
);

FILL FILL_2__7335_ (
);

FILL FILL_3__12168_ (
);

FILL SFILL59000x71050 (
);

OAI21X1 _12480_ (
    .A(_3385_),
    .B(vdd),
    .C(_3386_),
    .Y(_3360_[13])
);

FILL FILL_0__12195_ (
);

NAND3X1 _12060_ (
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [18]),
    .C(_3034__bF$buf4),
    .Y(_3091_)
);

FILL FILL_5__12915_ (
);

FILL FILL_4__8622_ (
);

FILL FILL_4__11908_ (
);

FILL FILL_4__8202_ (
);

FILL FILL_5_BUFX2_insert710 (
);

FILL FILL_5_BUFX2_insert711 (
);

FILL FILL_5__15387_ (
);

FILL FILL_5_BUFX2_insert712 (
);

FILL FILL_2__12522_ (
);

FILL FILL_2__12102_ (
);

FILL FILL_5_BUFX2_insert713 (
);

FILL FILL_5_BUFX2_insert714 (
);

DFFSR _9687_ (
    .Q(\datapath_1.regfile_1.regOut[22] [1]),
    .CLK(clk_bF$buf94),
    .R(rst_bF$buf94),
    .S(vdd),
    .D(_1368_[1])
);

FILL FILL_6__8128_ (
);

FILL FILL_5_BUFX2_insert715 (
);

NAND2X1 _9267_ (
    .A(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1213_)
);

FILL FILL_1_CLKBUF1_insert190 (
);

FILL FILL_5_BUFX2_insert716 (
);

FILL FILL_1_CLKBUF1_insert191 (
);

FILL FILL_5_BUFX2_insert717 (
);

FILL FILL_1_CLKBUF1_insert192 (
);

FILL FILL_1__11935_ (
);

FILL FILL_5_BUFX2_insert718 (
);

FILL FILL_1_CLKBUF1_insert193 (
);

FILL FILL_5_BUFX2_insert719 (
);

FILL FILL_1__11515_ (
);

FILL FILL_1_CLKBUF1_insert194 (
);

FILL FILL_1_CLKBUF1_insert195 (
);

FILL FILL_1_CLKBUF1_insert196 (
);

FILL SFILL104040x60050 (
);

FILL FILL_1_CLKBUF1_insert197 (
);

FILL FILL_1_CLKBUF1_insert198 (
);

FILL FILL_0__10928_ (
);

FILL FILL_1_CLKBUF1_insert199 (
);

FILL FILL_0__8522_ (
);

FILL FILL_0__10508_ (
);

FILL FILL_0__8102_ (
);

FILL FILL_5__6965_ (
);

FILL FILL_6__14707_ (
);

FILL FILL_4__15741_ (
);

FILL FILL_4__15321_ (
);

FILL FILL_3__9091_ (
);

NOR2X1 _13685_ (
    .A(_4182_),
    .B(_4192_),
    .Y(_4193_)
);

NOR2X1 _13265_ (
    .A(_3781_),
    .B(_3807_),
    .Y(\datapath_1.regfile_1.regEn [1])
);

FILL FILL_2__9901_ (
);

FILL FILL_3__14734_ (
);

FILL FILL_3__14314_ (
);

FILL SFILL3560x12050 (
);

FILL FILL_1__6957_ (
);

FILL FILL_4__9407_ (
);

FILL FILL_2__13727_ (
);

FILL FILL_2__13307_ (
);

FILL FILL_0__14761_ (
);

FILL FILL_0__14341_ (
);

FILL FILL_2__16199_ (
);

FILL FILL_0__9727_ (
);

FILL FILL_3__7824_ (
);

FILL FILL_2_BUFX2_insert840 (
);

FILL FILL_4__16106_ (
);

FILL FILL_2_BUFX2_insert841 (
);

FILL FILL_2_BUFX2_insert842 (
);

FILL FILL_2_BUFX2_insert843 (
);

FILL FILL_2_BUFX2_insert844 (
);

FILL FILL_4__11661_ (
);

FILL FILL_4__11241_ (
);

FILL FILL_2_BUFX2_insert845 (
);

FILL FILL_3__15939_ (
);

FILL FILL_2_BUFX2_insert846 (
);

FILL FILL_3__15519_ (
);

FILL FILL_2_BUFX2_insert847 (
);

FILL FILL_2_BUFX2_insert848 (
);

FILL FILL_2_BUFX2_insert849 (
);

FILL FILL_1__16133_ (
);

FILL FILL_3__10654_ (
);

FILL FILL_3__10234_ (
);

FILL SFILL12840x64050 (
);

FILL SFILL28920x11050 (
);

FILL FILL_0__15966_ (
);

FILL FILL_0__15546_ (
);

INVX1 _15831_ (
    .A(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_6292_)
);

NOR2X1 _15411_ (
    .A(_5879_),
    .B(_5882_),
    .Y(_5883_)
);

FILL FILL_0__15126_ (
);

FILL FILL_0__10681_ (
);

FILL FILL_0__10261_ (
);

FILL FILL_3__8609_ (
);

FILL FILL_5__13873_ (
);

FILL FILL_5__13453_ (
);

FILL FILL_5__13033_ (
);

OAI21X1 _7753_ (
    .A(_446_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .C(_447_),
    .Y(_393_[27])
);

OAI21X1 _7333_ (
    .A(_227_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_228_),
    .Y(_198_[15])
);

FILL SFILL79560x79050 (
);

FILL SFILL28840x18050 (
);

FILL FILL_4__12866_ (
);

FILL FILL_4__9160_ (
);

FILL FILL_4__12446_ (
);

FILL FILL_4__12026_ (
);

FILL FILL_2__13480_ (
);

FILL FILL_3__11859_ (
);

FILL FILL_1__12893_ (
);

FILL FILL_3__11439_ (
);

FILL FILL_1__12473_ (
);

FILL FILL_3__11019_ (
);

FILL FILL_1__12053_ (
);

FILL FILL_0__11886_ (
);

FILL FILL_0__9480_ (
);

FILL FILL_2__9498_ (
);

FILL SFILL79160x65050 (
);

FILL FILL_2__9078_ (
);

FILL FILL_0__11466_ (
);

OAI21X1 _11751_ (
    .A(_2376_),
    .B(_2503_),
    .C(_2470__bF$buf1),
    .Y(_2847_)
);

FILL FILL_0__11046_ (
);

OAI21X1 _11331_ (
    .A(_2437_),
    .B(_2445_),
    .C(_2449_),
    .Y(_2450_)
);

FILL FILL_6__15245_ (
);

FILL FILL_5__7083_ (
);

FILL FILL_5__14658_ (
);

FILL FILL_5__14238_ (
);

FILL FILL_3__15692_ (
);

FILL FILL_3__15272_ (
);

OAI21X1 _8958_ (
    .A(_1046_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .C(_1047_),
    .Y(_1043_[2])
);

DFFSR _8538_ (
    .Q(\datapath_1.regfile_1.regOut[13] [4]),
    .CLK(clk_bF$buf58),
    .R(rst_bF$buf1),
    .S(vdd),
    .D(_783_[4])
);

NAND2X1 _8118_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_630_)
);

FILL FILL_1__7495_ (
);

FILL FILL_1__7075_ (
);

FILL FILL_2__14685_ (
);

FILL FILL_2__14265_ (
);

FILL FILL_1__13678_ (
);

FILL FILL_1__13258_ (
);

FILL FILL_1_BUFX2_insert860 (
);

FILL FILL_3__8782_ (
);

FILL FILL_1_BUFX2_insert861 (
);

FILL FILL_1_BUFX2_insert862 (
);

FILL FILL_3__8362_ (
);

OAI21X1 _12956_ (
    .A(_3621_),
    .B(vdd),
    .C(_3622_),
    .Y(_3620_[1])
);

FILL FILL_1_BUFX2_insert863 (
);

DFFSR _12536_ (
    .Q(ALUOut[1]),
    .CLK(clk_bF$buf81),
    .R(rst_bF$buf65),
    .S(vdd),
    .D(_3360_[1])
);

FILL FILL_1_BUFX2_insert864 (
);

NAND2X1 _12116_ (
    .A(\datapath_1.a [0]),
    .B(ALUSrcA_bF$buf2),
    .Y(_3195_)
);

FILL FILL_1_BUFX2_insert865 (
);

FILL FILL_1_BUFX2_insert866 (
);

FILL FILL_1_BUFX2_insert867 (
);

FILL FILL_1_BUFX2_insert868 (
);

FILL FILL_1_BUFX2_insert869 (
);

FILL FILL_6__11165_ (
);

FILL FILL_0__13612_ (
);

FILL FILL_3__16057_ (
);

FILL FILL_5__10998_ (
);

FILL FILL_5__10578_ (
);

FILL FILL_5__10158_ (
);

FILL FILL_3__11192_ (
);

FILL FILL_0__16084_ (
);

FILL SFILL84360x83050 (
);

FILL FILL_2__10185_ (
);

FILL FILL_1__9641_ (
);

FILL FILL_1__9221_ (
);

FILL FILL_3__9987_ (
);

FILL FILL_2__16411_ (
);

FILL FILL_3__9147_ (
);

FILL FILL_4__10932_ (
);

FILL FILL_4__10512_ (
);

FILL FILL_1__15824_ (
);

FILL FILL_1__15404_ (
);

DFFSR _8291_ (
    .Q(\datapath_1.regfile_1.regOut[11] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_653_[13])
);

FILL FILL_0__14817_ (
);

FILL FILL111880x3050 (
);

FILL FILL_2__7984_ (
);

FILL FILL_2__7564_ (
);

BUFX2 BUFX2_insert530 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf77)
);

FILL FILL_3__12397_ (
);

BUFX2 BUFX2_insert531 (
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf76)
);

BUFX2 BUFX2_insert532 (
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf75)
);

BUFX2 BUFX2_insert533 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf74)
);

BUFX2 BUFX2_insert534 (
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf73)
);

BUFX2 BUFX2_insert535 (
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf72)
);

FILL FILL_6__13311_ (
);

BUFX2 BUFX2_insert536 (
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf71)
);

BUFX2 BUFX2_insert537 (
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf70)
);

BUFX2 BUFX2_insert538 (
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf69)
);

BUFX2 BUFX2_insert539 (
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf68)
);

FILL FILL_5__12724_ (
);

FILL FILL_5__12304_ (
);

FILL FILL_4__8851_ (
);

FILL FILL_4__8011_ (
);

FILL FILL_4__11717_ (
);

FILL FILL_2__12751_ (
);

FILL FILL_5__15196_ (
);

FILL FILL_2__12331_ (
);

NAND2X1 _9496_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1325_)
);

DFFSR _9076_ (
    .Q(\datapath_1.regfile_1.regOut[17] [30]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_1043_[30])
);

FILL FILL_1__11744_ (
);

FILL FILL_4__14189_ (
);

FILL FILL_1__11324_ (
);

FILL FILL_0__8751_ (
);

FILL FILL_2__8769_ (
);

FILL FILL_0__8331_ (
);

FILL FILL_2__8349_ (
);

FILL SFILL114520x64050 (
);

FILL FILL_0__10317_ (
);

DFFSR _10602_ (
    .Q(\datapath_1.regfile_1.regOut[29] [20]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf93),
    .S(vdd),
    .D(_1823_[20])
);

FILL FILL_0_BUFX2_insert50 (
);

FILL FILL_0_BUFX2_insert51 (
);

FILL FILL_4__15970_ (
);

FILL FILL_0_BUFX2_insert52 (
);

FILL FILL_0_BUFX2_insert53 (
);

FILL FILL_4__15550_ (
);

FILL FILL_0_BUFX2_insert54 (
);

FILL FILL_4__15130_ (
);

FILL SFILL3720x83050 (
);

FILL FILL_0_BUFX2_insert55 (
);

FILL FILL_0_BUFX2_insert56 (
);

FILL FILL_0_BUFX2_insert57 (
);

INVX8 _13494_ (
    .A(_3910_),
    .Y(_4005_)
);

DFFSR _13074_ (
    .Q(_2_[27]),
    .CLK(clk_bF$buf100),
    .R(rst_bF$buf112),
    .S(vdd),
    .D(_3620_[27])
);

FILL FILL_5__13929_ (
);

FILL FILL_0_BUFX2_insert58 (
);

FILL FILL_0_BUFX2_insert59 (
);

FILL FILL_3__14963_ (
);

FILL FILL_5__13509_ (
);

FILL FILL_3__14543_ (
);

OAI21X1 _7809_ (
    .A(_463_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .C(_464_),
    .Y(_458_[3])
);

FILL FILL_3__14123_ (
);

FILL FILL_4_BUFX2_insert370 (
);

FILL FILL_4__9636_ (
);

FILL FILL_4_BUFX2_insert371 (
);

FILL FILL_4_BUFX2_insert372 (
);

FILL FILL_4__9216_ (
);

FILL SFILL69080x25050 (
);

FILL FILL_4_BUFX2_insert373 (
);

FILL FILL_2__13956_ (
);

FILL FILL_0__14990_ (
);

FILL FILL_4_BUFX2_insert374 (
);

FILL FILL_2__13536_ (
);

FILL FILL_0__14570_ (
);

FILL FILL_2__13116_ (
);

FILL FILL_4_BUFX2_insert375 (
);

FILL FILL_0__14150_ (
);

FILL FILL_4_BUFX2_insert376 (
);

FILL FILL_4_BUFX2_insert377 (
);

FILL FILL_4_BUFX2_insert378 (
);

FILL FILL_4_BUFX2_insert379 (
);

FILL FILL_1__12529_ (
);

FILL FILL_1__12109_ (
);

FILL FILL_0__9536_ (
);

FILL FILL_3__7633_ (
);

FILL FILL_0__9116_ (
);

FILL FILL_3__7213_ (
);

OAI21X1 _11807_ (
    .A(_2368_),
    .B(_2363_),
    .C(_2898_),
    .Y(_2899_)
);

FILL FILL_5__7979_ (
);

FILL FILL_5__7559_ (
);

FILL FILL_4__16335_ (
);

FILL FILL_4__11890_ (
);

INVX1 _14699_ (
    .A(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_5185_)
);

FILL FILL_6__10016_ (
);

INVX1 _14279_ (
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_4774_)
);

FILL FILL_4__11470_ (
);

FILL FILL_4__11050_ (
);

FILL FILL_3__15748_ (
);

FILL FILL_3__15328_ (
);

FILL FILL_1__16362_ (
);

FILL FILL_3__10883_ (
);

FILL FILL_5__8500_ (
);

FILL FILL_3__10043_ (
);

FILL SFILL59080x68050 (
);

FILL FILL_0__15775_ (
);

FILL FILL_0__15355_ (
);

NOR2X1 _15640_ (
    .A(_6103_),
    .B(_6105_),
    .Y(_6106_)
);

NAND2X1 _15220_ (
    .A(\datapath_1.PCJump [23]),
    .B(_5475_),
    .Y(_5696_)
);

FILL FILL_0__10490_ (
);

FILL FILL_1__8912_ (
);

FILL SFILL83560x79050 (
);

FILL FILL_3__8838_ (
);

FILL SFILL3640x45050 (
);

FILL FILL_5__13682_ (
);

FILL FILL_5__13262_ (
);

OAI21X1 _7982_ (
    .A(_558_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .C(_559_),
    .Y(_523_[18])
);

OAI21X1 _7562_ (
    .A(_339_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .C(_340_),
    .Y(_328_[6])
);

DFFSR _7142_ (
    .Q(\datapath_1.regfile_1.regOut[2] [16]),
    .CLK(clk_bF$buf93),
    .R(rst_bF$buf51),
    .S(vdd),
    .D(_68_[16])
);

FILL SFILL43880x52050 (
);

FILL FILL_4__12255_ (
);

DFFSR _10199_ (
    .Q(\datapath_1.regfile_1.regOut[26] [1]),
    .CLK(clk_bF$buf65),
    .R(rst_bF$buf52),
    .S(vdd),
    .D(_1628_[1])
);

FILL FILL_3__11668_ (
);

FILL FILL_3__11248_ (
);

FILL SFILL59000x66050 (
);

FILL FILL_1__12282_ (
);

DFFSR _16425_ (
    .Q(\datapath_1.regfile_1.regOut[0] [8]),
    .CLK(clk_bF$buf112),
    .R(rst_bF$buf40),
    .S(vdd),
    .D(_6769_[8])
);

NOR3X1 _16005_ (
    .A(_6461_),
    .B(_6442_),
    .C(_6451_),
    .Y(_6462_)
);

FILL SFILL59080x23050 (
);

INVX1 _11980_ (
    .A(\datapath_1.PCJump [31]),
    .Y(_3028_)
);

FILL FILL_0__11695_ (
);

INVX1 _11560_ (
    .A(_2235_),
    .Y(_2669_)
);

FILL FILL_0__11275_ (
);

NOR2X1 _11140_ (
    .A(_2258_),
    .B(_2249_),
    .Y(_2259_)
);

FILL FILL_6__15894_ (
);

FILL SFILL104440x69050 (
);

FILL FILL_3_BUFX2_insert390 (
);

FILL FILL_4__7702_ (
);

FILL FILL_3_BUFX2_insert391 (
);

FILL FILL_3_BUFX2_insert392 (
);

FILL FILL_5__14887_ (
);

FILL FILL_5__14467_ (
);

FILL FILL_3_BUFX2_insert393 (
);

FILL FILL_2__11602_ (
);

FILL FILL_5__14047_ (
);

FILL FILL_3_BUFX2_insert394 (
);

NAND2X1 _8767_ (
    .A(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_961_)
);

FILL FILL_3__15081_ (
);

FILL FILL_3_BUFX2_insert395 (
);

FILL FILL_3_BUFX2_insert396 (
);

FILL FILL_6__7208_ (
);

NAND2X1 _8347_ (
    .A(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_742_)
);

FILL FILL_3_BUFX2_insert397 (
);

FILL FILL_3_BUFX2_insert398 (
);

FILL FILL_3_BUFX2_insert399 (
);

FILL FILL_2__14494_ (
);

FILL FILL_2__14074_ (
);

FILL FILL_0__7602_ (
);

FILL FILL_1__13487_ (
);

FILL FILL_4__14821_ (
);

FILL FILL_4__14401_ (
);

FILL SFILL59000x21050 (
);

FILL FILL_3__8591_ (
);

FILL SFILL49080x66050 (
);

NAND2X1 _12765_ (
    .A(IRWrite_bF$buf7),
    .B(memoryOutData[23]),
    .Y(_3536_)
);

OAI21X1 _12345_ (
    .A(_3358_),
    .B(MemToReg_bF$buf5),
    .C(_3359_),
    .Y(\datapath_1.mux_wd3.dout [0])
);

FILL FILL_3__13814_ (
);

FILL FILL_5__8097_ (
);

FILL FILL_4__8907_ (
);

FILL SFILL73560x77050 (
);

FILL SFILL104440x24050 (
);

FILL FILL_0__13841_ (
);

FILL FILL_0__13421_ (
);

FILL FILL_3__16286_ (
);

FILL FILL_0__13001_ (
);

FILL FILL_5__10387_ (
);

FILL FILL_1__8089_ (
);

FILL FILL_2__15699_ (
);

FILL FILL_2__15279_ (
);

FILL FILL_3__6904_ (
);

FILL FILL_1__9870_ (
);

FILL FILL_1__9030_ (
);

FILL FILL_4__15606_ (
);

FILL FILL_2__16220_ (
);

FILL FILL_3__9796_ (
);

FILL FILL_3__9376_ (
);

FILL SFILL113720x15050 (
);

FILL FILL_4__10321_ (
);

FILL FILL_1__15633_ (
);

FILL SFILL49080x21050 (
);

FILL FILL_1__15213_ (
);

FILL SFILL94440x73050 (
);

FILL FILL_0__14626_ (
);

INVX1 _14911_ (
    .A(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_5393_)
);

FILL FILL_0__14206_ (
);

FILL FILL_2__7373_ (
);

FILL FILL_4__7299_ (
);

FILL FILL_6__13120_ (
);

FILL FILL_2__11199_ (
);

FILL FILL_5__12953_ (
);

FILL FILL_5__12533_ (
);

FILL FILL_5__12113_ (
);

FILL FILL_4__8660_ (
);

FILL FILL_4__11946_ (
);

FILL FILL_4__8240_ (
);

FILL FILL_2__12980_ (
);

FILL FILL_4__11526_ (
);

FILL FILL_4__11106_ (
);

FILL FILL_2__12140_ (
);

FILL FILL_0__7199_ (
);

FILL FILL_3__10939_ (
);

FILL FILL_1__11973_ (
);

FILL FILL_3__10519_ (
);

FILL FILL_1__11553_ (
);

FILL FILL_1__11133_ (
);

FILL FILL_2__8998_ (
);

FILL FILL_0__8980_ (
);

FILL FILL_0__10966_ (
);

FILL FILL_2__8578_ (
);

OAI21X1 _10831_ (
    .A(_2010_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_2011_),
    .Y(_1953_[29])
);

FILL FILL_0__8140_ (
);

FILL FILL_0__10546_ (
);

FILL FILL_0__10126_ (
);

OAI21X1 _10411_ (
    .A(_1791_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1792_),
    .Y(_1758_[17])
);

FILL FILL_5__13738_ (
);

FILL FILL_5__13318_ (
);

FILL FILL_3__14772_ (
);

FILL FILL_3__14352_ (
);

NAND2X1 _7618_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_378_)
);

FILL FILL_1__6995_ (
);

FILL FILL_4__9865_ (
);

FILL FILL_4__9025_ (
);

FILL FILL_2__13765_ (
);

FILL FILL111800x64050 (
);

FILL FILL_2__13345_ (
);

FILL SFILL94360x35050 (
);

FILL FILL_1__12758_ (
);

FILL FILL_1__12338_ (
);

FILL FILL_3__7862_ (
);

FILL FILL_0__9765_ (
);

FILL FILL_0__9345_ (
);

FILL FILL_3__7442_ (
);

OAI21X1 _11616_ (
    .A(_2547_),
    .B(_2548_),
    .C(_2720_),
    .Y(_2721_)
);

FILL SFILL39400x3050 (
);

FILL FILL_5__7368_ (
);

FILL FILL_4__16144_ (
);

OAI22X1 _14088_ (
    .A(_4586_),
    .B(_3941_),
    .C(_3916_),
    .D(_4585_),
    .Y(_4587_)
);

FILL FILL_3__15977_ (
);

FILL FILL_3__15557_ (
);

FILL FILL_3__15137_ (
);

FILL FILL_1__16171_ (
);

FILL FILL_3__10692_ (
);

FILL FILL_3__10272_ (
);

FILL FILL_0__15584_ (
);

FILL FILL_0__15164_ (
);

FILL SFILL84360x78050 (
);

FILL SFILL79160x5050 (
);

FILL FILL_1__8721_ (
);

FILL SFILL53880x1050 (
);

FILL FILL_2__15911_ (
);

FILL FILL_3__8647_ (
);

FILL FILL_3__8227_ (
);

FILL FILL_5__13491_ (
);

FILL FILL_1__14904_ (
);

DFFSR _7791_ (
    .Q(\datapath_1.regfile_1.regOut[7] [25]),
    .CLK(clk_bF$buf111),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_393_[25])
);

NAND2X1 _7371_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_254_)
);

FILL FILL_4__12484_ (
);

FILL FILL_4__12064_ (
);

FILL SFILL8760x52050 (
);

FILL FILL_5__9934_ (
);

FILL FILL_3__11897_ (
);

FILL FILL_5__9514_ (
);

FILL FILL_3__11477_ (
);

FILL FILL_3__11057_ (
);

FILL FILL_1__12091_ (
);

FILL FILL_0__16369_ (
);

INVX1 _16234_ (
    .A(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_6685_)
);

FILL FILL_0__11084_ (
);

FILL SFILL114600x52050 (
);

FILL FILL_1__9926_ (
);

FILL FILL_5__11804_ (
);

FILL FILL_1__9506_ (
);

FILL FILL_4__7931_ (
);

FILL FILL_5__14696_ (
);

FILL FILL_2__11831_ (
);

FILL FILL_5__14276_ (
);

FILL FILL_2__11411_ (
);

NAND2X1 _8996_ (
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1073_)
);

NAND2X1 _8576_ (
    .A(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_854_)
);

DFFSR _8156_ (
    .Q(\datapath_1.regfile_1.regOut[10] [6]),
    .CLK(clk_bF$buf84),
    .R(rst_bF$buf45),
    .S(vdd),
    .D(_588_[6])
);

FILL FILL_1__10824_ (
);

FILL FILL_4__13689_ (
);

FILL FILL_4__13269_ (
);

FILL FILL_1__10404_ (
);

FILL FILL_0__7831_ (
);

FILL FILL_2__7849_ (
);

FILL FILL_2__7429_ (
);

FILL FILL_1__13296_ (
);

FILL FILL_4__14630_ (
);

FILL SFILL3720x78050 (
);

FILL FILL_4__14210_ (
);

NAND2X1 _12994_ (
    .A(vdd),
    .B(\datapath_1.rd2 [14]),
    .Y(_3648_)
);

NAND2X1 _12574_ (
    .A(vdd),
    .B(memoryOutData[2]),
    .Y(_3429_)
);

FILL FILL_0__12289_ (
);

INVX1 _12154_ (
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_3156_)
);

FILL FILL_3__13623_ (
);

FILL FILL_6__16068_ (
);

FILL FILL_4__8716_ (
);

FILL SFILL19080x60050 (
);

FILL FILL_2__12616_ (
);

FILL FILL_0__13650_ (
);

FILL FILL_0__13230_ (
);

FILL FILL_3__16095_ (
);

FILL FILL_5__10196_ (
);

FILL FILL_1__11609_ (
);

FILL FILL_2__15088_ (
);

FILL FILL_5__16002_ (
);

FILL FILL_0__8616_ (
);

FILL FILL_4__15835_ (
);

FILL FILL_4__15415_ (
);

FILL FILL_4__10970_ (
);

NOR2X1 _13779_ (
    .A(_4281_),
    .B(_4284_),
    .Y(_4285_)
);

FILL FILL_4__10550_ (
);

INVX1 _13359_ (
    .A(_3767_),
    .Y(_3875_)
);

FILL FILL_4__10130_ (
);

FILL SFILL3720x33050 (
);

FILL FILL_3__14828_ (
);

FILL FILL_3__14408_ (
);

FILL FILL_1__15862_ (
);

FILL FILL_1__15442_ (
);

FILL FILL_1__15022_ (
);

FILL SFILL38600x27050 (
);

FILL SFILL43960x40050 (
);

FILL FILL_0__14855_ (
);

INVX1 _14720_ (
    .A(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_5206_)
);

FILL FILL_0__14435_ (
);

FILL FILL_0__14015_ (
);

INVX1 _14300_ (
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_4795_)
);

BUFX2 BUFX2_insert910 (
    .A(IRWrite),
    .Y(IRWrite_bF$buf0)
);

FILL FILL_2__7182_ (
);

BUFX2 BUFX2_insert911 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf4 )
);

BUFX2 BUFX2_insert912 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf3 )
);

BUFX2 BUFX2_insert913 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf2 )
);

FILL SFILL49560x5050 (
);

BUFX2 BUFX2_insert914 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf1 )
);

BUFX2 BUFX2_insert915 (
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf0 )
);

BUFX2 BUFX2_insert916 (
    .A(_5549_),
    .Y(_5549__bF$buf4)
);

BUFX2 BUFX2_insert917 (
    .A(_5549_),
    .Y(_5549__bF$buf3)
);

BUFX2 BUFX2_insert918 (
    .A(_5549_),
    .Y(_5549__bF$buf2)
);

BUFX2 BUFX2_insert919 (
    .A(_5549_),
    .Y(_5549__bF$buf1)
);

FILL FILL_5__12762_ (
);

FILL FILL_5__12342_ (
);

FILL SFILL104520x57050 (
);

FILL SFILL43880x47050 (
);

FILL SFILL48920x2050 (
);

FILL FILL_4__11755_ (
);

FILL FILL_4__11335_ (
);

FILL FILL_1__16227_ (
);

FILL FILL_3__10748_ (
);

FILL FILL_1__11782_ (
);

FILL FILL_1__11362_ (
);

FILL SFILL108840x65050 (
);

OAI22X1 _15925_ (
    .A(_5463__bF$buf3),
    .B(_4943_),
    .C(_4942_),
    .D(_5504__bF$buf1),
    .Y(_6384_)
);

INVX1 _15505_ (
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_5974_)
);

FILL SFILL59080x18050 (
);

FILL FILL112280x51050 (
);

FILL FILL_0__10775_ (
);

FILL FILL_2__8387_ (
);

OAI21X1 _10640_ (
    .A(_1903_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .C(_1904_),
    .Y(_1888_[8])
);

DFFSR _10220_ (
    .Q(\datapath_1.regfile_1.regOut[26] [22]),
    .CLK(clk_bF$buf88),
    .R(rst_bF$buf14),
    .S(vdd),
    .D(_1628_[22])
);

FILL FILL_6__14554_ (
);

FILL FILL_6__14134_ (
);

FILL FILL_5__13967_ (
);

FILL FILL_5__13547_ (
);

FILL FILL_3__14581_ (
);

FILL FILL_5__13127_ (
);

NAND2X1 _7847_ (
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_490_)
);

FILL FILL_3__14161_ (
);

NAND2X1 _7427_ (
    .A(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_271_)
);

FILL FILL_4_BUFX2_insert750 (
);

DFFSR _7007_ (
    .Q(\datapath_1.regfile_1.regOut[1] [9]),
    .CLK(clk_bF$buf20),
    .R(rst_bF$buf5),
    .S(vdd),
    .D(_3_[9])
);

FILL FILL_4_BUFX2_insert751 (
);

FILL FILL_4__9674_ (
);

FILL FILL_4_BUFX2_insert752 (
);

FILL FILL_4__9254_ (
);

FILL FILL_2__13994_ (
);

FILL FILL_4_BUFX2_insert753 (
);

FILL FILL_4_BUFX2_insert754 (
);

FILL FILL_2__13574_ (
);

FILL SFILL104520x12050 (
);

FILL FILL_2__13154_ (
);

FILL FILL_4_BUFX2_insert755 (
);

FILL FILL_4_BUFX2_insert756 (
);

FILL FILL_4_BUFX2_insert757 (
);

FILL FILL_4_BUFX2_insert758 (
);

FILL FILL_4_BUFX2_insert759 (
);

FILL FILL_1__12987_ (
);

FILL FILL_1__12567_ (
);

FILL FILL_1__12147_ (
);

FILL FILL_4__13901_ (
);

FILL SFILL59000x16050 (
);

FILL FILL_0__9994_ (
);

FILL FILL_3__7671_ (
);

FILL FILL_3__7251_ (
);

OAI21X1 _11845_ (
    .A(_2926_),
    .B(_2930_),
    .C(_2932_),
    .Y(_2933_)
);

FILL FILL_0__9154_ (
);

NAND2X1 _11425_ (
    .A(_2132_),
    .B(_2133_),
    .Y(_2541_)
);

NAND2X1 _11005_ (
    .A(_2122_),
    .B(_2123_),
    .Y(_2124_)
);

FILL FILL_5__7597_ (
);

FILL FILL_5__7177_ (
);

FILL FILL_4__16373_ (
);

FILL FILL_6__10894_ (
);

FILL FILL_3__15786_ (
);

FILL FILL_3__15366_ (
);

FILL FILL_0__12501_ (
);

FILL FILL_1__7589_ (
);

FILL FILL_1__7169_ (
);

FILL FILL_2__14779_ (
);

FILL FILL_2__14359_ (
);

FILL FILL_0__15393_ (
);

FILL SFILL33880x45050 (
);

FILL FILL_1__8950_ (
);

FILL FILL_1__8530_ (
);

FILL FILL_1__8110_ (
);

FILL FILL_2__15720_ (
);

FILL FILL_2__15300_ (
);

FILL FILL_3__8876_ (
);

FILL FILL_3__8456_ (
);

FILL SFILL49080x16050 (
);

FILL FILL_1__14713_ (
);

NAND2X1 _7180_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_147_)
);

FILL SFILL94440x68050 (
);

FILL FILL_4__12293_ (
);

FILL FILL_0__13706_ (
);

FILL FILL_2__6873_ (
);

FILL FILL_5__9743_ (
);

FILL FILL_3__11286_ (
);

FILL SFILL49400x28050 (
);

FILL FILL_0__16178_ (
);

NOR2X1 _16043_ (
    .A(_6497_),
    .B(_6498_),
    .Y(_6499_)
);

FILL FILL_2__10699_ (
);

FILL FILL_2__10279_ (
);

FILL FILL_5__11613_ (
);

FILL FILL_1__9735_ (
);

FILL FILL_4__7740_ (
);

FILL FILL_3_BUFX2_insert770 (
);

FILL FILL_4__7320_ (
);

FILL FILL_3_BUFX2_insert771 (
);

FILL FILL_3_BUFX2_insert772 (
);

FILL FILL_3_BUFX2_insert773 (
);

FILL FILL_2__11640_ (
);

FILL SFILL18600x23050 (
);

FILL FILL_3_BUFX2_insert774 (
);

FILL FILL_2__11220_ (
);

FILL FILL_5__14085_ (
);

FILL SFILL49000x14050 (
);

FILL FILL_1__15918_ (
);

FILL FILL_3_BUFX2_insert775 (
);

FILL FILL_3_BUFX2_insert776 (
);

INVX1 _8385_ (
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_767_)
);

FILL FILL_3_BUFX2_insert777 (
);

FILL FILL_3_BUFX2_insert778 (
);

FILL FILL_3_BUFX2_insert779 (
);

FILL FILL_1__10633_ (
);

FILL FILL_4__13498_ (
);

FILL FILL_2__7238_ (
);

FILL FILL_0__7220_ (
);

FILL SFILL18840x6050 (
);

NAND2X1 _12383_ (
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [13]),
    .Y(_3321_)
);

FILL FILL_0__12098_ (
);

FILL FILL_3__13852_ (
);

FILL SFILL54280x34050 (
);

FILL FILL_3__13432_ (
);

FILL FILL_3__13012_ (
);

FILL FILL_4__8525_ (
);

FILL FILL_4__8105_ (
);

FILL FILL_2__12845_ (
);

FILL FILL_2__12425_ (
);

FILL FILL_2__12005_ (
);

FILL SFILL23400x72050 (
);

FILL SFILL39000x57050 (
);

FILL FILL_1__11838_ (
);

FILL FILL_1__11418_ (
);

FILL FILL_0__8845_ (
);

FILL FILL_5__16231_ (
);

FILL FILL_3__6942_ (
);

FILL FILL_0__8005_ (
);

FILL FILL_5__6868_ (
);

FILL FILL_4__15644_ (
);

FILL FILL_4__15224_ (
);

INVX1 _13588_ (
    .A(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_4097_)
);

OAI21X1 _13168_ (
    .A(_3742_),
    .B(PCEn_bF$buf6),
    .C(_3743_),
    .Y(_3685_[29])
);

FILL SFILL23800x41050 (
);

FILL FILL_2__9804_ (
);

FILL FILL_3__14637_ (
);

FILL FILL_1__15671_ (
);

FILL FILL_3__14217_ (
);

FILL SFILL88760x74050 (
);

FILL FILL_1__15251_ (
);

FILL FILL_0__14664_ (
);

FILL FILL_0__14244_ (
);

FILL SFILL84840x35050 (
);

FILL FILL111800x14050 (
);

FILL SFILL39000x12050 (
);

FILL FILL_1__7801_ (
);

FILL FILL_3__7727_ (
);

FILL FILL_3__7307_ (
);

FILL FILL_5__12991_ (
);

FILL FILL_5__12571_ (
);

FILL FILL_5__12151_ (
);

BUFX2 _6871_ (
    .A(_2_[1]),
    .Y(memoryWriteData[1])
);

FILL FILL_4__16009_ (
);

FILL FILL_4__11984_ (
);

FILL FILL_4__11564_ (
);

FILL SFILL8760x47050 (
);

FILL FILL_4__11144_ (
);

FILL FILL_1__16036_ (
);

FILL FILL_3__10977_ (
);

FILL FILL_3__10557_ (
);

FILL FILL_6_BUFX2_insert280 (
);

FILL FILL_3__10137_ (
);

FILL FILL_1__11591_ (
);

FILL FILL_1__11171_ (
);

FILL FILL_0__15869_ (
);

NAND2X1 _15734_ (
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .B(_5560_),
    .Y(_6197_)
);

FILL FILL_0__15449_ (
);

INVX1 _15314_ (
    .A(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_5788_)
);

FILL FILL_0__15029_ (
);

FILL FILL_6_BUFX2_insert285 (
);

FILL FILL_2__8196_ (
);

FILL FILL_0__10164_ (
);

FILL SFILL53960x37050 (
);

FILL SFILL84360x28050 (
);

BUFX2 BUFX2_insert60 (
    .A(_5463_),
    .Y(_5463__bF$buf2)
);

BUFX2 BUFX2_insert61 (
    .A(_5463_),
    .Y(_5463__bF$buf1)
);

BUFX2 BUFX2_insert62 (
    .A(_5463_),
    .Y(_5463__bF$buf0)
);

BUFX2 BUFX2_insert63 (
    .A(_3200_),
    .Y(_3200__bF$buf4)
);

BUFX2 BUFX2_insert64 (
    .A(_3200_),
    .Y(_3200__bF$buf3)
);

BUFX2 BUFX2_insert65 (
    .A(_3200_),
    .Y(_3200__bF$buf2)
);

BUFX2 BUFX2_insert66 (
    .A(_3200_),
    .Y(_3200__bF$buf1)
);

FILL FILL_2__10911_ (
);

FILL FILL_5__13776_ (
);

BUFX2 BUFX2_insert67 (
    .A(_3200_),
    .Y(_3200__bF$buf0)
);

FILL FILL_5__13356_ (
);

BUFX2 BUFX2_insert68 (
    .A(_3905_),
    .Y(_3905__bF$buf3)
);

BUFX2 BUFX2_insert69 (
    .A(_3905_),
    .Y(_3905__bF$buf2)
);

FILL FILL_3__14390_ (
);

DFFSR _7656_ (
    .Q(\datapath_1.regfile_1.regOut[6] [18]),
    .CLK(clk_bF$buf89),
    .R(rst_bF$buf111),
    .S(vdd),
    .D(_328_[18])
);

INVX1 _7236_ (
    .A(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_184_)
);

FILL FILL_4__9483_ (
);

FILL SFILL88680x36050 (
);

FILL FILL_4__12769_ (
);

FILL FILL_4__12349_ (
);

FILL FILL_2__13383_ (
);

FILL FILL_0__6911_ (
);

FILL FILL_2__6929_ (
);

FILL FILL_1__12376_ (
);

FILL FILL_4__13710_ (
);

FILL FILL_0__9383_ (
);

FILL FILL_3__7480_ (
);

FILL FILL_0__11789_ (
);

FILL FILL_0__11369_ (
);

FILL FILL_3__7060_ (
);

OAI21X1 _11654_ (
    .A(_2376_),
    .B(_2755_),
    .C(_2756_),
    .Y(_2757_)
);

NOR2X1 _11234_ (
    .A(_2352_),
    .B(_2351_),
    .Y(_2353_)
);

FILL FILL_3__12703_ (
);

FILL FILL_4__16182_ (
);

FILL FILL_0__12730_ (
);

FILL FILL_3__15595_ (
);

FILL FILL_3__15175_ (
);

FILL FILL_0__12310_ (
);

FILL FILL_2__14588_ (
);

FILL FILL_2__14168_ (
);

FILL FILL_5__15922_ (
);

FILL FILL_5__15502_ (
);

INVX1 _9802_ (
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_1488_)
);

FILL FILL_4__14915_ (
);

INVX1 _12859_ (
    .A(\datapath_1.a [12]),
    .Y(_3578_)
);

FILL FILL_3__8265_ (
);

INVX1 _12439_ (
    .A(ALUOut[0]),
    .Y(_3423_)
);

NAND3X1 _12019_ (
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[8]),
    .C(_3032__bF$buf4),
    .Y(_3060_)
);

FILL FILL_3__13908_ (
);

FILL FILL_1__14942_ (
);

FILL FILL_1__14522_ (
);

FILL FILL_1__14102_ (
);

FILL SFILL43960x35050 (
);

FILL FILL_0__13935_ (
);

NOR2X1 _13800_ (
    .A(_4304_),
    .B(_3910_),
    .Y(_4305_)
);

FILL FILL_0__13515_ (
);

FILL FILL_5_BUFX2_insert1090 (
);

FILL FILL_5__9552_ (
);

FILL FILL_5__9132_ (
);

FILL FILL_5_BUFX2_insert1091 (
);

FILL FILL_3__11095_ (
);

FILL FILL_5_BUFX2_insert1092 (
);

FILL FILL_5_BUFX2_insert1093 (
);

OAI22X1 _16272_ (
    .A(_5381_),
    .B(_5548__bF$buf1),
    .C(_5489__bF$buf0),
    .D(_5395_),
    .Y(_6722_)
);

FILL FILL_5__11842_ (
);

FILL FILL_1__9544_ (
);

FILL FILL_5__11422_ (
);

FILL FILL_1__9124_ (
);

FILL FILL_5__11002_ (
);

FILL FILL_2__16314_ (
);

FILL FILL_4__10835_ (
);

FILL FILL_4__10415_ (
);

FILL FILL_1__15727_ (
);

INVX1 _8194_ (
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_660_)
);

FILL FILL_1__15307_ (
);

FILL FILL_1__10442_ (
);

FILL FILL_1__10022_ (
);

FILL FILL112280x46050 (
);

FILL FILL_2__7887_ (
);

FILL FILL_2__7467_ (
);

FILL FILL_2__7047_ (
);

FILL FILL_6__13214_ (
);

FILL SFILL68680x77050 (
);

OAI21X1 _12192_ (
    .A(_3180_),
    .B(ALUSrcA_bF$buf3),
    .C(_3181_),
    .Y(\datapath_1.alu_1.ALUInA [25])
);

FILL FILL_5__12627_ (
);

FILL FILL_3__13661_ (
);

FILL FILL_5__12207_ (
);

FILL FILL_3__13241_ (
);

NAND2X1 _6927_ (
    .A(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_19_)
);

FILL FILL_4__8754_ (
);

FILL FILL_4__8334_ (
);

FILL FILL_2__12654_ (
);

FILL FILL_2__12234_ (
);

FILL FILL_5__15099_ (
);

OAI21X1 _9399_ (
    .A(_1279_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1280_),
    .Y(_1238_[21])
);

FILL FILL_1__11647_ (
);

FILL FILL_1__11227_ (
);

FILL FILL_0__8654_ (
);

FILL FILL_5__16040_ (
);

OR2X2 _10925_ (
    .A(_2062_),
    .B(_0_),
    .Y(IorD)
);

FILL FILL_0__8234_ (
);

NAND2X1 _10505_ (
    .A(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1835_)
);

FILL FILL_4__15873_ (
);

FILL FILL_4__15453_ (
);

FILL FILL_4__15033_ (
);

NAND3X1 _13397_ (
    .A(_3898_),
    .B(_3883_),
    .C(_3888_),
    .Y(_3909_)
);

FILL FILL_2__9613_ (
);

FILL FILL_3__14866_ (
);

FILL FILL_3__14446_ (
);

FILL FILL_3__14026_ (
);

FILL FILL_1__15480_ (
);

FILL FILL_1__15060_ (
);

FILL FILL_4__9539_ (
);

FILL FILL_4__9119_ (
);

FILL FILL_2__13859_ (
);

FILL FILL_2__13439_ (
);

FILL FILL_0__14893_ (
);

FILL FILL_0__14473_ (
);

FILL FILL_2__13019_ (
);

FILL FILL_0__14053_ (
);

FILL FILL_1__7610_ (
);

FILL FILL_2__14800_ (
);

FILL FILL_0__9859_ (
);

FILL FILL_3__7956_ (
);

FILL FILL_0__9019_ (
);

FILL FILL_3__7116_ (
);

FILL FILL_5__12380_ (
);

FILL SFILL115080x34050 (
);

FILL FILL_4__16238_ (
);

FILL FILL_4__11793_ (
);

FILL FILL_4__11373_ (
);

FILL FILL_1__16265_ (
);

FILL FILL_5__8823_ (
);

FILL FILL_3__10786_ (
);

FILL FILL_5__8403_ (
);

FILL FILL_3__10366_ (
);

FILL FILL_0__15678_ (
);

INVX1 _15963_ (
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_6421_)
);

FILL FILL_0__15258_ (
);

INVX1 _15543_ (
    .A(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_6011_)
);

OAI22X1 _15123_ (
    .A(_5485__bF$buf2),
    .B(_5601_),
    .C(_5483__bF$buf1),
    .D(_4034_),
    .Y(_5602_)
);

FILL FILL_0__10393_ (
);

FILL FILL_5__13585_ (
);

FILL FILL_2__10300_ (
);

FILL FILL_5__13165_ (
);

INVX1 _7885_ (
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_515_)
);

INVX1 _7465_ (
    .A(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_296_)
);

INVX1 _7045_ (
    .A(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_77_)
);

FILL FILL_4__12998_ (
);

FILL FILL_4__9292_ (
);

FILL FILL_4__12578_ (
);

FILL FILL_4__12158_ (
);

FILL SFILL94440x18050 (
);

FILL FILL_5__9608_ (
);

FILL FILL_1__12185_ (
);

NAND2X1 _16328_ (
    .A(gnd),
    .B(gnd),
    .Y(_6773_)
);

OAI21X1 _11883_ (
    .A(_2964_),
    .B(RegDst),
    .C(_2965_),
    .Y(\datapath_1.a3 [3])
);

FILL FILL_0__11598_ (
);

OAI21X1 _11463_ (
    .A(_2261_),
    .B(_2284_),
    .C(_2577_),
    .Y(_2578_)
);

FILL FILL_0__11178_ (
);

XOR2X1 _11043_ (
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2162_)
);

FILL FILL_6__15797_ (
);

FILL FILL_3__12512_ (
);

FILL FILL_4__7605_ (
);

FILL FILL_2__11925_ (
);

FILL FILL_2__11505_ (
);

FILL FILL_1__10918_ (
);

FILL FILL_2__14397_ (
);

FILL FILL_5__15731_ (
);

FILL FILL_5__15311_ (
);

FILL FILL_0__7505_ (
);

INVX1 _9611_ (
    .A(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_1381_)
);

FILL FILL_4__14724_ (
);

FILL FILL_4__14304_ (
);

FILL FILL_3__8494_ (
);

FILL FILL_3__8074_ (
);

DFFSR _12668_ (
    .Q(\datapath_1.Data [5]),
    .CLK(clk_bF$buf98),
    .R(rst_bF$buf41),
    .S(vdd),
    .D(_3425_[5])
);

FILL SFILL23800x36050 (
);

NAND3X1 _12248_ (
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [10]),
    .C(_3198__bF$buf3),
    .Y(_3225_)
);

FILL FILL_3__13717_ (
);

FILL FILL_1__14751_ (
);

FILL FILL_1__14331_ (
);

FILL FILL_0__13744_ (
);

FILL FILL_0__13324_ (
);

FILL FILL_3__16189_ (
);

FILL FILL_5__9781_ (
);

FILL FILL_5__9361_ (
);

FILL SFILL74120x83050 (
);

INVX1 _16081_ (
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_6536_)
);

FILL FILL_5__11651_ (
);

FILL FILL_1__9773_ (
);

FILL FILL_1__9353_ (
);

FILL FILL_5__11231_ (
);

FILL FILL_4__15929_ (
);

FILL FILL_4__15509_ (
);

FILL FILL_2__16123_ (
);

FILL FILL_3__9279_ (
);

FILL FILL_4__10644_ (
);

FILL FILL_1__15956_ (
);

FILL FILL_1__15536_ (
);

FILL FILL_1__15116_ (
);

FILL SFILL74520x52050 (
);

FILL FILL_1__10671_ (
);

FILL FILL_1__10251_ (
);

FILL FILL_0__14949_ (
);

INVX1 _14814_ (
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_5298_)
);

FILL FILL_0__14529_ (
);

FILL FILL_0__14109_ (
);

FILL FILL_2__7696_ (
);

FILL FILL_6__13863_ (
);

FILL FILL_5__12856_ (
);

FILL FILL_5__12436_ (
);

FILL FILL_3__13890_ (
);

FILL FILL_5__12016_ (
);

FILL FILL_3__13470_ (
);

FILL FILL_4__8983_ (
);

FILL FILL_4__8143_ (
);

FILL FILL_4__11849_ (
);

FILL FILL_2__12883_ (
);

FILL FILL_4__11429_ (
);

FILL FILL_2__12463_ (
);

FILL FILL_4__11009_ (
);

FILL FILL_2__12043_ (
);

FILL SFILL13800x34050 (
);

FILL FILL_1__11876_ (
);

FILL FILL_1__11456_ (
);

FILL FILL_1__11036_ (
);

FILL FILL_3__6980_ (
);

FILL FILL_0__8883_ (
);

FILL FILL_0__8463_ (
);

FILL FILL_6__9850_ (
);

DFFSR _10734_ (
    .Q(\datapath_1.regfile_1.regOut[30] [24]),
    .CLK(clk_bF$buf16),
    .R(rst_bF$buf54),
    .S(vdd),
    .D(_1888_[24])
);

FILL FILL_0__10449_ (
);

INVX1 _10314_ (
    .A(\datapath_1.regfile_1.regOut[27] [28]),
    .Y(_1748_)
);

FILL FILL_0__10029_ (
);

FILL FILL_4__15682_ (
);

FILL FILL_4__15262_ (
);

FILL SFILL64120x81050 (
);

FILL FILL_2__9422_ (
);

FILL FILL_0__11810_ (
);

FILL FILL_3__14675_ (
);

FILL FILL_3__14255_ (
);

FILL FILL_2__9002_ (
);

FILL FILL_1__6898_ (
);

FILL FILL_4__9768_ (
);

FILL FILL_4__9348_ (
);

FILL FILL_2__13668_ (
);

FILL FILL_2__13248_ (
);

FILL FILL_0__14282_ (
);

FILL FILL_0__9668_ (
);

FILL FILL_3__7765_ (
);

FILL FILL_0__9248_ (
);

NAND2X1 _11939_ (
    .A(IorD_bF$buf1),
    .B(ALUOut[17]),
    .Y(_3001_)
);

FILL FILL_3__7345_ (
);

OAI21X1 _11519_ (
    .A(_2507_),
    .B(_2518_),
    .C(_2259_),
    .Y(_2630_)
);

FILL FILL_1__13602_ (
);

FILL FILL_4__16047_ (
);

FILL FILL_6__10568_ (
);

FILL FILL_1_BUFX2_insert100 (
);

FILL FILL_4__11182_ (
);

FILL FILL_1_BUFX2_insert101 (
);

FILL FILL_1_BUFX2_insert102 (
);

FILL FILL_1_BUFX2_insert103 (
);

FILL FILL_1_BUFX2_insert104 (
);

FILL FILL_1__16074_ (
);

FILL FILL_1_BUFX2_insert105 (
);

FILL FILL_5__8632_ (
);

FILL FILL_1_BUFX2_insert106 (
);

FILL FILL_3__10175_ (
);

FILL FILL_1_BUFX2_insert107 (
);

FILL FILL_5__8212_ (
);

FILL FILL_1_BUFX2_insert108 (
);

FILL FILL_1_BUFX2_insert109 (
);

AOI22X1 _15772_ (
    .A(_5481_),
    .B(\datapath_1.regfile_1.regOut[30] [18]),
    .C(\datapath_1.regfile_1.regOut[6] [18]),
    .D(_5565__bF$buf2),
    .Y(_6234_)
);

FILL FILL_6_BUFX2_insert664 (
);

FILL FILL_0__15487_ (
);

OAI22X1 _15352_ (
    .A(_4316_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf0),
    .D(_4307_),
    .Y(_5825_)
);

FILL FILL_0__15067_ (
);

FILL FILL112360x34050 (
);

FILL FILL_3__16401_ (
);

FILL FILL_6_BUFX2_insert669 (
);

FILL FILL_5__10922_ (
);

FILL FILL_1__8624_ (
);

FILL FILL_5__10502_ (
);

FILL FILL_1__8204_ (
);

FILL FILL_2__15814_ (
);

FILL SFILL64040x43050 (
);

FILL FILL_5__13394_ (
);

FILL FILL_6__6975_ (
);

INVX1 _7694_ (
    .A(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_408_)
);

FILL FILL_1__14807_ (
);

DFFSR _7274_ (
    .Q(\datapath_1.regfile_1.regOut[3] [20]),
    .CLK(clk_bF$buf99),
    .R(rst_bF$buf8),
    .S(vdd),
    .D(_133_[20])
);

FILL FILL_4__12387_ (
);

FILL FILL_3__9911_ (
);

FILL FILL_2__6967_ (
);

FILL FILL_5__9417_ (
);

OAI22X1 _16137_ (
    .A(_6589_),
    .B(_5503__bF$buf1),
    .C(_5504__bF$buf2),
    .D(_6588_),
    .Y(_6590_)
);

AOI21X1 _11692_ (
    .A(_2165_),
    .B(_2764_),
    .C(_2791_),
    .Y(_2792_)
);

INVX1 _11272_ (
    .A(\datapath_1.alu_1.ALUInB [11]),
    .Y(_2391_)
);

FILL FILL_5__11707_ (
);

FILL FILL_3__12741_ (
);

FILL FILL_1__9409_ (
);

FILL FILL_3__12321_ (
);

FILL FILL_4__7834_ (
);

FILL FILL_4__7414_ (
);

FILL FILL_5__14599_ (
);

FILL FILL_2__11734_ (
);

FILL FILL_5__14179_ (
);

FILL FILL_2__11314_ (
);

OAI21X1 _8899_ (
    .A(_1027_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1028_),
    .Y(_978_[25])
);

OAI21X1 _8479_ (
    .A(_808_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_809_),
    .Y(_783_[13])
);

OAI21X1 _8059_ (
    .A(_589_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_590_),
    .Y(_588_[1])
);

FILL FILL_1__10307_ (
);

FILL FILL_5__15960_ (
);

FILL FILL_5__15540_ (
);

FILL FILL_0__7734_ (
);

FILL FILL_5__15120_ (
);

DFFSR _9840_ (
    .Q(\datapath_1.regfile_1.regOut[23] [26]),
    .CLK(clk_bF$buf108),
    .R(rst_bF$buf19),
    .S(vdd),
    .D(_1433_[26])
);

FILL FILL_0__7314_ (
);

OAI21X1 _9420_ (
    .A(_1293_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1294_),
    .Y(_1238_[28])
);

OAI21X1 _9000_ (
    .A(_1074_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1075_),
    .Y(_1043_[16])
);

FILL FILL_4__14953_ (
);

FILL FILL_4__14533_ (
);

FILL FILL_4__14113_ (
);

OAI21X1 _12897_ (
    .A(_3602_),
    .B(vdd),
    .C(_3603_),
    .Y(_3555_[24])
);

OAI21X1 _12477_ (
    .A(_3383_),
    .B(vdd),
    .C(_3384_),
    .Y(_3360_[12])
);

AOI22X1 _12057_ (
    .A(\datapath_1.ALUResult [17]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3089_)
);

FILL FILL_3__13946_ (
);

FILL FILL_1__14980_ (
);

FILL FILL_3__13526_ (
);

FILL FILL_1__14560_ (
);

FILL FILL_3__13106_ (
);

FILL FILL_1__14140_ (
);

FILL FILL_4__8619_ (
);

FILL FILL_5_BUFX2_insert680 (
);

FILL FILL_5_BUFX2_insert681 (
);

FILL FILL_2__12519_ (
);

FILL FILL_5_BUFX2_insert682 (
);

FILL FILL_0__13973_ (
);

FILL FILL_5_BUFX2_insert683 (
);

FILL FILL_0__13553_ (
);

FILL FILL_5_BUFX2_insert684 (
);

FILL FILL_0__13133_ (
);

FILL FILL_5_BUFX2_insert685 (
);

FILL FILL_5_BUFX2_insert686 (
);

FILL FILL_5_BUFX2_insert687 (
);

FILL FILL_5__9590_ (
);

FILL SFILL54040x41050 (
);

FILL FILL_5_BUFX2_insert688 (
);

FILL FILL_5__9170_ (
);

FILL FILL_5_BUFX2_insert689 (
);

FILL FILL_5__16325_ (
);

FILL FILL_0__8519_ (
);

FILL FILL_6__9906_ (
);

FILL FILL_5__11880_ (
);

FILL FILL_5__11460_ (
);

FILL FILL_1__9162_ (
);

FILL FILL_5__11040_ (
);

FILL FILL_4__15738_ (
);

FILL FILL_4__15318_ (
);

FILL FILL_2__16352_ (
);

FILL FILL_3__9088_ (
);

FILL FILL_4__10873_ (
);

FILL FILL_4__10453_ (
);

FILL FILL_4__10033_ (
);

FILL FILL_1__15765_ (
);

FILL FILL_1__15345_ (
);

FILL FILL_1__10060_ (
);

FILL FILL_0__14758_ (
);

INVX1 _14623_ (
    .A(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_5111_)
);

FILL FILL_0__14338_ (
);

OAI22X1 _14203_ (
    .A(_4698_),
    .B(_3955__bF$buf3),
    .C(_3954__bF$buf1),
    .D(_4699_),
    .Y(_4700_)
);

FILL FILL_2__7085_ (
);

FILL FILL_5__12245_ (
);

INVX1 _6965_ (
    .A(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_44_)
);

FILL FILL_4__8372_ (
);

FILL FILL_4__11658_ (
);

FILL FILL_4__11238_ (
);

FILL FILL_2__12272_ (
);

FILL FILL_1__11685_ (
);

FILL FILL_1__11265_ (
);

NAND3X1 _15828_ (
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf2),
    .Y(_6289_)
);

INVX1 _15408_ (
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_5880_)
);

FILL FILL_0__10678_ (
);

NOR2X1 _10963_ (
    .A(ALUOp[1]),
    .B(_2062_),
    .Y(_2095_)
);

FILL FILL_0__8272_ (
);

INVX1 _10543_ (
    .A(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_1860_)
);

FILL FILL_0__10258_ (
);

INVX1 _10123_ (
    .A(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_1641_)
);

FILL SFILL109400x71050 (
);

FILL FILL_6__14457_ (
);

FILL FILL_6__14037_ (
);

FILL FILL_4__15491_ (
);

FILL FILL_4__15071_ (
);

FILL FILL_2__9651_ (
);

FILL FILL_2__9231_ (
);

FILL FILL_3__14484_ (
);

FILL FILL_3__14064_ (
);

FILL FILL_4__9997_ (
);

FILL FILL_4__9157_ (
);

FILL FILL_2__13897_ (
);

FILL FILL_2__13477_ (
);

FILL FILL_0__14091_ (
);

FILL FILL_5__14811_ (
);

FILL FILL_4__13804_ (
);

FILL FILL_3__7994_ (
);

FILL FILL_0__9897_ (
);

FILL FILL_0__9477_ (
);

FILL FILL_3__7574_ (
);

OAI21X1 _11748_ (
    .A(_2344__bF$buf1),
    .B(_2389_),
    .C(_2347__bF$buf3),
    .Y(_2844_)
);

INVX1 _11328_ (
    .A(_2446_),
    .Y(_2447_)
);

FILL FILL_1__13831_ (
);

FILL FILL_1__13411_ (
);

FILL FILL_4__16276_ (
);

FILL FILL_3__15689_ (
);

FILL FILL_0__12824_ (
);

FILL FILL_0__12404_ (
);

FILL FILL_3__15269_ (
);

FILL FILL_5__8861_ (
);

FILL FILL_5__8441_ (
);

FILL FILL_5__8021_ (
);

FILL FILL_0__15296_ (
);

OAI22X1 _15581_ (
    .A(_4586_),
    .B(_5518__bF$buf0),
    .C(_5548__bF$buf4),
    .D(_4599_),
    .Y(_6048_)
);

INVX1 _15161_ (
    .A(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_5639_)
);

FILL FILL_3__16210_ (
);

FILL FILL_1__8853_ (
);

FILL FILL_5__10311_ (
);

FILL FILL_1__8013_ (
);

FILL FILL_2__15623_ (
);

FILL FILL_2__15203_ (
);

FILL FILL_3__8779_ (
);

FILL FILL_3__8359_ (
);

FILL FILL_1__14616_ (
);

OAI21X1 _7083_ (
    .A(_101_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_102_),
    .Y(_68_[17])
);

FILL FILL_4__12196_ (
);

FILL FILL_3__9720_ (
);

FILL SFILL69160x50050 (
);

FILL FILL_0__13609_ (
);

FILL FILL_3__9300_ (
);

FILL FILL_5__9646_ (
);

FILL FILL_5__9226_ (
);

FILL FILL_3__11189_ (
);

INVX1 _16366_ (
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_6798_)
);

FILL SFILL74120x33050 (
);

FILL FILL_5__11936_ (
);

AOI21X1 _11081_ (
    .A(_2194_),
    .B(_2199_),
    .C(_2196_),
    .Y(_2200_)
);

FILL FILL_1__9638_ (
);

FILL FILL_5__11516_ (
);

FILL FILL_3__12970_ (
);

FILL FILL_1__9218_ (
);

FILL FILL_3__12130_ (
);

FILL FILL_2__16408_ (
);

FILL SFILL99320x82050 (
);

FILL FILL_4__7223_ (
);

FILL FILL_4__10929_ (
);

FILL FILL_4__10509_ (
);

FILL FILL_2__11963_ (
);

FILL FILL_2__11543_ (
);

FILL FILL_6__7989_ (
);

FILL FILL_3_CLKBUF1_insert210 (
);

FILL FILL_2__11123_ (
);

FILL FILL_3_CLKBUF1_insert211 (
);

FILL FILL_3_CLKBUF1_insert212 (
);

DFFSR _8288_ (
    .Q(\datapath_1.regfile_1.regOut[11] [10]),
    .CLK(clk_bF$buf59),
    .R(rst_bF$buf103),
    .S(vdd),
    .D(_653_[10])
);

FILL FILL_3_CLKBUF1_insert213 (
);

FILL FILL_3_CLKBUF1_insert214 (
);

FILL FILL_1__10956_ (
);

FILL FILL_3_CLKBUF1_insert215 (
);

FILL FILL_3_CLKBUF1_insert216 (
);

FILL FILL_1__10536_ (
);

FILL FILL_3_CLKBUF1_insert217 (
);

FILL FILL_1__10116_ (
);

FILL FILL_3_CLKBUF1_insert218 (
);

FILL FILL_3_CLKBUF1_insert219 (
);

FILL FILL_0__7963_ (
);

FILL FILL_0__7543_ (
);

FILL FILL_6__8510_ (
);

FILL FILL_0__7123_ (
);

FILL FILL_4__14762_ (
);

FILL FILL_4__14342_ (
);

FILL SFILL64120x76050 (
);

NAND3X1 _12286_ (
    .A(_3251_),
    .B(_3252_),
    .C(_3253_),
    .Y(\datapath_1.alu_1.ALUInB [17])
);

FILL FILL_2__8502_ (
);

FILL FILL_3__13755_ (
);

FILL FILL_3__13335_ (
);

FILL FILL_4__8848_ (
);

FILL FILL_4__8008_ (
);

FILL FILL_2__12748_ (
);

FILL FILL_0__13782_ (
);

FILL FILL_2__12328_ (
);

FILL FILL_0__13362_ (
);

FILL FILL_3__6845_ (
);

FILL FILL_0__8748_ (
);

FILL FILL_5__16134_ (
);

FILL FILL_0__8328_ (
);

FILL FILL_1__9391_ (
);

FILL FILL_4__15967_ (
);

FILL FILL_4__15547_ (
);

FILL FILL_4__15127_ (
);

FILL FILL_2__16161_ (
);

FILL FILL_4__10682_ (
);

FILL FILL_4__10262_ (
);

FILL SFILL64120x31050 (
);

FILL FILL_1__15994_ (
);

FILL FILL_1__15574_ (
);

FILL FILL_1__15154_ (
);

FILL FILL_5__7712_ (
);

FILL FILL_0__14987_ (
);

INVX1 _14852_ (
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_5335_)
);

FILL FILL_0__14567_ (
);

FILL FILL_0__14147_ (
);

INVX1 _14432_ (
    .A(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_4924_)
);

FILL SFILL89320x80050 (
);

FILL FILL112360x29050 (
);

NAND3X1 _14012_ (
    .A(_4502_),
    .B(_4505_),
    .C(_4512_),
    .Y(_4513_)
);

FILL FILL_3__15901_ (
);

FILL FILL_1__7704_ (
);

FILL SFILL64040x38050 (
);

FILL FILL_5__12894_ (
);

FILL FILL_5__12474_ (
);

FILL FILL_5__12054_ (
);

FILL FILL_4__11887_ (
);

FILL FILL_4__11467_ (
);

FILL FILL_4__11047_ (
);

FILL FILL_2__12081_ (
);

FILL SFILL84120x3050 (
);

FILL FILL_1__16359_ (
);

FILL FILL_5__8917_ (
);

FILL FILL_1__11494_ (
);

FILL FILL_1__11074_ (
);

OAI21X1 _15637_ (
    .A(_6101_),
    .B(_5535__bF$buf4),
    .C(_6102_),
    .Y(_6103_)
);

INVX4 _15217_ (
    .A(_5535__bF$buf0),
    .Y(_5693_)
);

FILL FILL_2__8099_ (
);

FILL FILL_0__10487_ (
);

INVX1 _10772_ (
    .A(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_1972_)
);

FILL FILL_0__8081_ (
);

DFFSR _10352_ (
    .Q(\datapath_1.regfile_1.regOut[27] [26]),
    .CLK(clk_bF$buf14),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1693_[26])
);

FILL FILL_0__10067_ (
);

FILL FILL_1__8909_ (
);

FILL FILL_3__11821_ (
);

FILL FILL_3__11401_ (
);

FILL FILL_4__6914_ (
);

FILL FILL_2__10814_ (
);

FILL FILL_5__13679_ (
);

FILL FILL_2__9880_ (
);

FILL FILL_5__13259_ (
);

FILL SFILL113800x40050 (
);

FILL FILL_2__9040_ (
);

FILL FILL_3__14293_ (
);

OAI21X1 _7979_ (
    .A(_556_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_557_),
    .Y(_523_[17])
);

OAI21X1 _7559_ (
    .A(_337_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_338_),
    .Y(_328_[5])
);

DFFSR _7139_ (
    .Q(\datapath_1.regfile_1.regOut[2] [13]),
    .CLK(clk_bF$buf63),
    .R(rst_bF$buf110),
    .S(vdd),
    .D(_68_[13])
);

FILL FILL_4__9386_ (
);

FILL FILL_2__13286_ (
);

FILL FILL_5__14620_ (
);

FILL FILL_5__14200_ (
);

DFFSR _8920_ (
    .Q(\datapath_1.regfile_1.regOut[16] [2]),
    .CLK(clk_bF$buf52),
    .R(rst_bF$buf46),
    .S(vdd),
    .D(_978_[2])
);

FILL SFILL89240x42050 (
);

FILL FILL_1__12699_ (
);

OAI21X1 _8500_ (
    .A(_822_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .C(_823_),
    .Y(_783_[20])
);

FILL FILL_1__12279_ (
);

FILL FILL_4__13613_ (
);

INVX1 _11977_ (
    .A(\datapath_1.PCJump [30]),
    .Y(_3026_)
);

FILL FILL_0__9286_ (
);

AND2X2 _11557_ (
    .A(_2663_),
    .B(_2665_),
    .Y(_2666_)
);

NAND2X1 _11137_ (
    .A(_2254_),
    .B(_2255_),
    .Y(_2256_)
);

FILL FILL_3__12606_ (
);

FILL FILL_1__13640_ (
);

FILL FILL_1__13220_ (
);

FILL FILL_4__16085_ (
);

FILL FILL_6__10186_ (
);

FILL FILL_0__12633_ (
);

FILL FILL_3__15498_ (
);

FILL FILL_0__12213_ (
);

FILL FILL_3__15078_ (
);

FILL SFILL54040x36050 (
);

FILL FILL_5__8250_ (
);

NAND2X1 _15390_ (
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .B(_5649_),
    .Y(_5862_)
);

FILL FILL_5__15825_ (
);

FILL FILL_5__15405_ (
);

DFFSR _9705_ (
    .Q(\datapath_1.regfile_1.regOut[22] [19]),
    .CLK(clk_bF$buf41),
    .R(rst_bF$buf77),
    .S(vdd),
    .D(_1368_[19])
);

FILL FILL_5__10960_ (
);

FILL FILL_5__10540_ (
);

FILL FILL_5__10120_ (
);

FILL FILL_1__8242_ (
);

FILL FILL_4__14818_ (
);

FILL SFILL58360x44050 (
);

FILL FILL_2__15852_ (
);

FILL FILL_2__15432_ (
);

FILL FILL_3__8588_ (
);

FILL FILL_2__15012_ (
);

FILL FILL_1__14845_ (
);

FILL FILL_1__14425_ (
);

FILL FILL_1__14005_ (
);

FILL FILL_0__13838_ (
);

FILL FILL_0__13418_ (
);

INVX1 _13703_ (
    .A(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_4210_)
);

FILL FILL_5__9875_ (
);

FILL SFILL44040x79050 (
);

FILL FILL_5__9035_ (
);

AOI21X1 _16175_ (
    .A(\datapath_1.regfile_1.regOut[7] [28]),
    .B(_5490_),
    .C(_6626_),
    .Y(_6627_)
);

FILL FILL_1__9867_ (
);

FILL FILL_5__11745_ (
);

FILL FILL_5__11325_ (
);

FILL FILL_1__9027_ (
);

FILL SFILL79240x40050 (
);

FILL FILL_4__7872_ (
);

FILL FILL_2__16217_ (
);

FILL FILL_4__7452_ (
);

FILL FILL_4__7032_ (
);

FILL FILL_4__10318_ (
);

FILL FILL_2__11772_ (
);

FILL FILL_2__11352_ (
);

FILL FILL_6__7798_ (
);

FILL FILL_6__7378_ (
);

NAND2X1 _8097_ (
    .A(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_616_)
);

FILL FILL111880x53050 (
);

FILL FILL_1__10765_ (
);

FILL FILL_2_CLKBUF1_insert200 (
);

FILL FILL_2_CLKBUF1_insert201 (
);

AOI22X1 _14908_ (
    .A(\datapath_1.regfile_1.regOut[6] [30]),
    .B(_4001__bF$buf3),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_5390_)
);

FILL FILL_2_CLKBUF1_insert202 (
);

FILL FILL_2_CLKBUF1_insert203 (
);

FILL FILL_2_CLKBUF1_insert204 (
);

FILL FILL_2_CLKBUF1_insert205 (
);

FILL FILL_0__7352_ (
);

FILL FILL_2_CLKBUF1_insert206 (
);

FILL FILL_2_CLKBUF1_insert207 (
);

FILL FILL_2_CLKBUF1_insert208 (
);

FILL FILL_4__14991_ (
);

FILL FILL_2_CLKBUF1_insert209 (
);

FILL FILL_4__14571_ (
);

FILL FILL_4__14151_ (
);

NAND3X1 _12095_ (
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[27]),
    .C(_3032__bF$buf1),
    .Y(_3117_)
);

FILL FILL_3__13984_ (
);

FILL FILL_2__8731_ (
);

FILL FILL_2__8311_ (
);

FILL FILL_3__13564_ (
);

FILL SFILL94280x5050 (
);

FILL FILL_3__13144_ (
);

FILL SFILL69240x83050 (
);

FILL FILL_4__8657_ (
);

FILL FILL_4__8237_ (
);

FILL FILL_2__12977_ (
);

FILL SFILL109000x52050 (
);

FILL FILL_0__13591_ (
);

FILL FILL_2__12137_ (
);

FILL FILL_0__13171_ (
);

FILL FILL_5__16363_ (
);

FILL FILL_0__8977_ (
);

OAI21X1 _10828_ (
    .A(_2008_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_2009_),
    .Y(_1953_[28])
);

FILL FILL_0__8137_ (
);

FILL FILL_6__9524_ (
);

OAI21X1 _10408_ (
    .A(_1789_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .C(_1790_),
    .Y(_1758_[16])
);

FILL FILL_1__12911_ (
);

FILL FILL_4__15776_ (
);

FILL FILL_4__15356_ (
);

FILL FILL_2__16390_ (
);

FILL SFILL104440x8050 (
);

FILL FILL_4__10491_ (
);

FILL FILL_2__9936_ (
);

FILL FILL_0__11904_ (
);

FILL FILL_2__9516_ (
);

FILL FILL_3__14769_ (
);

FILL FILL_3__14349_ (
);

FILL FILL_1__15383_ (
);

FILL FILL_5__7941_ (
);

FILL FILL_5__7101_ (
);

FILL FILL_0__14796_ (
);

FILL FILL_0__14376_ (
);

INVX1 _14661_ (
    .A(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_5148_)
);

NOR2X1 _14241_ (
    .A(_4733_),
    .B(_4736_),
    .Y(_4737_)
);

FILL FILL_3__15710_ (
);

FILL FILL_1__7933_ (
);

FILL FILL_6__13290_ (
);

FILL FILL_2__14703_ (
);

FILL FILL_3__7859_ (
);

FILL FILL_3__7439_ (
);

FILL FILL_5__12283_ (
);

FILL SFILL99400x70050 (
);

FILL FILL_4__11696_ (
);

FILL FILL_4__11276_ (
);

FILL SFILL69160x45050 (
);

FILL FILL_1__16168_ (
);

FILL FILL_3__10689_ (
);

FILL FILL_5__8726_ (
);

FILL FILL_3__10269_ (
);

NOR3X1 _15866_ (
    .A(_6320_),
    .B(_6316_),
    .C(_6325_),
    .Y(_6326_)
);

FILL SFILL74120x28050 (
);

NOR2X1 _15446_ (
    .A(_5916_),
    .B(_5915_),
    .Y(_5917_)
);

NOR2X1 _15026_ (
    .A(_5505_),
    .B(_5502_),
    .Y(_5506_)
);

FILL FILL_0__10296_ (
);

OAI21X1 _10581_ (
    .A(_1884_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .C(_1885_),
    .Y(_1823_[31])
);

FILL SFILL38360x40050 (
);

OAI21X1 _10161_ (
    .A(_1665_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1666_),
    .Y(_1628_[19])
);

FILL FILL_1__8718_ (
);

FILL FILL_3__11630_ (
);

FILL FILL_3__11210_ (
);

FILL FILL_2__15908_ (
);

FILL FILL_0__16102_ (
);

FILL FILL_2__10623_ (
);

FILL FILL_5__13488_ (
);

DFFSR _7788_ (
    .Q(\datapath_1.regfile_1.regOut[7] [22]),
    .CLK(clk_bF$buf74),
    .R(rst_bF$buf88),
    .S(vdd),
    .D(_393_[22])
);

NAND2X1 _7368_ (
    .A(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_252_)
);

FILL FILL_2__13095_ (
);

FILL FILL_5_BUFX2_insert70 (
);

FILL FILL_5_BUFX2_insert71 (
);

FILL FILL_5_BUFX2_insert72 (
);

FILL FILL_5_BUFX2_insert73 (
);

FILL FILL_5_BUFX2_insert74 (
);

FILL FILL_1__12088_ (
);

FILL FILL_5_BUFX2_insert75 (
);

FILL FILL_4__13842_ (
);

FILL FILL_5_BUFX2_insert76 (
);

FILL FILL_4__13422_ (
);

FILL FILL_5_BUFX2_insert77 (
);

FILL FILL_5_BUFX2_insert78 (
);

FILL FILL_4__13002_ (
);

FILL FILL_5_BUFX2_insert79 (
);

FILL FILL_3__7192_ (
);

OAI21X1 _11786_ (
    .A(_2494_),
    .B(_2488_),
    .C(_2560_),
    .Y(_2879_)
);

FILL FILL_0__9095_ (
);

OAI21X1 _11366_ (
    .A(_2479_),
    .B(_2480_),
    .C(_2482_),
    .Y(_2483_)
);

FILL FILL_3__12835_ (
);

FILL FILL_3__12415_ (
);

FILL FILL_4__7928_ (
);

FILL FILL_4__7508_ (
);

FILL FILL_2__11828_ (
);

FILL FILL_0__12862_ (
);

FILL FILL_2__11408_ (
);

FILL SFILL99320x32050 (
);

FILL FILL_0__12442_ (
);

FILL FILL_0__12022_ (
);

FILL SFILL89320x6050 (
);

FILL SFILL23800x4050 (
);

FILL SFILL23720x9050 (
);

FILL SFILL63960x7050 (
);

FILL FILL_5__15634_ (
);

FILL FILL_5__15214_ (
);

FILL FILL_0__7828_ (
);

FILL SFILL28760x52050 (
);

NAND2X1 _9934_ (
    .A(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_1556_)
);

NAND2X1 _9514_ (
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1337_)
);

FILL FILL_1__8891_ (
);

FILL FILL_1__8471_ (
);

FILL FILL_4__14627_ (
);

FILL FILL_2__15661_ (
);

FILL FILL_4__14207_ (
);

FILL FILL_2__15241_ (
);

FILL FILL_3__8397_ (
);

FILL SFILL99240x39050 (
);

FILL SFILL64120x26050 (
);

FILL SFILL3640x5050 (
);

FILL FILL_1__14654_ (
);

FILL FILL_1__14234_ (
);

FILL FILL_0__13647_ (
);

INVX1 _13932_ (
    .A(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_4434_)
);

FILL FILL_0__13227_ (
);

INVX1 _13512_ (
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_4023_)
);

FILL FILL_5__9684_ (
);

FILL FILL_5__9264_ (
);

FILL FILL_6__12981_ (
);

FILL FILL_5__11974_ (
);

FILL FILL_1__9676_ (
);

FILL FILL_5__11554_ (
);

FILL FILL_1__9256_ (
);

FILL FILL_5__11134_ (
);

BUFX2 BUFX2_insert1060 (
    .A(_5531_),
    .Y(_5531__bF$buf1)
);

BUFX2 BUFX2_insert1061 (
    .A(_5531_),
    .Y(_5531__bF$buf0)
);

FILL FILL_4__7681_ (
);

FILL FILL_2__16026_ (
);

BUFX2 BUFX2_insert1062 (
    .A(_5472_),
    .Y(_5472__bF$buf3)
);

FILL FILL_4__10967_ (
);

BUFX2 BUFX2_insert1063 (
    .A(_5472_),
    .Y(_5472__bF$buf2)
);

BUFX2 BUFX2_insert1064 (
    .A(_5472_),
    .Y(_5472__bF$buf1)
);

FILL FILL_4__10547_ (
);

FILL FILL_4__10127_ (
);

BUFX2 BUFX2_insert1065 (
    .A(_5472_),
    .Y(_5472__bF$buf0)
);

FILL FILL_2__11581_ (
);

FILL SFILL54120x69050 (
);

BUFX2 BUFX2_insert1066 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf7 )
);

FILL FILL_2__11161_ (
);

FILL SFILL85000x22050 (
);

FILL FILL_1__15859_ (
);

BUFX2 BUFX2_insert1067 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf6 )
);

BUFX2 BUFX2_insert1068 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf5 )
);

FILL FILL_1__15439_ (
);

FILL FILL_1__15019_ (
);

BUFX2 BUFX2_insert1069 (
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf4 )
);

FILL FILL_1__10994_ (
);

FILL FILL_1__10574_ (
);

FILL FILL_1__10154_ (
);

INVX1 _14717_ (
    .A(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_5203_)
);

FILL SFILL33960x70050 (
);

BUFX2 BUFX2_insert880 (
    .A(_3201_),
    .Y(_3201__bF$buf4)
);

FILL FILL_2__7599_ (
);

FILL FILL_0__7581_ (
);

FILL FILL_2__7179_ (
);

BUFX2 BUFX2_insert881 (
    .A(_3201_),
    .Y(_3201__bF$buf3)
);

FILL FILL_0__7161_ (
);

BUFX2 BUFX2_insert882 (
    .A(_3201_),
    .Y(_3201__bF$buf2)
);

BUFX2 BUFX2_insert883 (
    .A(_3201_),
    .Y(_3201__bF$buf1)
);

FILL SFILL28680x14050 (
);

FILL FILL_3__10901_ (
);

FILL FILL_6__13766_ (
);

BUFX2 BUFX2_insert884 (
    .A(_3201_),
    .Y(_3201__bF$buf0)
);

BUFX2 BUFX2_insert885 (
    .A(_3944_),
    .Y(_3944__bF$buf4)
);

BUFX2 BUFX2_insert886 (
    .A(_3944_),
    .Y(_3944__bF$buf3)
);

FILL FILL_4__14380_ (
);

BUFX2 BUFX2_insert887 (
    .A(_3944_),
    .Y(_3944__bF$buf2)
);

BUFX2 BUFX2_insert888 (
    .A(_3944_),
    .Y(_3944__bF$buf1)
);

BUFX2 BUFX2_insert889 (
    .A(_3944_),
    .Y(_3944__bF$buf0)
);

FILL FILL_2__8960_ (
);

FILL FILL_5__12759_ (
);

FILL FILL_3__13793_ (
);

FILL FILL_5__12339_ (
);

FILL FILL_2__8120_ (
);

FILL FILL_3__13373_ (
);

FILL SFILL18760x50050 (
);

FILL FILL_4__8886_ (
);

FILL FILL_4__8466_ (
);

FILL FILL_2__12786_ (
);

FILL FILL_2__12366_ (
);

FILL FILL_5__13700_ (
);

FILL SFILL89240x37050 (
);

FILL FILL_1__11779_ (
);

FILL FILL_1__11359_ (
);

FILL FILL_5__16172_ (
);

FILL FILL_0__8786_ (
);

FILL FILL_3__6883_ (
);

FILL FILL_0__8366_ (
);

OAI21X1 _10637_ (
    .A(_1901_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1902_),
    .Y(_1888_[7])
);

DFFSR _10217_ (
    .Q(\datapath_1.regfile_1.regOut[26] [19]),
    .CLK(clk_bF$buf78),
    .R(rst_bF$buf113),
    .S(vdd),
    .D(_1628_[19])
);

FILL SFILL79320x73050 (
);

FILL SFILL18680x57050 (
);

FILL FILL_1__12720_ (
);

FILL FILL_4__15585_ (
);

FILL FILL_1__12300_ (
);

FILL FILL_4__15165_ (
);

FILL FILL_3__14998_ (
);

FILL FILL_2__9745_ (
);

FILL FILL_3__14578_ (
);

FILL FILL_0__11713_ (
);

FILL FILL_3__14158_ (
);

FILL FILL_1__15192_ (
);

FILL FILL_5__7750_ (
);

FILL FILL_5__7330_ (
);

AOI22X1 _14890_ (
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .B(_3942__bF$buf2),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_5372_)
);

AOI21X1 _14470_ (
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .B(_4038__bF$buf2),
    .C(_4960_),
    .Y(_4961_)
);

FILL FILL_0__14185_ (
);

FILL SFILL34680x4050 (
);

INVX1 _14050_ (
    .A(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_4550_)
);

FILL FILL_5__14905_ (
);

FILL FILL_1__7742_ (
);

FILL FILL_1__7322_ (
);

FILL FILL_2__14932_ (
);

FILL FILL_2__14512_ (
);

FILL FILL_3__7248_ (
);

FILL FILL_5__12092_ (
);

FILL FILL_1__13925_ (
);

FILL SFILL39560x53050 (
);

FILL FILL_1__13505_ (
);

FILL SFILL33960x6050 (
);

FILL SFILL18680x12050 (
);

FILL FILL_4__11085_ (
);

FILL FILL_0__12918_ (
);

FILL FILL_1__16397_ (
);

FILL SFILL79640x49050 (
);

FILL FILL_5__8955_ (
);

FILL FILL_3__10498_ (
);

FILL FILL_5__8115_ (
);

NOR2X1 _15675_ (
    .A(_6139_),
    .B(_6137_),
    .Y(_6140_)
);

OAI22X1 _15255_ (
    .A(_5463__bF$buf1),
    .B(_4168_),
    .C(_5730_),
    .D(_5504__bF$buf3),
    .Y(_5731_)
);

FILL FILL_3__16304_ (
);

OAI21X1 _10390_ (
    .A(_1777_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1778_),
    .Y(_1758_[10])
);

FILL FILL_5__10825_ (
);

FILL FILL_1__8527_ (
);

FILL FILL_5__10405_ (
);

FILL FILL_1__8107_ (
);

FILL FILL_2__15717_ (
);

FILL FILL_4__6952_ (
);

FILL FILL_0__16331_ (
);

FILL FILL_5__13297_ (
);

FILL FILL_2__10432_ (
);

FILL FILL_2__10012_ (
);

FILL FILL_6__6878_ (
);

NAND2X1 _7597_ (
    .A(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_364_)
);

NAND2X1 _7177_ (
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_145_)
);

FILL FILL111880x48050 (
);

FILL FILL_0__6852_ (
);

FILL SFILL44040x29050 (
);

FILL FILL_4__13651_ (
);

FILL FILL_4__13231_ (
);

NAND3X1 _11595_ (
    .A(_2240_),
    .B(_2248_),
    .C(_2701_),
    .Y(_2702_)
);

AND2X2 _11175_ (
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2294_)
);

FILL FILL_2__7811_ (
);

FILL FILL_3__12644_ (
);

FILL FILL_3__12224_ (
);

FILL FILL_4__7737_ (
);

FILL FILL_4__7317_ (
);

FILL FILL_2__11637_ (
);

FILL FILL_2__11217_ (
);

FILL FILL_0__12251_ (
);

FILL FILL_5__15863_ (
);

FILL FILL_5__15443_ (
);

FILL FILL_5__15023_ (
);

FILL FILL_0__7637_ (
);

NAND2X1 _9743_ (
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1449_)
);

FILL FILL_6__8604_ (
);

FILL FILL_0__7217_ (
);

DFFSR _9323_ (
    .Q(\datapath_1.regfile_1.regOut[19] [21]),
    .CLK(clk_bF$buf18),
    .R(rst_bF$buf24),
    .S(vdd),
    .D(_1173_[21])
);

FILL FILL_4__14856_ (
);

FILL FILL_2__15890_ (
);

FILL FILL_4__14436_ (
);

FILL FILL_4__14016_ (
);

FILL FILL_2__15470_ (
);

FILL FILL_2__15050_ (
);

FILL FILL_3__13849_ (
);

FILL FILL_3__13429_ (
);

FILL FILL_1__14883_ (
);

FILL FILL_1__14463_ (
);

FILL FILL_3__13009_ (
);

FILL FILL_1__14043_ (
);

FILL FILL_0__13876_ (
);

AOI22X1 _13741_ (
    .A(_4246_),
    .B(\datapath_1.regfile_1.regOut[19] [6]),
    .C(\datapath_1.regfile_1.regOut[12] [6]),
    .D(_4005__bF$buf3),
    .Y(_4247_)
);

FILL FILL_0__13456_ (
);

NOR2X1 _13321_ (
    .A(\datapath_1.a3 [1]),
    .B(_3753_),
    .Y(_3851_)
);

FILL FILL_0__13036_ (
);

FILL FILL_5__9493_ (
);

FILL FILL_5__16228_ (
);

FILL FILL_3__6939_ (
);

FILL FILL_5__11783_ (
);

FILL FILL_1__9485_ (
);

FILL FILL_5__11363_ (
);

FILL FILL_2__16255_ (
);

FILL SFILL99400x65050 (
);

FILL FILL_4__7490_ (
);

FILL FILL_4__10776_ (
);

FILL FILL_4__7070_ (
);

FILL FILL_2__11390_ (
);

FILL FILL_1__15668_ (
);

FILL FILL_1__15248_ (
);

FILL FILL_5__7806_ (
);

FILL FILL_1__10383_ (
);

OAI22X1 _14946_ (
    .A(_3884__bF$buf3),
    .B(_5425_),
    .C(_5426_),
    .D(_3916_),
    .Y(_5427_)
);

NAND3X1 _14526_ (
    .A(_5012_),
    .B(_5015_),
    .C(_5009_),
    .Y(_5016_)
);

NAND3X1 _14106_ (
    .A(_4604_),
    .B(_4596_),
    .C(_4597_),
    .Y(_4605_)
);

FILL FILL_0__15602_ (
);

FILL SFILL69160x1050 (
);

FILL FILL_5__12988_ (
);

FILL FILL_5__12568_ (
);

FILL FILL_5__12148_ (
);

BUFX2 _6868_ (
    .A(_1_[30]),
    .Y(memoryAddress[30])
);

FILL FILL_4__8695_ (
);

FILL FILL_4__8275_ (
);

FILL FILL_2__12595_ (
);

FILL FILL_2__12175_ (
);

FILL SFILL99400x20050 (
);

FILL FILL_1__11588_ (
);

FILL FILL_1__11168_ (
);

FILL FILL_4__12502_ (
);

FILL FILL_0__8595_ (
);

DFFSR _10866_ (
    .Q(\datapath_1.regfile_1.regOut[31] [28]),
    .CLK(clk_bF$buf83),
    .R(rst_bF$buf42),
    .S(vdd),
    .D(_1953_[28])
);

NAND2X1 _10446_ (
    .A(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1816_)
);

FILL SFILL59240x31050 (
);

NAND2X1 _10026_ (
    .A(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1597_)
);

FILL FILL_3__11915_ (
);

FILL FILL_4__15394_ (
);

FILL FILL_2__10908_ (
);

FILL FILL_2__9974_ (
);

FILL SFILL99320x27050 (
);

FILL FILL_0__11942_ (
);

FILL FILL_2__9554_ (
);

FILL FILL_2__9134_ (
);

FILL FILL_3__14387_ (
);

FILL FILL_0__11522_ (
);

FILL FILL_0__11102_ (
);

FILL FILL_6__15301_ (
);

FILL FILL_5__14714_ (
);

FILL SFILL28760x47050 (
);

FILL FILL_0__6908_ (
);

FILL FILL_1__7971_ (
);

FILL FILL_1__7551_ (
);

FILL FILL_4__13707_ (
);

FILL FILL_2__14741_ (
);

FILL FILL_2__14321_ (
);

FILL FILL_3__7477_ (
);

FILL SFILL83640x49050 (
);

FILL FILL_3__7057_ (
);

FILL FILL_1__13734_ (
);

FILL FILL_1__13314_ (
);

FILL FILL_4__16179_ (
);

FILL FILL_0__12727_ (
);

FILL FILL_0__12307_ (
);

FILL FILL_5__8764_ (
);

FILL FILL_5__8344_ (
);

FILL FILL_0__15199_ (
);

FILL FILL_6__11221_ (
);

INVX1 _15484_ (
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_5954_)
);

FILL FILL_5__15919_ (
);

NAND3X1 _15064_ (
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5513_),
    .C(_5462_),
    .Y(_5544_)
);

FILL FILL_3__16113_ (
);

FILL FILL_5__10634_ (
);

FILL FILL_1__8756_ (
);

FILL FILL_1__8336_ (
);

FILL FILL_2__15946_ (
);

FILL FILL_2__15526_ (
);

FILL FILL_2__15106_ (
);

FILL FILL_0__16140_ (
);

FILL FILL_2__10661_ (
);

FILL FILL_2__10241_ (
);

FILL FILL_1__14939_ (
);

FILL FILL_1__14519_ (
);

FILL FILL_4__12099_ (
);

FILL FILL_3__9623_ (
);

FILL FILL_5__9549_ (
);

FILL SFILL89320x25050 (
);

FILL FILL_5__9129_ (
);

FILL FILL_6__12846_ (
);

FILL FILL_4__13880_ (
);

FILL FILL_4__13460_ (
);

INVX1 _16269_ (
    .A(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_6719_)
);

FILL FILL_4__13040_ (
);

FILL FILL_5__11839_ (
);

FILL FILL_3__12873_ (
);

FILL FILL_2__7620_ (
);

FILL FILL_5__11419_ (
);

FILL FILL_2__7200_ (
);

FILL FILL_3__12453_ (
);

FILL SFILL18760x45050 (
);

FILL FILL_3__12033_ (
);

FILL FILL_4__7966_ (
);

FILL FILL_4__7546_ (
);

FILL FILL_2__11866_ (
);

FILL FILL_2__11446_ (
);

FILL FILL_0__12480_ (
);

FILL FILL_2__11026_ (
);

FILL FILL_0__12060_ (
);

FILL FILL_1__10439_ (
);

FILL FILL_1__10019_ (
);

FILL FILL_5__15672_ (
);

FILL SFILL39080x5050 (
);

FILL FILL_5__15252_ (
);

FILL FILL_0__7866_ (
);

DFFSR _9972_ (
    .Q(\datapath_1.regfile_1.regOut[24] [30]),
    .CLK(clk_bF$buf85),
    .R(rst_bF$buf64),
    .S(vdd),
    .D(_1498_[30])
);

FILL FILL_0__7446_ (
);

INVX1 _9552_ (
    .A(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_1362_)
);

FILL SFILL79320x68050 (
);

INVX1 _9132_ (
    .A(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_1143_)
);

FILL FILL_1__11800_ (
);

FILL FILL_4__14665_ (
);

FILL FILL_4__14245_ (
);

OAI21X1 _12189_ (
    .A(_3178_),
    .B(ALUSrcA_bF$buf6),
    .C(_3179_),
    .Y(\datapath_1.alu_1.ALUInA [24])
);

FILL FILL_2__8825_ (
);

FILL FILL_3__13658_ (
);

FILL FILL_2__8405_ (
);

FILL FILL_3__13238_ (
);

FILL FILL_1__14692_ (
);

FILL FILL_1__14272_ (
);

FILL FILL_0_BUFX2_insert520 (
);

FILL FILL_0_BUFX2_insert521 (
);

FILL FILL_0_BUFX2_insert522 (
);

FILL FILL_0_BUFX2_insert523 (
);

FILL FILL_0__13685_ (
);

FILL FILL_0_BUFX2_insert524 (
);

NOR2X1 _13970_ (
    .A(_4471_),
    .B(_4468_),
    .Y(_4472_)
);

FILL FILL_0__13265_ (
);

FILL FILL_0_BUFX2_insert525 (
);

OAI22X1 _13550_ (
    .A(_4058_),
    .B(_3930__bF$buf2),
    .C(_3954__bF$buf2),
    .D(_4059_),
    .Y(_4060_)
);

INVX1 _13130_ (
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3718_)
);

FILL FILL_0_BUFX2_insert526 (
);

FILL FILL_0_BUFX2_insert527 (
);

FILL FILL_0_BUFX2_insert528 (
);

FILL FILL_0_BUFX2_insert529 (
);

FILL SFILL23960x50 (
);

FILL FILL_5__16037_ (
);

FILL FILL_5__11592_ (
);

FILL FILL_1__9294_ (
);

FILL FILL_5__11172_ (
);

FILL SFILL79320x23050 (
);

FILL FILL_2__16064_ (
);

FILL FILL_4__10165_ (
);

FILL FILL_1__15897_ (
);

FILL FILL_1__15477_ (
);

FILL FILL_1__15057_ (
);

FILL FILL_5__7615_ (
);

FILL FILL111960x36050 (
);

FILL FILL_1__10192_ (
);

INVX1 _14755_ (
    .A(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_5240_)
);

INVX1 _14335_ (
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_4829_)
);

FILL FILL_3__15804_ (
);

FILL FILL_1__7607_ (
);

FILL FILL_0__15831_ (
);

FILL FILL_0__15411_ (
);

FILL FILL_5__12377_ (
);

FILL FILL_4__8084_ (
);

FILL FILL_1__11397_ (
);

FILL SFILL114760x69050 (
);

FILL FILL_4__12731_ (
);

FILL FILL_4__12311_ (
);

NAND2X1 _10675_ (
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1928_)
);

NAND2X1 _10255_ (
    .A(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1709_)
);

FILL FILL_3__11724_ (
);

FILL FILL_3__11304_ (
);

FILL FILL_2__9783_ (
);

FILL FILL_0__11751_ (
);

FILL FILL_2__9363_ (
);

FILL FILL_3__14196_ (
);

FILL FILL_0__11331_ (
);

FILL FILL_4__9289_ (
);

FILL SFILL69320x21050 (
);

FILL FILL_5__14943_ (
);

FILL FILL_5__14523_ (
);

FILL FILL_5__14103_ (
);

NAND2X1 _8823_ (
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .Y(_1042_)
);

INVX1 _8403_ (
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_779_)
);

FILL FILL_1__7360_ (
);

FILL FILL_4__13936_ (
);

FILL FILL_2__14970_ (
);

FILL FILL_4__13516_ (
);

FILL FILL_2__14550_ (
);

FILL FILL_2__14130_ (
);

FILL FILL_3__7286_ (
);

FILL FILL_3__12509_ (
);

FILL FILL_1__13963_ (
);

FILL FILL_1__13543_ (
);

FILL FILL_1__13123_ (
);

FILL SFILL69240x28050 (
);

FILL FILL_0__12956_ (
);

DFFSR _12821_ (
    .Q(\control_1.op [4]),
    .CLK(clk_bF$buf30),
    .R(rst_bF$buf4),
    .S(vdd),
    .D(_3490_[30])
);

NAND2X1 _12401_ (
    .A(MemToReg_bF$buf6),
    .B(\datapath_1.Data [19]),
    .Y(_3333_)
);

FILL FILL_0__12116_ (
);

FILL FILL_5__8993_ (
);

FILL FILL_5__8573_ (
);

NOR2X1 _15293_ (
    .A(_5766_),
    .B(_5767_),
    .Y(_5768_)
);

FILL FILL_5__15728_ (
);

FILL FILL_5__15308_ (
);

FILL FILL_3__16342_ (
);

INVX1 _9608_ (
    .A(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_1379_)
);

FILL FILL_1__8985_ (
);

FILL FILL_5__10443_ (
);

FILL FILL_5__10023_ (
);

FILL FILL_1__8145_ (
);

FILL FILL_2__15755_ (
);

FILL FILL_4__6990_ (
);

FILL FILL_2__15335_ (
);

FILL FILL_2__10890_ (
);

FILL FILL_2__10050_ (
);

FILL FILL_1__14748_ (
);

FILL FILL_1__14328_ (
);

FILL FILL_3__9852_ (
);

INVX4 _13606_ (
    .A(_3902__bF$buf1),
    .Y(_4115_)
);

FILL FILL_3__9012_ (
);

FILL FILL_0__6890_ (
);

FILL FILL_5__9778_ (
);

FILL FILL_5__9358_ (
);

FILL FILL_6__12655_ (
);

OAI22X1 _16078_ (
    .A(_6532_),
    .B(_5518__bF$buf0),
    .C(_5478__bF$buf3),
    .D(_5136_),
    .Y(_6533_)
);

FILL FILL_5__11648_ (
);

FILL FILL_5__11228_ (
);

FILL FILL_3__12262_ (
);

FILL FILL_4__7355_ (
);

FILL FILL_2__11675_ (
);

FILL FILL_2__11255_ (
);

FILL SFILL99400x15050 (
);

FILL FILL_1__10668_ (
);

FILL FILL_1__10248_ (
);

FILL FILL_5__15481_ (
);

FILL FILL_5__15061_ (
);

FILL FILL_0__7675_ (
);

INVX1 _9781_ (
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_1474_)
);

INVX1 _9361_ (
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_1255_)
);

FILL FILL_4__14894_ (
);

FILL FILL_4__14474_ (
);

FILL FILL_4__14054_ (
);

FILL FILL_3__13887_ (
);

FILL FILL_2__8634_ (
);

FILL FILL_3__13467_ (
);

FILL FILL_2__8214_ (
);

FILL FILL_1__14081_ (
);

FILL FILL_0__13494_ (
);

FILL SFILL89400x58050 (
);

FILL FILL_4__9921_ (
);

FILL FILL_4__9501_ (
);

FILL FILL_2__13821_ (
);

FILL FILL_2__13401_ (
);

FILL FILL_5__16266_ (
);

FILL FILL_3__6977_ (
);

FILL FILL_6__9007_ (
);

FILL FILL_4__15679_ (
);

FILL FILL_4__15259_ (
);

FILL FILL_2__16293_ (
);

FILL FILL_4__10394_ (
);

FILL FILL_2__9419_ (
);

FILL FILL_0__9401_ (
);

FILL FILL_0__11807_ (
);

FILL FILL_1__15286_ (
);

FILL FILL_5__7844_ (
);

FILL FILL_5__7424_ (
);

FILL FILL_4__16200_ (
);

INVX1 _14984_ (
    .A(\datapath_1.PCJump [26]),
    .Y(_5464_)
);

FILL FILL_0__14699_ (
);

OAI22X1 _14564_ (
    .A(_5051_),
    .B(_3930__bF$buf3),
    .C(_3931__bF$buf0),
    .D(_5052_),
    .Y(_5053_)
);

FILL FILL_0__14279_ (
);

NOR2X1 _14144_ (
    .A(_4641_),
    .B(_4631_),
    .Y(_4642_)
);

FILL FILL_3__15613_ (
);

FILL SFILL89400x13050 (
);

FILL FILL_1__7836_ (
);

FILL FILL_1__7416_ (
);

FILL SFILL94280x64050 (
);

FILL FILL_2__14606_ (
);

FILL FILL_0__15640_ (
);

FILL FILL_0__15220_ (
);

FILL FILL_5__12186_ (
);

FILL FILL_4__11599_ (
);

FILL FILL_4__11179_ (
);

FILL FILL_3__8703_ (
);

FILL FILL_5__8629_ (
);

FILL FILL_5__8209_ (
);

FILL FILL_4__12960_ (
);

NOR3X1 _15769_ (
    .A(_6231_),
    .B(_6211_),
    .C(_6221_),
    .Y(_6232_)
);

AOI22X1 _15349_ (
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_5822_)
);

FILL FILL_4__12120_ (
);

DFFSR _10484_ (
    .Q(\datapath_1.regfile_1.regOut[28] [30]),
    .CLK(clk_bF$buf76),
    .R(rst_bF$buf20),
    .S(vdd),
    .D(_1758_[30])
);

FILL FILL_5__10919_ (
);

INVX1 _10064_ (
    .A(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_1622_)
);

FILL FILL_3__11953_ (
);

FILL FILL_3__11533_ (
);

FILL FILL_3__11113_ (
);

FILL FILL_0__16005_ (
);

FILL FILL_2__10946_ (
);

FILL FILL_2__9592_ (
);

FILL FILL_0__11980_ (
);

FILL FILL_2__10526_ (
);

FILL FILL_2__9172_ (
);

FILL FILL_0__11560_ (
);

FILL FILL_2__10106_ (
);

FILL FILL_0__11140_ (
);

FILL FILL_4__9098_ (
);

FILL FILL_3__9908_ (
);

FILL FILL_5__14752_ (
);

FILL FILL_0__6946_ (
);

FILL FILL_5__14332_ (
);

INVX1 _8632_ (
    .A(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_891_)
);

FILL SFILL8680x81050 (
);

INVX1 _8212_ (
    .A(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_672_)
);

endmodule
