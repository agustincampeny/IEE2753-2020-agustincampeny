* NGSPICE file created from mips.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

.subckt mips gnd vdd MemRead MemWrite clk memoryAddress[31] memoryAddress[30] memoryAddress[29]
+ memoryAddress[28] memoryAddress[27] memoryAddress[26] memoryAddress[25] memoryAddress[24]
+ memoryAddress[23] memoryAddress[22] memoryAddress[21] memoryAddress[20] memoryAddress[19]
+ memoryAddress[18] memoryAddress[17] memoryAddress[16] memoryAddress[15] memoryAddress[14]
+ memoryAddress[13] memoryAddress[12] memoryAddress[11] memoryAddress[10] memoryAddress[9]
+ memoryAddress[8] memoryAddress[7] memoryAddress[6] memoryAddress[5] memoryAddress[4]
+ memoryAddress[3] memoryAddress[2] memoryAddress[1] memoryAddress[0] memoryOutData[31]
+ memoryOutData[30] memoryOutData[29] memoryOutData[28] memoryOutData[27] memoryOutData[26]
+ memoryOutData[25] memoryOutData[24] memoryOutData[23] memoryOutData[22] memoryOutData[21]
+ memoryOutData[20] memoryOutData[19] memoryOutData[18] memoryOutData[17] memoryOutData[16]
+ memoryOutData[15] memoryOutData[14] memoryOutData[13] memoryOutData[12] memoryOutData[11]
+ memoryOutData[10] memoryOutData[9] memoryOutData[8] memoryOutData[7] memoryOutData[6]
+ memoryOutData[5] memoryOutData[4] memoryOutData[3] memoryOutData[2] memoryOutData[1]
+ memoryOutData[0] memoryWriteData[31] memoryWriteData[30] memoryWriteData[29] memoryWriteData[28]
+ memoryWriteData[27] memoryWriteData[26] memoryWriteData[25] memoryWriteData[24]
+ memoryWriteData[23] memoryWriteData[22] memoryWriteData[21] memoryWriteData[20]
+ memoryWriteData[19] memoryWriteData[18] memoryWriteData[17] memoryWriteData[16]
+ memoryWriteData[15] memoryWriteData[14] memoryWriteData[13] memoryWriteData[12]
+ memoryWriteData[11] memoryWriteData[10] memoryWriteData[9] memoryWriteData[8] memoryWriteData[7]
+ memoryWriteData[6] memoryWriteData[5] memoryWriteData[4] memoryWriteData[3] memoryWriteData[2]
+ memoryWriteData[1] memoryWriteData[0] rst
XFILL_5__15675_ gnd vdd FILL
XFILL_5__12887_ gnd vdd FILL
XFILL_2__14515_ gnd vdd FILL
XFILL_4__10548_ gnd vdd FILL
XFILL_2__9369_ gnd vdd FILL
XFILL_1__13156_ gnd vdd FILL
XFILL_0__12906_ gnd vdd FILL
XFILL_2__11727_ gnd vdd FILL
XFILL_1__10368_ gnd vdd FILL
XSFILL54840x78050 gnd vdd FILL
XSFILL54040x59050 gnd vdd FILL
XFILL_2__15495_ gnd vdd FILL
XFILL_6__11108_ gnd vdd FILL
XFILL_0__13886_ gnd vdd FILL
XFILL_5__9078_ gnd vdd FILL
XFILL_5__14626_ gnd vdd FILL
XFILL_0__8384_ gnd vdd FILL
XSFILL94440x64050 gnd vdd FILL
XFILL_3__15805_ gnd vdd FILL
XFILL_4__16055_ gnd vdd FILL
XFILL_5__11838_ gnd vdd FILL
XFILL_4__13267_ gnd vdd FILL
XFILL_1__12107_ gnd vdd FILL
XFILL_3__7113_ gnd vdd FILL
XFILL_2__14446_ gnd vdd FILL
XFILL_0__15625_ gnd vdd FILL
XFILL_0__12837_ gnd vdd FILL
XFILL_1__13087_ gnd vdd FILL
XFILL_3__13997_ gnd vdd FILL
XFILL_2__11658_ gnd vdd FILL
XFILL_3__8093_ gnd vdd FILL
XFILL_1__10299_ gnd vdd FILL
XFILL_4__15006_ gnd vdd FILL
XSFILL95080x30050 gnd vdd FILL
XFILL_6__9891_ gnd vdd FILL
XFILL_0__7335_ gnd vdd FILL
XFILL_4__12218_ gnd vdd FILL
XFILL_5__14557_ gnd vdd FILL
X_7963_ _7972_/A _7451_/B gnd _7963_/Y vdd NAND2X1
XSFILL69240x40050 gnd vdd FILL
XFILL_5__11769_ gnd vdd FILL
XFILL_3__15736_ gnd vdd FILL
XFILL_3__7044_ gnd vdd FILL
XFILL_1__12038_ gnd vdd FILL
XSFILL33880x17050 gnd vdd FILL
XFILL_0__15556_ gnd vdd FILL
XFILL_2__14377_ gnd vdd FILL
XFILL_2__11589_ gnd vdd FILL
XFILL_6__8842_ gnd vdd FILL
XFILL_0__12768_ gnd vdd FILL
X_9702_ _9702_/Q _7021_/CLK _9062_/R vdd _9702_/D gnd vdd DFFSR
X_6914_ _7002_/Q gnd _6916_/A vdd INVX1
XFILL_5__13508_ gnd vdd FILL
XFILL_5__14488_ gnd vdd FILL
XFILL_2__16116_ gnd vdd FILL
XFILL_4__12149_ gnd vdd FILL
XFILL_2__13328_ gnd vdd FILL
XFILL_3__15667_ gnd vdd FILL
X_7894_ _7894_/Q _9436_/CLK _9454_/R vdd _7894_/D gnd vdd DFFSR
XFILL_0__14507_ gnd vdd FILL
XSFILL48920x39050 gnd vdd FILL
XFILL_3__12879_ gnd vdd FILL
XFILL_0__11719_ gnd vdd FILL
XFILL_0__9005_ gnd vdd FILL
XFILL_0__15487_ gnd vdd FILL
XFILL_0__12699_ gnd vdd FILL
XFILL_5__16227_ gnd vdd FILL
XFILL_3__14618_ gnd vdd FILL
X_6845_ _6845_/A gnd memoryAddress[7] vdd BUFX2
X_9633_ _9613_/B _9633_/B gnd _9633_/Y vdd NAND2X1
XFILL_5__13439_ gnd vdd FILL
XFILL_0__7197_ gnd vdd FILL
XFILL_2__16047_ gnd vdd FILL
XFILL_2__13259_ gnd vdd FILL
XFILL_3__15598_ gnd vdd FILL
XFILL_0__14438_ gnd vdd FILL
XFILL_3__8995_ gnd vdd FILL
XSFILL89960x10050 gnd vdd FILL
XSFILL49000x48050 gnd vdd FILL
XFILL_1__13989_ gnd vdd FILL
XFILL_4__15908_ gnd vdd FILL
X_9564_ _9564_/Q _8022_/CLK _9046_/R vdd _9564_/D gnd vdd DFFSR
XFILL_5__16158_ gnd vdd FILL
XFILL_3__14549_ gnd vdd FILL
XFILL_3__7946_ gnd vdd FILL
XFILL_1__15728_ gnd vdd FILL
XFILL_5_BUFX2_insert403 gnd vdd FILL
XFILL_0__14369_ gnd vdd FILL
XFILL_5_BUFX2_insert414 gnd vdd FILL
X_8515_ _8513_/Y _8469_/A _8515_/C gnd _8559_/D vdd OAI21X1
XFILL_5__15109_ gnd vdd FILL
XSFILL109560x59050 gnd vdd FILL
XFILL_5_BUFX2_insert425 gnd vdd FILL
XFILL_5__16089_ gnd vdd FILL
X_9495_ _9569_/Q gnd _9495_/Y vdd INVX1
XFILL_1__6961_ gnd vdd FILL
XFILL_4__15839_ gnd vdd FILL
XFILL_0__16108_ gnd vdd FILL
XFILL_5_BUFX2_insert436 gnd vdd FILL
XFILL_1__15659_ gnd vdd FILL
XFILL_3__7877_ gnd vdd FILL
XFILL_5_BUFX2_insert447 gnd vdd FILL
XFILL_5_BUFX2_insert458 gnd vdd FILL
XFILL_0__9907_ gnd vdd FILL
XFILL_1__8700_ gnd vdd FILL
XFILL_3__16219_ gnd vdd FILL
XFILL_6__7586_ gnd vdd FILL
X_8446_ _8444_/Y _8494_/B _8446_/C gnd _8446_/Y vdd OAI21X1
XFILL_5_BUFX2_insert469 gnd vdd FILL
XFILL_3__9616_ gnd vdd FILL
XFILL_1__9680_ gnd vdd FILL
XFILL_0__16039_ gnd vdd FILL
XFILL_1__6892_ gnd vdd FILL
XFILL_1__8631_ gnd vdd FILL
X_8377_ _8360_/B _8377_/B gnd _8377_/Y vdd NAND2X1
XFILL_3__9547_ gnd vdd FILL
XFILL_4__8340_ gnd vdd FILL
X_7328_ _7328_/A gnd _7330_/A vdd INVX1
XFILL_0__9769_ gnd vdd FILL
XFILL_4__8271_ gnd vdd FILL
XFILL_3__9478_ gnd vdd FILL
XSFILL18760x58050 gnd vdd FILL
X_7259_ _7173_/A _7143_/CLK _7015_/R vdd _7259_/D gnd vdd DFFSR
XFILL_4__7222_ gnd vdd FILL
XSFILL8600x68050 gnd vdd FILL
XFILL_1__8493_ gnd vdd FILL
XSFILL58360x44050 gnd vdd FILL
XFILL_6__8138_ gnd vdd FILL
XSFILL33800x61050 gnd vdd FILL
XFILL_1__7444_ gnd vdd FILL
XFILL_2_BUFX2_insert304 gnd vdd FILL
XFILL_2_BUFX2_insert315 gnd vdd FILL
XFILL_1__7375_ gnd vdd FILL
XSFILL23880x49050 gnd vdd FILL
XFILL_2_BUFX2_insert326 gnd vdd FILL
X_11900_ _11900_/A _12355_/A gnd _11901_/C vdd NAND2X1
XFILL_4__7084_ gnd vdd FILL
XFILL_2_BUFX2_insert337 gnd vdd FILL
XFILL_1__9114_ gnd vdd FILL
XFILL_2_BUFX2_insert348 gnd vdd FILL
X_12880_ _12938_/Q gnd _12880_/Y vdd INVX1
XFILL_2_BUFX2_insert359 gnd vdd FILL
XFILL111960x71050 gnd vdd FILL
XFILL112440x78050 gnd vdd FILL
X_11831_ _11238_/Y _11374_/Y gnd _11835_/A vdd NOR2X1
XFILL_1__9045_ gnd vdd FILL
X_14550_ _9965_/Q gnd _14550_/Y vdd INVX1
X_11762_ _11761_/Y _11762_/B gnd _11763_/C vdd OR2X2
X_13501_ _15095_/D _14068_/C _14342_/B _13499_/Y gnd _13502_/B vdd OAI22X1
X_10713_ _10623_/A _8921_/CLK _8942_/R vdd _10713_/D gnd vdd DFFSR
XBUFX2_insert303 _12414_/Y gnd _9788_/B vdd BUFX2
XFILL_4__7986_ gnd vdd FILL
X_14481_ _10859_/Q _14877_/D _14481_/C _7019_/Q gnd _14483_/A vdd AOI22X1
XBUFX2_insert314 _13454_/Y gnd _14030_/C vdd BUFX2
X_11693_ _11066_/Y _11366_/B gnd _11693_/Y vdd NAND2X1
XFILL_6_BUFX2_insert270 gnd vdd FILL
XFILL_4__9725_ gnd vdd FILL
XBUFX2_insert325 _13345_/Y gnd _9941_/B vdd BUFX2
X_16220_ _16220_/A _16220_/B gnd _16244_/A vdd NOR2X1
XFILL_4__6937_ gnd vdd FILL
XSFILL18840x38050 gnd vdd FILL
XBUFX2_insert336 _13494_/Y gnd _14037_/B vdd BUFX2
X_13432_ _13381_/A _13423_/B _13407_/Y gnd _13432_/Y vdd NAND3X1
XBUFX2_insert347 _10927_/Y gnd _12255_/A vdd BUFX2
XSFILL84280x14050 gnd vdd FILL
XBUFX2_insert358 _13306_/Y gnd _8006_/B vdd BUFX2
X_10644_ _10720_/Q gnd _10646_/A vdd INVX1
XFILL_2__8740_ gnd vdd FILL
XBUFX2_insert369 _13338_/Y gnd _9535_/A vdd BUFX2
XFILL_4__9656_ gnd vdd FILL
XFILL_5_CLKBUF1_insert204 gnd vdd FILL
XFILL_5_CLKBUF1_insert215 gnd vdd FILL
XFILL_4__6868_ gnd vdd FILL
X_16151_ _16150_/Y _16151_/B _16309_/A _16151_/D gnd _16151_/Y vdd OAI22X1
X_10575_ _10575_/A _10535_/A _10575_/C gnd _10575_/Y vdd OAI21X1
X_13363_ _13220_/A _13363_/B gnd _13363_/Y vdd NAND2X1
XSFILL69080x75050 gnd vdd FILL
XFILL_5_BUFX2_insert970 gnd vdd FILL
XFILL_1__9878_ gnd vdd FILL
XFILL_4__8607_ gnd vdd FILL
XSFILL85160x42050 gnd vdd FILL
X_15102_ _15102_/A _15102_/B _15099_/Y gnd _15103_/A vdd NAND3X1
XFILL_5__8380_ gnd vdd FILL
X_12314_ _12311_/Y _12312_/Y _12314_/C gnd _12314_/Y vdd NAND3X1
XFILL_5_BUFX2_insert981 gnd vdd FILL
XFILL_5_BUFX2_insert992 gnd vdd FILL
XFILL_3__10230_ gnd vdd FILL
XFILL_6__11390_ gnd vdd FILL
X_16082_ _16082_/A _15527_/C _15449_/C _14683_/A gnd _16084_/A vdd OAI22X1
X_13294_ _13294_/A gnd _13294_/Y vdd INVX1
XFILL_2__7622_ gnd vdd FILL
XFILL_1__8829_ gnd vdd FILL
XSFILL22920x65050 gnd vdd FILL
XFILL_2__10960_ gnd vdd FILL
XFILL_5__7331_ gnd vdd FILL
XFILL_0__10050_ gnd vdd FILL
X_15033_ _12813_/Q _12812_/Q gnd _15212_/B vdd NOR2X1
X_12245_ _6877_/A _12249_/B _12249_/C _12710_/A gnd _12246_/C vdd AOI22X1
XSFILL64840x4050 gnd vdd FILL
XFILL_4__11520_ gnd vdd FILL
XFILL_3__10161_ gnd vdd FILL
XFILL_2__7553_ gnd vdd FILL
XFILL_1__11340_ gnd vdd FILL
XFILL_2__10891_ gnd vdd FILL
XFILL_4__8469_ gnd vdd FILL
X_12176_ _12123_/B _12176_/B gnd _12176_/Y vdd NAND2X1
XFILL_5__13790_ gnd vdd FILL
XFILL_4__11451_ gnd vdd FILL
XFILL_2__12630_ gnd vdd FILL
XFILL_5__9001_ gnd vdd FILL
XFILL_2__7484_ gnd vdd FILL
XFILL_1__11271_ gnd vdd FILL
XFILL_5__12741_ gnd vdd FILL
XFILL_4__10402_ gnd vdd FILL
XFILL_5__7193_ gnd vdd FILL
X_11127_ _12174_/Y _12294_/Y gnd _11591_/A vdd NOR2X1
XFILL_4__14170_ gnd vdd FILL
XFILL_1__13010_ gnd vdd FILL
XFILL_3__13920_ gnd vdd FILL
XFILL_2__9223_ gnd vdd FILL
XFILL_4__11382_ gnd vdd FILL
XFILL_0__13740_ gnd vdd FILL
XFILL_0__10952_ gnd vdd FILL
X_15935_ _8376_/A _15978_/B _16293_/A _7148_/Q gnd _15936_/B vdd AOI22X1
XFILL_4__13121_ gnd vdd FILL
X_11058_ _12278_/Y _12162_/Y gnd _11061_/C vdd XNOR2X1
XSFILL114440x12050 gnd vdd FILL
XFILL_2__14300_ gnd vdd FILL
XFILL_5__15460_ gnd vdd FILL
XFILL_3__13851_ gnd vdd FILL
XFILL_2__9154_ gnd vdd FILL
XFILL_2__11512_ gnd vdd FILL
XFILL_2__12492_ gnd vdd FILL
XFILL_1__10153_ gnd vdd FILL
XFILL_2__15280_ gnd vdd FILL
XSFILL94360x79050 gnd vdd FILL
XFILL_0__13671_ gnd vdd FILL
X_10009_ _10007_/Y _10024_/B _10008_/Y gnd _10009_/Y vdd OAI21X1
XFILL_0__10883_ gnd vdd FILL
XFILL_5__14411_ gnd vdd FILL
XFILL_5__11623_ gnd vdd FILL
XFILL_5__15391_ gnd vdd FILL
XFILL_2__8105_ gnd vdd FILL
X_15866_ _15860_/Y _15866_/B _15866_/C gnd _15891_/A vdd NOR3X1
XFILL_0__15410_ gnd vdd FILL
XFILL_2__14231_ gnd vdd FILL
XFILL_4__10264_ gnd vdd FILL
XFILL_2__11443_ gnd vdd FILL
XFILL_0__12622_ gnd vdd FILL
XFILL_2_BUFX2_insert860 gnd vdd FILL
XFILL_3__13782_ gnd vdd FILL
XFILL_2__9085_ gnd vdd FILL
XFILL_0__16390_ gnd vdd FILL
XFILL_2_BUFX2_insert871 gnd vdd FILL
XFILL_1__14961_ gnd vdd FILL
XFILL_5__9903_ gnd vdd FILL
XSFILL99400x16050 gnd vdd FILL
XFILL_0__7120_ gnd vdd FILL
XFILL_3__10994_ gnd vdd FILL
XSFILL69160x55050 gnd vdd FILL
X_14817_ _9418_/A gnd _14818_/D vdd INVX1
XFILL_4__12003_ gnd vdd FILL
XFILL_5__14342_ gnd vdd FILL
XFILL_6__12913_ gnd vdd FILL
XFILL_3__15521_ gnd vdd FILL
XFILL_2_BUFX2_insert882 gnd vdd FILL
XFILL_5__11554_ gnd vdd FILL
XFILL_2_BUFX2_insert893 gnd vdd FILL
XFILL_3__12733_ gnd vdd FILL
X_15797_ _15797_/A gnd _15798_/D vdd INVX1
XFILL_0__15341_ gnd vdd FILL
XFILL_2__14162_ gnd vdd FILL
XFILL_4__10195_ gnd vdd FILL
XFILL_1__13912_ gnd vdd FILL
XFILL_2__11374_ gnd vdd FILL
XFILL_0__7051_ gnd vdd FILL
XFILL_5__10505_ gnd vdd FILL
XFILL_1__14892_ gnd vdd FILL
X_14748_ _8945_/Q gnd _14748_/Y vdd INVX1
XFILL_5__14273_ gnd vdd FILL
XFILL_2__13113_ gnd vdd FILL
XFILL_3__15452_ gnd vdd FILL
XFILL_5__11485_ gnd vdd FILL
XFILL_2__10325_ gnd vdd FILL
XFILL_2__14093_ gnd vdd FILL
XFILL_0__11504_ gnd vdd FILL
XFILL_1__13843_ gnd vdd FILL
XFILL_0__15272_ gnd vdd FILL
XFILL_5__9765_ gnd vdd FILL
XFILL_5__13224_ gnd vdd FILL
XFILL_5__16012_ gnd vdd FILL
XFILL_0__12484_ gnd vdd FILL
XSFILL74280x46050 gnd vdd FILL
XFILL_5__10436_ gnd vdd FILL
XFILL_4_BUFX2_insert3 gnd vdd FILL
XFILL_5__6977_ gnd vdd FILL
XFILL_3__14403_ gnd vdd FILL
XFILL_3__7800_ gnd vdd FILL
XFILL_2__13044_ gnd vdd FILL
XFILL_4__13954_ gnd vdd FILL
XFILL_3__11615_ gnd vdd FILL
X_14679_ _14678_/Y _14679_/B gnd _14680_/C vdd NOR2X1
XFILL_2__10256_ gnd vdd FILL
XFILL_3__15383_ gnd vdd FILL
XFILL_0__14223_ gnd vdd FILL
XFILL_3__12595_ gnd vdd FILL
XFILL_5__8716_ gnd vdd FILL
XFILL_2__9987_ gnd vdd FILL
XFILL_3__8780_ gnd vdd FILL
XFILL_0__11435_ gnd vdd FILL
XFILL_1__13774_ gnd vdd FILL
X_16418_ _16324_/A _8679_/CLK _7131_/R vdd _16326_/Y gnd vdd DFFSR
XFILL_5__13155_ gnd vdd FILL
XSFILL49080x22050 gnd vdd FILL
XFILL_5__10367_ gnd vdd FILL
XSFILL89320x68050 gnd vdd FILL
XFILL_3__14334_ gnd vdd FILL
XFILL_4__12905_ gnd vdd FILL
XFILL_4__13885_ gnd vdd FILL
XFILL_1__15513_ gnd vdd FILL
XFILL_3__7731_ gnd vdd FILL
XFILL_3__11546_ gnd vdd FILL
XFILL_1__12725_ gnd vdd FILL
XFILL_2__10187_ gnd vdd FILL
XFILL_0__14154_ gnd vdd FILL
X_8300_ _8248_/A _7661_/CLK _8819_/R vdd _8250_/Y gnd vdd DFFSR
XFILL_5__12106_ gnd vdd FILL
XBUFX2_insert870 _13379_/Y gnd _14738_/A vdd BUFX2
XFILL_5__8647_ gnd vdd FILL
XFILL_0__11366_ gnd vdd FILL
XBUFX2_insert881 _12216_/Y gnd _12269_/C vdd BUFX2
X_16349_ gnd gnd gnd _16349_/Y vdd NAND2X1
X_9280_ _9278_/Y _9232_/B _9279_/Y gnd _9326_/D vdd OAI21X1
XBUFX2_insert892 _12369_/Y gnd _9487_/B vdd BUFX2
XFILL_4__15624_ gnd vdd FILL
XFILL_4__12836_ gnd vdd FILL
XFILL_5__13086_ gnd vdd FILL
XFILL_0__7953_ gnd vdd FILL
XFILL_3__14265_ gnd vdd FILL
XFILL_0__13105_ gnd vdd FILL
XFILL_5__10298_ gnd vdd FILL
XFILL_1__12656_ gnd vdd FILL
XFILL_2__8869_ gnd vdd FILL
XFILL_0__10317_ gnd vdd FILL
XFILL_3__11477_ gnd vdd FILL
XFILL_1__15444_ gnd vdd FILL
XFILL_2__14995_ gnd vdd FILL
XFILL_0__14085_ gnd vdd FILL
XFILL_3__16004_ gnd vdd FILL
XFILL_5__8578_ gnd vdd FILL
X_8231_ _8232_/B _7079_/B gnd _8231_/Y vdd NAND2X1
XFILL_0__6904_ gnd vdd FILL
XFILL_5__12037_ gnd vdd FILL
XFILL_0__11297_ gnd vdd FILL
XFILL_3__13216_ gnd vdd FILL
XFILL_4__15555_ gnd vdd FILL
XFILL_3__9401_ gnd vdd FILL
XFILL_3__10428_ gnd vdd FILL
XFILL_4__12767_ gnd vdd FILL
XFILL_0__7884_ gnd vdd FILL
XFILL_3__14196_ gnd vdd FILL
XFILL_0__13036_ gnd vdd FILL
XFILL_1__11607_ gnd vdd FILL
XFILL_6__9110_ gnd vdd FILL
XFILL_2__13946_ gnd vdd FILL
XFILL_0__10248_ gnd vdd FILL
XFILL_1__12587_ gnd vdd FILL
XFILL_1__15375_ gnd vdd FILL
XFILL_3__7593_ gnd vdd FILL
XFILL_0__9623_ gnd vdd FILL
XFILL_4__14506_ gnd vdd FILL
XFILL_4__11718_ gnd vdd FILL
X_8162_ _8090_/A _7382_/CLK _8674_/R vdd _8162_/D gnd vdd DFFSR
XFILL_3__13147_ gnd vdd FILL
XFILL_4__15486_ gnd vdd FILL
XFILL_4__12698_ gnd vdd FILL
XFILL_3__10359_ gnd vdd FILL
XFILL_1__14326_ gnd vdd FILL
XFILL_1__11538_ gnd vdd FILL
XFILL_2__13877_ gnd vdd FILL
X_7113_ _7113_/A _7124_/A _7113_/C gnd _7153_/D vdd OAI21X1
XFILL_0__10179_ gnd vdd FILL
XFILL_0__9554_ gnd vdd FILL
XFILL_4__14437_ gnd vdd FILL
XFILL_2__15616_ gnd vdd FILL
XFILL_4__11649_ gnd vdd FILL
X_8093_ _8163_/Q gnd _8095_/A vdd INVX1
XFILL_5__13988_ gnd vdd FILL
XFILL_3__9263_ gnd vdd FILL
XFILL_2__12828_ gnd vdd FILL
XFILL_1__14257_ gnd vdd FILL
XFILL_1__11469_ gnd vdd FILL
XFILL_0__8505_ gnd vdd FILL
XSFILL104440x44050 gnd vdd FILL
XFILL_5__15727_ gnd vdd FILL
X_7044_ _7044_/A _7095_/B _7044_/C gnd _7130_/D vdd OAI21X1
XFILL_0__14987_ gnd vdd FILL
XFILL_0__9485_ gnd vdd FILL
XFILL_3__12029_ gnd vdd FILL
XFILL_4__14368_ gnd vdd FILL
XFILL_3__8214_ gnd vdd FILL
XFILL_1__13208_ gnd vdd FILL
XFILL_2__15547_ gnd vdd FILL
XSFILL33720x76050 gnd vdd FILL
XFILL_2__12759_ gnd vdd FILL
XFILL_1__14188_ gnd vdd FILL
XFILL_0__13938_ gnd vdd FILL
XFILL_4__13319_ gnd vdd FILL
XFILL_4__16107_ gnd vdd FILL
XFILL_5__15658_ gnd vdd FILL
XFILL_1__13139_ gnd vdd FILL
XFILL_4__14299_ gnd vdd FILL
XFILL_3__8145_ gnd vdd FILL
XSFILL89400x48050 gnd vdd FILL
XFILL_2__15478_ gnd vdd FILL
XFILL_0__13869_ gnd vdd FILL
XFILL_5__14609_ gnd vdd FILL
XFILL_4__16038_ gnd vdd FILL
XFILL_1__7160_ gnd vdd FILL
XSFILL99320x4050 gnd vdd FILL
XFILL_0__8367_ gnd vdd FILL
XFILL_5__15589_ gnd vdd FILL
XFILL_2__14429_ gnd vdd FILL
XFILL_3__8076_ gnd vdd FILL
X_8995_ _8995_/A gnd _8997_/A vdd INVX1
XFILL_0__15608_ gnd vdd FILL
XFILL_0__7318_ gnd vdd FILL
XFILL_1__7091_ gnd vdd FILL
X_7946_ _7944_/Y _7937_/B _7946_/C gnd _8028_/D vdd OAI21X1
XFILL_3__15719_ gnd vdd FILL
XFILL_0__15539_ gnd vdd FILL
XSFILL13640x43050 gnd vdd FILL
XFILL_0__7249_ gnd vdd FILL
X_7877_ _7821_/B _7877_/B gnd _7878_/C vdd NAND2X1
XSFILL59640x5050 gnd vdd FILL
XFILL_4__7840_ gnd vdd FILL
XSFILL13720x8050 gnd vdd FILL
X_9616_ _9616_/A _9615_/A _9616_/C gnd _9616_/Y vdd OAI21X1
XFILL_3__8978_ gnd vdd FILL
XFILL_1__9801_ gnd vdd FILL
X_9547_ _9548_/B _7499_/B gnd _9548_/C vdd NAND2X1
XFILL_4__9510_ gnd vdd FILL
XFILL_1__7993_ gnd vdd FILL
XFILL_3__7929_ gnd vdd FILL
XSFILL104520x24050 gnd vdd FILL
XFILL_5_BUFX2_insert233 gnd vdd FILL
XFILL_5_BUFX2_insert244 gnd vdd FILL
XSFILL33800x56050 gnd vdd FILL
XFILL_1__9732_ gnd vdd FILL
XFILL_5_BUFX2_insert255 gnd vdd FILL
XSFILL8760x22050 gnd vdd FILL
XFILL_1__6944_ gnd vdd FILL
XSFILL98760x44050 gnd vdd FILL
X_9478_ _9514_/A _9478_/B gnd _9479_/C vdd NAND2X1
XFILL_5_BUFX2_insert266 gnd vdd FILL
XFILL_5_BUFX2_insert277 gnd vdd FILL
X_10360_ _10360_/A _10405_/B _10360_/C gnd _10454_/D vdd OAI21X1
XFILL_5_BUFX2_insert288 gnd vdd FILL
XFILL_5_BUFX2_insert299 gnd vdd FILL
XFILL_4_BUFX2_insert900 gnd vdd FILL
X_8429_ _8379_/A _8429_/CLK _9203_/R vdd _8429_/D gnd vdd DFFSR
XFILL_1__9663_ gnd vdd FILL
XFILL_4_BUFX2_insert911 gnd vdd FILL
XFILL_4_BUFX2_insert922 gnd vdd FILL
XFILL_1__6875_ gnd vdd FILL
XFILL_4__9372_ gnd vdd FILL
XFILL_4_BUFX2_insert933 gnd vdd FILL
XFILL_1__8614_ gnd vdd FILL
X_10291_ _10325_/B _9779_/B gnd _10292_/C vdd NAND2X1
XFILL_4_BUFX2_insert944 gnd vdd FILL
XFILL_4_BUFX2_insert955 gnd vdd FILL
XFILL_4_BUFX2_insert966 gnd vdd FILL
XFILL_4__8323_ gnd vdd FILL
XFILL_1__9594_ gnd vdd FILL
XFILL111960x66050 gnd vdd FILL
XFILL_4_BUFX2_insert977 gnd vdd FILL
X_12030_ _12027_/Y _12030_/B _12029_/Y gnd _13110_/B vdd NAND3X1
XFILL_4_BUFX2_insert988 gnd vdd FILL
XFILL_4_BUFX2_insert999 gnd vdd FILL
XSFILL109240x36050 gnd vdd FILL
XSFILL13720x23050 gnd vdd FILL
XFILL_4__8254_ gnd vdd FILL
XSFILL79160x18050 gnd vdd FILL
XFILL112040x75050 gnd vdd FILL
XFILL_4__7205_ gnd vdd FILL
XFILL_1__8476_ gnd vdd FILL
XFILL_4__8185_ gnd vdd FILL
XFILL_1__7427_ gnd vdd FILL
X_13981_ _7447_/A gnd _15514_/B vdd INVX1
XFILL_2_BUFX2_insert101 gnd vdd FILL
X_15720_ _15720_/A _15720_/B gnd _15731_/B vdd NAND2X1
X_12932_ _12932_/Q _8180_/CLK _7391_/R vdd _12864_/Y gnd vdd DFFSR
XFILL_1__7358_ gnd vdd FILL
XFILL_4__7067_ gnd vdd FILL
X_15651_ _15651_/A _15651_/B _15651_/C gnd _12866_/B vdd AOI21X1
X_12863_ vdd _15610_/Y gnd _12864_/C vdd NAND2X1
XFILL_1_BUFX2_insert801 gnd vdd FILL
XFILL_1_BUFX2_insert812 gnd vdd FILL
XFILL_1__7289_ gnd vdd FILL
XFILL_5__6900_ gnd vdd FILL
X_14602_ _8126_/A gnd _14602_/Y vdd INVX1
XFILL_1_BUFX2_insert823 gnd vdd FILL
X_11814_ _11003_/Y _11484_/B _11349_/B _11236_/Y gnd _11815_/A vdd OAI22X1
XFILL_5__7880_ gnd vdd FILL
XFILL_2__9910_ gnd vdd FILL
XFILL_1_BUFX2_insert834 gnd vdd FILL
XFILL_1__9028_ gnd vdd FILL
X_15582_ _7709_/A _15969_/C _15581_/Y gnd _15582_/Y vdd AOI21X1
X_12794_ _12704_/A _12809_/CLK _12809_/R vdd _12794_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert845 gnd vdd FILL
XFILL_1_BUFX2_insert856 gnd vdd FILL
XFILL_1_BUFX2_insert867 gnd vdd FILL
X_14533_ _8248_/A gnd _14533_/Y vdd INVX1
XFILL_1_BUFX2_insert878 gnd vdd FILL
XFILL_2__10110_ gnd vdd FILL
XFILL_5__11270_ gnd vdd FILL
X_11745_ _11078_/Y _11270_/B gnd _11745_/Y vdd NAND2X1
XBUFX2_insert100 _15009_/Y gnd _15922_/C vdd BUFX2
XFILL_1_BUFX2_insert889 gnd vdd FILL
XFILL_2__11090_ gnd vdd FILL
XFILL_5__9550_ gnd vdd FILL
XFILL_4__7969_ gnd vdd FILL
X_14464_ _10219_/Q gnd _14464_/Y vdd INVX1
XFILL_3__11400_ gnd vdd FILL
XFILL_4__10951_ gnd vdd FILL
XFILL_2__10041_ gnd vdd FILL
X_11676_ _11046_/Y _11676_/B gnd _11677_/C vdd NAND2X1
XFILL_2__9772_ gnd vdd FILL
XFILL_5__8501_ gnd vdd FILL
XFILL_3__12380_ gnd vdd FILL
XFILL_0__11220_ gnd vdd FILL
X_16203_ _16203_/A _16203_/B _15338_/C gnd _12908_/B vdd AOI21X1
XFILL_1__10771_ gnd vdd FILL
XFILL_2__6984_ gnd vdd FILL
XFILL112120x55050 gnd vdd FILL
XFILL_5__9481_ gnd vdd FILL
X_13415_ _13414_/Y _13415_/B gnd _13427_/B vdd NOR2X1
XFILL_5__10152_ gnd vdd FILL
X_10627_ _10658_/B _7555_/B gnd _10627_/Y vdd NAND2X1
XFILL_4__13670_ gnd vdd FILL
XFILL_1__12510_ gnd vdd FILL
X_14395_ _9065_/Q gnd _15845_/B vdd INVX1
XFILL_2__8723_ gnd vdd FILL
XFILL_3__11331_ gnd vdd FILL
XSFILL64040x40050 gnd vdd FILL
XFILL_4__10882_ gnd vdd FILL
XFILL_4__9639_ gnd vdd FILL
XFILL_1__13490_ gnd vdd FILL
XFILL_0__11151_ gnd vdd FILL
X_16134_ _16225_/C _14750_/Y _16306_/C _14779_/Y gnd _16138_/B vdd OAI22X1
XFILL_4__12621_ gnd vdd FILL
X_13346_ _13312_/A gnd _13352_/B vdd INVX1
X_10558_ _10606_/Q gnd _10560_/A vdd INVX1
XFILL_2__13800_ gnd vdd FILL
XFILL_3__14050_ gnd vdd FILL
XFILL_5__14960_ gnd vdd FILL
XFILL_2__8654_ gnd vdd FILL
XFILL_1__12441_ gnd vdd FILL
XFILL_0__10102_ gnd vdd FILL
XFILL_3__11262_ gnd vdd FILL
XFILL_2__14780_ gnd vdd FILL
XFILL_2__11992_ gnd vdd FILL
XFILL_5__8363_ gnd vdd FILL
XFILL_0__11082_ gnd vdd FILL
XFILL_4__15340_ gnd vdd FILL
XFILL_3__13001_ gnd vdd FILL
X_16065_ _16064_/Y _16065_/B gnd _16065_/Y vdd NOR2X1
XFILL_5__13911_ gnd vdd FILL
X_13277_ _13326_/A _13262_/B gnd _13285_/B vdd NOR2X1
XFILL_2__7605_ gnd vdd FILL
X_10489_ _15122_/A gnd _10489_/Y vdd INVX1
XFILL_2__13731_ gnd vdd FILL
XFILL_1__15160_ gnd vdd FILL
XFILL_3__11193_ gnd vdd FILL
XFILL_5__14891_ gnd vdd FILL
XFILL_2__10943_ gnd vdd FILL
XFILL_2__8585_ gnd vdd FILL
XFILL_1__12372_ gnd vdd FILL
XFILL_0__10033_ gnd vdd FILL
XFILL_5__7314_ gnd vdd FILL
XFILL_0__14910_ gnd vdd FILL
X_15016_ _15644_/D gnd _16014_/C vdd INVX8
X_12228_ _12224_/A _12704_/A _12224_/C gnd _12228_/Y vdd NAND3X1
XFILL_4__11503_ gnd vdd FILL
XFILL_0__15890_ gnd vdd FILL
XFILL_5__13842_ gnd vdd FILL
XFILL_4__15271_ gnd vdd FILL
XFILL_2__16450_ gnd vdd FILL
XFILL_3__10144_ gnd vdd FILL
XFILL_4__12483_ gnd vdd FILL
XFILL_1__11323_ gnd vdd FILL
XFILL_1__14111_ gnd vdd FILL
XFILL_2__13662_ gnd vdd FILL
XFILL_1__15091_ gnd vdd FILL
XFILL_5__7245_ gnd vdd FILL
XFILL_0__14841_ gnd vdd FILL
XSFILL84200x53050 gnd vdd FILL
XFILL_2__10874_ gnd vdd FILL
XFILL_4__14222_ gnd vdd FILL
XFILL_2__15401_ gnd vdd FILL
X_12159_ _12159_/A _12134_/A _12159_/C gnd _12159_/Y vdd OAI21X1
XFILL_4__11434_ gnd vdd FILL
XFILL_5__13773_ gnd vdd FILL
XFILL_2__12613_ gnd vdd FILL
XSFILL104360x59050 gnd vdd FILL
XFILL_1__14042_ gnd vdd FILL
XFILL_3__14952_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1078 gnd vdd FILL
XFILL_2__7467_ gnd vdd FILL
XFILL_2__16381_ gnd vdd FILL
XFILL_1__11254_ gnd vdd FILL
XFILL_2__13593_ gnd vdd FILL
XFILL_0__14772_ gnd vdd FILL
XFILL_5__7176_ gnd vdd FILL
XFILL_0__11984_ gnd vdd FILL
XFILL_5__15512_ gnd vdd FILL
XFILL_0__9270_ gnd vdd FILL
XFILL_5__12724_ gnd vdd FILL
XFILL_6__10186_ gnd vdd FILL
XFILL_4__14153_ gnd vdd FILL
XFILL_2__9206_ gnd vdd FILL
XFILL_3__13903_ gnd vdd FILL
XFILL_2__15332_ gnd vdd FILL
XFILL_4__11365_ gnd vdd FILL
XFILL_3__14883_ gnd vdd FILL
XFILL_0__10935_ gnd vdd FILL
XFILL_0__13723_ gnd vdd FILL
XFILL_1__11185_ gnd vdd FILL
XFILL_4__13104_ gnd vdd FILL
XFILL_0__8221_ gnd vdd FILL
XFILL_4__10316_ gnd vdd FILL
X_15918_ _16438_/Q _15680_/B _15680_/C gnd _15927_/C vdd NAND3X1
XFILL_5__15443_ gnd vdd FILL
XFILL_5__12655_ gnd vdd FILL
XFILL_3__13834_ gnd vdd FILL
XFILL_6__14994_ gnd vdd FILL
XFILL_2__9137_ gnd vdd FILL
XFILL_4__14084_ gnd vdd FILL
XSFILL49080x17050 gnd vdd FILL
XFILL_1__10136_ gnd vdd FILL
XFILL_4__11296_ gnd vdd FILL
XFILL_2__15263_ gnd vdd FILL
XFILL_0__13654_ gnd vdd FILL
XFILL_2__12475_ gnd vdd FILL
XSFILL24520x34050 gnd vdd FILL
XSFILL23720x3050 gnd vdd FILL
XFILL_1__15993_ gnd vdd FILL
XFILL_6__6940_ gnd vdd FILL
X_7800_ _7798_/Y _7800_/B _7800_/C gnd _7894_/D vdd OAI21X1
XFILL_4__13035_ gnd vdd FILL
X_15849_ _15848_/Y _15849_/B gnd _15850_/B vdd NOR2X1
XFILL_5__11606_ gnd vdd FILL
XFILL_6__13945_ gnd vdd FILL
XSFILL64120x20050 gnd vdd FILL
XFILL_5__12586_ gnd vdd FILL
XFILL_5__15374_ gnd vdd FILL
XFILL_2__14214_ gnd vdd FILL
X_8780_ _8778_/Y _8714_/B _8779_/Y gnd _8818_/D vdd OAI21X1
XFILL_4__10247_ gnd vdd FILL
XFILL_0__12605_ gnd vdd FILL
XFILL_3__13765_ gnd vdd FILL
XFILL_2_BUFX2_insert690 gnd vdd FILL
XFILL_2__11426_ gnd vdd FILL
XFILL_3__10977_ gnd vdd FILL
XFILL_2__15194_ gnd vdd FILL
XFILL_1__10067_ gnd vdd FILL
XFILL_1__14944_ gnd vdd FILL
XFILL_0__16373_ gnd vdd FILL
XFILL_0__7103_ gnd vdd FILL
XFILL_0__13585_ gnd vdd FILL
XFILL_3__15504_ gnd vdd FILL
X_7731_ _7684_/B _9907_/B gnd _7732_/C vdd NAND2X1
XFILL_0__10797_ gnd vdd FILL
XFILL_5__14325_ gnd vdd FILL
XFILL_0__8083_ gnd vdd FILL
XFILL_5__11537_ gnd vdd FILL
XFILL_3__12716_ gnd vdd FILL
XFILL_2__8019_ gnd vdd FILL
XFILL112200x7050 gnd vdd FILL
XFILL_3__8901_ gnd vdd FILL
XSFILL13560x58050 gnd vdd FILL
XFILL_2__14145_ gnd vdd FILL
XFILL_4__10178_ gnd vdd FILL
XFILL_0__15324_ gnd vdd FILL
XFILL_3__9881_ gnd vdd FILL
XFILL_3__13696_ gnd vdd FILL
XFILL_2__11357_ gnd vdd FILL
XFILL_1__14875_ gnd vdd FILL
XFILL_0__7034_ gnd vdd FILL
XSFILL53960x63050 gnd vdd FILL
X_7662_ _7662_/Q _7662_/CLK _8430_/R vdd _7662_/D gnd vdd DFFSR
XFILL_5__14256_ gnd vdd FILL
XFILL_3__15435_ gnd vdd FILL
XFILL_5__11468_ gnd vdd FILL
XSFILL68760x23050 gnd vdd FILL
XFILL_3__8832_ gnd vdd FILL
XFILL_3__12647_ gnd vdd FILL
XFILL_2__10308_ gnd vdd FILL
XFILL_1__13826_ gnd vdd FILL
XFILL_0__15255_ gnd vdd FILL
XFILL_4__14986_ gnd vdd FILL
XFILL_2__11288_ gnd vdd FILL
XFILL_2__14076_ gnd vdd FILL
XFILL_0__12467_ gnd vdd FILL
XFILL_5_BUFX2_insert50 gnd vdd FILL
XFILL_5__13207_ gnd vdd FILL
XFILL_5_BUFX2_insert61 gnd vdd FILL
XFILL_6__15546_ gnd vdd FILL
X_9401_ _9401_/A _9657_/B gnd _9402_/C vdd NAND2X1
XFILL_5__10419_ gnd vdd FILL
XFILL_5__9748_ gnd vdd FILL
XFILL_6__12758_ gnd vdd FILL
XFILL_5_BUFX2_insert72 gnd vdd FILL
XFILL_5__14187_ gnd vdd FILL
XFILL_2__10239_ gnd vdd FILL
XFILL_3__15366_ gnd vdd FILL
XFILL_0__14206_ gnd vdd FILL
XFILL_5_BUFX2_insert83 gnd vdd FILL
X_7593_ _7593_/A gnd _7595_/A vdd INVX1
XFILL_2__13027_ gnd vdd FILL
XFILL_5__11399_ gnd vdd FILL
XFILL_4__13937_ gnd vdd FILL
XFILL_3__12578_ gnd vdd FILL
XFILL_3__8763_ gnd vdd FILL
XFILL_5_BUFX2_insert94 gnd vdd FILL
XFILL_0__11418_ gnd vdd FILL
XFILL_0__15186_ gnd vdd FILL
XFILL_1__13757_ gnd vdd FILL
XFILL_1__10969_ gnd vdd FILL
XFILL_5__9679_ gnd vdd FILL
XFILL_0__12398_ gnd vdd FILL
XFILL_5__13138_ gnd vdd FILL
XSFILL104440x39050 gnd vdd FILL
XFILL_3__14317_ gnd vdd FILL
X_9332_ _9332_/Q _7007_/CLK _9332_/R vdd _9332_/D gnd vdd DFFSR
XFILL_0__8985_ gnd vdd FILL
XFILL_3__7714_ gnd vdd FILL
XFILL_3__11529_ gnd vdd FILL
XFILL_1__12708_ gnd vdd FILL
XFILL_4__13868_ gnd vdd FILL
XFILL_3__15297_ gnd vdd FILL
XFILL_0__14137_ gnd vdd FILL
XSFILL8680x37050 gnd vdd FILL
XFILL_3__8694_ gnd vdd FILL
XFILL_0__11349_ gnd vdd FILL
XFILL_1__13688_ gnd vdd FILL
XFILL_0__7936_ gnd vdd FILL
X_9263_ _9321_/Q gnd _9263_/Y vdd INVX1
XFILL_4__15607_ gnd vdd FILL
XFILL_3__14248_ gnd vdd FILL
XFILL_4__13799_ gnd vdd FILL
XFILL_1__15427_ gnd vdd FILL
XFILL_4_BUFX2_insert229 gnd vdd FILL
XFILL_1__12639_ gnd vdd FILL
XFILL_0__14068_ gnd vdd FILL
XFILL_2__14978_ gnd vdd FILL
X_8214_ _8212_/Y _8244_/B _8214_/C gnd _8214_/Y vdd OAI21X1
XFILL_0__7867_ gnd vdd FILL
XSFILL48920x52050 gnd vdd FILL
XFILL_4__15538_ gnd vdd FILL
X_9194_ _9194_/Q _9194_/CLK _7914_/R vdd _9140_/Y gnd vdd DFFSR
XFILL_3__14179_ gnd vdd FILL
XFILL_0__13019_ gnd vdd FILL
XFILL_2__13929_ gnd vdd FILL
XFILL_1__15358_ gnd vdd FILL
XFILL_3__7576_ gnd vdd FILL
XFILL_0__9606_ gnd vdd FILL
X_8145_ _8133_/A _9041_/B gnd _8146_/C vdd NAND2X1
XFILL_3_BUFX2_insert907 gnd vdd FILL
XFILL_3_BUFX2_insert918 gnd vdd FILL
XFILL_0__7798_ gnd vdd FILL
XFILL_1__14309_ gnd vdd FILL
XFILL_4__15469_ gnd vdd FILL
XFILL_3_BUFX2_insert929 gnd vdd FILL
XSFILL49000x61050 gnd vdd FILL
XFILL_1__15289_ gnd vdd FILL
XFILL_1__8330_ gnd vdd FILL
XSFILL13640x38050 gnd vdd FILL
XFILL_0__9537_ gnd vdd FILL
X_8076_ _8118_/A _6924_/B gnd _8077_/C vdd NAND2X1
XFILL_3__9246_ gnd vdd FILL
X_7027_ _7027_/Q _7021_/CLK _9069_/R vdd _7027_/D gnd vdd DFFSR
XFILL_1__8261_ gnd vdd FILL
XFILL_0__9468_ gnd vdd FILL
XSFILL54120x52050 gnd vdd FILL
XFILL_1__7212_ gnd vdd FILL
XFILL_1__8192_ gnd vdd FILL
XFILL_3__8128_ gnd vdd FILL
XFILL_0__9399_ gnd vdd FILL
XFILL_4__9990_ gnd vdd FILL
XSFILL8760x17050 gnd vdd FILL
XFILL_1_BUFX2_insert108 gnd vdd FILL
XFILL_3__8059_ gnd vdd FILL
X_8978_ _9011_/A _7954_/B gnd _8979_/C vdd NAND2X1
XSFILL33960x10050 gnd vdd FILL
XFILL_1__7074_ gnd vdd FILL
X_7929_ _8023_/Q gnd _7929_/Y vdd INVX1
XFILL_4__8872_ gnd vdd FILL
XFILL_0_CLKBUF1_insert201 gnd vdd FILL
XSFILL18760x71050 gnd vdd FILL
XFILL_0_CLKBUF1_insert212 gnd vdd FILL
XSFILL23880x9050 gnd vdd FILL
XFILL_0_CLKBUF1_insert223 gnd vdd FILL
XSFILL8600x81050 gnd vdd FILL
XSFILL19240x78050 gnd vdd FILL
XFILL_4__7823_ gnd vdd FILL
XFILL_0_BUFX2_insert808 gnd vdd FILL
XFILL_0_BUFX2_insert819 gnd vdd FILL
X_11530_ _11527_/C _11574_/B _11529_/Y gnd _11530_/Y vdd OAI21X1
XFILL_1_BUFX2_insert1005 gnd vdd FILL
XFILL_1_BUFX2_insert1016 gnd vdd FILL
XFILL_4__7754_ gnd vdd FILL
XSFILL13720x18050 gnd vdd FILL
XFILL_1_BUFX2_insert1027 gnd vdd FILL
XFILL_1_BUFX2_insert1038 gnd vdd FILL
X_11461_ _11461_/A _11461_/B _11461_/C gnd _11466_/B vdd NAND3X1
XFILL_1_BUFX2_insert1049 gnd vdd FILL
XFILL_1__7976_ gnd vdd FILL
X_13200_ _13200_/Q _13180_/CLK _13180_/R vdd _13200_/D gnd vdd DFFSR
X_10412_ _10412_/A gnd _10414_/A vdd INVX1
XFILL_4__7685_ gnd vdd FILL
X_14180_ _10853_/Q _13884_/C _14180_/C _10531_/A gnd _14182_/A vdd AOI22X1
X_11392_ _11731_/B _11079_/Y _11392_/C gnd _11392_/Y vdd OAI21X1
XFILL_1__6927_ gnd vdd FILL
XFILL_4__9424_ gnd vdd FILL
XSFILL69240x8050 gnd vdd FILL
X_13131_ _13173_/A _13131_/B gnd _13132_/C vdd NAND2X1
XFILL_4_BUFX2_insert730 gnd vdd FILL
X_10343_ _10343_/Q _7400_/CLK _9704_/R vdd _10343_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert741 gnd vdd FILL
XFILL_1__9646_ gnd vdd FILL
XFILL_1__6858_ gnd vdd FILL
XFILL_4__9355_ gnd vdd FILL
XFILL_4_BUFX2_insert752 gnd vdd FILL
XFILL_4_BUFX2_insert763 gnd vdd FILL
XFILL_4_BUFX2_insert774 gnd vdd FILL
X_13062_ _6885_/A _8171_/CLK _8171_/R vdd _13062_/D gnd vdd DFFSR
X_10274_ _10272_/Y _10294_/A _10274_/C gnd _10340_/D vdd OAI21X1
XFILL_4_BUFX2_insert785 gnd vdd FILL
XFILL_2__8370_ gnd vdd FILL
XFILL_4_BUFX2_insert796 gnd vdd FILL
X_12013_ _12458_/B _12105_/B _12001_/C gnd gnd _12014_/C vdd AOI22X1
XFILL_4__9286_ gnd vdd FILL
XFILL_2__7321_ gnd vdd FILL
XFILL_1__8528_ gnd vdd FILL
XSFILL84120x68050 gnd vdd FILL
XSFILL43960x50 gnd vdd FILL
XSFILL18840x51050 gnd vdd FILL
XFILL_5__7030_ gnd vdd FILL
XFILL_4__8237_ gnd vdd FILL
XFILL_5__10770_ gnd vdd FILL
XFILL_1__8459_ gnd vdd FILL
XFILL_2__7252_ gnd vdd FILL
XFILL_3__10900_ gnd vdd FILL
XFILL_4__11150_ gnd vdd FILL
X_13964_ _9748_/A gnd _13966_/A vdd INVX1
XFILL_2__7183_ gnd vdd FILL
XFILL_4__7119_ gnd vdd FILL
XFILL_3__11880_ gnd vdd FILL
X_15703_ _7206_/A _15177_/B _16293_/A _7142_/Q gnd _15705_/A vdd AOI22X1
XFILL_4__8099_ gnd vdd FILL
XFILL_5__12440_ gnd vdd FILL
X_12915_ _12913_/Y vdd _12914_/Y gnd _12949_/D vdd OAI21X1
XFILL_5__8981_ gnd vdd FILL
XFILL_3__10831_ gnd vdd FILL
XFILL_4__11081_ gnd vdd FILL
X_13895_ _9311_/Q _13854_/B _13853_/B _8799_/Q gnd _13895_/Y vdd AOI22X1
XFILL_2__12260_ gnd vdd FILL
XFILL_0__10651_ gnd vdd FILL
XSFILL64040x35050 gnd vdd FILL
XFILL_5__7932_ gnd vdd FILL
X_15634_ _15634_/A _15633_/Y gnd _15641_/A vdd NOR2X1
XFILL_1__12990_ gnd vdd FILL
XFILL_6__13730_ gnd vdd FILL
X_12846_ _12844_/Y vdd _12846_/C gnd _12926_/D vdd OAI21X1
XFILL_5__12371_ gnd vdd FILL
XFILL_1_BUFX2_insert620 gnd vdd FILL
XFILL_4__10032_ gnd vdd FILL
XFILL_1_BUFX2_insert631 gnd vdd FILL
XFILL_3__13550_ gnd vdd FILL
XFILL_2__11211_ gnd vdd FILL
XFILL_3__10762_ gnd vdd FILL
XFILL_1_BUFX2_insert642 gnd vdd FILL
XFILL_2__12191_ gnd vdd FILL
XFILL_1__11941_ gnd vdd FILL
XFILL_0__13370_ gnd vdd FILL
XFILL_5__7863_ gnd vdd FILL
XFILL_1_BUFX2_insert653 gnd vdd FILL
XFILL_5__14110_ gnd vdd FILL
XFILL_5__11322_ gnd vdd FILL
XFILL_3__12501_ gnd vdd FILL
XFILL_5__15090_ gnd vdd FILL
X_15565_ _14068_/A _15565_/B gnd _15565_/Y vdd NOR2X1
XFILL_1_BUFX2_insert664 gnd vdd FILL
X_12777_ _12777_/A memoryOutData[27] gnd _12778_/C vdd NAND2X1
XFILL_4__14840_ gnd vdd FILL
XFILL_1_BUFX2_insert675 gnd vdd FILL
XFILL_2__11142_ gnd vdd FILL
XFILL_1_BUFX2_insert686 gnd vdd FILL
XFILL_0__12321_ gnd vdd FILL
XFILL_3__13481_ gnd vdd FILL
XFILL_1__11872_ gnd vdd FILL
XFILL_5__9602_ gnd vdd FILL
XFILL_3__10693_ gnd vdd FILL
XFILL_1__14660_ gnd vdd FILL
X_14516_ _9272_/A gnd _14518_/A vdd INVX1
XFILL_5__14041_ gnd vdd FILL
XFILL_1_BUFX2_insert697 gnd vdd FILL
XFILL_3__15220_ gnd vdd FILL
XFILL_6__16380_ gnd vdd FILL
X_11728_ _11447_/Y _11256_/Y _11050_/Y gnd _11728_/Y vdd OAI21X1
XFILL_5__11253_ gnd vdd FILL
XFILL_3__12432_ gnd vdd FILL
XFILL_6__13592_ gnd vdd FILL
X_15496_ _15496_/A _15495_/Y gnd _15496_/Y vdd NOR2X1
XFILL_1__13611_ gnd vdd FILL
XFILL_4__11983_ gnd vdd FILL
XFILL_0__15040_ gnd vdd FILL
XFILL_2__15950_ gnd vdd FILL
XFILL_2__11073_ gnd vdd FILL
XFILL_4__14771_ gnd vdd FILL
XFILL_5__9533_ gnd vdd FILL
XFILL_0__12252_ gnd vdd FILL
XFILL_1__10823_ gnd vdd FILL
XFILL_1__14591_ gnd vdd FILL
XSFILL84200x48050 gnd vdd FILL
X_14447_ _9194_/Q _14868_/D _14739_/C _15878_/A gnd _14447_/Y vdd AOI22X1
XFILL_4__10934_ gnd vdd FILL
XFILL_2__10024_ gnd vdd FILL
XSFILL18920x31050 gnd vdd FILL
X_11659_ _11656_/Y _11059_/Y _11044_/A gnd _11660_/B vdd OAI21X1
XFILL_5__11184_ gnd vdd FILL
XFILL_3__15151_ gnd vdd FILL
XFILL_4__13722_ gnd vdd FILL
XFILL_2__14901_ gnd vdd FILL
XFILL_3__12363_ gnd vdd FILL
XFILL_1__16330_ gnd vdd FILL
XFILL_2__9755_ gnd vdd FILL
XFILL_0__11203_ gnd vdd FILL
XFILL_2__6967_ gnd vdd FILL
XFILL_1__10754_ gnd vdd FILL
XFILL_1__13542_ gnd vdd FILL
XFILL_2__15881_ gnd vdd FILL
XFILL_5__9464_ gnd vdd FILL
XFILL_0__12183_ gnd vdd FILL
XFILL_5__10135_ gnd vdd FILL
XFILL_3__14102_ gnd vdd FILL
XSFILL59000x24050 gnd vdd FILL
XFILL_4__13653_ gnd vdd FILL
XFILL_2__8706_ gnd vdd FILL
XFILL_6__12474_ gnd vdd FILL
X_14378_ _9449_/Q _13883_/B _14378_/C gnd _14379_/B vdd AOI21X1
XFILL_3__11314_ gnd vdd FILL
XFILL_0__8770_ gnd vdd FILL
XFILL_5__15992_ gnd vdd FILL
XFILL_2__14832_ gnd vdd FILL
XFILL_3__15082_ gnd vdd FILL
XFILL_3__12294_ gnd vdd FILL
XFILL_0__11134_ gnd vdd FILL
XFILL_1__16261_ gnd vdd FILL
XFILL_1__10685_ gnd vdd FILL
XFILL_1__13473_ gnd vdd FILL
X_16117_ _14708_/A _15924_/B _15644_/D _16117_/D gnd _16121_/A vdd OAI22X1
XFILL_2__6898_ gnd vdd FILL
X_13329_ _13259_/C _13328_/Y gnd _13329_/Y vdd NOR2X1
XFILL_4__12604_ gnd vdd FILL
XFILL_5__9395_ gnd vdd FILL
XFILL_6__11425_ gnd vdd FILL
XFILL_0__7721_ gnd vdd FILL
XFILL_6__15193_ gnd vdd FILL
XFILL_3__14033_ gnd vdd FILL
XFILL_5__14943_ gnd vdd FILL
XFILL_5__10066_ gnd vdd FILL
XFILL_2__8637_ gnd vdd FILL
XFILL_1__15212_ gnd vdd FILL
XFILL_4__16372_ gnd vdd FILL
XFILL_3__7430_ gnd vdd FILL
XFILL_4__13584_ gnd vdd FILL
XFILL_3__11245_ gnd vdd FILL
XFILL_1__12424_ gnd vdd FILL
XFILL_4__10796_ gnd vdd FILL
XFILL_2__14763_ gnd vdd FILL
XFILL_2__11975_ gnd vdd FILL
XFILL_1__16192_ gnd vdd FILL
XFILL_0__15942_ gnd vdd FILL
XFILL_5__8346_ gnd vdd FILL
XFILL_0__11065_ gnd vdd FILL
X_16048_ _16048_/A _16089_/B gnd _16048_/Y vdd NOR2X1
XFILL_4__15323_ gnd vdd FILL
XSFILL64120x15050 gnd vdd FILL
XFILL_5__14874_ gnd vdd FILL
XFILL_2__13714_ gnd vdd FILL
XFILL_2__10926_ gnd vdd FILL
XFILL_0__10016_ gnd vdd FILL
XFILL_2__8568_ gnd vdd FILL
XFILL_1__12355_ gnd vdd FILL
XFILL_3__7361_ gnd vdd FILL
XFILL_1__15143_ gnd vdd FILL
XFILL_3__11176_ gnd vdd FILL
XFILL_2__14694_ gnd vdd FILL
XSFILL24120x31050 gnd vdd FILL
XFILL_5__8277_ gnd vdd FILL
XFILL_0__15873_ gnd vdd FILL
XFILL_3__9100_ gnd vdd FILL
XFILL_5__13825_ gnd vdd FILL
XFILL_4__15254_ gnd vdd FILL
XFILL_6__11287_ gnd vdd FILL
XFILL_3__10127_ gnd vdd FILL
XFILL_4__12466_ gnd vdd FILL
XFILL_0__7583_ gnd vdd FILL
XFILL_1__11306_ gnd vdd FILL
XSFILL39720x10050 gnd vdd FILL
XFILL_2__13645_ gnd vdd FILL
XFILL_5__7228_ gnd vdd FILL
XFILL_3__15984_ gnd vdd FILL
XFILL_0__14824_ gnd vdd FILL
XFILL_1__15074_ gnd vdd FILL
XFILL_3__7292_ gnd vdd FILL
XFILL_2__8499_ gnd vdd FILL
XFILL_1__12286_ gnd vdd FILL
XSFILL89320x81050 gnd vdd FILL
XFILL_4__14205_ gnd vdd FILL
XFILL_6__10238_ gnd vdd FILL
XSFILL53960x58050 gnd vdd FILL
XFILL_4__11417_ gnd vdd FILL
X_9950_ _9870_/A _7902_/CLK _7150_/R vdd _9950_/D gnd vdd DFFSR
XFILL_4__15185_ gnd vdd FILL
XFILL_5__13756_ gnd vdd FILL
XFILL_3__9031_ gnd vdd FILL
XSFILL3560x22050 gnd vdd FILL
XFILL_5__10968_ gnd vdd FILL
XFILL_3__10058_ gnd vdd FILL
XFILL_2__16364_ gnd vdd FILL
XFILL_4__12397_ gnd vdd FILL
XFILL_1__14025_ gnd vdd FILL
XFILL_3__14935_ gnd vdd FILL
XFILL_1__11237_ gnd vdd FILL
XFILL_2__13576_ gnd vdd FILL
XFILL_2__10788_ gnd vdd FILL
XFILL_0__11967_ gnd vdd FILL
XFILL_5__7159_ gnd vdd FILL
XFILL_0__14755_ gnd vdd FILL
XFILL_5__12707_ gnd vdd FILL
XFILL_0__9253_ gnd vdd FILL
XFILL_4__14136_ gnd vdd FILL
X_8901_ _8902_/B _9797_/B gnd _8901_/Y vdd NAND2X1
XFILL_2__15315_ gnd vdd FILL
XSFILL28760x34050 gnd vdd FILL
XFILL_4__11348_ gnd vdd FILL
XFILL_3__14866_ gnd vdd FILL
XFILL_5__10899_ gnd vdd FILL
XFILL_2__12527_ gnd vdd FILL
X_9881_ _9881_/A _9868_/A _9881_/C gnd _9953_/D vdd OAI21X1
XFILL_5__13687_ gnd vdd FILL
XFILL_0__10918_ gnd vdd FILL
XSFILL54040x67050 gnd vdd FILL
XFILL_2__16295_ gnd vdd FILL
XFILL_0__13706_ gnd vdd FILL
XFILL_1__11168_ gnd vdd FILL
XFILL_0__8204_ gnd vdd FILL
XFILL_0__11898_ gnd vdd FILL
XFILL_0__14686_ gnd vdd FILL
XFILL_5__15426_ gnd vdd FILL
X_8832_ _8896_/B _8832_/B gnd _8832_/Y vdd NAND2X1
XFILL_5__12638_ gnd vdd FILL
XSFILL94440x72050 gnd vdd FILL
XFILL_3__13817_ gnd vdd FILL
XBUFX2_insert0 _12381_/Y gnd _8091_/B vdd BUFX2
XFILL_4__14067_ gnd vdd FILL
XFILL_2__15246_ gnd vdd FILL
XFILL_1__10119_ gnd vdd FILL
XFILL_4__11279_ gnd vdd FILL
XFILL_3__14797_ gnd vdd FILL
XFILL_2__12458_ gnd vdd FILL
XFILL_1__15976_ gnd vdd FILL
XFILL_0__13637_ gnd vdd FILL
XFILL_1__11099_ gnd vdd FILL
XFILL_4__13018_ gnd vdd FILL
XFILL_0__8135_ gnd vdd FILL
XFILL_5__15357_ gnd vdd FILL
XFILL_5__12569_ gnd vdd FILL
X_8763_ _8813_/Q gnd _8765_/A vdd INVX1
XFILL_3__13748_ gnd vdd FILL
XFILL_2__11409_ gnd vdd FILL
XSFILL33880x25050 gnd vdd FILL
XFILL_3__9933_ gnd vdd FILL
XFILL_2__15177_ gnd vdd FILL
XFILL_1__14927_ gnd vdd FILL
XFILL_2__12389_ gnd vdd FILL
XFILL_0__16356_ gnd vdd FILL
XFILL_0__13568_ gnd vdd FILL
XFILL_5__14308_ gnd vdd FILL
XFILL_0__8066_ gnd vdd FILL
X_7714_ _7714_/A _7684_/B _7713_/Y gnd _7714_/Y vdd OAI21X1
XFILL_2__14128_ gnd vdd FILL
XFILL_5__15288_ gnd vdd FILL
XFILL_6_BUFX2_insert858 gnd vdd FILL
XFILL_0__15307_ gnd vdd FILL
XFILL_3__13679_ gnd vdd FILL
XFILL_3__9864_ gnd vdd FILL
XFILL_0__12519_ gnd vdd FILL
XSFILL48920x47050 gnd vdd FILL
X_8694_ _8790_/Q gnd _8694_/Y vdd INVX1
XFILL_1__14858_ gnd vdd FILL
XFILL_0__16287_ gnd vdd FILL
XFILL_0__13499_ gnd vdd FILL
XFILL_5__14239_ gnd vdd FILL
XFILL_3__15418_ gnd vdd FILL
X_7645_ _7645_/Q _7261_/CLK _8669_/R vdd _7645_/D gnd vdd DFFSR
XFILL_1__13809_ gnd vdd FILL
XFILL_2__14059_ gnd vdd FILL
XFILL_4__14969_ gnd vdd FILL
XFILL_3__16398_ gnd vdd FILL
XFILL_0__15238_ gnd vdd FILL
XFILL_3__9795_ gnd vdd FILL
XFILL_1__14789_ gnd vdd FILL
XSFILL49000x56050 gnd vdd FILL
XFILL_1__7830_ gnd vdd FILL
XFILL_3__15349_ gnd vdd FILL
X_7576_ _7577_/B _8600_/B gnd _7576_/Y vdd NAND2X1
XSFILL89400x61050 gnd vdd FILL
XFILL_3__8746_ gnd vdd FILL
XFILL_0__15169_ gnd vdd FILL
X_9315_ _9245_/A _7791_/CLK _9711_/R vdd _9315_/D gnd vdd DFFSR
XSFILL93640x24050 gnd vdd FILL
XFILL_0__8968_ gnd vdd FILL
XFILL_1__7761_ gnd vdd FILL
XFILL_4__7470_ gnd vdd FILL
XSFILL28840x14050 gnd vdd FILL
XFILL_1__9500_ gnd vdd FILL
XFILL_6__8386_ gnd vdd FILL
X_9246_ _9282_/A _9246_/B gnd _9246_/Y vdd NAND2X1
XFILL_1__7692_ gnd vdd FILL
XFILL_3__7628_ gnd vdd FILL
XFILL_0__8899_ gnd vdd FILL
XFILL_6__7337_ gnd vdd FILL
X_9177_ _9177_/Q _7129_/CLK _8542_/R vdd _9089_/Y gnd vdd DFFSR
XFILL_4__9140_ gnd vdd FILL
XFILL_3_BUFX2_insert704 gnd vdd FILL
XFILL_3__7559_ gnd vdd FILL
XFILL_3_BUFX2_insert715 gnd vdd FILL
X_8128_ _8128_/A _8079_/A _8127_/Y gnd _8174_/D vdd OAI21X1
XFILL_3_BUFX2_insert726 gnd vdd FILL
XFILL_3_BUFX2_insert737 gnd vdd FILL
XFILL_1__9362_ gnd vdd FILL
XFILL_3_BUFX2_insert748 gnd vdd FILL
XFILL_6__9007_ gnd vdd FILL
XFILL_3_BUFX2_insert759 gnd vdd FILL
XFILL_1__8313_ gnd vdd FILL
X_8059_ _8057_/Y _8107_/B _8059_/C gnd _8151_/D vdd OAI21X1
XFILL_1__9293_ gnd vdd FILL
XSFILL8600x76050 gnd vdd FILL
XFILL_3__9229_ gnd vdd FILL
XFILL_1_BUFX2_insert70 gnd vdd FILL
XSFILL39000x6050 gnd vdd FILL
XSFILL33000x50050 gnd vdd FILL
XFILL_1_BUFX2_insert81 gnd vdd FILL
XFILL_1_BUFX2_insert92 gnd vdd FILL
XFILL_1__8244_ gnd vdd FILL
X_10961_ _12773_/A _10969_/C gnd _10962_/B vdd NOR2X1
XSFILL23880x57050 gnd vdd FILL
X_12700_ _12700_/A _10944_/C _12700_/C gnd _12700_/Y vdd OAI21X1
X_13680_ _13678_/Y _13680_/B _14496_/A _13679_/Y gnd _13680_/Y vdd OAI22X1
X_10892_ _12695_/A _10883_/Y _10892_/C gnd _10895_/A vdd NOR3X1
X_12631_ vdd memoryOutData[21] gnd _12632_/C vdd NAND2X1
XSFILL13640x50 gnd vdd FILL
XFILL_1__7057_ gnd vdd FILL
XFILL_4__8855_ gnd vdd FILL
XFILL_0_BUFX2_insert605 gnd vdd FILL
X_15350_ _15383_/A _7645_/Q _7435_/A _15383_/D gnd _15354_/B vdd AOI22X1
XSFILL79960x50050 gnd vdd FILL
XSFILL79160x31050 gnd vdd FILL
XFILL_0_BUFX2_insert616 gnd vdd FILL
X_12562_ _11969_/B _13180_/CLK _13180_/R vdd _12522_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert627 gnd vdd FILL
XFILL_2__7870_ gnd vdd FILL
XFILL_0_BUFX2_insert638 gnd vdd FILL
XFILL_4__7806_ gnd vdd FILL
X_14301_ _14301_/A _13775_/B _13456_/A _14299_/Y gnd _14305_/A vdd OAI22X1
XFILL_0_BUFX2_insert649 gnd vdd FILL
X_11513_ _11513_/A _11513_/B _11553_/C gnd _11514_/A vdd OAI21X1
XFILL_4__8786_ gnd vdd FILL
X_15281_ _9435_/Q _15114_/C _15764_/C gnd _15282_/C vdd NAND3X1
X_12493_ _12553_/Q gnd _12493_/Y vdd INVX1
XFILL_4__7737_ gnd vdd FILL
X_14232_ _7014_/Q gnd _14232_/Y vdd INVX1
XSFILL18840x46050 gnd vdd FILL
X_11444_ _11025_/A _12129_/Y gnd _11444_/Y vdd XNOR2X1
XFILL_2__9540_ gnd vdd FILL
XFILL_1__7959_ gnd vdd FILL
X_14163_ _7456_/A gnd _14164_/D vdd INVX1
XSFILL69080x83050 gnd vdd FILL
XFILL_4__10650_ gnd vdd FILL
X_11375_ _11373_/Y _12117_/Y _11374_/Y _11238_/Y gnd _11839_/A vdd OAI22X1
XFILL_2__9471_ gnd vdd FILL
XFILL_4__9407_ gnd vdd FILL
XFILL_5__8200_ gnd vdd FILL
X_13114_ _13114_/A _13108_/B _13113_/Y gnd _13114_/Y vdd OAI21X1
X_10326_ _13452_/A _8818_/CLK _7270_/R vdd _10232_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert560 gnd vdd FILL
XFILL_4__7599_ gnd vdd FILL
XFILL_5__11940_ gnd vdd FILL
XFILL_4_BUFX2_insert571 gnd vdd FILL
XFILL_1__9629_ gnd vdd FILL
X_14094_ _15590_/A _14868_/A _14283_/C _9955_/Q gnd _14095_/B vdd AOI22X1
XFILL_3__11030_ gnd vdd FILL
XFILL_4__10581_ gnd vdd FILL
XFILL_4_BUFX2_insert582 gnd vdd FILL
XFILL_5__8131_ gnd vdd FILL
XFILL_4__9338_ gnd vdd FILL
XFILL_2__11760_ gnd vdd FILL
XFILL_4_BUFX2_insert593 gnd vdd FILL
X_13045_ vdd _13045_/B gnd _13045_/Y vdd NAND2X1
XFILL_4__12320_ gnd vdd FILL
X_10257_ _13920_/A gnd _10259_/A vdd INVX1
XFILL_2__8353_ gnd vdd FILL
XFILL_1__12140_ gnd vdd FILL
XFILL_5__11871_ gnd vdd FILL
XFILL_4__9269_ gnd vdd FILL
XFILL_0__12870_ gnd vdd FILL
XFILL_5__8062_ gnd vdd FILL
XFILL_2__11691_ gnd vdd FILL
XFILL_5__13610_ gnd vdd FILL
XFILL_6__11072_ gnd vdd FILL
XFILL_2__7304_ gnd vdd FILL
X_10188_ _10188_/A _10166_/A _10188_/C gnd _10226_/D vdd OAI21X1
XFILL_5__10822_ gnd vdd FILL
XFILL_4__12251_ gnd vdd FILL
XFILL_5__14590_ gnd vdd FILL
XFILL_2__13430_ gnd vdd FILL
XSFILL79240x11050 gnd vdd FILL
XFILL_1__12071_ gnd vdd FILL
XFILL_3__12981_ gnd vdd FILL
XFILL_2__10642_ gnd vdd FILL
XFILL_0__11821_ gnd vdd FILL
XSFILL3480x37050 gnd vdd FILL
XFILL_4__11202_ gnd vdd FILL
XFILL_5__10753_ gnd vdd FILL
XFILL_5__13541_ gnd vdd FILL
XFILL_3__14720_ gnd vdd FILL
XFILL_3__11932_ gnd vdd FILL
X_14996_ _12812_/Q _15220_/B gnd _15024_/C vdd NOR2X1
XFILL_4__12182_ gnd vdd FILL
XFILL_2__7235_ gnd vdd FILL
XFILL_1__11022_ gnd vdd FILL
XFILL_2__13361_ gnd vdd FILL
XFILL_2__10573_ gnd vdd FILL
XFILL_0__14540_ gnd vdd FILL
XSFILL28680x49050 gnd vdd FILL
XFILL_0__11752_ gnd vdd FILL
XSFILL114440x20050 gnd vdd FILL
XFILL_2__15100_ gnd vdd FILL
X_13947_ _9184_/Q gnd _15461_/A vdd INVX1
XFILL_4__11133_ gnd vdd FILL
XFILL_5__16260_ gnd vdd FILL
XFILL_5__10684_ gnd vdd FILL
XFILL_5__13472_ gnd vdd FILL
XFILL_2__12312_ gnd vdd FILL
XFILL_3__14651_ gnd vdd FILL
XFILL_0__10703_ gnd vdd FILL
XFILL_1__15830_ gnd vdd FILL
XFILL_3__11863_ gnd vdd FILL
XFILL_2__16080_ gnd vdd FILL
XFILL_2__7166_ gnd vdd FILL
XSFILL18920x26050 gnd vdd FILL
XFILL_2__13292_ gnd vdd FILL
XFILL_0__14471_ gnd vdd FILL
XFILL_5__15211_ gnd vdd FILL
XFILL_0__11683_ gnd vdd FILL
XFILL_3__13602_ gnd vdd FILL
XFILL_5__8964_ gnd vdd FILL
XFILL_5__12423_ gnd vdd FILL
XFILL_3__10814_ gnd vdd FILL
X_13878_ _9742_/A gnd _13879_/A vdd INVX1
XFILL_5__16191_ gnd vdd FILL
XFILL_2__15031_ gnd vdd FILL
XFILL_4__15941_ gnd vdd FILL
XSFILL59800x38050 gnd vdd FILL
XFILL_4__11064_ gnd vdd FILL
XSFILL59000x19050 gnd vdd FILL
XFILL_3__14582_ gnd vdd FILL
XFILL_0__16210_ gnd vdd FILL
XFILL_0__13422_ gnd vdd FILL
XFILL_2__12243_ gnd vdd FILL
XFILL_0__10634_ gnd vdd FILL
XFILL_2__7097_ gnd vdd FILL
XFILL_3__11794_ gnd vdd FILL
XSFILL99400x24050 gnd vdd FILL
XFILL_1__15761_ gnd vdd FILL
XFILL_1__12973_ gnd vdd FILL
XSFILL69160x63050 gnd vdd FILL
X_15617_ _8420_/Q _15978_/B _15380_/C _9888_/A gnd _15618_/B vdd AOI22X1
XFILL_5__8895_ gnd vdd FILL
XFILL_5__12354_ gnd vdd FILL
XFILL_6__10925_ gnd vdd FILL
XFILL_3__16321_ gnd vdd FILL
XFILL_1_BUFX2_insert450 gnd vdd FILL
XFILL_4__10015_ gnd vdd FILL
XFILL_5__15142_ gnd vdd FILL
X_12829_ _12829_/A gnd _12831_/A vdd INVX1
XFILL_1_BUFX2_insert461 gnd vdd FILL
XFILL_3__13533_ gnd vdd FILL
XFILL_1__14712_ gnd vdd FILL
XFILL_4__15872_ gnd vdd FILL
XFILL_3__6930_ gnd vdd FILL
XFILL_3__10745_ gnd vdd FILL
XFILL_0__13353_ gnd vdd FILL
XFILL_1__11924_ gnd vdd FILL
XFILL_1_BUFX2_insert472 gnd vdd FILL
XFILL_2__12174_ gnd vdd FILL
XFILL_0__16141_ gnd vdd FILL
XFILL_5__7846_ gnd vdd FILL
XFILL_1__15692_ gnd vdd FILL
XFILL_1_BUFX2_insert483 gnd vdd FILL
XFILL_0__10565_ gnd vdd FILL
XFILL_5__11305_ gnd vdd FILL
X_15548_ _15546_/Y _15548_/B _15548_/C gnd _15549_/A vdd NAND3X1
XFILL_1_BUFX2_insert494 gnd vdd FILL
XFILL_0__9940_ gnd vdd FILL
XSFILL104360x72050 gnd vdd FILL
XFILL_4__14823_ gnd vdd FILL
XFILL_5__15073_ gnd vdd FILL
XFILL_3__16252_ gnd vdd FILL
XFILL_5__12285_ gnd vdd FILL
XFILL_3__13464_ gnd vdd FILL
XFILL_0__12304_ gnd vdd FILL
XFILL_2__11125_ gnd vdd FILL
XFILL_1__14643_ gnd vdd FILL
XFILL_3__6861_ gnd vdd FILL
XFILL_0__16072_ gnd vdd FILL
XFILL_3__10676_ gnd vdd FILL
XFILL_0__13284_ gnd vdd FILL
XFILL_1__11855_ gnd vdd FILL
XFILL_0__10496_ gnd vdd FILL
XFILL_3__15203_ gnd vdd FILL
XSFILL74280x54050 gnd vdd FILL
XFILL_5__14024_ gnd vdd FILL
X_7430_ _7430_/A _7558_/B gnd _7431_/C vdd NAND2X1
XFILL_5__11236_ gnd vdd FILL
XFILL_0__9871_ gnd vdd FILL
XFILL_3__12415_ gnd vdd FILL
XFILL_3__8600_ gnd vdd FILL
XBUFX2_insert1007 _10928_/Y gnd _12216_/B vdd BUFX2
X_15479_ _15479_/A _16151_/B _16247_/C _15479_/D gnd _15480_/C vdd OAI22X1
XFILL_2__9807_ gnd vdd FILL
XFILL_3__16183_ gnd vdd FILL
XBUFX2_insert1018 _15054_/Y gnd _15646_/D vdd BUFX2
XFILL_4__11966_ gnd vdd FILL
XFILL_2__15933_ gnd vdd FILL
XFILL_0__15023_ gnd vdd FILL
XFILL_2__11056_ gnd vdd FILL
XFILL_4__14754_ gnd vdd FILL
XFILL_1__10806_ gnd vdd FILL
XBUFX2_insert1029 _13333_/Y gnd _9228_/A vdd BUFX2
XFILL_3__13395_ gnd vdd FILL
XFILL_0__12235_ gnd vdd FILL
XFILL_2__7999_ gnd vdd FILL
XFILL_1__14574_ gnd vdd FILL
XFILL_5__9516_ gnd vdd FILL
XFILL_0__8822_ gnd vdd FILL
XFILL_1__11786_ gnd vdd FILL
XSFILL89320x76050 gnd vdd FILL
XFILL_4__10917_ gnd vdd FILL
XSFILL49080x30050 gnd vdd FILL
X_7361_ _7361_/A gnd _7361_/Y vdd INVX1
XFILL_3__15134_ gnd vdd FILL
XFILL_4__13705_ gnd vdd FILL
XFILL_5__11167_ gnd vdd FILL
XFILL_2__9738_ gnd vdd FILL
XFILL_2__10007_ gnd vdd FILL
XFILL_3__8531_ gnd vdd FILL
XFILL_3__12346_ gnd vdd FILL
XFILL_1__16313_ gnd vdd FILL
XSFILL3560x17050 gnd vdd FILL
XFILL_4__11897_ gnd vdd FILL
XFILL_2__15864_ gnd vdd FILL
XFILL_4__14685_ gnd vdd FILL
XFILL_1__13525_ gnd vdd FILL
XFILL_0__12166_ gnd vdd FILL
X_9100_ _9101_/B _9100_/B gnd _9100_/Y vdd NAND2X1
XFILL_6__15245_ gnd vdd FILL
XFILL_5__10118_ gnd vdd FILL
XFILL_0__8753_ gnd vdd FILL
XFILL_4__13636_ gnd vdd FILL
XFILL_5__15975_ gnd vdd FILL
XFILL_2__14815_ gnd vdd FILL
XFILL_3__15065_ gnd vdd FILL
XFILL_5__11098_ gnd vdd FILL
X_7292_ _7292_/A gnd _7292_/Y vdd INVX1
XFILL_3__8462_ gnd vdd FILL
XFILL_1__16244_ gnd vdd FILL
XFILL_2__9669_ gnd vdd FILL
XFILL_3__12277_ gnd vdd FILL
XFILL_0__11117_ gnd vdd FILL
XFILL_1__13456_ gnd vdd FILL
XFILL_2__15795_ gnd vdd FILL
XFILL_1__10668_ gnd vdd FILL
XFILL_5__9378_ gnd vdd FILL
XFILL_0__7704_ gnd vdd FILL
XFILL_0__12097_ gnd vdd FILL
X_9031_ _9031_/A gnd _9033_/A vdd INVX1
XFILL_3__14016_ gnd vdd FILL
XFILL_5__10049_ gnd vdd FILL
XFILL_5__14926_ gnd vdd FILL
XSFILL94440x67050 gnd vdd FILL
XFILL_4__16355_ gnd vdd FILL
XFILL_4__13567_ gnd vdd FILL
XFILL_3__11228_ gnd vdd FILL
XFILL_1__12407_ gnd vdd FILL
XFILL_4__10779_ gnd vdd FILL
XSFILL49000x1050 gnd vdd FILL
XFILL_2__14746_ gnd vdd FILL
XFILL_0__15925_ gnd vdd FILL
XFILL_5__8329_ gnd vdd FILL
XFILL_1__16175_ gnd vdd FILL
XFILL_2__11958_ gnd vdd FILL
XFILL_0__11048_ gnd vdd FILL
XFILL_3__8393_ gnd vdd FILL
XFILL_1__13387_ gnd vdd FILL
XFILL_4__15306_ gnd vdd FILL
XFILL_0__7635_ gnd vdd FILL
XFILL_5__14857_ gnd vdd FILL
XFILL_4__12518_ gnd vdd FILL
XFILL_2__10909_ gnd vdd FILL
XSFILL69240x43050 gnd vdd FILL
XFILL_4__16286_ gnd vdd FILL
XFILL_3__7344_ gnd vdd FILL
XFILL_4__13498_ gnd vdd FILL
XFILL_3__11159_ gnd vdd FILL
XFILL_1__15126_ gnd vdd FILL
XFILL_1__12338_ gnd vdd FILL
XFILL_2__14677_ gnd vdd FILL
XFILL_6__7053_ gnd vdd FILL
XFILL_2__11889_ gnd vdd FILL
XFILL_0__15856_ gnd vdd FILL
XFILL_5__13808_ gnd vdd FILL
XFILL_6__14058_ gnd vdd FILL
XFILL_0__7566_ gnd vdd FILL
XFILL_4__12449_ gnd vdd FILL
XFILL_4__15237_ gnd vdd FILL
XFILL_2__16416_ gnd vdd FILL
XFILL_2__13628_ gnd vdd FILL
XFILL_5__14788_ gnd vdd FILL
XFILL_0__14807_ gnd vdd FILL
XFILL_1__15057_ gnd vdd FILL
XFILL_3__15967_ gnd vdd FILL
XFILL_1__12269_ gnd vdd FILL
XSFILL104440x52050 gnd vdd FILL
XFILL_0__15787_ gnd vdd FILL
X_9933_ _9933_/A gnd _9933_/Y vdd INVX1
XFILL_3__9014_ gnd vdd FILL
XFILL_0__12999_ gnd vdd FILL
XSFILL88520x28050 gnd vdd FILL
XFILL_5__13739_ gnd vdd FILL
XFILL_4__15168_ gnd vdd FILL
XFILL_2__16347_ gnd vdd FILL
XFILL_1__14008_ gnd vdd FILL
XFILL_0__7497_ gnd vdd FILL
XFILL_3__14918_ gnd vdd FILL
XSFILL9160x57050 gnd vdd FILL
XFILL_2__13559_ gnd vdd FILL
XSFILL98680x72050 gnd vdd FILL
XFILL_3__15898_ gnd vdd FILL
XFILL_0__14738_ gnd vdd FILL
XFILL_0__9236_ gnd vdd FILL
XFILL_4__14119_ gnd vdd FILL
X_9864_ _9864_/A gnd _9864_/Y vdd INVX1
XFILL_4__15099_ gnd vdd FILL
XFILL_3__14849_ gnd vdd FILL
XFILL_2__16278_ gnd vdd FILL
XSFILL89400x56050 gnd vdd FILL
XFILL_5__15409_ gnd vdd FILL
XFILL_0__14669_ gnd vdd FILL
XFILL_0__9167_ gnd vdd FILL
X_8815_ _8815_/Q _8815_/CLK _8047_/R vdd _8815_/D gnd vdd DFFSR
XFILL_5__16389_ gnd vdd FILL
XFILL_2__15229_ gnd vdd FILL
XFILL_0__16408_ gnd vdd FILL
X_9795_ _9793_/Y _9798_/B _9795_/C gnd _9839_/D vdd OAI21X1
XFILL_1__15959_ gnd vdd FILL
XFILL_4__6970_ gnd vdd FILL
XFILL_0__8118_ gnd vdd FILL
XFILL_6_BUFX2_insert633 gnd vdd FILL
XFILL_0__9098_ gnd vdd FILL
X_8746_ _8695_/B _7594_/B gnd _8747_/C vdd NAND2X1
XFILL_1__9980_ gnd vdd FILL
XFILL_3__9916_ gnd vdd FILL
XFILL_0__16339_ gnd vdd FILL
XFILL_6__6837_ gnd vdd FILL
XSFILL13640x51050 gnd vdd FILL
XSFILL94520x47050 gnd vdd FILL
XFILL_4__8640_ gnd vdd FILL
X_8677_ _8611_/A _8165_/CLK _9046_/R vdd _8677_/D gnd vdd DFFSR
XFILL_3__9847_ gnd vdd FILL
X_7628_ _7626_/Y _7562_/B _7627_/Y gnd _7666_/D vdd OAI21X1
XFILL_1__8862_ gnd vdd FILL
XSFILL114280x55050 gnd vdd FILL
XFILL_4__8571_ gnd vdd FILL
XFILL_3__9778_ gnd vdd FILL
XFILL_1__7813_ gnd vdd FILL
XFILL_1_CLKBUF1_insert115 gnd vdd FILL
XFILL_1_CLKBUF1_insert126 gnd vdd FILL
XFILL_3__8729_ gnd vdd FILL
XSFILL104520x32050 gnd vdd FILL
X_7559_ _7557_/Y _7598_/B _7558_/Y gnd _7643_/D vdd OAI21X1
XFILL_1_CLKBUF1_insert137 gnd vdd FILL
XFILL_1_CLKBUF1_insert148 gnd vdd FILL
XSFILL8760x30050 gnd vdd FILL
XFILL_1_CLKBUF1_insert159 gnd vdd FILL
XFILL_1__7744_ gnd vdd FILL
XSFILL33800x64050 gnd vdd FILL
XSFILL98760x52050 gnd vdd FILL
XFILL_4__7453_ gnd vdd FILL
X_11160_ _12183_/Y gnd _11160_/Y vdd INVX1
X_9229_ _9227_/Y _9228_/A _9229_/C gnd _9309_/D vdd OAI21X1
XFILL_1__7675_ gnd vdd FILL
XFILL_3_BUFX2_insert501 gnd vdd FILL
X_10111_ _10201_/Q gnd _10111_/Y vdd INVX1
XFILL_1__9414_ gnd vdd FILL
X_11091_ _12159_/Y gnd _11092_/B vdd INVX1
XFILL_3_BUFX2_insert512 gnd vdd FILL
XFILL_3_BUFX2_insert523 gnd vdd FILL
XFILL_4__9123_ gnd vdd FILL
XFILL_3_BUFX2_insert534 gnd vdd FILL
XFILL_3_BUFX2_insert545 gnd vdd FILL
X_10042_ _10042_/A _10024_/B _10041_/Y gnd _10042_/Y vdd OAI21X1
XFILL_3_BUFX2_insert556 gnd vdd FILL
XFILL_1__9345_ gnd vdd FILL
XFILL_3_BUFX2_insert567 gnd vdd FILL
XSFILL13720x31050 gnd vdd FILL
XFILL_3_BUFX2_insert578 gnd vdd FILL
XFILL_3_BUFX2_insert589 gnd vdd FILL
X_14850_ _9459_/Q _13883_/B _14850_/C gnd _14850_/Y vdd AOI21X1
XSFILL79160x26050 gnd vdd FILL
XFILL_1__9276_ gnd vdd FILL
XFILL_4__8005_ gnd vdd FILL
X_13801_ _9309_/Q gnd _13801_/Y vdd INVX1
XFILL_1__8227_ gnd vdd FILL
X_14781_ _13587_/C _16127_/D _14779_/Y _13574_/C gnd _14781_/Y vdd OAI22X1
X_11993_ _11993_/A _12113_/B _12113_/C gnd gnd _11994_/C vdd AOI22X1
X_13732_ _8837_/A gnd _13733_/A vdd INVX1
X_10944_ _10944_/A _10944_/B _10944_/C gnd _10944_/Y vdd AOI21X1
X_16451_ _16451_/A _16450_/B _16451_/C gnd _16451_/Y vdd OAI21X1
XSFILL44280x33050 gnd vdd FILL
X_13663_ _13663_/A _13663_/B gnd _13664_/A vdd NAND2X1
XFILL_1__7109_ gnd vdd FILL
XSFILL53800x2050 gnd vdd FILL
XSFILL99320x39050 gnd vdd FILL
X_10875_ _10887_/A gnd _10882_/A vdd INVX1
XFILL_2__8971_ gnd vdd FILL
XFILL_1__8089_ gnd vdd FILL
XFILL_5__7700_ gnd vdd FILL
X_15402_ _7902_/Q gnd _15404_/A vdd INVX1
XFILL_4__8907_ gnd vdd FILL
X_12614_ _12614_/A vdd _12613_/Y gnd _12678_/D vdd OAI21X1
X_16382_ gnd gnd gnd _16382_/Y vdd NAND2X1
XFILL_0_BUFX2_insert402 gnd vdd FILL
XFILL_4__9887_ gnd vdd FILL
X_13594_ _13594_/A _14344_/B _13853_/C _6911_/A gnd _13595_/B vdd AOI22X1
XFILL_3__10530_ gnd vdd FILL
XFILL_0_BUFX2_insert413 gnd vdd FILL
XFILL_5__7631_ gnd vdd FILL
XFILL_0_BUFX2_insert424 gnd vdd FILL
X_15333_ _8540_/Q gnd _15334_/B vdd INVX1
XFILL_4__8838_ gnd vdd FILL
XFILL_0_BUFX2_insert435 gnd vdd FILL
XFILL_0_BUFX2_insert446 gnd vdd FILL
XFILL_5__12070_ gnd vdd FILL
X_12545_ _12027_/B _13184_/CLK _8176_/R vdd _12471_/Y gnd vdd DFFSR
XFILL_6__10641_ gnd vdd FILL
XFILL_4__11820_ gnd vdd FILL
XFILL_0_BUFX2_insert457 gnd vdd FILL
XFILL_2__7853_ gnd vdd FILL
XFILL_0_BUFX2_insert468 gnd vdd FILL
XFILL_1__11640_ gnd vdd FILL
XFILL_5__7562_ gnd vdd FILL
XFILL_0_BUFX2_insert479 gnd vdd FILL
XFILL_0__10281_ gnd vdd FILL
XFILL_4__8769_ gnd vdd FILL
XFILL_5__11021_ gnd vdd FILL
XFILL_3__12200_ gnd vdd FILL
XSFILL13800x11050 gnd vdd FILL
X_15264_ _15264_/A _15264_/B gnd _15265_/C vdd NOR2X1
X_12476_ vdd _12476_/B gnd _12476_/Y vdd NAND2X1
XFILL_4__11751_ gnd vdd FILL
XFILL_0__12020_ gnd vdd FILL
XFILL_5__9301_ gnd vdd FILL
XFILL_3__10392_ gnd vdd FILL
XFILL_1__11571_ gnd vdd FILL
X_14215_ _14215_/A _14215_/B _14212_/Y gnd _14216_/B vdd NAND3X1
XFILL112120x63050 gnd vdd FILL
XFILL_4__10702_ gnd vdd FILL
XFILL_5__7493_ gnd vdd FILL
X_11427_ _11427_/A _11011_/Y _11374_/Y gnd _11428_/C vdd AOI21X1
XFILL_4__14470_ gnd vdd FILL
X_15195_ _15195_/A _15195_/B gnd _15196_/B vdd NOR2X1
XFILL_2__9523_ gnd vdd FILL
XFILL_3__12131_ gnd vdd FILL
XFILL_1__13310_ gnd vdd FILL
XFILL_1__10522_ gnd vdd FILL
XFILL_4__11682_ gnd vdd FILL
XFILL_5__9232_ gnd vdd FILL
XFILL_2__12861_ gnd vdd FILL
XFILL_6__15030_ gnd vdd FILL
XFILL_1__14290_ gnd vdd FILL
XFILL_4__13421_ gnd vdd FILL
X_14146_ _14389_/B _14146_/B _7268_/Q _14458_/C gnd _14146_/Y vdd AOI22X1
XFILL_2__14600_ gnd vdd FILL
XFILL_4__10633_ gnd vdd FILL
XFILL_5__15760_ gnd vdd FILL
X_11358_ _11358_/A _11358_/B _11202_/Y gnd _11359_/A vdd AOI21X1
XFILL_5__12972_ gnd vdd FILL
XFILL_3__12062_ gnd vdd FILL
XSFILL109640x1050 gnd vdd FILL
XFILL_2__11812_ gnd vdd FILL
XFILL_1__13241_ gnd vdd FILL
XFILL_1__10453_ gnd vdd FILL
XFILL_2__15580_ gnd vdd FILL
XCLKBUF1_insert114 CLKBUF1_insert216/A gnd _8046_/CLK vdd CLKBUF1
XFILL_5__9163_ gnd vdd FILL
XSFILL43720x47050 gnd vdd FILL
XFILL_4_BUFX2_insert390 gnd vdd FILL
X_10309_ _10264_/A _7877_/B gnd _10310_/C vdd NAND2X1
XFILL_5__14711_ gnd vdd FILL
XCLKBUF1_insert125 CLKBUF1_insert182/A gnd _7274_/CLK vdd CLKBUF1
XFILL_0__13971_ gnd vdd FILL
XFILL_4__13352_ gnd vdd FILL
XCLKBUF1_insert136 CLKBUF1_insert206/A gnd _8560_/CLK vdd CLKBUF1
XFILL_5__11923_ gnd vdd FILL
XFILL_2__8405_ gnd vdd FILL
X_14077_ _14909_/C _7139_/Q _14077_/C _13621_/B gnd _14085_/B vdd AOI22X1
XFILL_3__11013_ gnd vdd FILL
XFILL_4__16140_ gnd vdd FILL
XFILL_5__15691_ gnd vdd FILL
XFILL_2__14531_ gnd vdd FILL
XFILL_4__10564_ gnd vdd FILL
X_11289_ _11257_/Y _11431_/C _11289_/C gnd _11637_/B vdd OAI21X1
XFILL_0__15710_ gnd vdd FILL
XFILL_1__13172_ gnd vdd FILL
XFILL_5__8114_ gnd vdd FILL
XFILL_2__9385_ gnd vdd FILL
XCLKBUF1_insert147 CLKBUF1_insert193/A gnd _8151_/CLK vdd CLKBUF1
XFILL_2__11743_ gnd vdd FILL
XFILL_1__10384_ gnd vdd FILL
XCLKBUF1_insert158 CLKBUF1_insert206/A gnd _9306_/CLK vdd CLKBUF1
XSFILL69160x58050 gnd vdd FILL
XCLKBUF1_insert169 CLKBUF1_insert169/A gnd _8289_/CLK vdd CLKBUF1
XFILL_4__12303_ gnd vdd FILL
X_13028_ _13026_/Y vdd _13028_/C gnd _13072_/D vdd OAI21X1
XFILL_6__11124_ gnd vdd FILL
XFILL_5__9094_ gnd vdd FILL
XFILL_0__7420_ gnd vdd FILL
XSFILL99400x19050 gnd vdd FILL
XFILL_5__14642_ gnd vdd FILL
XFILL_4__16071_ gnd vdd FILL
XFILL_4__13283_ gnd vdd FILL
XFILL_2__8336_ gnd vdd FILL
XFILL_3__15821_ gnd vdd FILL
XFILL_1__12123_ gnd vdd FILL
XFILL_5__11854_ gnd vdd FILL
XFILL_4__10495_ gnd vdd FILL
XFILL_2__14462_ gnd vdd FILL
XFILL_0__15641_ gnd vdd FILL
XFILL_2__11674_ gnd vdd FILL
XFILL_0__12853_ gnd vdd FILL
XFILL_5__10805_ gnd vdd FILL
XFILL_0__7351_ gnd vdd FILL
XSFILL103880x60050 gnd vdd FILL
XFILL_2__16201_ gnd vdd FILL
XFILL_4__15022_ gnd vdd FILL
XFILL_4__12234_ gnd vdd FILL
XFILL_5__14573_ gnd vdd FILL
XSFILL104360x67050 gnd vdd FILL
XFILL_2__13413_ gnd vdd FILL
XFILL_2__10625_ gnd vdd FILL
XFILL_2__8267_ gnd vdd FILL
XFILL_3__12964_ gnd vdd FILL
XFILL_1__12054_ gnd vdd FILL
XFILL_5__11785_ gnd vdd FILL
XFILL_3__7060_ gnd vdd FILL
XFILL_3__15752_ gnd vdd FILL
XFILL_2__14393_ gnd vdd FILL
XFILL_0__11804_ gnd vdd FILL
XFILL_0__12784_ gnd vdd FILL
XFILL_0__15572_ gnd vdd FILL
XFILL_5__16312_ gnd vdd FILL
XSFILL74280x49050 gnd vdd FILL
XSFILL23640x14050 gnd vdd FILL
XFILL_5__13524_ gnd vdd FILL
XFILL_3__11915_ gnd vdd FILL
XFILL_3__14703_ gnd vdd FILL
XFILL_4__12165_ gnd vdd FILL
X_6930_ _6982_/B _7186_/B gnd _6930_/Y vdd NAND2X1
XFILL_2__7218_ gnd vdd FILL
XFILL_1__11005_ gnd vdd FILL
XFILL_2__16132_ gnd vdd FILL
XFILL_2__13344_ gnd vdd FILL
XFILL_3__15683_ gnd vdd FILL
X_14979_ _12770_/A gnd _14979_/Y vdd INVX8
XFILL_3__12895_ gnd vdd FILL
XFILL_2__10556_ gnd vdd FILL
XFILL_0__14523_ gnd vdd FILL
XFILL_0__11735_ gnd vdd FILL
XFILL_2__8198_ gnd vdd FILL
XFILL_0__9021_ gnd vdd FILL
XFILL_5__16243_ gnd vdd FILL
XFILL_4__11116_ gnd vdd FILL
XFILL_5__9996_ gnd vdd FILL
XFILL_5__13455_ gnd vdd FILL
XSFILL49080x25050 gnd vdd FILL
XFILL_3__14634_ gnd vdd FILL
X_6861_ _6861_/A gnd memoryAddress[23] vdd BUFX2
XFILL112200x43050 gnd vdd FILL
XFILL_4__12096_ gnd vdd FILL
XFILL_5__10667_ gnd vdd FILL
XFILL_1__15813_ gnd vdd FILL
XFILL_2__16063_ gnd vdd FILL
XFILL_3__11846_ gnd vdd FILL
XFILL_2__13275_ gnd vdd FILL
XFILL_6__7740_ gnd vdd FILL
XFILL_0__14454_ gnd vdd FILL
XFILL_2__10487_ gnd vdd FILL
XFILL_0__11666_ gnd vdd FILL
XFILL_5__12406_ gnd vdd FILL
X_8600_ _8609_/A _8600_/B gnd _8600_/Y vdd NAND2X1
XFILL_4__15924_ gnd vdd FILL
XFILL_5__16174_ gnd vdd FILL
XFILL_6__11957_ gnd vdd FILL
XFILL_2__15014_ gnd vdd FILL
XFILL_4__11047_ gnd vdd FILL
XFILL_3__14565_ gnd vdd FILL
XFILL_5__13386_ gnd vdd FILL
X_9580_ _9580_/Q _7020_/CLK _9580_/R vdd _9530_/Y gnd vdd DFFSR
XFILL_2__12226_ gnd vdd FILL
XFILL_0__13405_ gnd vdd FILL
XFILL_3__7962_ gnd vdd FILL
XFILL_0__10617_ gnd vdd FILL
XFILL_3__11777_ gnd vdd FILL
XFILL_1__15744_ gnd vdd FILL
XFILL_0__14385_ gnd vdd FILL
XFILL_1__12956_ gnd vdd FILL
XFILL_1_BUFX2_insert280 gnd vdd FILL
XFILL_0__11597_ gnd vdd FILL
XFILL_5__15125_ gnd vdd FILL
X_8531_ _8531_/A gnd _8533_/A vdd INVX1
XFILL_3__16304_ gnd vdd FILL
XFILL_5__8878_ gnd vdd FILL
XFILL_3__13516_ gnd vdd FILL
XFILL_5__12337_ gnd vdd FILL
XFILL_3__6913_ gnd vdd FILL
XFILL_4__15855_ gnd vdd FILL
XSFILL43800x27050 gnd vdd FILL
XFILL_1_BUFX2_insert291 gnd vdd FILL
XFILL_3__14496_ gnd vdd FILL
XFILL_1__11907_ gnd vdd FILL
XFILL_2__12157_ gnd vdd FILL
XFILL_0__16124_ gnd vdd FILL
XFILL_0__13336_ gnd vdd FILL
XFILL_1__15675_ gnd vdd FILL
XFILL_5_BUFX2_insert607 gnd vdd FILL
XFILL_3__7893_ gnd vdd FILL
XFILL_6__9410_ gnd vdd FILL
XFILL_0__10548_ gnd vdd FILL
XSFILL53960x71050 gnd vdd FILL
XFILL_1__12887_ gnd vdd FILL
XFILL_5__7829_ gnd vdd FILL
XFILL_0__9923_ gnd vdd FILL
XFILL_5_BUFX2_insert618 gnd vdd FILL
XFILL_4__14806_ gnd vdd FILL
XFILL_5__15056_ gnd vdd FILL
XFILL_5_BUFX2_insert629 gnd vdd FILL
X_8462_ _8542_/Q gnd _8464_/A vdd INVX1
XFILL_3__16235_ gnd vdd FILL
XFILL_3__9632_ gnd vdd FILL
XFILL_3__13447_ gnd vdd FILL
XFILL_5__12268_ gnd vdd FILL
XFILL_2__11108_ gnd vdd FILL
XFILL_3__10659_ gnd vdd FILL
XFILL_1__14626_ gnd vdd FILL
XFILL_3__6844_ gnd vdd FILL
XFILL_4__15786_ gnd vdd FILL
XSFILL53960x8050 gnd vdd FILL
XFILL_0__13267_ gnd vdd FILL
XFILL_4__12998_ gnd vdd FILL
XFILL_2__12088_ gnd vdd FILL
XFILL_0__16055_ gnd vdd FILL
XFILL_1__11838_ gnd vdd FILL
XFILL_5__14007_ gnd vdd FILL
XFILL_0_BUFX2_insert980 gnd vdd FILL
X_7413_ _7413_/Q _9589_/CLK _7413_/R vdd _7381_/Y gnd vdd DFFSR
XFILL_0__9854_ gnd vdd FILL
XFILL_5__11219_ gnd vdd FILL
XFILL_0_BUFX2_insert991 gnd vdd FILL
XFILL_3__16166_ gnd vdd FILL
XFILL_4__14737_ gnd vdd FILL
XFILL_5__12199_ gnd vdd FILL
X_8393_ _8391_/Y _8365_/A _8393_/C gnd _8433_/D vdd OAI21X1
XSFILL54040x80050 gnd vdd FILL
XFILL_2__15916_ gnd vdd FILL
XFILL_3__13378_ gnd vdd FILL
XFILL_4__11949_ gnd vdd FILL
XFILL_0__15006_ gnd vdd FILL
XFILL_0__12218_ gnd vdd FILL
XFILL_2__11039_ gnd vdd FILL
XFILL_1__14557_ gnd vdd FILL
XSFILL104440x47050 gnd vdd FILL
XFILL_1__11769_ gnd vdd FILL
X_7344_ _7366_/B _9008_/B gnd _7344_/Y vdd NAND2X1
XFILL_3__15117_ gnd vdd FILL
XFILL_0__9785_ gnd vdd FILL
XFILL_3__12329_ gnd vdd FILL
XFILL_3__8514_ gnd vdd FILL
XFILL_0__6997_ gnd vdd FILL
XFILL_3__16097_ gnd vdd FILL
XFILL_4__14668_ gnd vdd FILL
XFILL_1__13508_ gnd vdd FILL
XFILL_0__12149_ gnd vdd FILL
XFILL_2__15847_ gnd vdd FILL
XSFILL74360x29050 gnd vdd FILL
XFILL_3__9494_ gnd vdd FILL
XFILL_1__14488_ gnd vdd FILL
XFILL_0__8736_ gnd vdd FILL
XFILL_4__16407_ gnd vdd FILL
X_7275_ _7275_/Q _7261_/CLK _8669_/R vdd _7223_/Y gnd vdd DFFSR
XFILL_4__13619_ gnd vdd FILL
XFILL_3__15048_ gnd vdd FILL
XFILL_5__15958_ gnd vdd FILL
XFILL_1__16227_ gnd vdd FILL
XFILL_3__8445_ gnd vdd FILL
XFILL_4__14599_ gnd vdd FILL
XFILL_1__13439_ gnd vdd FILL
XFILL_2__15778_ gnd vdd FILL
XSFILL59160x2050 gnd vdd FILL
X_9014_ _9014_/A _7094_/B gnd _9014_/Y vdd NAND2X1
XFILL_5__14909_ gnd vdd FILL
XFILL_1__7460_ gnd vdd FILL
XFILL_4__16338_ gnd vdd FILL
XSFILL48920x60050 gnd vdd FILL
XFILL_2__14729_ gnd vdd FILL
XFILL_5__15889_ gnd vdd FILL
XFILL_3__8376_ gnd vdd FILL
XFILL_0__15908_ gnd vdd FILL
XFILL_6__7105_ gnd vdd FILL
XFILL_1__16158_ gnd vdd FILL
XFILL_0__7618_ gnd vdd FILL
XFILL_0__8598_ gnd vdd FILL
XFILL_3__7327_ gnd vdd FILL
XFILL_1__15109_ gnd vdd FILL
XFILL_4__16269_ gnd vdd FILL
XFILL_1__16089_ gnd vdd FILL
XFILL_0__15839_ gnd vdd FILL
XFILL_2_BUFX2_insert508 gnd vdd FILL
XSFILL13640x46050 gnd vdd FILL
XFILL_1__9130_ gnd vdd FILL
XFILL_2_BUFX2_insert519 gnd vdd FILL
XFILL_0__7549_ gnd vdd FILL
XSFILL109560x80050 gnd vdd FILL
X_9916_ _9917_/B _9532_/B gnd _9917_/C vdd NAND2X1
XSFILL39080x57050 gnd vdd FILL
XFILL_3__7189_ gnd vdd FILL
XFILL_0__9219_ gnd vdd FILL
XFILL_1__8012_ gnd vdd FILL
XSFILL54120x60050 gnd vdd FILL
X_9847_ _6903_/A _9865_/A gnd _9847_/Y vdd NAND2X1
XFILL_6_BUFX2_insert1027 gnd vdd FILL
XFILL_4__9810_ gnd vdd FILL
XSFILL8760x25050 gnd vdd FILL
XSFILL33800x59050 gnd vdd FILL
X_9778_ _9778_/A gnd _9780_/A vdd INVX1
XFILL_4__9741_ gnd vdd FILL
XSFILL94440x50 gnd vdd FILL
XFILL_4__6953_ gnd vdd FILL
XBUFX2_insert507 BUFX2_insert570/A gnd _12689_/R vdd BUFX2
X_10660_ _10661_/B _8228_/B gnd _10660_/Y vdd NAND2X1
XBUFX2_insert518 BUFX2_insert518/A gnd _8038_/R vdd BUFX2
X_8729_ _8727_/Y _8765_/B _8729_/C gnd _8801_/D vdd OAI21X1
XBUFX2_insert529 BUFX2_insert518/A gnd _7789_/R vdd BUFX2
XFILL_6_BUFX2_insert474 gnd vdd FILL
XFILL_4__9672_ gnd vdd FILL
XFILL_6_BUFX2_insert485 gnd vdd FILL
XFILL_4__6884_ gnd vdd FILL
XFILL_1__8914_ gnd vdd FILL
X_10591_ _13919_/A _7156_/CLK _7775_/R vdd _10515_/Y gnd vdd DFFSR
XFILL_1__9894_ gnd vdd FILL
XFILL_4__8623_ gnd vdd FILL
XFILL111960x69050 gnd vdd FILL
XFILL_4_BUFX2_insert1020 gnd vdd FILL
X_12330_ _12330_/A _12328_/Y _12330_/C gnd _12330_/Y vdd NAND3X1
XFILL_6__9539_ gnd vdd FILL
XFILL_1__8845_ gnd vdd FILL
XFILL_4_BUFX2_insert1031 gnd vdd FILL
XFILL_4_BUFX2_insert1042 gnd vdd FILL
XFILL_4_BUFX2_insert1053 gnd vdd FILL
XSFILL13720x26050 gnd vdd FILL
XFILL_4_BUFX2_insert1064 gnd vdd FILL
X_12261_ _6881_/A _12249_/B _12249_/C _12800_/Q gnd _12262_/C vdd AOI22X1
XFILL112040x78050 gnd vdd FILL
XSFILL23880x70050 gnd vdd FILL
XFILL_4_BUFX2_insert1086 gnd vdd FILL
XFILL_4__7505_ gnd vdd FILL
XFILL_1__8776_ gnd vdd FILL
X_14000_ _13999_/Y _14545_/B gnd _14000_/Y vdd NOR2X1
XFILL_4__8485_ gnd vdd FILL
X_11212_ _11212_/A _11211_/Y _11348_/A gnd _11212_/Y vdd OAI21X1
XFILL_1__7727_ gnd vdd FILL
X_12192_ _12192_/A _12123_/B _12192_/C gnd _12192_/Y vdd OAI21X1
XFILL_4__7436_ gnd vdd FILL
X_11143_ _11143_/A _11118_/Y gnd _11404_/A vdd NAND2X1
XFILL_3_BUFX2_insert320 gnd vdd FILL
XFILL_4__7367_ gnd vdd FILL
XFILL_3_BUFX2_insert331 gnd vdd FILL
XFILL_3_BUFX2_insert342 gnd vdd FILL
X_15951_ _14518_/A _15342_/B _15950_/Y gnd _15954_/A vdd OAI21X1
X_11074_ _11713_/C _11073_/Y _11074_/C gnd _11388_/B vdd OAI21X1
XFILL_3_BUFX2_insert353 gnd vdd FILL
XFILL_4__9106_ gnd vdd FILL
XFILL_2__9170_ gnd vdd FILL
XFILL_1__7589_ gnd vdd FILL
XFILL_3_BUFX2_insert364 gnd vdd FILL
XFILL_3_BUFX2_insert375 gnd vdd FILL
XFILL_4__7298_ gnd vdd FILL
XFILL_3_BUFX2_insert386 gnd vdd FILL
XSFILL58840x43050 gnd vdd FILL
XFILL_2_BUFX2_insert1090 gnd vdd FILL
X_14902_ _8912_/A gnd _14904_/A vdd INVX1
X_10025_ _10087_/Q gnd _10025_/Y vdd INVX1
XFILL_2__8121_ gnd vdd FILL
X_15882_ _15881_/Y _15879_/Y gnd _15882_/Y vdd NOR2X1
XFILL_3_BUFX2_insert397 gnd vdd FILL
XFILL_4__10280_ gnd vdd FILL
XFILL_4__9037_ gnd vdd FILL
XSFILL19320x66050 gnd vdd FILL
X_14833_ _14833_/A _14833_/B gnd _14833_/Y vdd NOR2X1
XFILL_5__11570_ gnd vdd FILL
XFILL_2__10410_ gnd vdd FILL
XFILL_1__9259_ gnd vdd FILL
XSFILL23560x29050 gnd vdd FILL
XFILL_2__11390_ gnd vdd FILL
XFILL_5__9850_ gnd vdd FILL
XFILL_5__10521_ gnd vdd FILL
XFILL_3__11700_ gnd vdd FILL
X_14764_ _14764_/A _14764_/B _14764_/C gnd _14764_/Y vdd NAND3X1
X_11976_ _11976_/A _11975_/A _11976_/C gnd _6867_/A vdd OAI21X1
XFILL_0__11520_ gnd vdd FILL
XFILL112120x58050 gnd vdd FILL
X_13715_ _7941_/A gnd _15286_/C vdd INVX1
XFILL_5__9781_ gnd vdd FILL
XFILL_5__13240_ gnd vdd FILL
X_10927_ _10911_/A _10938_/B gnd _10927_/Y vdd NOR2X1
XFILL_5__10452_ gnd vdd FILL
XFILL_5__6993_ gnd vdd FILL
X_14695_ _9284_/A gnd _16090_/A vdd INVX1
XFILL_3__11631_ gnd vdd FILL
XFILL_2__10272_ gnd vdd FILL
XFILL_4__13970_ gnd vdd FILL
XSFILL64840x62050 gnd vdd FILL
XSFILL64040x43050 gnd vdd FILL
XFILL_4_CLKBUF1_insert121 gnd vdd FILL
XFILL_0__11451_ gnd vdd FILL
XFILL_1__13790_ gnd vdd FILL
XFILL_4_CLKBUF1_insert132 gnd vdd FILL
XFILL_5__8732_ gnd vdd FILL
XFILL_4__9939_ gnd vdd FILL
X_13646_ _14643_/B gnd _13864_/B vdd INVX8
XFILL_4_CLKBUF1_insert143 gnd vdd FILL
X_16434_ _15747_/A _8792_/CLK _9048_/R vdd _16434_/D gnd vdd DFFSR
XFILL_5__10383_ gnd vdd FILL
XFILL_2__12011_ gnd vdd FILL
XFILL_5__13171_ gnd vdd FILL
XFILL_3__14350_ gnd vdd FILL
XFILL_4_CLKBUF1_insert154 gnd vdd FILL
X_10858_ _10802_/A _8297_/CLK _7796_/R vdd _10858_/D gnd vdd DFFSR
XFILL_0__10402_ gnd vdd FILL
XFILL_2__8954_ gnd vdd FILL
XFILL_3__11562_ gnd vdd FILL
XFILL_1__12741_ gnd vdd FILL
XFILL_0__14170_ gnd vdd FILL
XFILL_4_CLKBUF1_insert165 gnd vdd FILL
XFILL_4_CLKBUF1_insert176 gnd vdd FILL
XFILL_0__11382_ gnd vdd FILL
XFILL_3__13301_ gnd vdd FILL
XFILL_4_CLKBUF1_insert187 gnd vdd FILL
X_16365_ _16363_/Y gnd _16365_/C gnd _16431_/D vdd OAI21X1
XFILL_0_BUFX2_insert232 gnd vdd FILL
XFILL_5__12122_ gnd vdd FILL
XFILL_4__15640_ gnd vdd FILL
XFILL_4_CLKBUF1_insert198 gnd vdd FILL
X_13577_ _13479_/C _13577_/B _14744_/B _13576_/Y gnd _13578_/B vdd OAI22X1
XFILL_3__10513_ gnd vdd FILL
X_10789_ _10787_/Y _10789_/B _10788_/Y gnd _10789_/Y vdd OAI21X1
XFILL_0__13121_ gnd vdd FILL
XFILL_0_BUFX2_insert243 gnd vdd FILL
XFILL_4__12852_ gnd vdd FILL
XFILL_3__14281_ gnd vdd FILL
XFILL_0_BUFX2_insert254 gnd vdd FILL
XFILL_2__8885_ gnd vdd FILL
XFILL_3__11493_ gnd vdd FILL
XFILL_1__15460_ gnd vdd FILL
XFILL_5__7614_ gnd vdd FILL
X_15316_ _9224_/A gnd _15317_/A vdd INVX1
XFILL_0_BUFX2_insert265 gnd vdd FILL
XFILL_3__16020_ gnd vdd FILL
XFILL_0__6920_ gnd vdd FILL
X_12528_ _12526_/Y vdd _12527_/Y gnd _12564_/D vdd OAI21X1
XFILL_5__12053_ gnd vdd FILL
XFILL_0_BUFX2_insert276 gnd vdd FILL
XFILL_5__8594_ gnd vdd FILL
XFILL_3__13232_ gnd vdd FILL
XFILL_0_BUFX2_insert287 gnd vdd FILL
X_16296_ _16296_/A _16296_/B _16295_/Y gnd _16320_/A vdd NOR3X1
XFILL_4__11803_ gnd vdd FILL
XFILL_3__10444_ gnd vdd FILL
XFILL_2__7836_ gnd vdd FILL
XFILL_4__15571_ gnd vdd FILL
XFILL_1__14411_ gnd vdd FILL
XFILL_4__12783_ gnd vdd FILL
XFILL_1__11623_ gnd vdd FILL
XFILL_2__13962_ gnd vdd FILL
XFILL_0_BUFX2_insert298 gnd vdd FILL
XSFILL58920x23050 gnd vdd FILL
XFILL_1__15391_ gnd vdd FILL
XFILL_0__10264_ gnd vdd FILL
XFILL_5__7545_ gnd vdd FILL
XFILL_5__11004_ gnd vdd FILL
X_15247_ _13668_/Y _15920_/B _15920_/C _13669_/D gnd _15247_/Y vdd OAI22X1
X_12459_ _12457_/Y vdd _12458_/Y gnd _12459_/Y vdd OAI21X1
XFILL_4__14522_ gnd vdd FILL
XFILL_0__6851_ gnd vdd FILL
XFILL_2__15701_ gnd vdd FILL
XFILL_3__13163_ gnd vdd FILL
XFILL_0__12003_ gnd vdd FILL
XFILL_2__12913_ gnd vdd FILL
XFILL_4__11734_ gnd vdd FILL
XFILL_1__14342_ gnd vdd FILL
XFILL_3__10375_ gnd vdd FILL
XFILL_2__13893_ gnd vdd FILL
XFILL_1__11554_ gnd vdd FILL
XFILL_5__15812_ gnd vdd FILL
XFILL_0__10195_ gnd vdd FILL
XFILL_5__7476_ gnd vdd FILL
X_15178_ _8793_/Q _15821_/B _15178_/C _10239_/A gnd _15178_/Y vdd AOI22X1
XFILL_3__12114_ gnd vdd FILL
XSFILL59000x32050 gnd vdd FILL
XFILL_4__14453_ gnd vdd FILL
XFILL_2__9506_ gnd vdd FILL
XFILL_2__15632_ gnd vdd FILL
XFILL_6__10486_ gnd vdd FILL
XFILL_2_BUFX2_insert14 gnd vdd FILL
XFILL_4__11665_ gnd vdd FILL
XFILL_2__12844_ gnd vdd FILL
XFILL_1__10505_ gnd vdd FILL
XFILL_3__13094_ gnd vdd FILL
XFILL_2_BUFX2_insert25 gnd vdd FILL
XSFILL104760x83050 gnd vdd FILL
XFILL_5__9215_ gnd vdd FILL
XFILL_2_BUFX2_insert36 gnd vdd FILL
XFILL_1__14273_ gnd vdd FILL
XFILL_2__7698_ gnd vdd FILL
X_14129_ _14129_/A _14128_/Y gnd _14133_/C vdd NOR2X1
XFILL_0__8521_ gnd vdd FILL
XFILL_2_BUFX2_insert47 gnd vdd FILL
XFILL_1__11485_ gnd vdd FILL
XFILL_4__13404_ gnd vdd FILL
XFILL_4__10616_ gnd vdd FILL
X_7060_ _7060_/A gnd _7060_/Y vdd INVX1
XFILL_5__15743_ gnd vdd FILL
XFILL_1__16012_ gnd vdd FILL
XFILL_3__8230_ gnd vdd FILL
XFILL_3__12045_ gnd vdd FILL
XFILL_2_BUFX2_insert58 gnd vdd FILL
XFILL_5__12955_ gnd vdd FILL
XFILL_1__13224_ gnd vdd FILL
XFILL_2_BUFX2_insert69 gnd vdd FILL
XFILL112200x38050 gnd vdd FILL
XFILL_2__15563_ gnd vdd FILL
XFILL_4__14384_ gnd vdd FILL
XFILL_4__11596_ gnd vdd FILL
XFILL_2__12775_ gnd vdd FILL
XFILL_5__9146_ gnd vdd FILL
XFILL_1__10436_ gnd vdd FILL
XSFILL23720x6050 gnd vdd FILL
XFILL_0__13954_ gnd vdd FILL
XFILL_0__8452_ gnd vdd FILL
XFILL_5__11906_ gnd vdd FILL
XFILL_4__16123_ gnd vdd FILL
XFILL_4__13335_ gnd vdd FILL
XFILL_5__15674_ gnd vdd FILL
XFILL_2__14514_ gnd vdd FILL
XFILL_4__10547_ gnd vdd FILL
XSFILL64120x23050 gnd vdd FILL
XFILL_5__12886_ gnd vdd FILL
XFILL_2__9368_ gnd vdd FILL
XFILL_2__11726_ gnd vdd FILL
XFILL_1__10367_ gnd vdd FILL
XFILL_1__13155_ gnd vdd FILL
XFILL_2__15494_ gnd vdd FILL
XFILL_0__12905_ gnd vdd FILL
XFILL_0__13885_ gnd vdd FILL
XFILL_5__14625_ gnd vdd FILL
XFILL_4__13266_ gnd vdd FILL
XFILL_2__8319_ gnd vdd FILL
XFILL_0__8383_ gnd vdd FILL
XFILL_3__15804_ gnd vdd FILL
XFILL_3__7112_ gnd vdd FILL
XFILL_4__16054_ gnd vdd FILL
XFILL_5__11837_ gnd vdd FILL
XFILL_1__12106_ gnd vdd FILL
XFILL_2__14445_ gnd vdd FILL
XFILL_3__8092_ gnd vdd FILL
XFILL_0__15624_ gnd vdd FILL
XFILL_2__9299_ gnd vdd FILL
XFILL_2__11657_ gnd vdd FILL
XFILL_0__12836_ gnd vdd FILL
XFILL_1__13086_ gnd vdd FILL
XFILL_3__13996_ gnd vdd FILL
XFILL_1__10298_ gnd vdd FILL
XFILL_6__15915_ gnd vdd FILL
XSFILL53960x66050 gnd vdd FILL
XFILL_0__7334_ gnd vdd FILL
XFILL_4__15005_ gnd vdd FILL
XFILL_4__12217_ gnd vdd FILL
XFILL_5__14556_ gnd vdd FILL
XSFILL3560x30050 gnd vdd FILL
XFILL_3__7043_ gnd vdd FILL
X_7962_ _8034_/Q gnd _7964_/A vdd INVX1
XFILL_5__11768_ gnd vdd FILL
XFILL_3__15735_ gnd vdd FILL
XFILL_1__12037_ gnd vdd FILL
XFILL_2__14376_ gnd vdd FILL
XFILL_0__15555_ gnd vdd FILL
XFILL_2__11588_ gnd vdd FILL
X_9701_ _9701_/Q _8926_/CLK _8670_/R vdd _9637_/Y gnd vdd DFFSR
XFILL_0__12767_ gnd vdd FILL
XFILL_5__13507_ gnd vdd FILL
X_6913_ _6913_/A _6951_/A _6912_/Y gnd _6913_/Y vdd OAI21X1
XFILL_4__12148_ gnd vdd FILL
XFILL_2__16115_ gnd vdd FILL
XFILL_2__13327_ gnd vdd FILL
XFILL_5__14487_ gnd vdd FILL
XSFILL54040x75050 gnd vdd FILL
XFILL_3__15666_ gnd vdd FILL
XFILL_2__10539_ gnd vdd FILL
XFILL_0__14506_ gnd vdd FILL
XFILL_3__12878_ gnd vdd FILL
X_7893_ _7893_/A _7800_/B _7892_/Y gnd _7925_/D vdd OAI21X1
XFILL_5__11699_ gnd vdd FILL
XFILL_0__11718_ gnd vdd FILL
XFILL_0__9004_ gnd vdd FILL
XFILL_5__16226_ gnd vdd FILL
XFILL_0__15486_ gnd vdd FILL
XFILL_0__12698_ gnd vdd FILL
X_9632_ _9700_/Q gnd _9632_/Y vdd INVX1
XFILL_6__15777_ gnd vdd FILL
XFILL_5__9979_ gnd vdd FILL
XFILL_5__13438_ gnd vdd FILL
XFILL_3__14617_ gnd vdd FILL
XFILL_2__16046_ gnd vdd FILL
XFILL_4__12079_ gnd vdd FILL
X_6844_ _6844_/A gnd memoryAddress[6] vdd BUFX2
XFILL_0__7196_ gnd vdd FILL
XFILL_3__11829_ gnd vdd FILL
XFILL_2__13258_ gnd vdd FILL
XFILL_3__8994_ gnd vdd FILL
XFILL_3__15597_ gnd vdd FILL
XFILL_0__14437_ gnd vdd FILL
XFILL_1__13988_ gnd vdd FILL
XFILL_6__14728_ gnd vdd FILL
XFILL_0__11649_ gnd vdd FILL
XFILL_4__15907_ gnd vdd FILL
XFILL_5__16157_ gnd vdd FILL
XFILL_5__13369_ gnd vdd FILL
XSFILL33880x33050 gnd vdd FILL
XFILL_2__12209_ gnd vdd FILL
X_9563_ _9477_/A _8151_/CLK _9944_/R vdd _9479_/Y gnd vdd DFFSR
XSFILL33080x14050 gnd vdd FILL
XFILL_1__15727_ gnd vdd FILL
XFILL_3__14548_ gnd vdd FILL
XFILL_3__7945_ gnd vdd FILL
XFILL_0__14368_ gnd vdd FILL
XFILL111800x11050 gnd vdd FILL
XFILL_5__15108_ gnd vdd FILL
XFILL_5_BUFX2_insert404 gnd vdd FILL
X_8514_ _8469_/A _8642_/B gnd _8515_/C vdd NAND2X1
XFILL_5_BUFX2_insert415 gnd vdd FILL
XFILL_1__6960_ gnd vdd FILL
XFILL_5__16088_ gnd vdd FILL
XFILL_4__15838_ gnd vdd FILL
XFILL_3__14479_ gnd vdd FILL
XSFILL48920x55050 gnd vdd FILL
XFILL_0__16107_ gnd vdd FILL
XFILL_5_BUFX2_insert426 gnd vdd FILL
X_9494_ _9494_/A _9554_/B _9493_/Y gnd _9494_/Y vdd OAI21X1
XFILL_0__13319_ gnd vdd FILL
XFILL_1__15658_ gnd vdd FILL
XFILL_5_BUFX2_insert437 gnd vdd FILL
XFILL_3__7876_ gnd vdd FILL
XSFILL88520x41050 gnd vdd FILL
XFILL_5_BUFX2_insert448 gnd vdd FILL
XFILL_5__15039_ gnd vdd FILL
XFILL_0__9906_ gnd vdd FILL
XFILL_0__14299_ gnd vdd FILL
XFILL_3__16218_ gnd vdd FILL
XFILL_5_BUFX2_insert459 gnd vdd FILL
X_8445_ _8494_/B _7293_/B gnd _8446_/C vdd NAND2X1
XFILL_3__9615_ gnd vdd FILL
XFILL_1__14609_ gnd vdd FILL
XFILL_1__6891_ gnd vdd FILL
XFILL_4__15769_ gnd vdd FILL
XFILL_0__16038_ gnd vdd FILL
XFILL_6__16329_ gnd vdd FILL
XFILL_1__15589_ gnd vdd FILL
XFILL_1__8630_ gnd vdd FILL
X_8376_ _8376_/A gnd _8378_/A vdd INVX1
XFILL_3__16149_ gnd vdd FILL
XFILL_3__9546_ gnd vdd FILL
XSFILL3640x10050 gnd vdd FILL
XSFILL109560x75050 gnd vdd FILL
XFILL_6__9255_ gnd vdd FILL
XFILL_0__9768_ gnd vdd FILL
XSFILL64120x50 gnd vdd FILL
X_7327_ _7327_/A _7369_/B _7326_/Y gnd _7395_/D vdd OAI21X1
XFILL_4__8270_ gnd vdd FILL
XFILL_3__9477_ gnd vdd FILL
XFILL_6__8206_ gnd vdd FILL
XSFILL28840x22050 gnd vdd FILL
XFILL_0__8719_ gnd vdd FILL
XSFILL54120x55050 gnd vdd FILL
XFILL_4__7221_ gnd vdd FILL
X_7258_ _7258_/Q _8541_/CLK _7258_/R vdd _7172_/Y gnd vdd DFFSR
XFILL_1__8492_ gnd vdd FILL
XFILL_1__7443_ gnd vdd FILL
X_7189_ _7250_/B _7317_/B gnd _7189_/Y vdd NAND2X1
XFILL_3__8359_ gnd vdd FILL
XFILL_1__7374_ gnd vdd FILL
XFILL_1_BUFX2_insert0 gnd vdd FILL
XFILL_2_BUFX2_insert305 gnd vdd FILL
XFILL_2_BUFX2_insert316 gnd vdd FILL
XFILL_4__7083_ gnd vdd FILL
XFILL_2_BUFX2_insert327 gnd vdd FILL
XFILL_2_BUFX2_insert338 gnd vdd FILL
XFILL_1__9113_ gnd vdd FILL
XSFILL18760x74050 gnd vdd FILL
XFILL_2_BUFX2_insert349 gnd vdd FILL
X_11830_ _11830_/A gnd _11997_/A vdd INVX1
XSFILL9240x50050 gnd vdd FILL
XFILL_1__9044_ gnd vdd FILL
X_11761_ _11761_/A _11760_/Y _11245_/Y gnd _11761_/Y vdd AOI21X1
X_13500_ _8791_/Q gnd _15095_/D vdd INVX1
X_10712_ _15130_/B _7640_/CLK _7515_/R vdd _10622_/Y gnd vdd DFFSR
X_14480_ _14480_/A _14480_/B gnd _14483_/C vdd NOR2X1
XFILL_4__7985_ gnd vdd FILL
XBUFX2_insert304 _11983_/Y gnd _12011_/C vdd BUFX2
X_11692_ _11046_/Y _11684_/B _11691_/Y gnd _11699_/A vdd AOI21X1
XSFILL113880x18050 gnd vdd FILL
XFILL_6_BUFX2_insert260 gnd vdd FILL
XBUFX2_insert315 _13454_/Y gnd _14894_/B vdd BUFX2
XBUFX2_insert326 _13345_/Y gnd _9868_/A vdd BUFX2
XFILL_4__9724_ gnd vdd FILL
X_13431_ _10198_/Q gnd _13433_/A vdd INVX1
XFILL_4__6936_ gnd vdd FILL
X_10643_ _10643_/A _10676_/B _10642_/Y gnd _10643_/Y vdd OAI21X1
XBUFX2_insert337 _13494_/Y gnd _14414_/B vdd BUFX2
XSFILL39560x53050 gnd vdd FILL
XBUFX2_insert348 _10927_/Y gnd _12327_/A vdd BUFX2
XBUFX2_insert359 _13306_/Y gnd _7931_/B vdd BUFX2
XFILL_4__6867_ gnd vdd FILL
XFILL_5_CLKBUF1_insert205 gnd vdd FILL
XFILL_4__9655_ gnd vdd FILL
X_16150_ _14774_/D gnd _16150_/Y vdd INVX1
XFILL_5_CLKBUF1_insert216 gnd vdd FILL
X_13362_ _13259_/C _13219_/B gnd _13362_/Y vdd NOR2X1
X_10574_ _10535_/A _8014_/B gnd _10575_/C vdd NAND2X1
XFILL_5_BUFX2_insert960 gnd vdd FILL
XFILL_1__9877_ gnd vdd FILL
XFILL_4__8606_ gnd vdd FILL
X_15101_ _7895_/Q _16204_/B _16014_/C _8185_/A gnd _15102_/B vdd AOI22X1
XFILL_5_BUFX2_insert971 gnd vdd FILL
X_12313_ _6894_/A _12301_/B _12301_/C _12313_/D gnd _12314_/C vdd AOI22X1
XFILL_5_BUFX2_insert982 gnd vdd FILL
X_16081_ _8385_/A gnd _16082_/A vdd INVX1
X_13293_ _13297_/C _13293_/B gnd _13293_/Y vdd NOR2X1
XFILL_5_BUFX2_insert993 gnd vdd FILL
XFILL_2__7621_ gnd vdd FILL
XSFILL84440x5050 gnd vdd FILL
XFILL_1__8828_ gnd vdd FILL
XFILL_5__7330_ gnd vdd FILL
XSFILL18840x54050 gnd vdd FILL
X_15032_ _15244_/C _15031_/Y gnd _15035_/C vdd NAND2X1
XSFILL84280x30050 gnd vdd FILL
X_12244_ _12248_/A _12716_/A _12248_/C gnd _12246_/B vdd NAND3X1
XFILL_2__7552_ gnd vdd FILL
XFILL_1__8759_ gnd vdd FILL
XFILL_3__10160_ gnd vdd FILL
XFILL_2__10890_ gnd vdd FILL
XFILL_4__8468_ gnd vdd FILL
X_12175_ _11947_/A gnd _12177_/A vdd INVX1
XSFILL63960x29050 gnd vdd FILL
XFILL_4__11450_ gnd vdd FILL
XFILL_5__9000_ gnd vdd FILL
XFILL_2__7483_ gnd vdd FILL
XFILL_1__11270_ gnd vdd FILL
XFILL_4__7419_ gnd vdd FILL
XFILL_4__8399_ gnd vdd FILL
XFILL_4__10401_ gnd vdd FILL
XFILL_5__7192_ gnd vdd FILL
X_11126_ _11126_/A gnd _11591_/C vdd INVX2
XFILL_5__12740_ gnd vdd FILL
XFILL_2__9222_ gnd vdd FILL
XFILL_4__11381_ gnd vdd FILL
XFILL112280x12050 gnd vdd FILL
XSFILL64040x38050 gnd vdd FILL
XFILL_0__10951_ gnd vdd FILL
XFILL_4__13120_ gnd vdd FILL
X_15934_ _7276_/Q _15177_/B _15969_/C _7736_/A gnd _15934_/Y vdd AOI22X1
X_11057_ _11028_/Y _11041_/Y _11056_/Y gnd _11057_/Y vdd OAI21X1
XFILL_2__9153_ gnd vdd FILL
XFILL_2__11511_ gnd vdd FILL
XFILL_1__10152_ gnd vdd FILL
XFILL_3__13850_ gnd vdd FILL
XFILL_2__12491_ gnd vdd FILL
XFILL_0__13670_ gnd vdd FILL
X_10008_ _10024_/B _6936_/B gnd _10008_/Y vdd NAND2X1
XFILL_0__10882_ gnd vdd FILL
XFILL_5__14410_ gnd vdd FILL
XFILL_2__8104_ gnd vdd FILL
XFILL_5__11622_ gnd vdd FILL
XFILL_6__13961_ gnd vdd FILL
XFILL_5__15390_ gnd vdd FILL
XFILL_2__14230_ gnd vdd FILL
XFILL_4__10263_ gnd vdd FILL
X_15865_ _15862_/Y _15865_/B _15865_/C gnd _15866_/C vdd NAND3X1
XFILL_3__13781_ gnd vdd FILL
XFILL_2__9084_ gnd vdd FILL
XFILL_2__11442_ gnd vdd FILL
XFILL_0__12621_ gnd vdd FILL
XSFILL3480x45050 gnd vdd FILL
XFILL_1__14960_ gnd vdd FILL
XFILL_2_BUFX2_insert850 gnd vdd FILL
XFILL_3__10993_ gnd vdd FILL
XFILL_5__9902_ gnd vdd FILL
XFILL_6__15700_ gnd vdd FILL
XFILL_4__12002_ gnd vdd FILL
XFILL_2_BUFX2_insert861 gnd vdd FILL
X_14816_ _14816_/A gnd _16180_/B vdd INVX1
XFILL_2_BUFX2_insert872 gnd vdd FILL
XFILL_5__14341_ gnd vdd FILL
XFILL_3__12732_ gnd vdd FILL
XFILL_3__15520_ gnd vdd FILL
XFILL_2_BUFX2_insert883 gnd vdd FILL
XFILL_5__11553_ gnd vdd FILL
XFILL_2__14161_ gnd vdd FILL
X_15796_ _10796_/A gnd _15796_/Y vdd INVX1
XFILL_4__10194_ gnd vdd FILL
XFILL_1__13911_ gnd vdd FILL
XFILL_2_BUFX2_insert894 gnd vdd FILL
XFILL_0__15340_ gnd vdd FILL
XFILL_2__11373_ gnd vdd FILL
XFILL_1__14891_ gnd vdd FILL
XFILL_0__7050_ gnd vdd FILL
XFILL_5__10504_ gnd vdd FILL
X_11959_ _11959_/A gnd _11961_/A vdd INVX1
XFILL_2__13112_ gnd vdd FILL
X_14747_ _9329_/Q gnd _14747_/Y vdd INVX1
XFILL_5__14272_ gnd vdd FILL
XFILL_3__15451_ gnd vdd FILL
XFILL_5__11484_ gnd vdd FILL
XFILL_2__10324_ gnd vdd FILL
XFILL_1__13842_ gnd vdd FILL
XFILL_2__14092_ gnd vdd FILL
XFILL_0__11503_ gnd vdd FILL
XFILL_5__16011_ gnd vdd FILL
XFILL_0__12483_ gnd vdd FILL
XFILL_0__15271_ gnd vdd FILL
XFILL_5__9764_ gnd vdd FILL
XFILL_5__13223_ gnd vdd FILL
XFILL_6__15562_ gnd vdd FILL
XFILL_6__12774_ gnd vdd FILL
XFILL_5__6976_ gnd vdd FILL
XFILL_3__14402_ gnd vdd FILL
XSFILL59000x27050 gnd vdd FILL
XFILL_5__10435_ gnd vdd FILL
X_14678_ _14410_/A _16079_/D _14711_/B _14678_/D gnd _14678_/Y vdd OAI22X1
XFILL_3__11614_ gnd vdd FILL
XFILL_3__15382_ gnd vdd FILL
XFILL_4_BUFX2_insert4 gnd vdd FILL
XFILL_4__13953_ gnd vdd FILL
XFILL_2__13043_ gnd vdd FILL
XFILL_0__14222_ gnd vdd FILL
XFILL_2__10255_ gnd vdd FILL
XFILL_3__12594_ gnd vdd FILL
XFILL_0__11434_ gnd vdd FILL
XFILL_1__13773_ gnd vdd FILL
XSFILL69160x71050 gnd vdd FILL
XFILL_5__8715_ gnd vdd FILL
XFILL_2__9986_ gnd vdd FILL
XFILL_6__14513_ gnd vdd FILL
XSFILL99400x32050 gnd vdd FILL
X_13629_ _10495_/A gnd _13629_/Y vdd INVX1
X_16417_ _16417_/Q _8022_/CLK _9046_/R vdd _16323_/Y gnd vdd DFFSR
XFILL_5__13154_ gnd vdd FILL
XFILL_3__14333_ gnd vdd FILL
XFILL_4__12904_ gnd vdd FILL
XFILL_5__10366_ gnd vdd FILL
XFILL_1__15512_ gnd vdd FILL
XFILL_3__7730_ gnd vdd FILL
XFILL_3__11545_ gnd vdd FILL
XFILL_4__13884_ gnd vdd FILL
XFILL_1__12724_ gnd vdd FILL
XBUFX2_insert860 _13314_/Y gnd _8249_/A vdd BUFX2
XFILL_2__10186_ gnd vdd FILL
XFILL_0__14153_ gnd vdd FILL
XFILL_0__11365_ gnd vdd FILL
XFILL_5__12105_ gnd vdd FILL
XBUFX2_insert871 _13379_/Y gnd _13818_/A vdd BUFX2
XFILL_5__8646_ gnd vdd FILL
XFILL_0__7952_ gnd vdd FILL
XFILL_4__15623_ gnd vdd FILL
XFILL_6__11656_ gnd vdd FILL
X_16348_ _13909_/A gnd _16350_/A vdd INVX1
XFILL_3__14264_ gnd vdd FILL
XFILL_4__12835_ gnd vdd FILL
XFILL_5__13085_ gnd vdd FILL
XFILL_5__10297_ gnd vdd FILL
XBUFX2_insert882 _12216_/Y gnd _12289_/C vdd BUFX2
XSFILL64120x18050 gnd vdd FILL
XBUFX2_insert893 _12369_/Y gnd _9615_/B vdd BUFX2
XFILL_0__10316_ gnd vdd FILL
XFILL_0__13104_ gnd vdd FILL
XFILL_3__11476_ gnd vdd FILL
XFILL_1__15443_ gnd vdd FILL
XFILL_1__12655_ gnd vdd FILL
XFILL_2__8868_ gnd vdd FILL
XFILL_2__14994_ gnd vdd FILL
XFILL_0__14084_ gnd vdd FILL
XSFILL74280x62050 gnd vdd FILL
XFILL_0__6903_ gnd vdd FILL
XFILL_0__11296_ gnd vdd FILL
XFILL_5__8577_ gnd vdd FILL
XFILL_3__13215_ gnd vdd FILL
XFILL_3__16003_ gnd vdd FILL
X_8230_ _8230_/A gnd _8232_/A vdd INVX1
XFILL_5__12036_ gnd vdd FILL
XFILL_6__14375_ gnd vdd FILL
X_16279_ _15842_/A _16279_/B _16277_/Y _16137_/C gnd _16280_/B vdd OAI22X1
XFILL_3__10427_ gnd vdd FILL
XFILL_0__7883_ gnd vdd FILL
XFILL_4__15554_ gnd vdd FILL
XFILL_3__9400_ gnd vdd FILL
XFILL_4__12766_ gnd vdd FILL
XFILL_2__7819_ gnd vdd FILL
XFILL_3__14195_ gnd vdd FILL
XFILL_0__13035_ gnd vdd FILL
XFILL_1__11606_ gnd vdd FILL
XFILL_2__13945_ gnd vdd FILL
XFILL_3__7592_ gnd vdd FILL
XFILL_1__15374_ gnd vdd FILL
XFILL_6__16114_ gnd vdd FILL
XFILL_0__10247_ gnd vdd FILL
XFILL_6__13326_ gnd vdd FILL
XFILL_1__12586_ gnd vdd FILL
XFILL_0__9622_ gnd vdd FILL
XFILL_4__14505_ gnd vdd FILL
XFILL_6__10538_ gnd vdd FILL
X_8161_ _8087_/A _8161_/CLK _7140_/R vdd _8161_/D gnd vdd DFFSR
XFILL_3__13146_ gnd vdd FILL
XFILL_4__11717_ gnd vdd FILL
XSFILL3560x25050 gnd vdd FILL
XFILL_3__10358_ gnd vdd FILL
XFILL_1__14325_ gnd vdd FILL
XFILL_4__15485_ gnd vdd FILL
XFILL_4__12697_ gnd vdd FILL
XFILL_2__13876_ gnd vdd FILL
XFILL_1__11537_ gnd vdd FILL
XFILL_5__7459_ gnd vdd FILL
XFILL_0__10178_ gnd vdd FILL
X_7112_ _7124_/A _8136_/B gnd _7113_/C vdd NAND2X1
XFILL_0__9553_ gnd vdd FILL
X_8092_ _8092_/A _8100_/A _8091_/Y gnd _8162_/D vdd OAI21X1
XSFILL28760x37050 gnd vdd FILL
XFILL_4__14436_ gnd vdd FILL
XFILL_2__15615_ gnd vdd FILL
XFILL_5__13987_ gnd vdd FILL
XFILL_3__9262_ gnd vdd FILL
XFILL_4__11648_ gnd vdd FILL
XFILL_2__12827_ gnd vdd FILL
XFILL_1__14256_ gnd vdd FILL
XFILL_3__10289_ gnd vdd FILL
XFILL_0__8504_ gnd vdd FILL
XFILL_6__12208_ gnd vdd FILL
XSFILL33880x7050 gnd vdd FILL
XFILL_1__11468_ gnd vdd FILL
XFILL_5__15726_ gnd vdd FILL
X_7043_ _7095_/B _8195_/B gnd _7044_/C vdd NAND2X1
XFILL_0__14986_ gnd vdd FILL
XFILL_0__9484_ gnd vdd FILL
XSFILL94440x75050 gnd vdd FILL
XFILL_3__12028_ gnd vdd FILL
XFILL_3__8213_ gnd vdd FILL
XFILL_1__13207_ gnd vdd FILL
XFILL_2__15546_ gnd vdd FILL
XFILL_4__14367_ gnd vdd FILL
XFILL_4__11579_ gnd vdd FILL
XFILL_2__12758_ gnd vdd FILL
XFILL_1__10419_ gnd vdd FILL
XFILL_1__14187_ gnd vdd FILL
XSFILL29640x65050 gnd vdd FILL
XFILL_0__13937_ gnd vdd FILL
XFILL_5__9129_ gnd vdd FILL
XFILL_4__16106_ gnd vdd FILL
XFILL_1__11399_ gnd vdd FILL
XFILL_4__13318_ gnd vdd FILL
XFILL_5__15657_ gnd vdd FILL
XFILL_5__12869_ gnd vdd FILL
XSFILL69240x51050 gnd vdd FILL
XFILL_2__11709_ gnd vdd FILL
XFILL_3__8144_ gnd vdd FILL
XFILL_1__13138_ gnd vdd FILL
XFILL_4__14298_ gnd vdd FILL
XFILL_2__15477_ gnd vdd FILL
XFILL_0__13868_ gnd vdd FILL
XFILL_5__14608_ gnd vdd FILL
XFILL_4__16037_ gnd vdd FILL
XFILL_0__8366_ gnd vdd FILL
XFILL_4__13249_ gnd vdd FILL
XFILL_5__15588_ gnd vdd FILL
XFILL_2__14428_ gnd vdd FILL
XFILL_3__8075_ gnd vdd FILL
X_8994_ _8994_/A _9014_/A _8993_/Y gnd _9060_/D vdd OAI21X1
XFILL_0__15607_ gnd vdd FILL
XFILL_3__13979_ gnd vdd FILL
XFILL_0__7317_ gnd vdd FILL
XFILL_0__13799_ gnd vdd FILL
XFILL_5__14539_ gnd vdd FILL
X_7945_ _7937_/B _7177_/B gnd _7946_/C vdd NAND2X1
XFILL_3__15718_ gnd vdd FILL
XFILL_1__7090_ gnd vdd FILL
XFILL_2__14359_ gnd vdd FILL
XFILL_0__15538_ gnd vdd FILL
XFILL_0__7248_ gnd vdd FILL
XFILL_3__15649_ gnd vdd FILL
X_7876_ _7876_/A gnd _7876_/Y vdd INVX1
XSFILL89400x64050 gnd vdd FILL
XFILL_5__16209_ gnd vdd FILL
XFILL_0__15469_ gnd vdd FILL
X_9615_ _9615_/A _9615_/B gnd _9616_/C vdd NAND2X1
XFILL_0__7179_ gnd vdd FILL
XFILL_2__16029_ gnd vdd FILL
XSFILL110040x58050 gnd vdd FILL
XFILL_3__8977_ gnd vdd FILL
XFILL_1__9800_ gnd vdd FILL
X_9546_ _9586_/Q gnd _9546_/Y vdd INVX1
XFILL_1__7992_ gnd vdd FILL
XFILL_3__7928_ gnd vdd FILL
XFILL_6__7637_ gnd vdd FILL
XFILL_5_BUFX2_insert234 gnd vdd FILL
XFILL_5_BUFX2_insert245 gnd vdd FILL
XFILL_1__9731_ gnd vdd FILL
XFILL_1__6943_ gnd vdd FILL
XFILL_5_BUFX2_insert256 gnd vdd FILL
X_9477_ _9477_/A gnd _9479_/A vdd INVX1
XFILL_5_BUFX2_insert267 gnd vdd FILL
XSFILL95160x21050 gnd vdd FILL
XFILL_3__7859_ gnd vdd FILL
XFILL_5_BUFX2_insert278 gnd vdd FILL
X_8428_ _8376_/A _7661_/CLK _9203_/R vdd _8428_/D gnd vdd DFFSR
XFILL_1__9662_ gnd vdd FILL
XFILL_5_BUFX2_insert289 gnd vdd FILL
XFILL_1__6874_ gnd vdd FILL
XFILL_4_BUFX2_insert901 gnd vdd FILL
XSFILL83560x79050 gnd vdd FILL
XFILL_4__9371_ gnd vdd FILL
XFILL_4_BUFX2_insert912 gnd vdd FILL
XFILL_4_BUFX2_insert923 gnd vdd FILL
XFILL_1__8613_ gnd vdd FILL
XFILL_4_BUFX2_insert934 gnd vdd FILL
XFILL_4_BUFX2_insert945 gnd vdd FILL
X_10290_ _15863_/B gnd _10290_/Y vdd INVX1
XSFILL8600x79050 gnd vdd FILL
X_8359_ _8360_/B _7975_/B gnd _8359_/Y vdd NAND2X1
XFILL_4__8322_ gnd vdd FILL
XSFILL104520x40050 gnd vdd FILL
XFILL_1__9593_ gnd vdd FILL
XFILL_4_BUFX2_insert956 gnd vdd FILL
XFILL_3__9529_ gnd vdd FILL
XFILL_4_BUFX2_insert967 gnd vdd FILL
XFILL_4_BUFX2_insert978 gnd vdd FILL
XSFILL33800x72050 gnd vdd FILL
XFILL_4_BUFX2_insert989 gnd vdd FILL
XFILL_4__8253_ gnd vdd FILL
XFILL_4__7204_ gnd vdd FILL
XFILL_1__8475_ gnd vdd FILL
XSFILL104360x2050 gnd vdd FILL
XFILL_4__8184_ gnd vdd FILL
XFILL_1__7426_ gnd vdd FILL
X_13980_ _13980_/A gnd _15512_/B vdd INVX1
XFILL_2_BUFX2_insert102 gnd vdd FILL
XSFILL23480x62050 gnd vdd FILL
X_12931_ _12859_/A _8176_/CLK _8816_/R vdd _12931_/D gnd vdd DFFSR
XFILL_1__7357_ gnd vdd FILL
XFILL_4__7066_ gnd vdd FILL
XSFILL79160x34050 gnd vdd FILL
X_15650_ _15650_/A _15650_/B _15650_/C gnd _15651_/B vdd NOR3X1
X_12862_ _12932_/Q gnd _12862_/Y vdd INVX1
XSFILL113720x77050 gnd vdd FILL
XFILL_1__7288_ gnd vdd FILL
XFILL_1_BUFX2_insert802 gnd vdd FILL
X_14601_ _8894_/A gnd _14601_/Y vdd INVX1
X_11813_ _11005_/Y _11778_/B _11366_/B _11015_/D gnd _11815_/B vdd OAI22X1
XFILL_1_BUFX2_insert813 gnd vdd FILL
XFILL_1__9027_ gnd vdd FILL
X_15581_ _14088_/A _16311_/A _15581_/C _14101_/D gnd _15581_/Y vdd OAI22X1
XFILL_1_BUFX2_insert824 gnd vdd FILL
XFILL_1_BUFX2_insert835 gnd vdd FILL
X_12793_ _12701_/A _12667_/CLK _12809_/R vdd _12793_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert846 gnd vdd FILL
XSFILL18840x49050 gnd vdd FILL
X_14532_ _14532_/A _13879_/B _14862_/C _14532_/D gnd _14536_/B vdd OAI22X1
XFILL_1_BUFX2_insert857 gnd vdd FILL
XFILL_1_BUFX2_insert868 gnd vdd FILL
X_11744_ _11744_/A _11050_/Y _11743_/Y gnd _11753_/B vdd AOI21X1
XSFILL84280x25050 gnd vdd FILL
XFILL_1_BUFX2_insert879 gnd vdd FILL
XBUFX2_insert101 _15009_/Y gnd _15683_/C vdd BUFX2
X_14463_ _13868_/B _14463_/B _14872_/C _14461_/Y gnd _14467_/B vdd OAI22X1
XFILL_4__7968_ gnd vdd FILL
XSFILL99320x47050 gnd vdd FILL
X_11675_ _11675_/A gnd _12482_/B vdd INVX1
XFILL_4__10950_ gnd vdd FILL
XFILL_2__10040_ gnd vdd FILL
XFILL_2__9771_ gnd vdd FILL
XFILL_2__6983_ gnd vdd FILL
XFILL_5__8500_ gnd vdd FILL
X_16202_ _16202_/A _16180_/Y _16202_/C gnd _16203_/B vdd NOR3X1
X_13414_ _13410_/Y _13630_/B _13633_/C _13411_/Y gnd _13414_/Y vdd OAI22X1
XFILL_1__10770_ gnd vdd FILL
XFILL_4__6919_ gnd vdd FILL
XFILL_5__10151_ gnd vdd FILL
XFILL_5__9480_ gnd vdd FILL
X_10626_ _15235_/A gnd _10626_/Y vdd INVX1
XFILL_6__12490_ gnd vdd FILL
X_14394_ _9577_/Q gnd _14394_/Y vdd INVX1
XFILL_3__11330_ gnd vdd FILL
XFILL_4__10881_ gnd vdd FILL
XFILL_2__8722_ gnd vdd FILL
XFILL_1__9929_ gnd vdd FILL
XFILL_0__11150_ gnd vdd FILL
XFILL_4__9638_ gnd vdd FILL
X_16133_ _7281_/Q _15177_/B _16014_/C _8305_/Q gnd _16139_/B vdd AOI22X1
X_13345_ _13259_/C _13294_/A gnd _13345_/Y vdd NOR2X1
XFILL_6__11441_ gnd vdd FILL
XFILL_4__12620_ gnd vdd FILL
X_10557_ _10557_/A _10557_/B _10556_/Y gnd _10557_/Y vdd OAI21X1
XFILL_2__8653_ gnd vdd FILL
XFILL_3__11261_ gnd vdd FILL
XFILL_1__12440_ gnd vdd FILL
XSFILL43880x2050 gnd vdd FILL
XFILL_5_BUFX2_insert790 gnd vdd FILL
XFILL_2__11991_ gnd vdd FILL
XFILL_5__8362_ gnd vdd FILL
XFILL_0__11081_ gnd vdd FILL
XFILL_3__13000_ gnd vdd FILL
XFILL_6__14160_ gnd vdd FILL
X_16064_ _16063_/Y _16099_/B _16099_/C _14665_/B gnd _16064_/Y vdd OAI22X1
XFILL_5__13910_ gnd vdd FILL
X_13276_ _13297_/C _13276_/B gnd _13276_/Y vdd NOR2X1
XFILL_2__7604_ gnd vdd FILL
X_10488_ _10486_/Y _10505_/A _10488_/C gnd _10582_/D vdd OAI21X1
XFILL_2__13730_ gnd vdd FILL
XFILL_5__14890_ gnd vdd FILL
XFILL_2__10942_ gnd vdd FILL
XFILL_2__8584_ gnd vdd FILL
XFILL_0__10032_ gnd vdd FILL
XSFILL79240x14050 gnd vdd FILL
XFILL_5__7313_ gnd vdd FILL
XFILL_3__11192_ gnd vdd FILL
XFILL112120x71050 gnd vdd FILL
XFILL_1__12371_ gnd vdd FILL
X_15015_ _14983_/A _15061_/C _16035_/B gnd _15015_/Y vdd NAND3X1
X_12227_ _12227_/A gnd _12239_/C gnd _12227_/Y vdd NAND3X1
XFILL_5__13841_ gnd vdd FILL
XFILL_4__11502_ gnd vdd FILL
XFILL_4__12482_ gnd vdd FILL
XFILL_1__14110_ gnd vdd FILL
XFILL_3__10143_ gnd vdd FILL
XFILL_4__15270_ gnd vdd FILL
XFILL_2__13661_ gnd vdd FILL
XFILL_1__11322_ gnd vdd FILL
XFILL_0__14840_ gnd vdd FILL
XFILL_5__7244_ gnd vdd FILL
XFILL_1__15090_ gnd vdd FILL
XFILL_2__10873_ gnd vdd FILL
XFILL_6__13042_ gnd vdd FILL
XSFILL114440x23050 gnd vdd FILL
XFILL_6__10254_ gnd vdd FILL
XFILL_2__15400_ gnd vdd FILL
XFILL_4__14221_ gnd vdd FILL
X_12158_ _12134_/A _12865_/A gnd _12159_/C vdd NAND2X1
XFILL_4__11433_ gnd vdd FILL
XFILL_2__12612_ gnd vdd FILL
XFILL_5__13772_ gnd vdd FILL
XFILL_1__14041_ gnd vdd FILL
XFILL_3__14951_ gnd vdd FILL
XFILL_2__16380_ gnd vdd FILL
XFILL_2__7466_ gnd vdd FILL
XFILL_2__13592_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1079 gnd vdd FILL
XFILL_1__11253_ gnd vdd FILL
XFILL_5__15511_ gnd vdd FILL
XFILL_5__7175_ gnd vdd FILL
X_11109_ _12302_/Y gnd _11109_/Y vdd INVX1
XFILL_0__14771_ gnd vdd FILL
XFILL_5__12723_ gnd vdd FILL
XFILL_0__11983_ gnd vdd FILL
XSFILL89240x1050 gnd vdd FILL
XFILL_2__15331_ gnd vdd FILL
XFILL_4__14152_ gnd vdd FILL
X_12089_ _12089_/A _12113_/B _12061_/C gnd gnd _12089_/Y vdd AOI22X1
XFILL_3__13902_ gnd vdd FILL
XFILL_4__11364_ gnd vdd FILL
XFILL_1__11184_ gnd vdd FILL
XFILL_0__13722_ gnd vdd FILL
XFILL_3__14882_ gnd vdd FILL
XFILL_0__10934_ gnd vdd FILL
XSFILL69160x66050 gnd vdd FILL
XFILL_0__8220_ gnd vdd FILL
XSFILL99400x27050 gnd vdd FILL
XFILL_4__10315_ gnd vdd FILL
X_15917_ _15917_/A _15917_/B _15917_/C gnd _15928_/A vdd NAND3X1
XFILL_4__13103_ gnd vdd FILL
XFILL_5__15442_ gnd vdd FILL
XFILL_5__12654_ gnd vdd FILL
XFILL_2__9136_ gnd vdd FILL
XFILL_4__14083_ gnd vdd FILL
XFILL_3__13833_ gnd vdd FILL
XFILL_1__10135_ gnd vdd FILL
XFILL_4__11295_ gnd vdd FILL
XFILL_2__15262_ gnd vdd FILL
XFILL_2__12474_ gnd vdd FILL
XFILL_0__13653_ gnd vdd FILL
XFILL_1__15992_ gnd vdd FILL
XFILL_4__13034_ gnd vdd FILL
XFILL_5__11605_ gnd vdd FILL
XFILL_2__14213_ gnd vdd FILL
XFILL_5__15373_ gnd vdd FILL
X_15848_ _15848_/A _15848_/B _15524_/A _15848_/D gnd _15848_/Y vdd OAI22X1
XFILL_4__10246_ gnd vdd FILL
XSFILL104360x75050 gnd vdd FILL
XFILL_5__12585_ gnd vdd FILL
XFILL_2__11425_ gnd vdd FILL
XFILL_3__10976_ gnd vdd FILL
XFILL_0__12604_ gnd vdd FILL
XFILL_2__15193_ gnd vdd FILL
XFILL_3__13764_ gnd vdd FILL
XFILL_2_BUFX2_insert680 gnd vdd FILL
XFILL_1__14943_ gnd vdd FILL
XFILL_1__10066_ gnd vdd FILL
XFILL_0__7102_ gnd vdd FILL
XFILL_0__16372_ gnd vdd FILL
XFILL_2_BUFX2_insert691 gnd vdd FILL
XSFILL74280x57050 gnd vdd FILL
XFILL_5__14324_ gnd vdd FILL
XFILL_0__10796_ gnd vdd FILL
XFILL_0__13584_ gnd vdd FILL
XFILL_3__15503_ gnd vdd FILL
X_7730_ _7786_/Q gnd _7730_/Y vdd INVX1
XFILL_0__8082_ gnd vdd FILL
XFILL_5__11536_ gnd vdd FILL
XFILL_2__8018_ gnd vdd FILL
XFILL_3__12715_ gnd vdd FILL
XFILL_2__14144_ gnd vdd FILL
X_15779_ _7212_/A _15177_/B _16014_/C _8236_/A gnd _15779_/Y vdd AOI22X1
XFILL_3__8900_ gnd vdd FILL
XFILL_4__10177_ gnd vdd FILL
XFILL_0__15323_ gnd vdd FILL
XFILL_2__11356_ gnd vdd FILL
XFILL_3__13695_ gnd vdd FILL
XFILL_1__14874_ gnd vdd FILL
XFILL_3__9880_ gnd vdd FILL
XFILL_0__7033_ gnd vdd FILL
XFILL_6__12826_ gnd vdd FILL
XFILL_5__14255_ gnd vdd FILL
XSFILL49080x33050 gnd vdd FILL
XFILL_3__12646_ gnd vdd FILL
X_7661_ _7611_/A _7661_/CLK _7789_/R vdd _7661_/D gnd vdd DFFSR
XFILL112200x51050 gnd vdd FILL
XFILL_2__10307_ gnd vdd FILL
XFILL_3__15434_ gnd vdd FILL
XFILL_5__11467_ gnd vdd FILL
XFILL_3__8831_ gnd vdd FILL
XFILL_1__13825_ gnd vdd FILL
XFILL_4__14985_ gnd vdd FILL
XFILL_2__14075_ gnd vdd FILL
XFILL_5_BUFX2_insert40 gnd vdd FILL
XFILL_0__15254_ gnd vdd FILL
XFILL_2__11287_ gnd vdd FILL
XFILL_5_BUFX2_insert51 gnd vdd FILL
XFILL_0__12466_ gnd vdd FILL
X_9400_ _9400_/A gnd _9400_/Y vdd INVX1
XFILL_5__9747_ gnd vdd FILL
XFILL_5_BUFX2_insert62 gnd vdd FILL
XFILL_5__6959_ gnd vdd FILL
XFILL_5__10418_ gnd vdd FILL
XFILL_5__14186_ gnd vdd FILL
XFILL_2__13026_ gnd vdd FILL
XFILL_4__13936_ gnd vdd FILL
X_7592_ _7592_/A _7592_/B _7591_/Y gnd _7592_/Y vdd OAI21X1
XFILL_5_BUFX2_insert73 gnd vdd FILL
XFILL_3__12577_ gnd vdd FILL
XFILL_3__15365_ gnd vdd FILL
XFILL_0__14205_ gnd vdd FILL
XFILL_5__11398_ gnd vdd FILL
XFILL_2__10238_ gnd vdd FILL
XFILL_1__13756_ gnd vdd FILL
XFILL_5_BUFX2_insert84 gnd vdd FILL
XFILL_3__8762_ gnd vdd FILL
XFILL_0__11417_ gnd vdd FILL
XFILL_1__10968_ gnd vdd FILL
XFILL_0__15185_ gnd vdd FILL
XFILL_5_BUFX2_insert95 gnd vdd FILL
XFILL_0__12397_ gnd vdd FILL
X_9331_ _9293_/A _7021_/CLK _9062_/R vdd _9331_/D gnd vdd DFFSR
XFILL_5__9678_ gnd vdd FILL
XSFILL4440x48050 gnd vdd FILL
XFILL_5__13137_ gnd vdd FILL
XSFILL13560x74050 gnd vdd FILL
XFILL_0__8984_ gnd vdd FILL
XFILL_3__14316_ gnd vdd FILL
XFILL_3__11528_ gnd vdd FILL
XFILL_4__13867_ gnd vdd FILL
XFILL_1__12707_ gnd vdd FILL
XFILL_3__7713_ gnd vdd FILL
XSFILL49000x4050 gnd vdd FILL
XFILL_3__15296_ gnd vdd FILL
XFILL_0__14136_ gnd vdd FILL
XFILL_2__10169_ gnd vdd FILL
XBUFX2_insert690 _13362_/Y gnd _10548_/B vdd BUFX2
XFILL_5__8629_ gnd vdd FILL
XFILL_1__13687_ gnd vdd FILL
XFILL_0__11348_ gnd vdd FILL
XFILL_0__7935_ gnd vdd FILL
XFILL_1__10899_ gnd vdd FILL
XFILL_4__15606_ gnd vdd FILL
X_9262_ _9262_/A _9208_/B _9261_/Y gnd _9262_/Y vdd OAI21X1
XFILL_3__14247_ gnd vdd FILL
XSFILL69240x46050 gnd vdd FILL
XFILL_3__11459_ gnd vdd FILL
XFILL_1__15426_ gnd vdd FILL
XFILL_1__12638_ gnd vdd FILL
XFILL_4__13798_ gnd vdd FILL
XFILL_0__14067_ gnd vdd FILL
XFILL_6__7353_ gnd vdd FILL
XFILL_2__14977_ gnd vdd FILL
XFILL_0__11279_ gnd vdd FILL
XFILL_5__12019_ gnd vdd FILL
X_8213_ _8244_/B _8853_/B gnd _8214_/C vdd NAND2X1
XFILL_0__7866_ gnd vdd FILL
XFILL_4__15537_ gnd vdd FILL
XFILL_4__12749_ gnd vdd FILL
XFILL_3__14178_ gnd vdd FILL
X_9193_ _9193_/Q _9705_/CLK _7649_/R vdd _9193_/D gnd vdd DFFSR
XFILL_1__15357_ gnd vdd FILL
XFILL_0__13018_ gnd vdd FILL
XFILL_3__7575_ gnd vdd FILL
XFILL_2__13928_ gnd vdd FILL
XFILL_1__12569_ gnd vdd FILL
XSFILL104440x55050 gnd vdd FILL
XSFILL8760x50 gnd vdd FILL
XFILL_0__9605_ gnd vdd FILL
XFILL_3__13129_ gnd vdd FILL
X_8144_ _8180_/Q gnd _8146_/A vdd INVX1
XFILL_1__14308_ gnd vdd FILL
XFILL_4__15468_ gnd vdd FILL
XFILL_3_BUFX2_insert908 gnd vdd FILL
XSFILL8680x53050 gnd vdd FILL
XFILL_2__13859_ gnd vdd FILL
XFILL_3_BUFX2_insert919 gnd vdd FILL
XFILL_1__15288_ gnd vdd FILL
XFILL_0__9536_ gnd vdd FILL
XFILL_4__14419_ gnd vdd FILL
X_8075_ _8157_/Q gnd _8077_/A vdd INVX1
XFILL_3__9245_ gnd vdd FILL
XFILL_4__15399_ gnd vdd FILL
XFILL_1__14239_ gnd vdd FILL
XSFILL89400x59050 gnd vdd FILL
XFILL_0__14969_ gnd vdd FILL
X_7026_ _6986_/A _8537_/CLK _8166_/R vdd _6988_/Y gnd vdd DFFSR
XFILL_5__15709_ gnd vdd FILL
XFILL_1__8260_ gnd vdd FILL
XFILL_0__9467_ gnd vdd FILL
XFILL_2__15529_ gnd vdd FILL
XFILL_1__7211_ gnd vdd FILL
XFILL_3__8127_ gnd vdd FILL
XFILL_1__8191_ gnd vdd FILL
XFILL_0__9398_ gnd vdd FILL
XSFILL13640x54050 gnd vdd FILL
XFILL_0__8349_ gnd vdd FILL
XFILL_3__8058_ gnd vdd FILL
X_8977_ _9055_/Q gnd _8979_/A vdd INVX1
XFILL_1_BUFX2_insert109 gnd vdd FILL
XSFILL69320x26050 gnd vdd FILL
XFILL_1__7073_ gnd vdd FILL
X_7928_ _7928_/A _7972_/A _7928_/C gnd _7928_/Y vdd OAI21X1
XFILL_4__8871_ gnd vdd FILL
XFILL_0_CLKBUF1_insert202 gnd vdd FILL
XFILL_6__9787_ gnd vdd FILL
XFILL_0_CLKBUF1_insert213 gnd vdd FILL
XSFILL104520x35050 gnd vdd FILL
X_7859_ _7892_/A _9779_/B gnd _7860_/C vdd NAND2X1
XFILL_0_CLKBUF1_insert224 gnd vdd FILL
XFILL_4__7822_ gnd vdd FILL
XFILL_0_BUFX2_insert809 gnd vdd FILL
XFILL_6__8738_ gnd vdd FILL
XSFILL8760x33050 gnd vdd FILL
XSFILL33800x67050 gnd vdd FILL
XFILL_1_BUFX2_insert1006 gnd vdd FILL
XFILL_1_BUFX2_insert1017 gnd vdd FILL
XFILL_4__7753_ gnd vdd FILL
XFILL_1_BUFX2_insert1028 gnd vdd FILL
X_11460_ _11502_/B _11189_/Y _11174_/C gnd _11461_/C vdd OAI21X1
XFILL_1_BUFX2_insert1039 gnd vdd FILL
X_9529_ _9529_/A _9785_/B gnd _9530_/C vdd NAND2X1
XFILL_1__7975_ gnd vdd FILL
XFILL_4__7684_ gnd vdd FILL
X_10411_ _10409_/Y _10395_/A _10411_/C gnd _10471_/D vdd OAI21X1
XFILL_1__6926_ gnd vdd FILL
X_11391_ _11081_/C gnd _11392_/C vdd INVX1
XFILL_4__9423_ gnd vdd FILL
X_13130_ _13192_/Q gnd _13130_/Y vdd INVX1
X_10342_ _14221_/A _8562_/CLK _7270_/R vdd _10342_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert720 gnd vdd FILL
XFILL_4_BUFX2_insert731 gnd vdd FILL
XFILL_1__6857_ gnd vdd FILL
XFILL_1__9645_ gnd vdd FILL
XFILL_4_BUFX2_insert742 gnd vdd FILL
XSFILL13720x34050 gnd vdd FILL
XFILL_4__9354_ gnd vdd FILL
XFILL_4_BUFX2_insert753 gnd vdd FILL
XFILL_4_BUFX2_insert764 gnd vdd FILL
X_13061_ _6884_/A _13184_/CLK _8033_/R vdd _13061_/D gnd vdd DFFSR
XSFILL79160x29050 gnd vdd FILL
XFILL_3_CLKBUF1_insert1074 gnd vdd FILL
X_10273_ _10294_/A _9889_/B gnd _10274_/C vdd NAND2X1
XFILL_4_BUFX2_insert775 gnd vdd FILL
XFILL_4_BUFX2_insert786 gnd vdd FILL
X_12012_ _12012_/A _12707_/A _11996_/C gnd _12012_/Y vdd NAND3X1
XFILL_4__9285_ gnd vdd FILL
XFILL_4_BUFX2_insert797 gnd vdd FILL
XFILL_1__8527_ gnd vdd FILL
XFILL_2__7320_ gnd vdd FILL
XFILL_4__8236_ gnd vdd FILL
XFILL_1__8458_ gnd vdd FILL
XFILL_2__7251_ gnd vdd FILL
X_13963_ _13963_/A _13963_/B _13960_/Y gnd _13974_/B vdd NAND3X1
XFILL_2__7182_ gnd vdd FILL
XFILL_4__7118_ gnd vdd FILL
XFILL_1__8389_ gnd vdd FILL
X_15702_ _15699_/Y _15702_/B _15702_/C gnd _15705_/C vdd NOR3X1
XFILL_4__8098_ gnd vdd FILL
X_12914_ vdd _16283_/Y gnd _12914_/Y vdd NAND2X1
XFILL_5__8980_ gnd vdd FILL
XFILL_3__10830_ gnd vdd FILL
XFILL_4__11080_ gnd vdd FILL
X_13894_ _13893_/Y _13894_/B gnd _13897_/C vdd NOR2X1
XFILL_4__7049_ gnd vdd FILL
XFILL_0__10650_ gnd vdd FILL
XFILL_5__7931_ gnd vdd FILL
XFILL_6__10941_ gnd vdd FILL
X_12845_ vdd _12845_/B gnd _12846_/C vdd NAND2X1
XFILL_1_BUFX2_insert610 gnd vdd FILL
X_15633_ _16235_/A _15633_/B _14137_/Y _15633_/D gnd _15633_/Y vdd OAI22X1
XFILL_4__10031_ gnd vdd FILL
XFILL_5__12370_ gnd vdd FILL
XFILL_2__11210_ gnd vdd FILL
XFILL_3__10761_ gnd vdd FILL
XFILL_1_BUFX2_insert621 gnd vdd FILL
XFILL_1_BUFX2_insert632 gnd vdd FILL
XFILL_1__11940_ gnd vdd FILL
XFILL_2__12190_ gnd vdd FILL
XFILL_1_BUFX2_insert643 gnd vdd FILL
XFILL_0__10581_ gnd vdd FILL
XFILL_5__7862_ gnd vdd FILL
XFILL_1_BUFX2_insert654 gnd vdd FILL
XFILL_3__12500_ gnd vdd FILL
XFILL_5__11321_ gnd vdd FILL
X_12776_ _12818_/Q gnd _12776_/Y vdd INVX1
X_15564_ _15564_/A _15564_/B gnd _15564_/Y vdd NOR2X1
XSFILL13800x14050 gnd vdd FILL
XFILL_3__13480_ gnd vdd FILL
XFILL_2__11141_ gnd vdd FILL
XFILL_1_BUFX2_insert665 gnd vdd FILL
XFILL_5__9601_ gnd vdd FILL
XFILL_3__10692_ gnd vdd FILL
XFILL_0__12320_ gnd vdd FILL
XFILL_1_BUFX2_insert676 gnd vdd FILL
XFILL112120x66050 gnd vdd FILL
XFILL_1_BUFX2_insert687 gnd vdd FILL
XFILL_1__11871_ gnd vdd FILL
X_14515_ _14515_/A _13813_/B _14160_/B _14513_/Y gnd _14519_/A vdd OAI22X1
XFILL_5__14040_ gnd vdd FILL
X_11727_ _11724_/Y _11726_/Y _11727_/C gnd _12029_/A vdd NAND3X1
XFILL_1_BUFX2_insert698 gnd vdd FILL
XFILL_3__12431_ gnd vdd FILL
X_15495_ _15495_/A _15495_/B _15482_/Y gnd _15495_/Y vdd NAND3X1
XFILL_5__11252_ gnd vdd FILL
XFILL_1__13610_ gnd vdd FILL
XFILL_4__14770_ gnd vdd FILL
XSFILL64040x51050 gnd vdd FILL
XFILL_4__11982_ gnd vdd FILL
XFILL_1__10822_ gnd vdd FILL
XFILL_0__12251_ gnd vdd FILL
XFILL_2__11072_ gnd vdd FILL
XFILL_5__9532_ gnd vdd FILL
XFILL_1__14590_ gnd vdd FILL
X_11658_ _11658_/A _11285_/A _11657_/Y gnd _11658_/Y vdd OAI21X1
XFILL_5__11183_ gnd vdd FILL
XFILL_3__15150_ gnd vdd FILL
XFILL_4__13721_ gnd vdd FILL
X_14446_ _14738_/A _7402_/Q _7914_/Q _13865_/B gnd _14448_/A vdd AOI22X1
XFILL_4__10933_ gnd vdd FILL
XFILL_3__12362_ gnd vdd FILL
XFILL_2__10023_ gnd vdd FILL
XFILL_2__14900_ gnd vdd FILL
XFILL_2__6966_ gnd vdd FILL
XFILL_2__9754_ gnd vdd FILL
XFILL_1__13541_ gnd vdd FILL
XFILL_0__11202_ gnd vdd FILL
XFILL_1__10753_ gnd vdd FILL
XFILL_0__12182_ gnd vdd FILL
XFILL_2__15880_ gnd vdd FILL
XFILL_5__9463_ gnd vdd FILL
X_10609_ _14763_/B _8433_/CLK _7921_/R vdd _10609_/D gnd vdd DFFSR
X_14377_ _14376_/Y _14377_/B gnd _14378_/C vdd NOR2X1
XFILL_3__11313_ gnd vdd FILL
XFILL_5__10134_ gnd vdd FILL
XFILL_3__14101_ gnd vdd FILL
XFILL_2__8705_ gnd vdd FILL
XFILL_4__13652_ gnd vdd FILL
XFILL_5__15991_ gnd vdd FILL
XFILL_3__15081_ gnd vdd FILL
X_11589_ _11571_/A _11589_/B _11589_/C gnd _11600_/A vdd NAND3X1
XFILL_2__14831_ gnd vdd FILL
XFILL_3__12293_ gnd vdd FILL
XFILL_0__11133_ gnd vdd FILL
XFILL_1__16260_ gnd vdd FILL
XFILL_1__13472_ gnd vdd FILL
XFILL_2__9685_ gnd vdd FILL
XFILL_2__6897_ gnd vdd FILL
XFILL_1__10684_ gnd vdd FILL
XFILL_0__7720_ gnd vdd FILL
X_13328_ _13235_/C _13209_/Y gnd _13328_/Y vdd NAND2X1
X_16116_ _16115_/Y _16116_/B gnd _16122_/A vdd NOR2X1
XFILL_4__12603_ gnd vdd FILL
XFILL_3__14032_ gnd vdd FILL
XFILL_5__14942_ gnd vdd FILL
XFILL_5__9394_ gnd vdd FILL
XFILL_5__10065_ gnd vdd FILL
XFILL_4__16371_ gnd vdd FILL
XFILL_1__15211_ gnd vdd FILL
XFILL_3__11244_ gnd vdd FILL
XFILL_2__8636_ gnd vdd FILL
XFILL_1__12423_ gnd vdd FILL
XFILL_4__10795_ gnd vdd FILL
XFILL_4__13583_ gnd vdd FILL
XFILL_2__14762_ gnd vdd FILL
XFILL_2__11974_ gnd vdd FILL
XFILL_1__16191_ gnd vdd FILL
XFILL_0__15941_ gnd vdd FILL
XFILL_0__11064_ gnd vdd FILL
XSFILL84200x64050 gnd vdd FILL
XFILL_5__8345_ gnd vdd FILL
X_13259_ _13258_/Y _13326_/A _13259_/C gnd _13263_/C vdd OAI21X1
XFILL_4__15322_ gnd vdd FILL
X_16047_ _9281_/A _15892_/B gnd _16047_/Y vdd NAND2X1
XFILL_5__14873_ gnd vdd FILL
XSFILL70040x70050 gnd vdd FILL
XFILL_4__12534_ gnd vdd FILL
XFILL_2__8567_ gnd vdd FILL
XFILL_2__10925_ gnd vdd FILL
XFILL_3__7360_ gnd vdd FILL
XFILL_0__10015_ gnd vdd FILL
XFILL_2__13713_ gnd vdd FILL
XFILL_1__15142_ gnd vdd FILL
XFILL_3__11175_ gnd vdd FILL
XFILL_1__12354_ gnd vdd FILL
XFILL_2__14693_ gnd vdd FILL
XFILL_5__8276_ gnd vdd FILL
XFILL_0__15872_ gnd vdd FILL
XFILL_5__13824_ gnd vdd FILL
XSFILL59000x40050 gnd vdd FILL
XFILL_3__10126_ gnd vdd FILL
XFILL_4__15253_ gnd vdd FILL
XFILL_0__7582_ gnd vdd FILL
XFILL_2__13644_ gnd vdd FILL
XFILL_4__12465_ gnd vdd FILL
XFILL_1__11305_ gnd vdd FILL
XFILL_3__15983_ gnd vdd FILL
XFILL_0__14823_ gnd vdd FILL
XFILL_1__15073_ gnd vdd FILL
XFILL_2__8498_ gnd vdd FILL
XFILL_3__7291_ gnd vdd FILL
XFILL_5__7227_ gnd vdd FILL
XFILL_1__12285_ gnd vdd FILL
XFILL_4__14204_ gnd vdd FILL
XFILL_5__13755_ gnd vdd FILL
XFILL_3__9030_ gnd vdd FILL
XFILL_4__11416_ gnd vdd FILL
XFILL_5__10967_ gnd vdd FILL
XFILL_4__15184_ gnd vdd FILL
XFILL_2__16363_ gnd vdd FILL
XFILL112200x46050 gnd vdd FILL
XFILL_2__7449_ gnd vdd FILL
XFILL_1__14024_ gnd vdd FILL
XFILL_3__14934_ gnd vdd FILL
XFILL_3__10057_ gnd vdd FILL
XFILL_4__12396_ gnd vdd FILL
XFILL_2__13575_ gnd vdd FILL
XFILL_1__11236_ gnd vdd FILL
XFILL_2__10787_ gnd vdd FILL
XFILL_2_CLKBUF1_insert190 gnd vdd FILL
XFILL_5__7158_ gnd vdd FILL
XSFILL89480x33050 gnd vdd FILL
XFILL_0__14754_ gnd vdd FILL
XFILL_5__12706_ gnd vdd FILL
XFILL_0__9252_ gnd vdd FILL
XFILL_0__11966_ gnd vdd FILL
X_8900_ _8900_/A gnd _8902_/A vdd INVX1
XFILL_4__14135_ gnd vdd FILL
XSFILL64120x31050 gnd vdd FILL
XFILL_5__13686_ gnd vdd FILL
XFILL_2__15314_ gnd vdd FILL
XFILL_2__12526_ gnd vdd FILL
X_9880_ _9896_/B _6936_/B gnd _9881_/C vdd NAND2X1
XFILL_4__11347_ gnd vdd FILL
XFILL_5__10898_ gnd vdd FILL
XFILL_3__14865_ gnd vdd FILL
XFILL_0__13705_ gnd vdd FILL
XFILL_2__16294_ gnd vdd FILL
XFILL_0__10917_ gnd vdd FILL
XFILL_0__8203_ gnd vdd FILL
XFILL_1__11167_ gnd vdd FILL
XFILL_5__7089_ gnd vdd FILL
XFILL_0__14685_ gnd vdd FILL
XFILL_5__15425_ gnd vdd FILL
X_8831_ _8831_/A gnd _8833_/A vdd INVX1
XFILL_5__12637_ gnd vdd FILL
XFILL_0__11897_ gnd vdd FILL
XFILL_3__13816_ gnd vdd FILL
XFILL_2__15245_ gnd vdd FILL
XFILL_4__14066_ gnd vdd FILL
XFILL_2__9119_ gnd vdd FILL
XFILL_4__11278_ gnd vdd FILL
XFILL_2__12457_ gnd vdd FILL
XBUFX2_insert1 _12381_/Y gnd _7451_/B vdd BUFX2
XFILL_1__10118_ gnd vdd FILL
XFILL_0__13636_ gnd vdd FILL
XFILL_1__15975_ gnd vdd FILL
XFILL_3__14796_ gnd vdd FILL
XFILL_0__8134_ gnd vdd FILL
XFILL_1__11098_ gnd vdd FILL
XFILL_5__15356_ gnd vdd FILL
XFILL_4__13017_ gnd vdd FILL
XFILL_5__12568_ gnd vdd FILL
X_8762_ _8760_/Y _8714_/B _8762_/C gnd _8812_/D vdd OAI21X1
XFILL_2__11408_ gnd vdd FILL
XFILL_2__15176_ gnd vdd FILL
XFILL_3__13747_ gnd vdd FILL
XFILL_3__9932_ gnd vdd FILL
XFILL_3__10959_ gnd vdd FILL
XFILL_2__12388_ gnd vdd FILL
XFILL_0__16355_ gnd vdd FILL
XSFILL43400x32050 gnd vdd FILL
XFILL_1__10049_ gnd vdd FILL
XFILL_1__14926_ gnd vdd FILL
XFILL_5__14307_ gnd vdd FILL
XFILL_0__13567_ gnd vdd FILL
XFILL_0__8065_ gnd vdd FILL
XFILL_6__6853_ gnd vdd FILL
X_7713_ _7684_/B _7713_/B gnd _7713_/Y vdd NAND2X1
XFILL_0__10779_ gnd vdd FILL
XFILL_5__11519_ gnd vdd FILL
XFILL_6__13858_ gnd vdd FILL
XFILL_2__14127_ gnd vdd FILL
XFILL_5__15287_ gnd vdd FILL
XSFILL54040x83050 gnd vdd FILL
XFILL_0__15306_ gnd vdd FILL
XFILL_5__12499_ gnd vdd FILL
XFILL_6_BUFX2_insert848 gnd vdd FILL
XFILL_2__11339_ gnd vdd FILL
X_8693_ _8659_/A _9205_/CLK _7285_/R vdd _8661_/Y gnd vdd DFFSR
XFILL_1__14857_ gnd vdd FILL
XFILL_3__13678_ gnd vdd FILL
XFILL_0__12518_ gnd vdd FILL
XFILL_3__9863_ gnd vdd FILL
XFILL_0__16286_ gnd vdd FILL
XFILL_5__14238_ gnd vdd FILL
XFILL_0__13498_ gnd vdd FILL
X_7644_ _7560_/A _9436_/CLK _7644_/R vdd _7562_/Y gnd vdd DFFSR
XFILL_3__15417_ gnd vdd FILL
XFILL_1__13808_ gnd vdd FILL
XFILL_3__12629_ gnd vdd FILL
XFILL_2__14058_ gnd vdd FILL
XFILL_4__14968_ gnd vdd FILL
XSFILL73880x25050 gnd vdd FILL
XFILL_0__15237_ gnd vdd FILL
XSFILL8680x48050 gnd vdd FILL
XFILL_3__16397_ gnd vdd FILL
XFILL_0__12449_ gnd vdd FILL
XFILL_3__9794_ gnd vdd FILL
XFILL_1__14788_ gnd vdd FILL
XFILL_5__14169_ gnd vdd FILL
XSFILL33880x41050 gnd vdd FILL
XFILL_2__13009_ gnd vdd FILL
XFILL_4__13919_ gnd vdd FILL
XFILL_3__15348_ gnd vdd FILL
X_7575_ _7575_/A gnd _7577_/A vdd INVX1
XFILL_3__8745_ gnd vdd FILL
XFILL_4__14899_ gnd vdd FILL
XFILL_1__13739_ gnd vdd FILL
XFILL_0__15168_ gnd vdd FILL
X_9314_ _9314_/Q _8818_/CLK _8278_/R vdd _9314_/D gnd vdd DFFSR
XFILL_6__8454_ gnd vdd FILL
XFILL_6__15459_ gnd vdd FILL
XFILL_1__7760_ gnd vdd FILL
XSFILL48920x63050 gnd vdd FILL
XFILL_0__8967_ gnd vdd FILL
XFILL_0__14119_ gnd vdd FILL
XFILL_3__15279_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1080 gnd vdd FILL
XSFILL64200x11050 gnd vdd FILL
XFILL_0__15099_ gnd vdd FILL
X_9245_ _9245_/A gnd _9247_/A vdd INVX1
XFILL_1__7691_ gnd vdd FILL
XFILL_1__15409_ gnd vdd FILL
XFILL_0__8898_ gnd vdd FILL
XFILL_3__7627_ gnd vdd FILL
XFILL_1__16389_ gnd vdd FILL
XSFILL49000x72050 gnd vdd FILL
XSFILL13640x49050 gnd vdd FILL
XFILL_0__7849_ gnd vdd FILL
X_9176_ _9176_/Q _7143_/CLK _7015_/R vdd _9176_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert705 gnd vdd FILL
XFILL_3__7558_ gnd vdd FILL
XFILL_3_BUFX2_insert716 gnd vdd FILL
XSFILL109560x83050 gnd vdd FILL
X_8127_ _8079_/A _7743_/B gnd _8127_/Y vdd NAND2X1
XFILL_1__9361_ gnd vdd FILL
XFILL_3_BUFX2_insert727 gnd vdd FILL
XFILL_3_BUFX2_insert738 gnd vdd FILL
XFILL_3_BUFX2_insert749 gnd vdd FILL
XSFILL28840x30050 gnd vdd FILL
XFILL_3__7489_ gnd vdd FILL
XFILL_1__8312_ gnd vdd FILL
XFILL_0__9519_ gnd vdd FILL
XFILL_6__7198_ gnd vdd FILL
XFILL_1__9292_ gnd vdd FILL
XFILL_4__8021_ gnd vdd FILL
X_8058_ _8107_/B _9978_/B gnd _8059_/C vdd NAND2X1
XFILL_3__9228_ gnd vdd FILL
XFILL_1_BUFX2_insert60 gnd vdd FILL
X_7009_ _6935_/A _7916_/CLK _7276_/R vdd _7009_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert71 gnd vdd FILL
XFILL_1__8243_ gnd vdd FILL
XFILL_1_BUFX2_insert82 gnd vdd FILL
XFILL_1_BUFX2_insert93 gnd vdd FILL
XFILL_3__9159_ gnd vdd FILL
XSFILL33960x21050 gnd vdd FILL
X_10960_ _10930_/Y _10952_/Y gnd _10969_/C vdd NAND2X1
XSFILL18760x82050 gnd vdd FILL
XFILL_1__7125_ gnd vdd FILL
X_10891_ _10871_/Y gnd _10891_/Y vdd INVX1
X_12630_ _12407_/B gnd _12632_/A vdd INVX1
XFILL_1__7056_ gnd vdd FILL
XSFILL13720x29050 gnd vdd FILL
XFILL_4__8854_ gnd vdd FILL
XFILL_0_BUFX2_insert606 gnd vdd FILL
X_12561_ _12091_/B _13175_/CLK _13199_/R vdd _12519_/Y gnd vdd DFFSR
XSFILL23880x73050 gnd vdd FILL
XSFILL23080x54050 gnd vdd FILL
XFILL_0_BUFX2_insert617 gnd vdd FILL
XFILL_0_BUFX2_insert628 gnd vdd FILL
XFILL_4__7805_ gnd vdd FILL
XFILL_0_BUFX2_insert639 gnd vdd FILL
X_14300_ _8873_/A gnd _14301_/A vdd INVX1
X_11512_ _11498_/A _11491_/B gnd _11512_/Y vdd NOR2X1
XFILL_4__8785_ gnd vdd FILL
X_15280_ _15280_/A _15280_/B gnd _15285_/A vdd NOR2X1
X_12492_ _12492_/A vdd _12491_/Y gnd _12492_/Y vdd OAI21X1
XSFILL28920x10050 gnd vdd FILL
X_14231_ _9574_/Q gnd _14231_/Y vdd INVX1
XFILL_4__7736_ gnd vdd FILL
X_11443_ _11035_/Y _11776_/A gnd _11446_/A vdd NOR2X1
XFILL_1__7958_ gnd vdd FILL
X_14162_ _8548_/Q gnd _14164_/B vdd INVX1
X_11374_ _12222_/Y _12120_/Y gnd _11374_/Y vdd AND2X2
XFILL_1__6909_ gnd vdd FILL
XFILL_2__9470_ gnd vdd FILL
XFILL_4__9406_ gnd vdd FILL
XSFILL84680x36050 gnd vdd FILL
XFILL_1__7889_ gnd vdd FILL
X_13113_ _13108_/B _12034_/Y gnd _13113_/Y vdd NAND2X1
X_10325_ _10323_/Y _10325_/B _10324_/Y gnd _10357_/D vdd OAI21X1
XFILL_4__7598_ gnd vdd FILL
X_14093_ _9117_/A _14868_/D _14037_/C _7011_/Q gnd _14095_/A vdd AOI22X1
XFILL_4_BUFX2_insert550 gnd vdd FILL
XFILL_1__9628_ gnd vdd FILL
XFILL_4_BUFX2_insert561 gnd vdd FILL
XFILL_4__10580_ gnd vdd FILL
XFILL_4_BUFX2_insert572 gnd vdd FILL
XFILL_5__8130_ gnd vdd FILL
XFILL_4_BUFX2_insert583 gnd vdd FILL
XFILL_4__9337_ gnd vdd FILL
X_13044_ _6901_/A gnd _13044_/Y vdd INVX1
X_10256_ _10254_/Y _10304_/B _10256_/C gnd _10256_/Y vdd OAI21X1
XFILL_4_BUFX2_insert594 gnd vdd FILL
XFILL_2__8352_ gnd vdd FILL
XFILL_5__11870_ gnd vdd FILL
XFILL_2__11690_ gnd vdd FILL
XFILL_5__8061_ gnd vdd FILL
XFILL_4__9268_ gnd vdd FILL
XSFILL99320x60050 gnd vdd FILL
XFILL_5__10821_ gnd vdd FILL
XFILL_2__7303_ gnd vdd FILL
X_10187_ _10166_/A _7243_/B gnd _10188_/C vdd NAND2X1
XFILL_4__12250_ gnd vdd FILL
XFILL_2__10641_ gnd vdd FILL
XFILL_1__12070_ gnd vdd FILL
XFILL_4__8219_ gnd vdd FILL
XFILL_3__12980_ gnd vdd FILL
XFILL_0__11820_ gnd vdd FILL
XFILL_5__13540_ gnd vdd FILL
XFILL_4__11201_ gnd vdd FILL
XFILL_5__10752_ gnd vdd FILL
XFILL_4__12181_ gnd vdd FILL
XFILL_2__7234_ gnd vdd FILL
XFILL_2__13360_ gnd vdd FILL
X_14995_ _12813_/Q gnd _15220_/B vdd INVX2
XFILL_3__11931_ gnd vdd FILL
XSFILL63960x6050 gnd vdd FILL
XFILL112280x20050 gnd vdd FILL
XFILL_1__11021_ gnd vdd FILL
XFILL_2__10572_ gnd vdd FILL
XSFILL64040x46050 gnd vdd FILL
XFILL_0__11751_ gnd vdd FILL
XFILL_6__14830_ gnd vdd FILL
XFILL_4__11132_ gnd vdd FILL
XFILL_5__13471_ gnd vdd FILL
XFILL_2__12311_ gnd vdd FILL
X_13946_ _9952_/Q gnd _13948_/D vdd INVX1
XFILL_5__10683_ gnd vdd FILL
XFILL_3__14650_ gnd vdd FILL
XFILL_2__7165_ gnd vdd FILL
XFILL_2__13291_ gnd vdd FILL
XFILL_0__10702_ gnd vdd FILL
XFILL112280x5050 gnd vdd FILL
XFILL_3__11862_ gnd vdd FILL
XFILL_0__14470_ gnd vdd FILL
XFILL_5__15210_ gnd vdd FILL
XFILL_5__12422_ gnd vdd FILL
XFILL_5__8963_ gnd vdd FILL
XFILL_0__11682_ gnd vdd FILL
XFILL_3__13601_ gnd vdd FILL
XFILL_6__11973_ gnd vdd FILL
XFILL_5__16190_ gnd vdd FILL
XFILL_2__15030_ gnd vdd FILL
XFILL_4__15940_ gnd vdd FILL
XFILL_4__11063_ gnd vdd FILL
XFILL_3__10813_ gnd vdd FILL
X_13877_ _10590_/Q gnd _13877_/Y vdd INVX1
XFILL_2__12242_ gnd vdd FILL
XFILL_3__14581_ gnd vdd FILL
XFILL_0__13421_ gnd vdd FILL
XFILL_2__7096_ gnd vdd FILL
XFILL_1__15760_ gnd vdd FILL
XFILL_3__11793_ gnd vdd FILL
XFILL_1__12972_ gnd vdd FILL
XFILL_0__10633_ gnd vdd FILL
XSFILL3480x53050 gnd vdd FILL
X_15616_ _7268_/Q _15177_/B _15969_/C _7780_/Q gnd _15616_/Y vdd AOI22X1
XFILL_4__10014_ gnd vdd FILL
XFILL_5__15141_ gnd vdd FILL
XFILL_5__8894_ gnd vdd FILL
XFILL_5__12353_ gnd vdd FILL
XFILL_3__16320_ gnd vdd FILL
XFILL_6__14692_ gnd vdd FILL
XFILL_1_BUFX2_insert440 gnd vdd FILL
X_12828_ _12826_/Y vdd _12827_/Y gnd _12920_/D vdd OAI21X1
XFILL_1_BUFX2_insert451 gnd vdd FILL
XFILL_3__10744_ gnd vdd FILL
XFILL_1__14711_ gnd vdd FILL
XFILL_3__13532_ gnd vdd FILL
XFILL_4__15871_ gnd vdd FILL
XFILL_1_BUFX2_insert462 gnd vdd FILL
XFILL_1__11923_ gnd vdd FILL
XFILL_2__12173_ gnd vdd FILL
XFILL_0__16140_ gnd vdd FILL
XFILL_0__13352_ gnd vdd FILL
XFILL_1__15691_ gnd vdd FILL
XFILL_1_BUFX2_insert473 gnd vdd FILL
XFILL_5__7845_ gnd vdd FILL
XFILL_6__13643_ gnd vdd FILL
XSFILL84200x59050 gnd vdd FILL
XFILL_0__10564_ gnd vdd FILL
XFILL_1_BUFX2_insert484 gnd vdd FILL
XFILL_5__11304_ gnd vdd FILL
XFILL_4__14822_ gnd vdd FILL
X_15547_ _15547_/A _15175_/B _16212_/A _8602_/A gnd _15548_/B vdd AOI22X1
XFILL_5__15072_ gnd vdd FILL
X_12759_ _12721_/B memoryOutData[21] gnd _12760_/C vdd NAND2X1
XFILL_5__12284_ gnd vdd FILL
XFILL_2__11124_ gnd vdd FILL
XFILL_1_BUFX2_insert495 gnd vdd FILL
XFILL_3__16251_ gnd vdd FILL
XFILL_1__14642_ gnd vdd FILL
XFILL_3__6860_ gnd vdd FILL
XFILL_3__13463_ gnd vdd FILL
XFILL_0__12303_ gnd vdd FILL
XFILL_3__10675_ gnd vdd FILL
XFILL_0__16071_ gnd vdd FILL
XFILL_1__11854_ gnd vdd FILL
XFILL_0__13283_ gnd vdd FILL
XFILL_0__10495_ gnd vdd FILL
XFILL_5__14023_ gnd vdd FILL
XFILL_3__15202_ gnd vdd FILL
XSFILL59800x54050 gnd vdd FILL
XFILL_5__11235_ gnd vdd FILL
XFILL_2__9806_ gnd vdd FILL
XFILL_3__12414_ gnd vdd FILL
XFILL_0__9870_ gnd vdd FILL
XFILL_6__10786_ gnd vdd FILL
XFILL_4__14753_ gnd vdd FILL
X_15478_ _10848_/Q gnd _15479_/A vdd INVX1
XFILL_1__10805_ gnd vdd FILL
XFILL_3__16182_ gnd vdd FILL
XFILL_4__11965_ gnd vdd FILL
XFILL_2__15932_ gnd vdd FILL
XFILL_0__15022_ gnd vdd FILL
XFILL_3__13394_ gnd vdd FILL
XBUFX2_insert1008 _10928_/Y gnd _12312_/A vdd BUFX2
XFILL_2__11055_ gnd vdd FILL
XFILL_1__14573_ gnd vdd FILL
XSFILL99400x40050 gnd vdd FILL
XFILL_0__12234_ gnd vdd FILL
XBUFX2_insert1019 _13340_/Y gnd _9597_/A vdd BUFX2
XFILL_5__9515_ gnd vdd FILL
XFILL_2__7998_ gnd vdd FILL
XFILL_6__12525_ gnd vdd FILL
XFILL_1__11785_ gnd vdd FILL
XFILL_6__16293_ gnd vdd FILL
XFILL_4__13704_ gnd vdd FILL
X_14429_ _14721_/A _15884_/B _14545_/B _15879_/D gnd _14429_/Y vdd OAI22X1
XFILL_4__10916_ gnd vdd FILL
X_7360_ _7358_/Y _7297_/B _7360_/C gnd _7360_/Y vdd OAI21X1
XFILL_3__12345_ gnd vdd FILL
XFILL_1__16312_ gnd vdd FILL
XFILL_2__10006_ gnd vdd FILL
XFILL_3__15133_ gnd vdd FILL
XFILL_5__11166_ gnd vdd FILL
XFILL_2__9737_ gnd vdd FILL
XFILL_4__14684_ gnd vdd FILL
XFILL_1__13524_ gnd vdd FILL
XFILL_3__8530_ gnd vdd FILL
XFILL_4__11896_ gnd vdd FILL
XFILL_2__6949_ gnd vdd FILL
XFILL_2__15863_ gnd vdd FILL
XFILL_0__12165_ gnd vdd FILL
XSFILL23720x9050 gnd vdd FILL
XFILL_5__10117_ gnd vdd FILL
XFILL_0__8752_ gnd vdd FILL
XFILL_4__13635_ gnd vdd FILL
XSFILL64120x26050 gnd vdd FILL
XFILL_5__15974_ gnd vdd FILL
XFILL_1__16243_ gnd vdd FILL
XFILL_3__8461_ gnd vdd FILL
XFILL_2__14814_ gnd vdd FILL
XFILL_3__15064_ gnd vdd FILL
XFILL_3__12276_ gnd vdd FILL
XFILL_5__11097_ gnd vdd FILL
X_7291_ _7289_/Y _7369_/B _7290_/Y gnd _7383_/D vdd OAI21X1
XFILL_1__13455_ gnd vdd FILL
XFILL_2__9668_ gnd vdd FILL
XFILL_0__11116_ gnd vdd FILL
XSFILL74280x70050 gnd vdd FILL
XFILL_0__7703_ gnd vdd FILL
XFILL_0__12096_ gnd vdd FILL
XFILL_2__15794_ gnd vdd FILL
XFILL_1__10667_ gnd vdd FILL
XFILL_5__9377_ gnd vdd FILL
X_9030_ _9030_/A _9017_/A _9030_/C gnd _9072_/D vdd OAI21X1
XFILL_5__10048_ gnd vdd FILL
XFILL_6__12387_ gnd vdd FILL
XFILL_3__14015_ gnd vdd FILL
XFILL_4__16354_ gnd vdd FILL
XFILL_5__14925_ gnd vdd FILL
XFILL_3__11227_ gnd vdd FILL
XFILL_1__12406_ gnd vdd FILL
XFILL_4__13566_ gnd vdd FILL
XFILL_2__8619_ gnd vdd FILL
XFILL_0__15924_ gnd vdd FILL
XFILL_1__16174_ gnd vdd FILL
XFILL_2__11957_ gnd vdd FILL
XFILL_4__10778_ gnd vdd FILL
XFILL_0__11047_ gnd vdd FILL
XFILL_3__8392_ gnd vdd FILL
XFILL_2__14745_ gnd vdd FILL
XFILL_2__9599_ gnd vdd FILL
XFILL_5__8328_ gnd vdd FILL
XFILL_1__13386_ gnd vdd FILL
XFILL_4__15305_ gnd vdd FILL
XSFILL114920x14050 gnd vdd FILL
XFILL_0__7634_ gnd vdd FILL
XFILL_6__11338_ gnd vdd FILL
XSFILL53960x69050 gnd vdd FILL
XFILL_5__14856_ gnd vdd FILL
XFILL_4__12517_ gnd vdd FILL
XFILL_2__10908_ gnd vdd FILL
XFILL_4__16285_ gnd vdd FILL
XSFILL3560x33050 gnd vdd FILL
XFILL_3__7343_ gnd vdd FILL
XFILL_3__11158_ gnd vdd FILL
XFILL_1__15125_ gnd vdd FILL
XFILL_4__13497_ gnd vdd FILL
XFILL_1__12337_ gnd vdd FILL
XFILL_2__11888_ gnd vdd FILL
XFILL_0__15855_ gnd vdd FILL
XFILL_2__14676_ gnd vdd FILL
XFILL_5__13807_ gnd vdd FILL
XFILL_5__8259_ gnd vdd FILL
XFILL_0__7565_ gnd vdd FILL
XFILL_4__15236_ gnd vdd FILL
XFILL_3__10109_ gnd vdd FILL
XFILL_4__12448_ gnd vdd FILL
XFILL_2__16415_ gnd vdd FILL
XFILL_5__14787_ gnd vdd FILL
XFILL_2__13627_ gnd vdd FILL
XFILL_0__14806_ gnd vdd FILL
XFILL_5__11999_ gnd vdd FILL
XFILL_1__15056_ gnd vdd FILL
XFILL_3__15966_ gnd vdd FILL
XFILL_3__11089_ gnd vdd FILL
XFILL_1__12268_ gnd vdd FILL
XFILL_0__15786_ gnd vdd FILL
XSFILL94440x83050 gnd vdd FILL
XFILL_0__12998_ gnd vdd FILL
X_9932_ _9932_/A _9865_/A _9932_/C gnd _9970_/D vdd OAI21X1
XFILL_5__13738_ gnd vdd FILL
XFILL_3__9013_ gnd vdd FILL
XFILL_1__14007_ gnd vdd FILL
XFILL_0__7496_ gnd vdd FILL
XFILL_4__15167_ gnd vdd FILL
XFILL_3__14917_ gnd vdd FILL
XFILL_2__16346_ gnd vdd FILL
XFILL_4__12379_ gnd vdd FILL
XFILL_2__13558_ gnd vdd FILL
XFILL_1__11219_ gnd vdd FILL
XFILL_3__15897_ gnd vdd FILL
XFILL_0__14737_ gnd vdd FILL
XFILL_0__11949_ gnd vdd FILL
XFILL_1__12199_ gnd vdd FILL
XFILL_0__9235_ gnd vdd FILL
XSFILL3560x2050 gnd vdd FILL
XFILL_4__14118_ gnd vdd FILL
XFILL_5__13669_ gnd vdd FILL
XFILL_2__12509_ gnd vdd FILL
XSFILL33880x36050 gnd vdd FILL
X_9863_ _9863_/A _9902_/B _9862_/Y gnd _9947_/D vdd OAI21X1
XFILL_3__14848_ gnd vdd FILL
XFILL_4__15098_ gnd vdd FILL
XFILL_2__13489_ gnd vdd FILL
XFILL_2__16277_ gnd vdd FILL
XFILL_5__15408_ gnd vdd FILL
XFILL_0__14668_ gnd vdd FILL
XFILL111800x14050 gnd vdd FILL
X_8814_ _8814_/Q _7790_/CLK _9566_/R vdd _8768_/Y gnd vdd DFFSR
XFILL_0__9166_ gnd vdd FILL
XFILL_5__16388_ gnd vdd FILL
XFILL_4__14049_ gnd vdd FILL
XFILL_2__15228_ gnd vdd FILL
XSFILL48920x58050 gnd vdd FILL
XFILL_0__16407_ gnd vdd FILL
X_9794_ _9798_/B _9794_/B gnd _9795_/C vdd NAND2X1
XFILL_0__13619_ gnd vdd FILL
XFILL_3__14779_ gnd vdd FILL
XFILL_0__8117_ gnd vdd FILL
XFILL_1__15958_ gnd vdd FILL
XFILL_0__14599_ gnd vdd FILL
XFILL_5__15339_ gnd vdd FILL
XFILL_6__7885_ gnd vdd FILL
XFILL_6_BUFX2_insert623 gnd vdd FILL
XFILL_0__9097_ gnd vdd FILL
X_8745_ _8745_/A gnd _8745_/Y vdd INVX1
XFILL_3__9915_ gnd vdd FILL
XFILL_2__15159_ gnd vdd FILL
XFILL_0__16338_ gnd vdd FILL
XFILL_1__14909_ gnd vdd FILL
XSFILL49000x67050 gnd vdd FILL
XSFILL44600x3050 gnd vdd FILL
XFILL_1__15889_ gnd vdd FILL
XFILL_3__16449_ gnd vdd FILL
X_8676_ _8608_/A _7642_/CLK _8676_/R vdd _8676_/D gnd vdd DFFSR
XFILL_6_BUFX2_insert689 gnd vdd FILL
XSFILL89400x72050 gnd vdd FILL
XFILL_3__9846_ gnd vdd FILL
XSFILL3640x13050 gnd vdd FILL
XFILL_0__16269_ gnd vdd FILL
XSFILL109560x78050 gnd vdd FILL
X_7627_ _7562_/B _9803_/B gnd _7627_/Y vdd NAND2X1
XFILL_1__8861_ gnd vdd FILL
XFILL_3__9777_ gnd vdd FILL
XFILL_4__8570_ gnd vdd FILL
XFILL_3__6989_ gnd vdd FILL
XFILL_1__7812_ gnd vdd FILL
XSFILL54120x58050 gnd vdd FILL
XFILL_1_CLKBUF1_insert116 gnd vdd FILL
X_7558_ _7598_/B _7558_/B gnd _7558_/Y vdd NAND2X1
XFILL_3__8728_ gnd vdd FILL
XFILL_1_CLKBUF1_insert127 gnd vdd FILL
XFILL_0__9999_ gnd vdd FILL
XFILL_1_CLKBUF1_insert138 gnd vdd FILL
XFILL_1__7743_ gnd vdd FILL
XFILL_1_CLKBUF1_insert149 gnd vdd FILL
X_7489_ _7535_/Q gnd _7489_/Y vdd INVX1
XFILL_4__7452_ gnd vdd FILL
XFILL_3__8659_ gnd vdd FILL
XSFILL33960x16050 gnd vdd FILL
X_9228_ _9228_/A _7180_/B gnd _9229_/C vdd NAND2X1
XFILL_1__7674_ gnd vdd FILL
X_10110_ _10108_/Y _10106_/A _10110_/C gnd _10110_/Y vdd OAI21X1
XSFILL18760x77050 gnd vdd FILL
XFILL_1__9413_ gnd vdd FILL
X_11090_ _11089_/Y _11062_/Y _11090_/C gnd _11663_/C vdd AOI21X1
XFILL_3_BUFX2_insert502 gnd vdd FILL
X_9159_ _9159_/A gnd _9161_/A vdd INVX1
XFILL_3_BUFX2_insert513 gnd vdd FILL
XFILL_4__9122_ gnd vdd FILL
XFILL_3_BUFX2_insert524 gnd vdd FILL
XFILL_3_BUFX2_insert535 gnd vdd FILL
X_10041_ _10024_/B _9785_/B gnd _10041_/Y vdd NAND2X1
XSFILL33800x80050 gnd vdd FILL
XFILL_3_BUFX2_insert546 gnd vdd FILL
XFILL_1__9344_ gnd vdd FILL
XFILL_3_BUFX2_insert557 gnd vdd FILL
XFILL_3_BUFX2_insert568 gnd vdd FILL
XSFILL48600x40050 gnd vdd FILL
XFILL_3_BUFX2_insert579 gnd vdd FILL
XFILL_1__9275_ gnd vdd FILL
XSFILL23880x68050 gnd vdd FILL
XFILL_4__8004_ gnd vdd FILL
X_13800_ _13799_/Y _14865_/B gnd _13800_/Y vdd NOR2X1
XFILL_1__8226_ gnd vdd FILL
X_11992_ _11988_/B gnd _12096_/C gnd _11994_/B vdd NAND3X1
X_14780_ _7623_/A gnd _16127_/D vdd INVX1
X_10943_ _10957_/B _10943_/B _10943_/C gnd _10945_/B vdd NAND3X1
X_13731_ _9179_/Q gnd _13733_/D vdd INVX1
X_16450_ _16450_/A _16450_/B _16450_/C gnd _16451_/C vdd AOI21X1
XFILL_1__7108_ gnd vdd FILL
X_13662_ _13661_/Y _13662_/B gnd _13663_/A vdd NOR2X1
X_10874_ _10871_/Y _10874_/B gnd _10887_/A vdd NOR2X1
XFILL_1__8088_ gnd vdd FILL
XFILL_2__8970_ gnd vdd FILL
XFILL_4__8906_ gnd vdd FILL
X_15401_ _13842_/Y _15681_/B _15681_/C _15401_/D gnd _15405_/B vdd OAI22X1
X_12613_ vdd memoryOutData[15] gnd _12613_/Y vdd NAND2X1
XFILL_4__9886_ gnd vdd FILL
XFILL_1__7039_ gnd vdd FILL
X_13593_ _13377_/Y _13418_/A gnd _14344_/B vdd AND2X2
X_16381_ _14418_/A gnd _16381_/Y vdd INVX1
XFILL_0_BUFX2_insert403 gnd vdd FILL
XFILL_0_BUFX2_insert414 gnd vdd FILL
XFILL_5__7630_ gnd vdd FILL
XSFILL18840x57050 gnd vdd FILL
XFILL_0_BUFX2_insert425 gnd vdd FILL
XFILL_4__8837_ gnd vdd FILL
X_15332_ _8668_/Q gnd _15334_/C vdd INVX1
X_12544_ _12023_/B _9060_/CLK _9060_/R vdd _12468_/Y gnd vdd DFFSR
XSFILL84280x33050 gnd vdd FILL
XFILL_0_BUFX2_insert436 gnd vdd FILL
XFILL_0_BUFX2_insert447 gnd vdd FILL
XFILL_0_BUFX2_insert458 gnd vdd FILL
XFILL_2__7852_ gnd vdd FILL
XFILL_0__10280_ gnd vdd FILL
XFILL_0_BUFX2_insert469 gnd vdd FILL
XFILL_4__8768_ gnd vdd FILL
XFILL_5__7561_ gnd vdd FILL
XFILL_5__11020_ gnd vdd FILL
XSFILL99320x55050 gnd vdd FILL
X_12475_ _12035_/B gnd _12477_/A vdd INVX1
X_15263_ _13733_/A _15565_/B _15801_/A _13691_/Y gnd _15264_/A vdd OAI22X1
XFILL_4__11750_ gnd vdd FILL
XFILL_3__10391_ gnd vdd FILL
XFILL_5__9300_ gnd vdd FILL
XFILL_4__7719_ gnd vdd FILL
XFILL_6__12310_ gnd vdd FILL
XFILL_1__11570_ gnd vdd FILL
X_14214_ _10659_/A _14868_/A _14214_/C _10019_/A gnd _14215_/B vdd AOI22X1
X_11426_ _12218_/Y _12117_/Y gnd _11427_/A vdd AND2X2
XFILL_6__13290_ gnd vdd FILL
XFILL_4__10701_ gnd vdd FILL
X_15194_ _15683_/C _13586_/Y _13612_/Y _15410_/D gnd _15195_/A vdd OAI22X1
XSFILL23960x48050 gnd vdd FILL
XFILL_5__7492_ gnd vdd FILL
XFILL_3__12130_ gnd vdd FILL
XFILL_4__8699_ gnd vdd FILL
XFILL_2__9522_ gnd vdd FILL
XFILL_1__10521_ gnd vdd FILL
XFILL_2__12860_ gnd vdd FILL
XSFILL63560x34050 gnd vdd FILL
XFILL_4__11681_ gnd vdd FILL
XFILL112280x15050 gnd vdd FILL
XFILL_5__9231_ gnd vdd FILL
X_14145_ _13865_/C _7780_/Q _7584_/A _14145_/D gnd _14145_/Y vdd AOI22X1
XFILL_4__13420_ gnd vdd FILL
X_11357_ _11203_/Y gnd _11358_/A vdd INVX1
XFILL_4__10632_ gnd vdd FILL
XFILL_3__12061_ gnd vdd FILL
XFILL_5__12971_ gnd vdd FILL
XFILL_2__11811_ gnd vdd FILL
XFILL_1__13240_ gnd vdd FILL
XSFILL109320x40050 gnd vdd FILL
XFILL_1__10452_ gnd vdd FILL
XFILL_5__9162_ gnd vdd FILL
X_10308_ _14703_/A gnd _10308_/Y vdd INVX1
XFILL_5__14710_ gnd vdd FILL
XFILL_0__13970_ gnd vdd FILL
XFILL_5__11922_ gnd vdd FILL
XFILL_6__12172_ gnd vdd FILL
XFILL_4_BUFX2_insert380 gnd vdd FILL
X_14076_ _8349_/A _14414_/B _13864_/B _8675_/Q gnd _14085_/A vdd AOI22X1
XFILL_3__11012_ gnd vdd FILL
XCLKBUF1_insert115 CLKBUF1_insert150/A gnd _9834_/CLK vdd CLKBUF1
XFILL_4__13351_ gnd vdd FILL
XFILL_5__15690_ gnd vdd FILL
XCLKBUF1_insert126 CLKBUF1_insert187/A gnd _12669_/CLK vdd CLKBUF1
XFILL_4_BUFX2_insert391 gnd vdd FILL
XFILL_2__8404_ gnd vdd FILL
X_11288_ _11448_/A _11653_/A _11288_/C gnd _11289_/C vdd AOI21X1
XFILL_2__14530_ gnd vdd FILL
XCLKBUF1_insert137 CLKBUF1_insert182/A gnd _9716_/CLK vdd CLKBUF1
XFILL_2__11742_ gnd vdd FILL
XFILL_4__10563_ gnd vdd FILL
XSFILL79240x22050 gnd vdd FILL
XFILL_2__9384_ gnd vdd FILL
XFILL_1__13171_ gnd vdd FILL
XFILL_5__8113_ gnd vdd FILL
XCLKBUF1_insert148 CLKBUF1_insert182/A gnd _8815_/CLK vdd CLKBUF1
XFILL_1__10383_ gnd vdd FILL
X_13027_ vdd _13027_/B gnd _13028_/C vdd NAND2X1
XCLKBUF1_insert159 CLKBUF1_insert193/A gnd _8152_/CLK vdd CLKBUF1
XFILL_5__14641_ gnd vdd FILL
X_10239_ _10239_/A gnd _10239_/Y vdd INVX1
XFILL_4__12302_ gnd vdd FILL
XFILL_5__9093_ gnd vdd FILL
XFILL_3__15820_ gnd vdd FILL
XFILL_4__16070_ gnd vdd FILL
XFILL_5__11853_ gnd vdd FILL
XFILL_4__13282_ gnd vdd FILL
XFILL_2__8335_ gnd vdd FILL
XFILL_2__14461_ gnd vdd FILL
XFILL_4__10494_ gnd vdd FILL
XFILL_1__12122_ gnd vdd FILL
XFILL_0__15640_ gnd vdd FILL
XFILL_2__11673_ gnd vdd FILL
XSFILL114440x31050 gnd vdd FILL
XFILL_0__12852_ gnd vdd FILL
XFILL_0__7350_ gnd vdd FILL
XFILL_4__15021_ gnd vdd FILL
XFILL_5__10804_ gnd vdd FILL
XFILL_5__14572_ gnd vdd FILL
XFILL_2__16200_ gnd vdd FILL
XFILL_2__13412_ gnd vdd FILL
XFILL_4__12233_ gnd vdd FILL
XFILL_2__10624_ gnd vdd FILL
XFILL_2__8266_ gnd vdd FILL
XFILL_3__15751_ gnd vdd FILL
XFILL_5__11784_ gnd vdd FILL
XFILL_3__12963_ gnd vdd FILL
XFILL_1__12053_ gnd vdd FILL
XFILL_2__14392_ gnd vdd FILL
XSFILL84360x13050 gnd vdd FILL
XFILL_0__11803_ gnd vdd FILL
XFILL_0__15571_ gnd vdd FILL
XFILL_5__16311_ gnd vdd FILL
XFILL_6__10005_ gnd vdd FILL
XFILL_0__12783_ gnd vdd FILL
XFILL_5__13523_ gnd vdd FILL
XFILL_2__7217_ gnd vdd FILL
XFILL_3__14702_ gnd vdd FILL
XFILL_2__13343_ gnd vdd FILL
XFILL_3__11914_ gnd vdd FILL
XFILL_4__12164_ gnd vdd FILL
X_14978_ _14978_/A _14978_/B _15812_/C gnd _13045_/B vdd AOI21X1
XFILL_2__16131_ gnd vdd FILL
XFILL_1__11004_ gnd vdd FILL
XFILL_3__15682_ gnd vdd FILL
XFILL_2__10555_ gnd vdd FILL
XFILL_0__14522_ gnd vdd FILL
XFILL_2__8197_ gnd vdd FILL
XFILL_0__9020_ gnd vdd FILL
XSFILL69160x74050 gnd vdd FILL
XFILL_3__12894_ gnd vdd FILL
XSFILL99400x35050 gnd vdd FILL
XFILL_0__11734_ gnd vdd FILL
XFILL_5__16242_ gnd vdd FILL
XFILL_5__9995_ gnd vdd FILL
XFILL_5__13454_ gnd vdd FILL
X_13929_ _13929_/A _13929_/B gnd _13930_/A vdd NOR2X1
XFILL_4__11115_ gnd vdd FILL
XFILL_3__14633_ gnd vdd FILL
X_6860_ _6860_/A gnd memoryAddress[22] vdd BUFX2
XFILL_4__12095_ gnd vdd FILL
XFILL_5__10666_ gnd vdd FILL
XFILL_2__16062_ gnd vdd FILL
XFILL_2__13274_ gnd vdd FILL
XFILL_1__15812_ gnd vdd FILL
XFILL_3__11845_ gnd vdd FILL
XFILL_0__14453_ gnd vdd FILL
XFILL_2__10486_ gnd vdd FILL
XFILL_5__12405_ gnd vdd FILL
XFILL_0__11665_ gnd vdd FILL
XFILL_4__15923_ gnd vdd FILL
XFILL_5__16173_ gnd vdd FILL
XFILL_2__15013_ gnd vdd FILL
XFILL_4__11046_ gnd vdd FILL
XFILL_5__13385_ gnd vdd FILL
XFILL_2__12225_ gnd vdd FILL
XFILL_3__14564_ gnd vdd FILL
XFILL_2__7079_ gnd vdd FILL
XFILL_0__13404_ gnd vdd FILL
XFILL_3__7961_ gnd vdd FILL
XFILL_0__10616_ gnd vdd FILL
XFILL_1__12955_ gnd vdd FILL
XFILL_3__11776_ gnd vdd FILL
XFILL_1__15743_ gnd vdd FILL
XSFILL23640x30050 gnd vdd FILL
XFILL_0__14384_ gnd vdd FILL
XFILL_5__15124_ gnd vdd FILL
XFILL_1_BUFX2_insert270 gnd vdd FILL
XSFILL74280x65050 gnd vdd FILL
XFILL_3__16303_ gnd vdd FILL
XFILL_5__8877_ gnd vdd FILL
XFILL_5__12336_ gnd vdd FILL
XFILL_0__11596_ gnd vdd FILL
X_8530_ _8528_/Y _8496_/A _8530_/C gnd _8564_/D vdd OAI21X1
XFILL_4__15854_ gnd vdd FILL
XFILL_1_BUFX2_insert281 gnd vdd FILL
XFILL_3__13515_ gnd vdd FILL
XSFILL109400x20050 gnd vdd FILL
XFILL_3__6912_ gnd vdd FILL
XFILL_1_BUFX2_insert292 gnd vdd FILL
XFILL_1__11906_ gnd vdd FILL
XFILL_0__16123_ gnd vdd FILL
XFILL_2__12156_ gnd vdd FILL
XFILL_0__13335_ gnd vdd FILL
XFILL_3__14495_ gnd vdd FILL
XFILL_1__15674_ gnd vdd FILL
XFILL_1__12886_ gnd vdd FILL
XFILL_5__7828_ gnd vdd FILL
XFILL_0__10547_ gnd vdd FILL
XFILL_3__7892_ gnd vdd FILL
XFILL_4__14805_ gnd vdd FILL
XFILL_5_BUFX2_insert608 gnd vdd FILL
XFILL_5__15055_ gnd vdd FILL
XSFILL49080x41050 gnd vdd FILL
XFILL_0__9922_ gnd vdd FILL
XFILL_3__16234_ gnd vdd FILL
X_8461_ _8461_/A _8460_/A _8461_/C gnd _8461_/Y vdd OAI21X1
XFILL_5_BUFX2_insert619 gnd vdd FILL
XFILL_5__12267_ gnd vdd FILL
XFILL_2__11107_ gnd vdd FILL
XFILL_1__14625_ gnd vdd FILL
XFILL_3__10658_ gnd vdd FILL
XFILL_3__13446_ gnd vdd FILL
XFILL_4__15785_ gnd vdd FILL
XSFILL3560x28050 gnd vdd FILL
XFILL_3__9631_ gnd vdd FILL
XFILL_4__12997_ gnd vdd FILL
XFILL_2__12087_ gnd vdd FILL
XFILL_3__6843_ gnd vdd FILL
XFILL_0__16054_ gnd vdd FILL
XFILL_1__11837_ gnd vdd FILL
XFILL_0__13266_ gnd vdd FILL
XFILL_5__14006_ gnd vdd FILL
XFILL_5__7759_ gnd vdd FILL
XFILL_6__16345_ gnd vdd FILL
XFILL_0_BUFX2_insert970 gnd vdd FILL
X_7412_ _7376_/A _8180_/CLK _7391_/R vdd _7412_/D gnd vdd DFFSR
XFILL_5__11218_ gnd vdd FILL
XFILL_4__14736_ gnd vdd FILL
XFILL_0_BUFX2_insert981 gnd vdd FILL
XFILL_0__9853_ gnd vdd FILL
XFILL_2__15915_ gnd vdd FILL
XFILL_3__16165_ gnd vdd FILL
XFILL_4__11948_ gnd vdd FILL
XFILL_0__15005_ gnd vdd FILL
XFILL_5__12198_ gnd vdd FILL
XSFILL114520x11050 gnd vdd FILL
X_8392_ _8365_/A _8008_/B gnd _8393_/C vdd NAND2X1
XFILL_2__11038_ gnd vdd FILL
XFILL_0_BUFX2_insert992 gnd vdd FILL
XFILL_1__14556_ gnd vdd FILL
XFILL_3__13377_ gnd vdd FILL
XFILL_0__12217_ gnd vdd FILL
XFILL_1__11768_ gnd vdd FILL
X_7343_ _7401_/Q gnd _7345_/A vdd INVX1
XFILL_5__11149_ gnd vdd FILL
XFILL_3__15116_ gnd vdd FILL
XFILL_0__6996_ gnd vdd FILL
XFILL_0__9784_ gnd vdd FILL
XFILL_3__12328_ gnd vdd FILL
XFILL_3__8513_ gnd vdd FILL
XFILL_4__14667_ gnd vdd FILL
XFILL_1__13507_ gnd vdd FILL
XFILL_4__11879_ gnd vdd FILL
XFILL_3__16096_ gnd vdd FILL
XFILL_2__15846_ gnd vdd FILL
XFILL_1__14487_ gnd vdd FILL
XFILL_5__9429_ gnd vdd FILL
XFILL_0__12148_ gnd vdd FILL
XFILL_3__9493_ gnd vdd FILL
XFILL_4__16406_ gnd vdd FILL
XFILL_1__11699_ gnd vdd FILL
XFILL_4__13618_ gnd vdd FILL
XFILL_0__8735_ gnd vdd FILL
XFILL_1__16226_ gnd vdd FILL
XSFILL69240x54050 gnd vdd FILL
XFILL_5__15957_ gnd vdd FILL
XFILL_3__15047_ gnd vdd FILL
X_7274_ _7274_/Q _7274_/CLK _7274_/R vdd _7274_/D gnd vdd DFFSR
XFILL_4__14598_ gnd vdd FILL
XFILL_3__12259_ gnd vdd FILL
XFILL_3__8444_ gnd vdd FILL
XFILL_1__13438_ gnd vdd FILL
XFILL_2__15777_ gnd vdd FILL
X_9013_ _9067_/Q gnd _9015_/A vdd INVX1
XFILL_0__12079_ gnd vdd FILL
XFILL_2__12989_ gnd vdd FILL
XFILL_4__16337_ gnd vdd FILL
XFILL_6__15158_ gnd vdd FILL
XFILL_5__14908_ gnd vdd FILL
XFILL_4__13549_ gnd vdd FILL
XFILL_2__14728_ gnd vdd FILL
XFILL_1__16157_ gnd vdd FILL
XFILL_5__15888_ gnd vdd FILL
XFILL_3__8375_ gnd vdd FILL
XFILL_0__15907_ gnd vdd FILL
XFILL_1__13369_ gnd vdd FILL
XSFILL104440x63050 gnd vdd FILL
XFILL_6__14109_ gnd vdd FILL
XFILL_0__7617_ gnd vdd FILL
XFILL_5__14839_ gnd vdd FILL
XFILL_0__8597_ gnd vdd FILL
XFILL_4__16268_ gnd vdd FILL
XFILL_1__15108_ gnd vdd FILL
XSFILL8680x61050 gnd vdd FILL
XSFILL79240x9050 gnd vdd FILL
XSFILL23720x10050 gnd vdd FILL
XFILL_3__7326_ gnd vdd FILL
XFILL_1__16088_ gnd vdd FILL
XFILL_0__15838_ gnd vdd FILL
XFILL_2__14659_ gnd vdd FILL
XSFILL89960x24050 gnd vdd FILL
XFILL_4__15219_ gnd vdd FILL
XFILL_0__7548_ gnd vdd FILL
XFILL_2_BUFX2_insert509 gnd vdd FILL
XFILL_4__16199_ gnd vdd FILL
XFILL_1__15039_ gnd vdd FILL
XFILL_3__15949_ gnd vdd FILL
XSFILL89400x67050 gnd vdd FILL
XFILL_0__15769_ gnd vdd FILL
X_9915_ _9965_/Q gnd _9915_/Y vdd INVX1
XFILL_0__7479_ gnd vdd FILL
XFILL_2__16329_ gnd vdd FILL
XFILL_3__7188_ gnd vdd FILL
XFILL_1__8011_ gnd vdd FILL
XSFILL94440x3050 gnd vdd FILL
XFILL_0__9218_ gnd vdd FILL
X_9846_ _9942_/Q gnd _9848_/A vdd INVX1
XFILL_6__8986_ gnd vdd FILL
XFILL_6_BUFX2_insert1017 gnd vdd FILL
XSFILL13640x62050 gnd vdd FILL
XFILL_6__7937_ gnd vdd FILL
XFILL_0__9149_ gnd vdd FILL
X_9777_ _9775_/Y _9798_/B _9777_/C gnd _9777_/Y vdd OAI21X1
X_6989_ _7027_/Q gnd _6989_/Y vdd INVX1
XFILL_4__9740_ gnd vdd FILL
XFILL_4__6952_ gnd vdd FILL
XBUFX2_insert508 BUFX2_insert570/A gnd _12799_/R vdd BUFX2
X_8728_ _8765_/B _8472_/B gnd _8729_/C vdd NAND2X1
XBUFX2_insert519 BUFX2_insert556/A gnd _7270_/R vdd BUFX2
XFILL_6_BUFX2_insert464 gnd vdd FILL
XFILL_4__9671_ gnd vdd FILL
XFILL_6__9607_ gnd vdd FILL
XFILL_4__6883_ gnd vdd FILL
X_10590_ _10590_/Q _8025_/CLK _8025_/R vdd _10590_/D gnd vdd DFFSR
XFILL_1__8913_ gnd vdd FILL
X_8659_ _8659_/A gnd _8661_/A vdd INVX1
XFILL_1__9893_ gnd vdd FILL
XFILL_4__8622_ gnd vdd FILL
XFILL_4_BUFX2_insert1010 gnd vdd FILL
XSFILL33800x75050 gnd vdd FILL
XSFILL8760x41050 gnd vdd FILL
XFILL_4_BUFX2_insert1021 gnd vdd FILL
XFILL_1__8844_ gnd vdd FILL
XFILL_4_BUFX2_insert1032 gnd vdd FILL
XFILL_4_BUFX2_insert1043 gnd vdd FILL
XSFILL48600x35050 gnd vdd FILL
XFILL_4_BUFX2_insert1054 gnd vdd FILL
X_12260_ _12248_/A _12802_/Q _12248_/C gnd _12260_/Y vdd NAND3X1
XFILL_4_BUFX2_insert1065 gnd vdd FILL
XFILL_4_BUFX2_insert1087 gnd vdd FILL
XSFILL104360x5050 gnd vdd FILL
XFILL_4__7504_ gnd vdd FILL
XFILL_1__8775_ gnd vdd FILL
X_11211_ _11198_/Y _12334_/Y _11210_/Y gnd _11211_/Y vdd OAI21X1
XFILL_4__8484_ gnd vdd FILL
X_12191_ _12122_/A _12898_/A gnd _12192_/C vdd NAND2X1
XFILL_1__7726_ gnd vdd FILL
XFILL_4__7435_ gnd vdd FILL
X_11142_ _11142_/A _11057_/Y _11141_/Y gnd _11185_/A vdd AOI21X1
XSFILL13720x42050 gnd vdd FILL
XFILL_3_BUFX2_insert310 gnd vdd FILL
XFILL_3_BUFX2_insert321 gnd vdd FILL
XSFILL79160x37050 gnd vdd FILL
XFILL_4__7366_ gnd vdd FILL
X_15950_ _9400_/A _15945_/C _16148_/C gnd _15950_/Y vdd NAND3X1
X_11073_ _12258_/Y _12147_/Y gnd _11073_/Y vdd NOR2X1
XFILL_3_BUFX2_insert332 gnd vdd FILL
XFILL_3_BUFX2_insert343 gnd vdd FILL
XFILL_3_BUFX2_insert354 gnd vdd FILL
XFILL_1__7588_ gnd vdd FILL
XFILL_4__9105_ gnd vdd FILL
XFILL_3_BUFX2_insert365 gnd vdd FILL
XFILL_4__7297_ gnd vdd FILL
X_10024_ _10024_/A _10024_/B _10023_/Y gnd _10086_/D vdd OAI21X1
XSFILL94200x40050 gnd vdd FILL
X_14901_ _16272_/A _14901_/B _14900_/Y gnd _14901_/Y vdd OAI21X1
XFILL_2__8120_ gnd vdd FILL
XFILL_3_BUFX2_insert376 gnd vdd FILL
XFILL_3_BUFX2_insert387 gnd vdd FILL
XFILL_2_BUFX2_insert1091 gnd vdd FILL
X_15881_ _15527_/A _14444_/A _15527_/C _15881_/D gnd _15881_/Y vdd OAI22X1
XFILL_3_BUFX2_insert398 gnd vdd FILL
XFILL_4__9036_ gnd vdd FILL
X_14832_ _14832_/A _14824_/Y _14831_/Y gnd _14833_/A vdd NAND3X1
XSFILL84280x28050 gnd vdd FILL
XFILL_1__9258_ gnd vdd FILL
XFILL_5__10520_ gnd vdd FILL
XFILL_1__8209_ gnd vdd FILL
X_14763_ _14065_/C _14763_/B _7025_/Q _14926_/C gnd _14764_/B vdd AOI22X1
XSFILL43240x80050 gnd vdd FILL
X_11975_ _11975_/A _12430_/A gnd _11976_/C vdd NAND2X1
X_13714_ _13713_/Y _13698_/Y gnd _13714_/Y vdd NOR2X1
XFILL_5__9780_ gnd vdd FILL
X_10926_ _10911_/A _10898_/Y gnd _10926_/Y vdd NOR2X1
XFILL_5__10451_ gnd vdd FILL
XFILL_5__6992_ gnd vdd FILL
X_14694_ _14358_/B _16107_/A _7620_/A _14145_/D gnd _14694_/Y vdd AOI22X1
XFILL_3__11630_ gnd vdd FILL
XFILL_2__10271_ gnd vdd FILL
XFILL_4_CLKBUF1_insert111 gnd vdd FILL
XFILL_4_CLKBUF1_insert122 gnd vdd FILL
XFILL_5__8731_ gnd vdd FILL
XFILL_0__11450_ gnd vdd FILL
XFILL_4__9938_ gnd vdd FILL
X_16433_ _14262_/A _7282_/CLK _8166_/R vdd _16433_/D gnd vdd DFFSR
X_13645_ _8282_/Q _14557_/C _13645_/C _9946_/Q gnd _13648_/A vdd AOI22X1
XFILL_4_CLKBUF1_insert133 gnd vdd FILL
XFILL_5__13170_ gnd vdd FILL
XFILL_2__12010_ gnd vdd FILL
X_10857_ _14358_/A _9328_/CLK _7408_/R vdd _10857_/D gnd vdd DFFSR
XFILL_5__10382_ gnd vdd FILL
XFILL_4_CLKBUF1_insert144 gnd vdd FILL
XFILL_3__11561_ gnd vdd FILL
XFILL_1__12740_ gnd vdd FILL
XFILL_0__10401_ gnd vdd FILL
XFILL_4_CLKBUF1_insert155 gnd vdd FILL
XFILL_2__8953_ gnd vdd FILL
XFILL_4_CLKBUF1_insert166 gnd vdd FILL
XSFILL43880x5050 gnd vdd FILL
XFILL_4__9869_ gnd vdd FILL
XFILL_5__12121_ gnd vdd FILL
XFILL_4_CLKBUF1_insert177 gnd vdd FILL
XFILL_0__11381_ gnd vdd FILL
XFILL_3__13300_ gnd vdd FILL
XFILL_3__10512_ gnd vdd FILL
X_16364_ gnd gnd gnd _16365_/C vdd NAND2X1
XSFILL13800x22050 gnd vdd FILL
X_10788_ _10789_/B _8228_/B gnd _10788_/Y vdd NAND2X1
XFILL_4_CLKBUF1_insert188 gnd vdd FILL
XFILL_4__12851_ gnd vdd FILL
X_13576_ _7420_/A gnd _13576_/Y vdd INVX1
XFILL_0_BUFX2_insert233 gnd vdd FILL
XFILL_4_CLKBUF1_insert199 gnd vdd FILL
XFILL_0_BUFX2_insert244 gnd vdd FILL
XFILL_0__13120_ gnd vdd FILL
XFILL_3__11492_ gnd vdd FILL
XFILL_3__14280_ gnd vdd FILL
XFILL_5__7613_ gnd vdd FILL
XFILL_0_BUFX2_insert255 gnd vdd FILL
XFILL_2__8884_ gnd vdd FILL
X_15315_ _15314_/Y _15169_/D gnd _15318_/C vdd NOR2X1
X_12527_ vdd _12105_/A gnd _12527_/Y vdd NAND2X1
XFILL_5__12052_ gnd vdd FILL
XFILL_5__8593_ gnd vdd FILL
XFILL_4__11802_ gnd vdd FILL
XFILL_0_BUFX2_insert266 gnd vdd FILL
XFILL_3__13231_ gnd vdd FILL
XFILL_3__10443_ gnd vdd FILL
XFILL_0_BUFX2_insert277 gnd vdd FILL
XFILL_4__15570_ gnd vdd FILL
X_16295_ _16292_/Y _16294_/Y _16295_/C gnd _16295_/Y vdd NAND3X1
XFILL_1__14410_ gnd vdd FILL
XFILL_4__12782_ gnd vdd FILL
XFILL_2__7835_ gnd vdd FILL
XFILL_0_BUFX2_insert288 gnd vdd FILL
XFILL_1__11622_ gnd vdd FILL
XFILL_1__15390_ gnd vdd FILL
XFILL_0_BUFX2_insert299 gnd vdd FILL
XFILL_0__10263_ gnd vdd FILL
XFILL_2__13961_ gnd vdd FILL
XFILL_5__7544_ gnd vdd FILL
XFILL_6__16130_ gnd vdd FILL
XFILL_5__11003_ gnd vdd FILL
X_15246_ _15246_/A _15680_/B _15680_/C gnd _15257_/C vdd NAND3X1
XFILL_4__14521_ gnd vdd FILL
XFILL_0__6850_ gnd vdd FILL
XSFILL114440x26050 gnd vdd FILL
XFILL_2__15700_ gnd vdd FILL
X_12458_ vdd _12458_/B gnd _12458_/Y vdd NAND2X1
XFILL_3__13162_ gnd vdd FILL
XFILL_4__11733_ gnd vdd FILL
XFILL_2__12912_ gnd vdd FILL
XFILL_0__12002_ gnd vdd FILL
XFILL_1__14341_ gnd vdd FILL
XFILL_3__10374_ gnd vdd FILL
XFILL_1__11553_ gnd vdd FILL
XFILL_2__13892_ gnd vdd FILL
XFILL_0__10194_ gnd vdd FILL
XFILL_5__15811_ gnd vdd FILL
X_11409_ _11141_/A _11562_/B _11409_/C gnd _11411_/A vdd AOI21X1
XFILL_5__7475_ gnd vdd FILL
X_15177_ _7167_/A _15177_/B gnd _15184_/A vdd NAND2X1
XFILL_4__14452_ gnd vdd FILL
X_12389_ _12422_/A _12612_/A gnd _12390_/C vdd NAND2X1
XFILL_2__9505_ gnd vdd FILL
XFILL_3__12113_ gnd vdd FILL
XFILL_1__10504_ gnd vdd FILL
XFILL_2__15631_ gnd vdd FILL
XFILL_2_BUFX2_insert15 gnd vdd FILL
XFILL_3__13093_ gnd vdd FILL
XFILL_4__11664_ gnd vdd FILL
XFILL_2__12843_ gnd vdd FILL
XFILL_5__9214_ gnd vdd FILL
XFILL_1__14272_ gnd vdd FILL
XFILL_2_BUFX2_insert26 gnd vdd FILL
XFILL_6__12224_ gnd vdd FILL
XFILL_1__11484_ gnd vdd FILL
XFILL_2__7697_ gnd vdd FILL
X_14128_ _14127_/Y _13795_/B _13876_/C _14128_/D gnd _14128_/Y vdd OAI22X1
XFILL_4__13403_ gnd vdd FILL
XFILL_0__8520_ gnd vdd FILL
XFILL_2_BUFX2_insert37 gnd vdd FILL
XFILL_1__16011_ gnd vdd FILL
XFILL_2_BUFX2_insert48 gnd vdd FILL
XFILL_3__12044_ gnd vdd FILL
XFILL_4__10615_ gnd vdd FILL
XFILL_5__12954_ gnd vdd FILL
XFILL_5__15742_ gnd vdd FILL
XFILL_1__13223_ gnd vdd FILL
XFILL_2_BUFX2_insert59 gnd vdd FILL
XFILL_4__14383_ gnd vdd FILL
XFILL_2__12774_ gnd vdd FILL
XFILL_2__15562_ gnd vdd FILL
XFILL_1__10435_ gnd vdd FILL
XFILL_4__11595_ gnd vdd FILL
XFILL_5__9145_ gnd vdd FILL
XFILL_0__13953_ gnd vdd FILL
XFILL_0__8451_ gnd vdd FILL
XFILL_5__11905_ gnd vdd FILL
XFILL_4__16122_ gnd vdd FILL
XFILL_4__13334_ gnd vdd FILL
XFILL_5__15673_ gnd vdd FILL
X_14059_ _9698_/Q gnd _14061_/A vdd INVX1
XSFILL104360x78050 gnd vdd FILL
XFILL_2__14513_ gnd vdd FILL
XFILL_2__11725_ gnd vdd FILL
XFILL_5__12885_ gnd vdd FILL
XFILL_4__10546_ gnd vdd FILL
XFILL_2__9367_ gnd vdd FILL
XFILL_1__13154_ gnd vdd FILL
XFILL_0__12904_ gnd vdd FILL
XSFILL49560x5050 gnd vdd FILL
XFILL_1__10366_ gnd vdd FILL
XFILL_2__15493_ gnd vdd FILL
XFILL_0__13884_ gnd vdd FILL
XFILL_0__8382_ gnd vdd FILL
XFILL_5__14624_ gnd vdd FILL
XFILL_3__15803_ gnd vdd FILL
XFILL_3__7111_ gnd vdd FILL
XFILL_4__16053_ gnd vdd FILL
XFILL_5__11836_ gnd vdd FILL
XFILL_4__13265_ gnd vdd FILL
XFILL_1__12105_ gnd vdd FILL
XFILL_2__8318_ gnd vdd FILL
XSFILL109400x15050 gnd vdd FILL
XFILL_0__15623_ gnd vdd FILL
XFILL_3__8091_ gnd vdd FILL
XFILL_2__11656_ gnd vdd FILL
XFILL_2__14444_ gnd vdd FILL
XFILL_0__12835_ gnd vdd FILL
XFILL_1__13085_ gnd vdd FILL
XFILL_3__13995_ gnd vdd FILL
XFILL_2__9298_ gnd vdd FILL
XSFILL88840x75050 gnd vdd FILL
XFILL_0__7333_ gnd vdd FILL
XFILL_1__10297_ gnd vdd FILL
XFILL_6__11037_ gnd vdd FILL
XFILL_4__15004_ gnd vdd FILL
XFILL_5__14555_ gnd vdd FILL
XFILL_4__12216_ gnd vdd FILL
XFILL_3__7042_ gnd vdd FILL
XFILL112200x54050 gnd vdd FILL
X_7961_ _7959_/Y _7970_/B _7961_/C gnd _8033_/D vdd OAI21X1
XSFILL49080x36050 gnd vdd FILL
XFILL_5__11767_ gnd vdd FILL
XFILL_3__15734_ gnd vdd FILL
XFILL_2__8249_ gnd vdd FILL
XFILL_1__12036_ gnd vdd FILL
XFILL_2__14375_ gnd vdd FILL
XFILL_0__15554_ gnd vdd FILL
XFILL_2__11587_ gnd vdd FILL
XFILL_0__12766_ gnd vdd FILL
X_9700_ _9700_/Q _9306_/CLK _8801_/R vdd _9700_/D gnd vdd DFFSR
XSFILL39320x13050 gnd vdd FILL
XFILL_5__13506_ gnd vdd FILL
X_6912_ _6951_/A _8832_/B gnd _6912_/Y vdd NAND2X1
XFILL_5__14486_ gnd vdd FILL
XFILL_2__16114_ gnd vdd FILL
XFILL_4__12147_ gnd vdd FILL
XFILL_2__13326_ gnd vdd FILL
XFILL_3__15665_ gnd vdd FILL
XFILL_0__14505_ gnd vdd FILL
XFILL_5__11698_ gnd vdd FILL
XFILL_2__10538_ gnd vdd FILL
X_7892_ _7892_/A _9940_/B gnd _7892_/Y vdd NAND2X1
XFILL_3__12877_ gnd vdd FILL
XFILL_0__11717_ gnd vdd FILL
XFILL_0__9003_ gnd vdd FILL
XSFILL3960x44050 gnd vdd FILL
XFILL_0__15485_ gnd vdd FILL
XFILL_0__12697_ gnd vdd FILL
XFILL_5__16225_ gnd vdd FILL
XFILL_5__13437_ gnd vdd FILL
X_9631_ _9629_/Y _9597_/A _9631_/C gnd _9699_/D vdd OAI21X1
XFILL_5__9978_ gnd vdd FILL
XFILL_3__14616_ gnd vdd FILL
XFILL_5__10649_ gnd vdd FILL
X_6843_ _6843_/A gnd memoryAddress[5] vdd BUFX2
XFILL_0__7195_ gnd vdd FILL
XFILL_2__13257_ gnd vdd FILL
XFILL_2__16045_ gnd vdd FILL
XFILL_4__12078_ gnd vdd FILL
XFILL_3__11828_ gnd vdd FILL
XSFILL49000x7050 gnd vdd FILL
XFILL_3__15596_ gnd vdd FILL
XFILL_0__14436_ gnd vdd FILL
XSFILL53960x82050 gnd vdd FILL
XFILL_3__8993_ gnd vdd FILL
XFILL_1__13987_ gnd vdd FILL
XFILL_0__11648_ gnd vdd FILL
XFILL_5__16156_ gnd vdd FILL
X_9562_ _9562_/Q _9195_/CLK _8051_/R vdd _9562_/D gnd vdd DFFSR
XFILL_4__15906_ gnd vdd FILL
XFILL_5__13368_ gnd vdd FILL
XFILL_2__12208_ gnd vdd FILL
XFILL_4__11029_ gnd vdd FILL
XFILL_3__14547_ gnd vdd FILL
XSFILL18600x14050 gnd vdd FILL
XFILL_3__7944_ gnd vdd FILL
XFILL_1__15726_ gnd vdd FILL
XSFILL69240x49050 gnd vdd FILL
XFILL_3__11759_ gnd vdd FILL
XFILL_0__14367_ gnd vdd FILL
XFILL_5__15107_ gnd vdd FILL
XFILL_5__12319_ gnd vdd FILL
X_8513_ _8559_/Q gnd _8513_/Y vdd INVX1
XFILL_0__11579_ gnd vdd FILL
XFILL_5_BUFX2_insert405 gnd vdd FILL
XFILL_5__16087_ gnd vdd FILL
XFILL_5__13299_ gnd vdd FILL
XFILL_5_BUFX2_insert416 gnd vdd FILL
XFILL_2__12139_ gnd vdd FILL
XFILL_0__16106_ gnd vdd FILL
XFILL_4__15837_ gnd vdd FILL
X_9493_ _9554_/B _8853_/B gnd _9493_/Y vdd NAND2X1
XFILL_3__14478_ gnd vdd FILL
XFILL_0__13318_ gnd vdd FILL
XFILL_1__15657_ gnd vdd FILL
XFILL_1__12869_ gnd vdd FILL
XFILL_5_BUFX2_insert427 gnd vdd FILL
XFILL_3__7875_ gnd vdd FILL
XSFILL104440x58050 gnd vdd FILL
XFILL_5_BUFX2_insert438 gnd vdd FILL
XFILL_5__15038_ gnd vdd FILL
XFILL_0__9905_ gnd vdd FILL
XFILL_0__14298_ gnd vdd FILL
XSFILL64200x1050 gnd vdd FILL
XFILL_3__16217_ gnd vdd FILL
XFILL_5_BUFX2_insert449 gnd vdd FILL
XSFILL103800x1050 gnd vdd FILL
X_8444_ _8536_/Q gnd _8444_/Y vdd INVX1
XFILL_3__9614_ gnd vdd FILL
XFILL_3__13429_ gnd vdd FILL
XFILL_4__15768_ gnd vdd FILL
XFILL_1__6890_ gnd vdd FILL
XFILL_0__16037_ gnd vdd FILL
XFILL_1__14608_ gnd vdd FILL
XSFILL8680x56050 gnd vdd FILL
XFILL_0__13249_ gnd vdd FILL
XFILL_1__15588_ gnd vdd FILL
XFILL_4__14719_ gnd vdd FILL
X_8375_ _8375_/A _8333_/B _8374_/Y gnd _8375_/Y vdd OAI21X1
XSFILL104040x60050 gnd vdd FILL
XFILL_3__16148_ gnd vdd FILL
XFILL_4__15699_ gnd vdd FILL
XFILL_3__9545_ gnd vdd FILL
XFILL_1__14539_ gnd vdd FILL
X_7326_ _7369_/B _7326_/B gnd _7326_/Y vdd NAND2X1
XFILL_0__9767_ gnd vdd FILL
XFILL_2__15829_ gnd vdd FILL
XFILL_0__6979_ gnd vdd FILL
XFILL_3__16079_ gnd vdd FILL
XFILL_3__9476_ gnd vdd FILL
XFILL_0__8718_ gnd vdd FILL
X_7257_ _7167_/A _7129_/CLK _8542_/R vdd _7257_/D gnd vdd DFFSR
XFILL_1__8491_ gnd vdd FILL
XFILL_1__16209_ gnd vdd FILL
XSFILL108680x63050 gnd vdd FILL
XFILL_4__7220_ gnd vdd FILL
XSFILL13640x57050 gnd vdd FILL
XFILL_1__7442_ gnd vdd FILL
XFILL_0__8649_ gnd vdd FILL
X_7188_ _7188_/A gnd _7190_/A vdd INVX1
XFILL_3__8358_ gnd vdd FILL
XFILL_6__8067_ gnd vdd FILL
XFILL_1__7373_ gnd vdd FILL
XFILL_3__7309_ gnd vdd FILL
XFILL_2_BUFX2_insert306 gnd vdd FILL
XFILL_1_BUFX2_insert1 gnd vdd FILL
XFILL_4__7082_ gnd vdd FILL
XFILL_2_BUFX2_insert317 gnd vdd FILL
XFILL_2_BUFX2_insert328 gnd vdd FILL
XFILL_1__9112_ gnd vdd FILL
XFILL_2_BUFX2_insert339 gnd vdd FILL
XSFILL104520x38050 gnd vdd FILL
XFILL_1__9043_ gnd vdd FILL
XSFILL8760x36050 gnd vdd FILL
XSFILL17880x62050 gnd vdd FILL
X_11760_ _11019_/Y _11020_/Y _11776_/B gnd _11760_/Y vdd OAI21X1
X_9829_ _9829_/Q _8025_/CLK _8025_/R vdd _9765_/Y gnd vdd DFFSR
X_10711_ _13530_/A _7640_/CLK _7515_/R vdd _10619_/Y gnd vdd DFFSR
XFILL_4__7984_ gnd vdd FILL
X_11691_ _11684_/B _11046_/Y _11743_/A gnd _11691_/Y vdd OAI21X1
XBUFX2_insert305 _11983_/Y gnd _12031_/C vdd BUFX2
XFILL_4__9723_ gnd vdd FILL
XBUFX2_insert316 _13454_/Y gnd _14872_/C vdd BUFX2
XFILL_4__6935_ gnd vdd FILL
X_13430_ _14045_/A gnd _13430_/Y vdd INVX8
X_10642_ _10676_/B _7954_/B gnd _10642_/Y vdd NAND2X1
XBUFX2_insert327 _13345_/Y gnd _9937_/A vdd BUFX2
XBUFX2_insert338 _12811_/Q gnd _11884_/A vdd BUFX2
XBUFX2_insert349 _10927_/Y gnd _12216_/A vdd BUFX2
XSFILL13720x37050 gnd vdd FILL
XFILL_4__9654_ gnd vdd FILL
X_13361_ _13361_/A _13360_/Y gnd _13361_/Y vdd NOR2X1
XFILL_4__6866_ gnd vdd FILL
X_10573_ _10573_/A gnd _10575_/A vdd INVX1
XFILL_5_CLKBUF1_insert206 gnd vdd FILL
XSFILL23880x81050 gnd vdd FILL
XFILL_5_CLKBUF1_insert217 gnd vdd FILL
XFILL_5_BUFX2_insert950 gnd vdd FILL
XFILL_1__9876_ gnd vdd FILL
XFILL_4__8605_ gnd vdd FILL
X_15100_ _15981_/B gnd _16204_/B vdd INVX4
XFILL_5_BUFX2_insert961 gnd vdd FILL
X_12312_ _12312_/A _12313_/D _12312_/C gnd _12312_/Y vdd NAND3X1
X_13292_ _13297_/A _13292_/B gnd _13293_/B vdd OR2X2
XFILL_5_BUFX2_insert972 gnd vdd FILL
X_16080_ _16079_/Y _16078_/Y gnd _16085_/A vdd NOR2X1
XFILL_5_BUFX2_insert983 gnd vdd FILL
XFILL_2__7620_ gnd vdd FILL
XFILL_1__8827_ gnd vdd FILL
XFILL_5_BUFX2_insert994 gnd vdd FILL
X_15031_ _15012_/Y _15031_/B _15656_/B gnd _15031_/Y vdd AOI21X1
X_12243_ _12239_/A gnd _12239_/C gnd _12246_/A vdd NAND3X1
XFILL_2__7551_ gnd vdd FILL
XFILL_1__8758_ gnd vdd FILL
XSFILL13640x3050 gnd vdd FILL
XFILL_4__8467_ gnd vdd FILL
X_12174_ _12174_/A _12117_/B _12174_/C gnd _12174_/Y vdd OAI21X1
XFILL_1__7709_ gnd vdd FILL
XFILL_2__7482_ gnd vdd FILL
XFILL_4__7418_ gnd vdd FILL
XFILL_5__7191_ gnd vdd FILL
X_11125_ _11125_/A _11125_/B gnd _11126_/A vdd NOR2X1
XFILL_4__8398_ gnd vdd FILL
XFILL_4__10400_ gnd vdd FILL
XFILL_2__9221_ gnd vdd FILL
XFILL_4__11380_ gnd vdd FILL
XFILL_0__10950_ gnd vdd FILL
XFILL_4__7349_ gnd vdd FILL
X_15933_ _15932_/Y _15930_/Y gnd _15936_/C vdd NOR2X1
X_11056_ _11056_/A _11055_/Y gnd _11056_/Y vdd NOR2X1
XFILL_2__11510_ gnd vdd FILL
XFILL_2__9152_ gnd vdd FILL
XFILL_1__10151_ gnd vdd FILL
XFILL_2__12490_ gnd vdd FILL
X_10007_ _14016_/A gnd _10007_/Y vdd INVX1
XFILL_0__10881_ gnd vdd FILL
XFILL_5__11621_ gnd vdd FILL
XFILL_2__8103_ gnd vdd FILL
X_15864_ _16293_/A _7090_/A _15380_/C _9906_/A gnd _15865_/C vdd AOI22X1
XFILL_4__10262_ gnd vdd FILL
XSFILL13800x17050 gnd vdd FILL
XFILL_2__11441_ gnd vdd FILL
XFILL_2__9083_ gnd vdd FILL
XFILL_4__9019_ gnd vdd FILL
XFILL_0__12620_ gnd vdd FILL
XFILL_3__13780_ gnd vdd FILL
XFILL_2_BUFX2_insert840 gnd vdd FILL
XFILL_5__9901_ gnd vdd FILL
XFILL_2_BUFX2_insert851 gnd vdd FILL
XFILL_3__10992_ gnd vdd FILL
XFILL112120x69050 gnd vdd FILL
XFILL_4__12001_ gnd vdd FILL
X_14815_ _14814_/Y _14615_/B _14815_/C _14813_/Y gnd _14815_/Y vdd OAI22X1
XFILL_5__14340_ gnd vdd FILL
XFILL_2_BUFX2_insert862 gnd vdd FILL
XFILL_5__11552_ gnd vdd FILL
XFILL_3__12731_ gnd vdd FILL
XFILL_2__14160_ gnd vdd FILL
X_15795_ _15795_/A _15795_/B _15795_/C gnd _15795_/Y vdd OAI21X1
XFILL_2_BUFX2_insert873 gnd vdd FILL
XFILL_4__10193_ gnd vdd FILL
XSFILL64040x54050 gnd vdd FILL
XFILL_2_BUFX2_insert884 gnd vdd FILL
XFILL_1__13910_ gnd vdd FILL
XFILL_2__11372_ gnd vdd FILL
XFILL_2_BUFX2_insert895 gnd vdd FILL
XFILL_1__14890_ gnd vdd FILL
XFILL_5__10503_ gnd vdd FILL
XFILL_2__13111_ gnd vdd FILL
XFILL_5__14271_ gnd vdd FILL
X_14746_ _10481_/Q _14389_/B _14273_/C _8519_/A gnd _14746_/Y vdd AOI22X1
X_11958_ _11956_/Y _11909_/A _11958_/C gnd _6861_/A vdd OAI21X1
XFILL_3__15450_ gnd vdd FILL
XFILL_5__11483_ gnd vdd FILL
XFILL_2__10323_ gnd vdd FILL
XFILL_3__12662_ gnd vdd FILL
XFILL_1__13841_ gnd vdd FILL
XFILL_2__14091_ gnd vdd FILL
XFILL_0__11502_ gnd vdd FILL
XFILL_5__16010_ gnd vdd FILL
XFILL_0__15270_ gnd vdd FILL
XFILL_5__13222_ gnd vdd FILL
XFILL_5__9763_ gnd vdd FILL
XFILL_0__12482_ gnd vdd FILL
XFILL_5__6975_ gnd vdd FILL
X_10909_ _10938_/A gnd _10944_/A vdd INVX2
XFILL_3__14401_ gnd vdd FILL
XFILL_5__10434_ gnd vdd FILL
XFILL_3__11613_ gnd vdd FILL
X_14677_ _7535_/Q gnd _14678_/D vdd INVX1
XSFILL43880x12050 gnd vdd FILL
XFILL_4__13952_ gnd vdd FILL
XFILL_2__13042_ gnd vdd FILL
XFILL_2__10254_ gnd vdd FILL
XFILL_3__15381_ gnd vdd FILL
X_11889_ _11889_/A _11975_/A _11889_/C gnd _6838_/A vdd OAI21X1
XFILL_0__14221_ gnd vdd FILL
XFILL_4_BUFX2_insert5 gnd vdd FILL
XFILL_3__12593_ gnd vdd FILL
XFILL_2__9985_ gnd vdd FILL
XSFILL3480x61050 gnd vdd FILL
XFILL_5__8714_ gnd vdd FILL
XFILL_1__13772_ gnd vdd FILL
XFILL_0__11433_ gnd vdd FILL
X_16416_ _16414_/Y gnd _16416_/C gnd _16448_/D vdd OAI21X1
X_13628_ _10751_/A gnd _13628_/Y vdd INVX1
XFILL_5__13153_ gnd vdd FILL
XFILL_4__12903_ gnd vdd FILL
XFILL_3__14332_ gnd vdd FILL
XFILL_5__10365_ gnd vdd FILL
XFILL_1__12723_ gnd vdd FILL
XFILL_4__13883_ gnd vdd FILL
XFILL_1__15511_ gnd vdd FILL
XFILL_3__11544_ gnd vdd FILL
XFILL_0__14152_ gnd vdd FILL
XFILL_2__10185_ gnd vdd FILL
XSFILL84200x67050 gnd vdd FILL
XFILL_5__12104_ gnd vdd FILL
XFILL_5__8645_ gnd vdd FILL
XBUFX2_insert850 _13269_/Y gnd _7064_/A vdd BUFX2
XFILL_0__11364_ gnd vdd FILL
X_16347_ _16345_/Y gnd _16347_/C gnd _16425_/D vdd OAI21X1
XFILL_4__15622_ gnd vdd FILL
XBUFX2_insert861 _13314_/Y gnd _8244_/B vdd BUFX2
XFILL_0__7951_ gnd vdd FILL
XFILL_4__12834_ gnd vdd FILL
XBUFX2_insert872 _13435_/Y gnd _14211_/A vdd BUFX2
XFILL_5__13084_ gnd vdd FILL
X_13559_ _13559_/A _13558_/Y gnd _13559_/Y vdd NAND2X1
XFILL_3__14263_ gnd vdd FILL
XFILL_0__13103_ gnd vdd FILL
XFILL_5__10296_ gnd vdd FILL
XBUFX2_insert883 _12216_/Y gnd _12249_/C vdd BUFX2
XFILL_1__12654_ gnd vdd FILL
XBUFX2_insert894 _12369_/Y gnd _8207_/B vdd BUFX2
XFILL_0__10315_ gnd vdd FILL
XFILL_3__11475_ gnd vdd FILL
XFILL_2__8867_ gnd vdd FILL
XFILL_1__15442_ gnd vdd FILL
XFILL_2__14993_ gnd vdd FILL
XFILL_0__14083_ gnd vdd FILL
XFILL_5__8576_ gnd vdd FILL
XFILL_3__16002_ gnd vdd FILL
XFILL_0__6902_ gnd vdd FILL
XFILL_5__12035_ gnd vdd FILL
XFILL_0__11295_ gnd vdd FILL
XFILL_3__13214_ gnd vdd FILL
XFILL_4__15553_ gnd vdd FILL
X_16278_ _8564_/Q gnd _16279_/B vdd INVX1
XFILL_4__12765_ gnd vdd FILL
XFILL_0__7882_ gnd vdd FILL
XFILL_2__7818_ gnd vdd FILL
XFILL_3__10426_ gnd vdd FILL
XFILL_1__11605_ gnd vdd FILL
XFILL_1__15373_ gnd vdd FILL
XFILL_3__14194_ gnd vdd FILL
XFILL_0__13034_ gnd vdd FILL
XFILL_2__13944_ gnd vdd FILL
XFILL_3__7591_ gnd vdd FILL
XFILL_1__12585_ gnd vdd FILL
XFILL_0__10246_ gnd vdd FILL
X_15229_ _15223_/Y _15225_/Y _15229_/C gnd _15229_/Y vdd NAND3X1
XFILL_4__14504_ gnd vdd FILL
XFILL_0__9621_ gnd vdd FILL
XFILL_4__11716_ gnd vdd FILL
X_8160_ _8160_/Q _7007_/CLK _9332_/R vdd _8160_/D gnd vdd DFFSR
XFILL_3__13145_ gnd vdd FILL
XFILL_1__14324_ gnd vdd FILL
XFILL_4__15484_ gnd vdd FILL
XFILL_4__12696_ gnd vdd FILL
XFILL112200x49050 gnd vdd FILL
XFILL_1__11536_ gnd vdd FILL
XFILL_2__7749_ gnd vdd FILL
XFILL_2__13875_ gnd vdd FILL
XFILL_5__7458_ gnd vdd FILL
X_7111_ _7153_/Q gnd _7113_/A vdd INVX1
XFILL_0__10177_ gnd vdd FILL
XFILL_4__14435_ gnd vdd FILL
XFILL_0__9552_ gnd vdd FILL
XFILL_2__15614_ gnd vdd FILL
X_8091_ _8100_/A _8091_/B gnd _8091_/Y vdd NAND2X1
XFILL_4__11647_ gnd vdd FILL
XFILL_1__14255_ gnd vdd FILL
XFILL_5__13986_ gnd vdd FILL
XFILL_3__10288_ gnd vdd FILL
XFILL_3__9261_ gnd vdd FILL
XFILL_2__12826_ gnd vdd FILL
XFILL_1__11467_ gnd vdd FILL
XFILL_0__8503_ gnd vdd FILL
XFILL_0__14985_ gnd vdd FILL
XFILL_5__15725_ gnd vdd FILL
X_7042_ _7130_/Q gnd _7044_/A vdd INVX1
XFILL_0__9483_ gnd vdd FILL
XFILL_2__9419_ gnd vdd FILL
XFILL_3__12027_ gnd vdd FILL
XFILL_4__14366_ gnd vdd FILL
XFILL_3__8212_ gnd vdd FILL
XFILL_2__15545_ gnd vdd FILL
XFILL_1__10418_ gnd vdd FILL
XFILL_4__11578_ gnd vdd FILL
XFILL_1__14186_ gnd vdd FILL
XFILL_2__12757_ gnd vdd FILL
XFILL_5__9128_ gnd vdd FILL
XFILL_0__13936_ gnd vdd FILL
XFILL_4__16105_ gnd vdd FILL
XFILL_1__11398_ gnd vdd FILL
XFILL_4__13317_ gnd vdd FILL
XSFILL53960x77050 gnd vdd FILL
XFILL_5__15656_ gnd vdd FILL
XFILL_4__10529_ gnd vdd FILL
XFILL_5__12868_ gnd vdd FILL
XSFILL3560x41050 gnd vdd FILL
XFILL_3__8143_ gnd vdd FILL
XFILL_1__13137_ gnd vdd FILL
XFILL_2__11708_ gnd vdd FILL
XFILL_4__14297_ gnd vdd FILL
XFILL_2__15476_ gnd vdd FILL
XFILL_0__13867_ gnd vdd FILL
XFILL_5__14607_ gnd vdd FILL
XFILL_4__16036_ gnd vdd FILL
XSFILL28760x53050 gnd vdd FILL
XFILL_0__8365_ gnd vdd FILL
XFILL_5__11819_ gnd vdd FILL
XFILL_4__13248_ gnd vdd FILL
XFILL_3__8074_ gnd vdd FILL
X_8993_ _9014_/A _8225_/B gnd _8993_/Y vdd NAND2X1
XFILL_5__15587_ gnd vdd FILL
XFILL_2__14427_ gnd vdd FILL
XFILL_3__13978_ gnd vdd FILL
XFILL_2__11639_ gnd vdd FILL
XFILL_0__15606_ gnd vdd FILL
XFILL_0__13798_ gnd vdd FILL
XFILL_0__7316_ gnd vdd FILL
X_7944_ _7944_/A gnd _7944_/Y vdd INVX1
XFILL_3__15717_ gnd vdd FILL
XFILL_5__14538_ gnd vdd FILL
XFILL_1__12019_ gnd vdd FILL
XFILL_0__15537_ gnd vdd FILL
XFILL_2__14358_ gnd vdd FILL
XFILL_0__12749_ gnd vdd FILL
XFILL_0__7247_ gnd vdd FILL
XFILL_6__15828_ gnd vdd FILL
XFILL_5__14469_ gnd vdd FILL
XFILL_2__13309_ gnd vdd FILL
XFILL_3__15648_ gnd vdd FILL
X_7875_ _7873_/Y _7892_/A _7875_/C gnd _7875_/Y vdd OAI21X1
XFILL_2__14289_ gnd vdd FILL
XFILL_0__15468_ gnd vdd FILL
XFILL111800x22050 gnd vdd FILL
XFILL_5__16208_ gnd vdd FILL
XFILL_6__8754_ gnd vdd FILL
XFILL_0__7178_ gnd vdd FILL
X_9614_ _9694_/Q gnd _9616_/A vdd INVX1
XSFILL48920x66050 gnd vdd FILL
XFILL_2__16028_ gnd vdd FILL
XFILL_0__14419_ gnd vdd FILL
XFILL_3__15579_ gnd vdd FILL
XSFILL89560x16050 gnd vdd FILL
XFILL_3__8976_ gnd vdd FILL
XFILL_6__7705_ gnd vdd FILL
XSFILL64200x14050 gnd vdd FILL
XFILL_0__15399_ gnd vdd FILL
X_9545_ _9543_/Y _9466_/A _9545_/C gnd _9585_/D vdd OAI21X1
XSFILL48920x50 gnd vdd FILL
XFILL_5__16139_ gnd vdd FILL
XFILL_1__7991_ gnd vdd FILL
XFILL_1__15709_ gnd vdd FILL
XFILL_3__7927_ gnd vdd FILL
XSFILL49000x75050 gnd vdd FILL
XFILL_1__9730_ gnd vdd FILL
XFILL_5_BUFX2_insert235 gnd vdd FILL
X_9476_ _9476_/A _9551_/B _9475_/Y gnd _9562_/D vdd OAI21X1
XFILL_1__6942_ gnd vdd FILL
XSFILL89400x80050 gnd vdd FILL
XFILL_5_BUFX2_insert246 gnd vdd FILL
XFILL_5_BUFX2_insert257 gnd vdd FILL
XFILL_3__7858_ gnd vdd FILL
XFILL_5_BUFX2_insert268 gnd vdd FILL
XSFILL3640x21050 gnd vdd FILL
X_8427_ _8427_/Q _7915_/CLK _7915_/R vdd _8375_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert279 gnd vdd FILL
XFILL_1__9661_ gnd vdd FILL
XFILL_1__6873_ gnd vdd FILL
XFILL_4_BUFX2_insert902 gnd vdd FILL
XFILL_4__9370_ gnd vdd FILL
XSFILL28840x33050 gnd vdd FILL
XFILL_4_BUFX2_insert913 gnd vdd FILL
XSFILL79480x68050 gnd vdd FILL
XFILL_1__8612_ gnd vdd FILL
XFILL_4_BUFX2_insert924 gnd vdd FILL
X_8358_ _8422_/Q gnd _8360_/A vdd INVX1
XFILL_4_BUFX2_insert935 gnd vdd FILL
XFILL_4__8321_ gnd vdd FILL
XFILL_1__9592_ gnd vdd FILL
XFILL_4_BUFX2_insert946 gnd vdd FILL
XFILL_3__9528_ gnd vdd FILL
XFILL_4_BUFX2_insert957 gnd vdd FILL
XFILL_4_BUFX2_insert968 gnd vdd FILL
X_7309_ _7307_/Y _7308_/A _7309_/C gnd _7389_/D vdd OAI21X1
XSFILL79080x70050 gnd vdd FILL
XFILL_4_BUFX2_insert979 gnd vdd FILL
X_8289_ _8215_/A _8289_/CLK _8688_/R vdd _8289_/D gnd vdd DFFSR
XFILL_4__8252_ gnd vdd FILL
XSFILL33960x24050 gnd vdd FILL
XFILL_4__7203_ gnd vdd FILL
XFILL_1__8474_ gnd vdd FILL
XFILL_4__8183_ gnd vdd FILL
XSFILL74840x36050 gnd vdd FILL
XFILL_1__7425_ gnd vdd FILL
XFILL_2_BUFX2_insert103 gnd vdd FILL
X_12930_ _12856_/A _7532_/CLK _8816_/R vdd _12930_/D gnd vdd DFFSR
XFILL_1__7356_ gnd vdd FILL
XFILL_4__7065_ gnd vdd FILL
X_12861_ _12859_/Y vdd _12861_/C gnd _12931_/D vdd OAI21X1
XSFILL23880x76050 gnd vdd FILL
XFILL_1__7287_ gnd vdd FILL
X_14600_ _14598_/Y _13871_/A _14456_/C _14599_/Y gnd _14600_/Y vdd OAI22X1
XFILL_1_BUFX2_insert803 gnd vdd FILL
X_11812_ _11810_/Y _11005_/Y _11802_/A gnd _11812_/Y vdd OAI21X1
XFILL_1_BUFX2_insert814 gnd vdd FILL
XFILL_1__9026_ gnd vdd FILL
X_15580_ _15580_/A _15580_/B _15579_/Y gnd _15586_/B vdd NAND3X1
XFILL_1_BUFX2_insert825 gnd vdd FILL
X_12792_ _12792_/Q _7005_/CLK _12799_/R vdd _12700_/Y gnd vdd DFFSR
XSFILL28920x13050 gnd vdd FILL
XFILL_1_BUFX2_insert836 gnd vdd FILL
XFILL_1_BUFX2_insert847 gnd vdd FILL
X_14531_ _9016_/A gnd _14532_/D vdd INVX1
XFILL_1_BUFX2_insert858 gnd vdd FILL
X_11743_ _11743_/A _11737_/C gnd _11743_/Y vdd NAND2X1
XFILL_1_BUFX2_insert869 gnd vdd FILL
XBUFX2_insert102 _15009_/Y gnd _15010_/A vdd BUFX2
XFILL_4__7967_ gnd vdd FILL
X_14462_ _8299_/Q gnd _14463_/B vdd INVX1
X_11674_ _11673_/Y _11674_/B gnd _11675_/A vdd NOR2X1
XFILL_2__9770_ gnd vdd FILL
X_16201_ _16201_/A _16201_/B gnd _16202_/A vdd NAND2X1
XFILL_2__6982_ gnd vdd FILL
XFILL_4__6918_ gnd vdd FILL
X_13413_ _11884_/A _13390_/B gnd _13630_/B vdd NAND2X1
X_10625_ _10623_/Y _10661_/B _10625_/C gnd _10713_/D vdd OAI21X1
XFILL_5__10150_ gnd vdd FILL
XSFILL58840x49050 gnd vdd FILL
X_14393_ _14700_/A _14393_/B _13587_/C _15815_/D gnd _14393_/Y vdd OAI22X1
XFILL_2__8721_ gnd vdd FILL
XFILL_1__9928_ gnd vdd FILL
XFILL_4__10880_ gnd vdd FILL
XFILL_4__9637_ gnd vdd FILL
XSFILL18840x65050 gnd vdd FILL
XFILL_4__6849_ gnd vdd FILL
X_16132_ _7751_/A _15969_/C gnd _16132_/Y vdd NAND2X1
X_13344_ _13343_/Y _13335_/A gnd _13344_/Y vdd AND2X2
X_10556_ _10557_/B _8764_/B gnd _10556_/Y vdd NAND2X1
XSFILL84280x41050 gnd vdd FILL
XSFILL34120x13050 gnd vdd FILL
XFILL_3__11260_ gnd vdd FILL
XFILL_2__8652_ gnd vdd FILL
XFILL_1__9859_ gnd vdd FILL
XFILL_5_BUFX2_insert780 gnd vdd FILL
XFILL_2__11990_ gnd vdd FILL
XFILL_0__11080_ gnd vdd FILL
XFILL_5__8361_ gnd vdd FILL
XFILL_5_BUFX2_insert791 gnd vdd FILL
XSFILL99320x63050 gnd vdd FILL
X_16063_ _8943_/Q gnd _16063_/Y vdd INVX1
X_13275_ _13297_/A _13275_/B gnd _13276_/B vdd OR2X2
X_10487_ _6903_/A _10505_/A gnd _10488_/C vdd NAND2X1
XFILL_2__7603_ gnd vdd FILL
XFILL_3__11191_ gnd vdd FILL
XFILL_2__10941_ gnd vdd FILL
XFILL_5__7312_ gnd vdd FILL
XFILL_1__12370_ gnd vdd FILL
XFILL_6__13110_ gnd vdd FILL
XFILL_4__8519_ gnd vdd FILL
XFILL_0__10031_ gnd vdd FILL
XFILL_2__8583_ gnd vdd FILL
X_15014_ _15036_/A _15012_/Y _15014_/C gnd _15177_/B vdd NOR3X1
XFILL_4__9499_ gnd vdd FILL
X_12226_ _12226_/A _12226_/B _12226_/C gnd _12226_/Y vdd NAND3X1
XFILL_4__11501_ gnd vdd FILL
XFILL_5__13840_ gnd vdd FILL
XFILL_3__10142_ gnd vdd FILL
XFILL_4__12481_ gnd vdd FILL
XSFILL63960x9050 gnd vdd FILL
XFILL_1__11321_ gnd vdd FILL
XFILL_2__13660_ gnd vdd FILL
XFILL_2__10872_ gnd vdd FILL
XFILL_5__7243_ gnd vdd FILL
XSFILL64040x49050 gnd vdd FILL
XFILL_4__14220_ gnd vdd FILL
X_12157_ _11929_/A gnd _12159_/A vdd INVX1
XFILL_5__13771_ gnd vdd FILL
XFILL_4__11432_ gnd vdd FILL
XFILL_5__10983_ gnd vdd FILL
XFILL_2__12611_ gnd vdd FILL
XFILL_1__14040_ gnd vdd FILL
XFILL_3__14950_ gnd vdd FILL
XFILL_2__7465_ gnd vdd FILL
XFILL_1__11252_ gnd vdd FILL
XFILL_2__13591_ gnd vdd FILL
XFILL_0__14770_ gnd vdd FILL
X_11108_ _12180_/Y gnd _11108_/Y vdd INVX1
XFILL_5__12722_ gnd vdd FILL
XFILL_5__15510_ gnd vdd FILL
XFILL_0__11982_ gnd vdd FILL
XFILL_5__7174_ gnd vdd FILL
XFILL_4__14151_ gnd vdd FILL
X_12088_ _12012_/A _12764_/A _11996_/C gnd _12090_/B vdd NAND3X1
XFILL_3__13901_ gnd vdd FILL
XFILL_2__15330_ gnd vdd FILL
XSFILL79240x30050 gnd vdd FILL
XFILL_4__11363_ gnd vdd FILL
XFILL_3__14881_ gnd vdd FILL
XFILL_0__13721_ gnd vdd FILL
XFILL_0__10933_ gnd vdd FILL
XFILL_1__11183_ gnd vdd FILL
X_15916_ _10677_/A _15916_/B _15915_/Y gnd _15917_/B vdd AOI21X1
XFILL_4__13102_ gnd vdd FILL
X_11039_ _11384_/A _11038_/Y gnd _11040_/C vdd NOR2X1
XFILL_5__12653_ gnd vdd FILL
XSFILL93480x78050 gnd vdd FILL
XFILL_4__10314_ gnd vdd FILL
XFILL_5__15441_ gnd vdd FILL
XFILL_3__13832_ gnd vdd FILL
XFILL_2__9135_ gnd vdd FILL
XFILL_4__14082_ gnd vdd FILL
XFILL_2__12473_ gnd vdd FILL
XSFILL69160x3050 gnd vdd FILL
XFILL_1__10134_ gnd vdd FILL
XFILL_4__11294_ gnd vdd FILL
XFILL_2__15261_ gnd vdd FILL
XSFILL28680x68050 gnd vdd FILL
XFILL_0__13652_ gnd vdd FILL
XFILL_1__15991_ gnd vdd FILL
XFILL_5__11604_ gnd vdd FILL
XFILL_5__15372_ gnd vdd FILL
X_15847_ _9193_/Q gnd _15848_/B vdd INVX1
XFILL_4__13033_ gnd vdd FILL
XFILL_2__14212_ gnd vdd FILL
XFILL_5__12584_ gnd vdd FILL
XFILL_4__10245_ gnd vdd FILL
XFILL_2__11424_ gnd vdd FILL
XFILL_0__12603_ gnd vdd FILL
XFILL_2_BUFX2_insert670 gnd vdd FILL
XFILL_3__13763_ gnd vdd FILL
XFILL_0__7101_ gnd vdd FILL
XFILL_3__10975_ gnd vdd FILL
XFILL_2__15192_ gnd vdd FILL
XFILL_0__16371_ gnd vdd FILL
XFILL_1__14942_ gnd vdd FILL
XFILL_2_BUFX2_insert681 gnd vdd FILL
XFILL_1__10065_ gnd vdd FILL
XFILL_5__14323_ gnd vdd FILL
XFILL_0__13583_ gnd vdd FILL
XFILL_0__10795_ gnd vdd FILL
XFILL_0__8081_ gnd vdd FILL
XFILL_5__11535_ gnd vdd FILL
XFILL_3__15502_ gnd vdd FILL
XFILL_2_BUFX2_insert692 gnd vdd FILL
XFILL_3__12714_ gnd vdd FILL
XFILL_6__13874_ gnd vdd FILL
X_15778_ _7724_/A _15969_/C gnd _15778_/Y vdd NAND2X1
XFILL_2__8017_ gnd vdd FILL
XFILL_4__10176_ gnd vdd FILL
XFILL_2__14143_ gnd vdd FILL
XFILL_0__15322_ gnd vdd FILL
XFILL_2__11355_ gnd vdd FILL
XFILL_0__12534_ gnd vdd FILL
XFILL_3__13694_ gnd vdd FILL
XFILL_1__14873_ gnd vdd FILL
XFILL_6__15613_ gnd vdd FILL
XFILL_0__7032_ gnd vdd FILL
XFILL_5__14254_ gnd vdd FILL
X_14729_ _14729_/A _14728_/Y gnd _14730_/A vdd NOR2X1
X_7660_ _7608_/A _7661_/CLK _9203_/R vdd _7660_/D gnd vdd DFFSR
XFILL_2__10306_ gnd vdd FILL
XFILL_3__15433_ gnd vdd FILL
XFILL_5__11466_ gnd vdd FILL
XFILL_3__12645_ gnd vdd FILL
XFILL_4__14984_ gnd vdd FILL
XFILL_2__14074_ gnd vdd FILL
XFILL_3__8830_ gnd vdd FILL
XFILL_1__13824_ gnd vdd FILL
XFILL_0__15253_ gnd vdd FILL
XFILL_5_BUFX2_insert30 gnd vdd FILL
XFILL_2__11286_ gnd vdd FILL
XFILL_0__12465_ gnd vdd FILL
XFILL_5__9746_ gnd vdd FILL
XFILL_5_BUFX2_insert41 gnd vdd FILL
XFILL_5__6958_ gnd vdd FILL
XFILL_5__10417_ gnd vdd FILL
XFILL_5__14185_ gnd vdd FILL
XFILL_2__13025_ gnd vdd FILL
XFILL_5_BUFX2_insert52 gnd vdd FILL
XFILL_4__13935_ gnd vdd FILL
X_7591_ _7592_/B _7975_/B gnd _7591_/Y vdd NAND2X1
XFILL_0__14204_ gnd vdd FILL
XFILL_3__15364_ gnd vdd FILL
XSFILL64120x29050 gnd vdd FILL
XFILL_5_BUFX2_insert63 gnd vdd FILL
XFILL_5__11397_ gnd vdd FILL
XFILL_2__10237_ gnd vdd FILL
XFILL_5_BUFX2_insert74 gnd vdd FILL
XFILL_3__12576_ gnd vdd FILL
XFILL_3__8761_ gnd vdd FILL
XFILL_0__11416_ gnd vdd FILL
XFILL_1__10967_ gnd vdd FILL
XFILL_0__15184_ gnd vdd FILL
XFILL_1__13755_ gnd vdd FILL
XFILL_5_BUFX2_insert85 gnd vdd FILL
XFILL_5__9677_ gnd vdd FILL
XFILL_5__13136_ gnd vdd FILL
X_9330_ _9290_/A _8818_/CLK _8278_/R vdd _9292_/Y gnd vdd DFFSR
XFILL_0__12396_ gnd vdd FILL
XFILL_6__11707_ gnd vdd FILL
XFILL_6__8470_ gnd vdd FILL
XFILL_5_BUFX2_insert96 gnd vdd FILL
XFILL_3__14315_ gnd vdd FILL
XFILL_5__6889_ gnd vdd FILL
XFILL_6__15475_ gnd vdd FILL
XFILL_4__13866_ gnd vdd FILL
XFILL_0__8983_ gnd vdd FILL
XSFILL89880x52050 gnd vdd FILL
XFILL_3__7712_ gnd vdd FILL
XFILL_3__11527_ gnd vdd FILL
XFILL_1__12706_ gnd vdd FILL
XFILL_0__14135_ gnd vdd FILL
XFILL_2__10168_ gnd vdd FILL
XFILL_3__15295_ gnd vdd FILL
XFILL_1__13686_ gnd vdd FILL
XBUFX2_insert680 _15005_/Y gnd _15915_/C vdd BUFX2
XFILL_6__7421_ gnd vdd FILL
XFILL_5__8628_ gnd vdd FILL
XFILL_2__9899_ gnd vdd FILL
XFILL_0__11347_ gnd vdd FILL
XFILL_1__10898_ gnd vdd FILL
XBUFX2_insert691 _13362_/Y gnd _10581_/B vdd BUFX2
XFILL_6__14426_ gnd vdd FILL
X_9261_ _9208_/B _7853_/B gnd _9261_/Y vdd NAND2X1
XFILL_0__7934_ gnd vdd FILL
XFILL_4__15605_ gnd vdd FILL
XFILL_3__14246_ gnd vdd FILL
XFILL_5__10279_ gnd vdd FILL
XSFILL3560x36050 gnd vdd FILL
XFILL_1__12637_ gnd vdd FILL
XFILL_4__13797_ gnd vdd FILL
XFILL_3__11458_ gnd vdd FILL
XFILL_1__15425_ gnd vdd FILL
XFILL_0__14066_ gnd vdd FILL
XFILL_2__14976_ gnd vdd FILL
XFILL_5__12018_ gnd vdd FILL
X_8212_ _8212_/A gnd _8212_/Y vdd INVX1
XFILL_0__11278_ gnd vdd FILL
XFILL_4__15536_ gnd vdd FILL
XFILL_6__11569_ gnd vdd FILL
XFILL_4__12748_ gnd vdd FILL
XFILL_0__7865_ gnd vdd FILL
X_9192_ _9192_/Q _7016_/CLK _8424_/R vdd _9134_/Y gnd vdd DFFSR
XFILL_3__10409_ gnd vdd FILL
XSFILL53560x74050 gnd vdd FILL
XFILL_3__14177_ gnd vdd FILL
XFILL_0__13017_ gnd vdd FILL
XFILL_2__13927_ gnd vdd FILL
XFILL_1__12568_ gnd vdd FILL
XFILL_1__15356_ gnd vdd FILL
XFILL_3__7574_ gnd vdd FILL
XFILL_3__11389_ gnd vdd FILL
XFILL_0__9604_ gnd vdd FILL
X_8143_ _8143_/A _8142_/A _8143_/C gnd _8143_/Y vdd OAI21X1
XFILL_3__13128_ gnd vdd FILL
XFILL_4__15467_ gnd vdd FILL
XFILL_6__14288_ gnd vdd FILL
XFILL_1__14307_ gnd vdd FILL
XFILL_1__11519_ gnd vdd FILL
XFILL_3_BUFX2_insert909 gnd vdd FILL
XFILL_2__13858_ gnd vdd FILL
XFILL_6__9022_ gnd vdd FILL
XFILL_1__15287_ gnd vdd FILL
XFILL_6__16027_ gnd vdd FILL
XFILL_1__12499_ gnd vdd FILL
XFILL_6__13239_ gnd vdd FILL
XFILL_0__9535_ gnd vdd FILL
XFILL_4__14418_ gnd vdd FILL
X_8074_ _8074_/A _8142_/A _8074_/C gnd _8156_/D vdd OAI21X1
XSFILL3560x5050 gnd vdd FILL
XFILL_4__15398_ gnd vdd FILL
XSFILL69240x62050 gnd vdd FILL
XFILL_1__14238_ gnd vdd FILL
XFILL_3__9244_ gnd vdd FILL
XSFILL33880x39050 gnd vdd FILL
XFILL_5__13969_ gnd vdd FILL
XFILL_2__13789_ gnd vdd FILL
XFILL_5__15708_ gnd vdd FILL
XFILL_0__14968_ gnd vdd FILL
X_7025_ _7025_/Q _8433_/CLK _7921_/R vdd _7025_/D gnd vdd DFFSR
XFILL_4__14349_ gnd vdd FILL
XFILL_0__9466_ gnd vdd FILL
XFILL_2__15528_ gnd vdd FILL
XFILL_1__14169_ gnd vdd FILL
XSFILL104440x71050 gnd vdd FILL
XFILL_0__13919_ gnd vdd FILL
XFILL_0__14899_ gnd vdd FILL
XFILL_1__7210_ gnd vdd FILL
XFILL_5__15639_ gnd vdd FILL
XFILL_1__8190_ gnd vdd FILL
XFILL_3__8126_ gnd vdd FILL
XFILL_0__9397_ gnd vdd FILL
XFILL_2__15459_ gnd vdd FILL
XFILL_4__16019_ gnd vdd FILL
XFILL_0__8348_ gnd vdd FILL
X_8976_ _8976_/A _8969_/A _8975_/Y gnd _9054_/D vdd OAI21X1
XFILL_3__8057_ gnd vdd FILL
XFILL_6__9855_ gnd vdd FILL
XSFILL3640x16050 gnd vdd FILL
XFILL_1__7072_ gnd vdd FILL
X_7927_ _8951_/A _7972_/A gnd _7928_/C vdd NAND2X1
XFILL_4__8870_ gnd vdd FILL
XSFILL28840x28050 gnd vdd FILL
XFILL_0_CLKBUF1_insert203 gnd vdd FILL
X_7858_ _7914_/Q gnd _7860_/A vdd INVX1
XFILL_4__7821_ gnd vdd FILL
XFILL_0_CLKBUF1_insert214 gnd vdd FILL
XSFILL13640x70050 gnd vdd FILL
XSFILL54280x20050 gnd vdd FILL
X_7789_ _7739_/A _8051_/CLK _7789_/R vdd _7789_/D gnd vdd DFFSR
XFILL_3__8959_ gnd vdd FILL
XFILL_1_BUFX2_insert1007 gnd vdd FILL
XFILL_4__7752_ gnd vdd FILL
XSFILL69320x42050 gnd vdd FILL
XFILL_1_BUFX2_insert1018 gnd vdd FILL
XSFILL33960x19050 gnd vdd FILL
XFILL_1_BUFX2_insert1029 gnd vdd FILL
X_9528_ _9580_/Q gnd _9530_/A vdd INVX1
XFILL_1__7974_ gnd vdd FILL
X_10410_ _10395_/A _9258_/B gnd _10411_/C vdd NAND2X1
XFILL_4__7683_ gnd vdd FILL
X_11390_ _11379_/Y _11385_/Y _11390_/C gnd _11623_/A vdd AOI21X1
XFILL_1__6925_ gnd vdd FILL
X_9459_ _9459_/Q _9453_/CLK _9453_/R vdd _9459_/D gnd vdd DFFSR
XFILL_6__8599_ gnd vdd FILL
XFILL_4__9422_ gnd vdd FILL
XSFILL104520x51050 gnd vdd FILL
X_10341_ _10341_/Q _7781_/CLK _8670_/R vdd _10277_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert710 gnd vdd FILL
XFILL_4_BUFX2_insert721 gnd vdd FILL
XFILL_1__9644_ gnd vdd FILL
XFILL_4_BUFX2_insert732 gnd vdd FILL
XFILL_1__6856_ gnd vdd FILL
XFILL_4__9353_ gnd vdd FILL
XFILL_4_BUFX2_insert743 gnd vdd FILL
X_13060_ _6883_/A _9823_/CLK _9056_/R vdd _13060_/D gnd vdd DFFSR
X_10272_ _14135_/C gnd _10272_/Y vdd INVX1
XFILL_4_BUFX2_insert754 gnd vdd FILL
XFILL_4_BUFX2_insert765 gnd vdd FILL
XFILL_3_CLKBUF1_insert1075 gnd vdd FILL
XFILL_4_BUFX2_insert776 gnd vdd FILL
X_12011_ _12047_/A _12361_/A _12011_/C gnd _12014_/A vdd NAND3X1
XFILL_4_BUFX2_insert787 gnd vdd FILL
XFILL_4__9284_ gnd vdd FILL
XFILL_4_BUFX2_insert798 gnd vdd FILL
XFILL_1__8526_ gnd vdd FILL
XFILL_4__8235_ gnd vdd FILL
XFILL_1__8457_ gnd vdd FILL
XSFILL13720x50050 gnd vdd FILL
XFILL_2__7250_ gnd vdd FILL
XSFILL79960x64050 gnd vdd FILL
XSFILL79160x45050 gnd vdd FILL
X_13962_ _8340_/A _14414_/B _14926_/C _7008_/Q gnd _13963_/B vdd AOI22X1
XFILL_2__7181_ gnd vdd FILL
XFILL_4__7117_ gnd vdd FILL
XFILL_1__8388_ gnd vdd FILL
X_15701_ _14240_/D _15656_/B _15656_/C gnd _15702_/B vdd NOR3X1
XFILL_4__8097_ gnd vdd FILL
X_12913_ _12949_/Q gnd _12913_/Y vdd INVX1
XFILL_1__7339_ gnd vdd FILL
X_13893_ _13891_/Y _14441_/B _14377_/B _15436_/C gnd _13893_/Y vdd OAI22X1
XFILL_4__7048_ gnd vdd FILL
XFILL_5__7930_ gnd vdd FILL
X_15632_ _15632_/A _14164_/D _15632_/C gnd _15634_/A vdd OAI21X1
X_12844_ _12844_/A gnd _12844_/Y vdd INVX1
XFILL_1_BUFX2_insert600 gnd vdd FILL
XFILL_4__10030_ gnd vdd FILL
XFILL_1_BUFX2_insert611 gnd vdd FILL
XFILL_1_BUFX2_insert622 gnd vdd FILL
XFILL_3__10760_ gnd vdd FILL
XFILL_1_BUFX2_insert633 gnd vdd FILL
XFILL_5__7861_ gnd vdd FILL
XFILL_5__11320_ gnd vdd FILL
XFILL_0__10580_ gnd vdd FILL
XFILL_1_BUFX2_insert644 gnd vdd FILL
X_15563_ _15563_/A _14039_/Y _15563_/C _14061_/A gnd _15564_/B vdd OAI22X1
XFILL_1__9009_ gnd vdd FILL
X_12775_ _12773_/Y _12789_/A _12775_/C gnd _12817_/D vdd OAI21X1
XSFILL99320x58050 gnd vdd FILL
XFILL_1_BUFX2_insert655 gnd vdd FILL
XFILL_2__11140_ gnd vdd FILL
XSFILL59080x12050 gnd vdd FILL
XFILL_5__9600_ gnd vdd FILL
XFILL_1_BUFX2_insert666 gnd vdd FILL
XFILL_1_BUFX2_insert677 gnd vdd FILL
XFILL_1__11870_ gnd vdd FILL
XFILL_3__10691_ gnd vdd FILL
X_14514_ _8888_/A gnd _14515_/A vdd INVX1
XFILL_4__8999_ gnd vdd FILL
XFILL_1_BUFX2_insert688 gnd vdd FILL
X_11726_ _11720_/A _11726_/B _11725_/Y gnd _11726_/Y vdd OAI21X1
XFILL_5__11251_ gnd vdd FILL
XFILL_3__12430_ gnd vdd FILL
XFILL_1_BUFX2_insert699 gnd vdd FILL
X_15494_ _15490_/Y _15494_/B gnd _15495_/B vdd NOR2X1
XFILL_4__11981_ gnd vdd FILL
XFILL_1__10821_ gnd vdd FILL
XFILL_2__11071_ gnd vdd FILL
XFILL_5__9531_ gnd vdd FILL
XFILL_0__12250_ gnd vdd FILL
XFILL112280x18050 gnd vdd FILL
XFILL_4__13720_ gnd vdd FILL
X_14445_ _14445_/A _14444_/Y gnd _14445_/Y vdd NOR2X1
XFILL_4__10932_ gnd vdd FILL
XFILL_2__10022_ gnd vdd FILL
X_11657_ _11059_/Y _11656_/Y gnd _11657_/Y vdd NOR2X1
XFILL_5__11182_ gnd vdd FILL
XFILL_3__12361_ gnd vdd FILL
XFILL_2__9753_ gnd vdd FILL
XFILL_1__13540_ gnd vdd FILL
XFILL_0__11201_ gnd vdd FILL
XFILL_1__10752_ gnd vdd FILL
XFILL_2__6965_ gnd vdd FILL
XFILL_5__9462_ gnd vdd FILL
XFILL_0__12181_ gnd vdd FILL
X_10608_ _10608_/Q _8289_/CLK _7152_/R vdd _10566_/Y gnd vdd DFFSR
XSFILL13800x30050 gnd vdd FILL
XFILL_5__10133_ gnd vdd FILL
XFILL_3__14100_ gnd vdd FILL
XFILL_6__15260_ gnd vdd FILL
XFILL_2__8704_ gnd vdd FILL
XFILL_4__13651_ gnd vdd FILL
X_14376_ _10159_/A gnd _14376_/Y vdd INVX1
XFILL_3__11312_ gnd vdd FILL
XFILL_5__15990_ gnd vdd FILL
XFILL_2__14830_ gnd vdd FILL
X_11588_ _11146_/B _11588_/B _11587_/Y gnd _11589_/B vdd NAND3X1
XFILL_3__15080_ gnd vdd FILL
XFILL_1__13471_ gnd vdd FILL
XFILL_2__9684_ gnd vdd FILL
XFILL_3__12292_ gnd vdd FILL
XFILL_0__11132_ gnd vdd FILL
XSFILL79240x25050 gnd vdd FILL
XFILL_1__10683_ gnd vdd FILL
XFILL_6__14211_ gnd vdd FILL
XFILL_2__6896_ gnd vdd FILL
X_16115_ _16114_/Y _15958_/B _15010_/A _14700_/B gnd _16115_/Y vdd OAI22X1
XFILL_4__12602_ gnd vdd FILL
X_13327_ _13241_/Y _13274_/A gnd _13327_/Y vdd AND2X2
XFILL_5__9393_ gnd vdd FILL
XFILL_4__16370_ gnd vdd FILL
X_10539_ _10537_/Y _10539_/B _10538_/Y gnd _10599_/D vdd OAI21X1
XFILL_3__14031_ gnd vdd FILL
XFILL_5__14941_ gnd vdd FILL
XFILL_5__10064_ gnd vdd FILL
XFILL_2__8635_ gnd vdd FILL
XFILL_1__12422_ gnd vdd FILL
XFILL_1__15210_ gnd vdd FILL
XFILL_4__13582_ gnd vdd FILL
XFILL_3__11243_ gnd vdd FILL
XFILL_1__16190_ gnd vdd FILL
XFILL_2__14761_ gnd vdd FILL
XFILL_4__10794_ gnd vdd FILL
XFILL_2__11973_ gnd vdd FILL
XFILL_0__15940_ gnd vdd FILL
XFILL_5__8344_ gnd vdd FILL
XFILL_0__11063_ gnd vdd FILL
X_16046_ _16046_/A _16046_/B _14265_/C gnd _12896_/B vdd AOI21X1
XFILL_4__15321_ gnd vdd FILL
XFILL_6__11354_ gnd vdd FILL
X_13258_ _13281_/B _13337_/A _13270_/A gnd _13258_/Y vdd OAI21X1
XFILL_4__12533_ gnd vdd FILL
XFILL_5__14872_ gnd vdd FILL
XFILL_2__13712_ gnd vdd FILL
XFILL_1__15141_ gnd vdd FILL
XFILL_3__11174_ gnd vdd FILL
XFILL_1__12353_ gnd vdd FILL
XFILL_2__10924_ gnd vdd FILL
XFILL_2__8566_ gnd vdd FILL
XFILL_0__10014_ gnd vdd FILL
XFILL_6__10305_ gnd vdd FILL
XFILL_2__14692_ gnd vdd FILL
XSFILL84360x16050 gnd vdd FILL
XFILL_6__14073_ gnd vdd FILL
X_12209_ _12117_/B _12950_/Q gnd _12210_/C vdd NAND2X1
XFILL_5__8275_ gnd vdd FILL
XFILL_0__15871_ gnd vdd FILL
XFILL_5__13823_ gnd vdd FILL
XFILL_3__10125_ gnd vdd FILL
XFILL_4__15252_ gnd vdd FILL
XFILL_0__7581_ gnd vdd FILL
XFILL_4__12464_ gnd vdd FILL
X_13189_ _11929_/A _12537_/CLK _12536_/R vdd _13123_/Y gnd vdd DFFSR
XFILL_1__11304_ gnd vdd FILL
XFILL_3__15982_ gnd vdd FILL
XFILL_2__13643_ gnd vdd FILL
XFILL_1__15072_ gnd vdd FILL
XFILL_0__14822_ gnd vdd FILL
XFILL_5__7226_ gnd vdd FILL
XFILL_2__8497_ gnd vdd FILL
XFILL_1__12284_ gnd vdd FILL
XFILL_3__7290_ gnd vdd FILL
XFILL_4__14203_ gnd vdd FILL
XSFILL99400x38050 gnd vdd FILL
XFILL_4__11415_ gnd vdd FILL
XFILL_5__10966_ gnd vdd FILL
XFILL_4__15183_ gnd vdd FILL
XFILL_5__13754_ gnd vdd FILL
XFILL_1__14023_ gnd vdd FILL
XFILL_3__10056_ gnd vdd FILL
XFILL_3__14933_ gnd vdd FILL
XFILL_2__7448_ gnd vdd FILL
XFILL_4__12395_ gnd vdd FILL
XFILL_2__16362_ gnd vdd FILL
XFILL_1__11235_ gnd vdd FILL
XSFILL84200x80050 gnd vdd FILL
XFILL_2_CLKBUF1_insert180 gnd vdd FILL
XFILL_2__10786_ gnd vdd FILL
XFILL_0__14753_ gnd vdd FILL
XFILL_2__13574_ gnd vdd FILL
XFILL_2_CLKBUF1_insert191 gnd vdd FILL
XFILL_0__11965_ gnd vdd FILL
XFILL_5__12705_ gnd vdd FILL
XFILL_0__9251_ gnd vdd FILL
XFILL_4__14134_ gnd vdd FILL
XFILL_5__13685_ gnd vdd FILL
XFILL_2__15313_ gnd vdd FILL
XFILL_4__11346_ gnd vdd FILL
XFILL_3__14864_ gnd vdd FILL
XFILL_5__10897_ gnd vdd FILL
XFILL_2__12525_ gnd vdd FILL
XFILL_0__13704_ gnd vdd FILL
XFILL_0__10916_ gnd vdd FILL
XFILL_2__16293_ gnd vdd FILL
XFILL_2__7379_ gnd vdd FILL
XFILL_1__11166_ gnd vdd FILL
XFILL_0__8202_ gnd vdd FILL
XFILL_0__14684_ gnd vdd FILL
XFILL_5__12636_ gnd vdd FILL
XSFILL74280x68050 gnd vdd FILL
XFILL_0__11896_ gnd vdd FILL
XFILL_5__7088_ gnd vdd FILL
XFILL_5__15424_ gnd vdd FILL
XFILL_3__13815_ gnd vdd FILL
XFILL_4__14065_ gnd vdd FILL
XFILL_2__9118_ gnd vdd FILL
X_8830_ _8830_/A _8916_/A _8829_/Y gnd _8830_/Y vdd OAI21X1
XFILL_2__15244_ gnd vdd FILL
XFILL_1__10117_ gnd vdd FILL
XFILL_4__11277_ gnd vdd FILL
XSFILL109400x23050 gnd vdd FILL
XFILL_0__13635_ gnd vdd FILL
XFILL_3__14795_ gnd vdd FILL
XBUFX2_insert2 _12381_/Y gnd _7579_/B vdd BUFX2
XFILL_2__12456_ gnd vdd FILL
XFILL_1__15974_ gnd vdd FILL
XFILL_1__11097_ gnd vdd FILL
XFILL_4__13016_ gnd vdd FILL
XFILL_0__8133_ gnd vdd FILL
XFILL_5__12567_ gnd vdd FILL
XFILL_5__15355_ gnd vdd FILL
X_8761_ _8714_/B _8889_/B gnd _8762_/C vdd NAND2X1
XSFILL49080x44050 gnd vdd FILL
XFILL112200x62050 gnd vdd FILL
XFILL_3__13746_ gnd vdd FILL
XFILL_3__9931_ gnd vdd FILL
XFILL_2__11407_ gnd vdd FILL
XFILL_3__10958_ gnd vdd FILL
XFILL_2__15175_ gnd vdd FILL
XFILL_1__10048_ gnd vdd FILL
XFILL_2__12387_ gnd vdd FILL
XFILL_0__16354_ gnd vdd FILL
XFILL_1__14925_ gnd vdd FILL
XFILL_0__13566_ gnd vdd FILL
XFILL_0__8064_ gnd vdd FILL
X_7712_ _7780_/Q gnd _7714_/A vdd INVX1
XFILL_0__10778_ gnd vdd FILL
XFILL_5__11518_ gnd vdd FILL
XFILL_5__14306_ gnd vdd FILL
XFILL_6_BUFX2_insert827 gnd vdd FILL
XFILL_5__15286_ gnd vdd FILL
XFILL_6_BUFX2_insert838 gnd vdd FILL
XFILL_0__15305_ gnd vdd FILL
XFILL_2__14126_ gnd vdd FILL
XFILL_5__12498_ gnd vdd FILL
XFILL_4__10159_ gnd vdd FILL
X_8692_ _8656_/A _9578_/CLK _9460_/R vdd _8658_/Y gnd vdd DFFSR
XFILL_3__13677_ gnd vdd FILL
XFILL_0__12517_ gnd vdd FILL
XFILL_3__9862_ gnd vdd FILL
XFILL_2__11338_ gnd vdd FILL
XFILL_1__14856_ gnd vdd FILL
XFILL_0__16285_ gnd vdd FILL
XFILL_3__10889_ gnd vdd FILL
XSFILL4440x59050 gnd vdd FILL
XFILL_0__13497_ gnd vdd FILL
XFILL_5__14237_ gnd vdd FILL
XSFILL43800x46050 gnd vdd FILL
XSFILL115240x7050 gnd vdd FILL
XFILL_5__11449_ gnd vdd FILL
XFILL_3__15416_ gnd vdd FILL
X_7643_ _7643_/Q _7143_/CLK _7015_/R vdd _7643_/D gnd vdd DFFSR
XFILL_3__12628_ gnd vdd FILL
XFILL_1__13807_ gnd vdd FILL
XFILL_0__15236_ gnd vdd FILL
XFILL_2__14057_ gnd vdd FILL
XFILL_4__14967_ gnd vdd FILL
XFILL_3__16396_ gnd vdd FILL
XFILL_2__11269_ gnd vdd FILL
XFILL_0__12448_ gnd vdd FILL
XFILL_3__9793_ gnd vdd FILL
XFILL_5__9729_ gnd vdd FILL
XFILL_1__11999_ gnd vdd FILL
XFILL_1__14787_ gnd vdd FILL
XFILL_5__14168_ gnd vdd FILL
XFILL_3__15347_ gnd vdd FILL
XFILL_2__13008_ gnd vdd FILL
X_7574_ _7572_/Y _7570_/A _7574_/C gnd _7574_/Y vdd OAI21X1
XFILL_4__13918_ gnd vdd FILL
XFILL_3__8744_ gnd vdd FILL
XSFILL69240x57050 gnd vdd FILL
XFILL_4__14898_ gnd vdd FILL
XFILL_0__15167_ gnd vdd FILL
XFILL_1__13738_ gnd vdd FILL
X_9313_ _9313_/Q _8560_/CLK _9313_/R vdd _9313_/D gnd vdd DFFSR
XFILL_0__12379_ gnd vdd FILL
XFILL_5__13119_ gnd vdd FILL
XFILL_5__14099_ gnd vdd FILL
XFILL_0__8966_ gnd vdd FILL
XFILL_4__13849_ gnd vdd FILL
XFILL_0__14118_ gnd vdd FILL
XFILL_3__15278_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1081 gnd vdd FILL
XSFILL104440x66050 gnd vdd FILL
XFILL_1__13669_ gnd vdd FILL
XFILL_0__15098_ gnd vdd FILL
X_9244_ _9244_/A _9208_/B _9243_/Y gnd _9314_/D vdd OAI21X1
XFILL_3__14229_ gnd vdd FILL
XFILL_1__7690_ gnd vdd FILL
XFILL_1__15408_ gnd vdd FILL
XSFILL8680x64050 gnd vdd FILL
XFILL_3__7626_ gnd vdd FILL
XFILL_0__8897_ gnd vdd FILL
XFILL_0__14049_ gnd vdd FILL
XFILL_2__14959_ gnd vdd FILL
XFILL_1__16388_ gnd vdd FILL
XFILL_0__7848_ gnd vdd FILL
XFILL_4__15519_ gnd vdd FILL
X_9175_ _9175_/Q _8551_/CLK _9959_/R vdd _9083_/Y gnd vdd DFFSR
XFILL_1__15339_ gnd vdd FILL
XFILL_3__7557_ gnd vdd FILL
X_8126_ _8126_/A gnd _8128_/A vdd INVX1
XFILL_3_BUFX2_insert706 gnd vdd FILL
XFILL_1__9360_ gnd vdd FILL
XFILL_3_BUFX2_insert717 gnd vdd FILL
XFILL_3_BUFX2_insert728 gnd vdd FILL
XFILL_3_BUFX2_insert739 gnd vdd FILL
XFILL_3__7488_ gnd vdd FILL
XFILL_1__8311_ gnd vdd FILL
XFILL_0__9518_ gnd vdd FILL
XSFILL94440x6050 gnd vdd FILL
X_8057_ _8057_/A gnd _8057_/Y vdd INVX1
XFILL_3__9227_ gnd vdd FILL
XFILL_1__9291_ gnd vdd FILL
XFILL_4__8020_ gnd vdd FILL
XFILL_1_BUFX2_insert50 gnd vdd FILL
XFILL_1_BUFX2_insert61 gnd vdd FILL
X_7008_ _7008_/Q _7791_/CLK _7648_/R vdd _7008_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert72 gnd vdd FILL
XFILL_1__8242_ gnd vdd FILL
XFILL_1_BUFX2_insert83 gnd vdd FILL
XFILL_3__9158_ gnd vdd FILL
XFILL_1_BUFX2_insert94 gnd vdd FILL
XSFILL39080x76050 gnd vdd FILL
XFILL_3__8109_ gnd vdd FILL
XFILL_3__9089_ gnd vdd FILL
XFILL_1__7124_ gnd vdd FILL
X_10890_ _10963_/A gnd _10890_/Y vdd INVX1
X_8959_ _8959_/A gnd _8961_/A vdd INVX1
XFILL_1__7055_ gnd vdd FILL
XSFILL33800x78050 gnd vdd FILL
XFILL_4__8853_ gnd vdd FILL
X_12560_ _12418_/A _13201_/CLK _13201_/R vdd _12516_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert607 gnd vdd FILL
XFILL_4__7804_ gnd vdd FILL
XFILL_0_BUFX2_insert618 gnd vdd FILL
XFILL_0_BUFX2_insert629 gnd vdd FILL
XSFILL104360x8050 gnd vdd FILL
X_11511_ _11511_/A _11846_/C _11510_/Y gnd _11514_/C vdd AOI21X1
XFILL_4__8784_ gnd vdd FILL
X_12491_ vdd _12057_/A gnd _12491_/Y vdd NAND2X1
XFILL_4__7735_ gnd vdd FILL
X_14230_ _13614_/C _14228_/Y _13882_/B _14229_/Y gnd _14234_/A vdd OAI22X1
X_11442_ _12242_/Y _12135_/Y gnd _11776_/A vdd XNOR2X1
XFILL_1__7957_ gnd vdd FILL
XSFILL13720x45050 gnd vdd FILL
X_14161_ _14157_/Y _14161_/B gnd _14169_/A vdd NOR2X1
X_11373_ _12218_/Y gnd _11373_/Y vdd INVX1
XFILL_1__6908_ gnd vdd FILL
XFILL_4__9405_ gnd vdd FILL
XSFILL54600x57050 gnd vdd FILL
XFILL_1__7888_ gnd vdd FILL
X_13112_ _13186_/Q gnd _13114_/A vdd INVX1
X_10324_ _10325_/B _9172_/B gnd _10324_/Y vdd NAND2X1
XFILL_4__7597_ gnd vdd FILL
XFILL_4_BUFX2_insert540 gnd vdd FILL
XFILL_1__9627_ gnd vdd FILL
XFILL_4_BUFX2_insert551 gnd vdd FILL
X_14092_ _14092_/A _14092_/B gnd _14092_/Y vdd NOR2X1
XFILL_4_BUFX2_insert562 gnd vdd FILL
XFILL_1__6839_ gnd vdd FILL
XFILL_4__9336_ gnd vdd FILL
XFILL_4_BUFX2_insert573 gnd vdd FILL
X_10255_ _10304_/B _8719_/B gnd _10256_/C vdd NAND2X1
XFILL_4_BUFX2_insert584 gnd vdd FILL
X_13043_ _13041_/Y vdd _13042_/Y gnd _13077_/D vdd OAI21X1
XFILL_4_BUFX2_insert595 gnd vdd FILL
XFILL_2__8351_ gnd vdd FILL
XFILL_4__9267_ gnd vdd FILL
XFILL_5__8060_ gnd vdd FILL
XFILL_5__10820_ gnd vdd FILL
XFILL_1__8509_ gnd vdd FILL
X_10186_ _10186_/A gnd _10188_/A vdd INVX1
XFILL_2__7302_ gnd vdd FILL
XFILL_2__10640_ gnd vdd FILL
XFILL_4__8218_ gnd vdd FILL
XFILL_1__9489_ gnd vdd FILL
XFILL_6__10021_ gnd vdd FILL
XSFILL58840x62050 gnd vdd FILL
XSFILL99480x12050 gnd vdd FILL
XFILL_4__11200_ gnd vdd FILL
XFILL_5__10751_ gnd vdd FILL
XSFILL74120x10050 gnd vdd FILL
XFILL_4__12180_ gnd vdd FILL
X_14994_ _14994_/A _14987_/Y gnd _15008_/C vdd NOR2X1
XFILL_3__11930_ gnd vdd FILL
XFILL_2__7233_ gnd vdd FILL
XFILL_1__11020_ gnd vdd FILL
XFILL_2__10571_ gnd vdd FILL
XFILL_4__8149_ gnd vdd FILL
XFILL_0__11750_ gnd vdd FILL
XFILL_5__13470_ gnd vdd FILL
XFILL_3_CLKBUF1_insert220 gnd vdd FILL
XFILL_4__11131_ gnd vdd FILL
X_13945_ _13944_/Y _13587_/C _14456_/C _15479_/D gnd _13949_/A vdd OAI22X1
XFILL_5__10682_ gnd vdd FILL
XFILL_2__12310_ gnd vdd FILL
XFILL_2__13290_ gnd vdd FILL
XFILL_0__10701_ gnd vdd FILL
XFILL_3__11861_ gnd vdd FILL
XFILL_2__7164_ gnd vdd FILL
XSFILL43880x8050 gnd vdd FILL
XFILL_5__8962_ gnd vdd FILL
XFILL_5__12421_ gnd vdd FILL
XSFILL109320x38050 gnd vdd FILL
XFILL_0__11681_ gnd vdd FILL
XFILL_3__13600_ gnd vdd FILL
XSFILL63960x53050 gnd vdd FILL
XSFILL13800x25050 gnd vdd FILL
XFILL_3__10812_ gnd vdd FILL
X_13876_ _13875_/Y _13876_/B _13876_/C _13874_/Y gnd _13876_/Y vdd OAI22X1
XFILL_2__12241_ gnd vdd FILL
XFILL_4__11062_ gnd vdd FILL
XFILL_2__7095_ gnd vdd FILL
XFILL_3__14580_ gnd vdd FILL
XFILL_0__13420_ gnd vdd FILL
XFILL_0__10632_ gnd vdd FILL
XFILL_3__11792_ gnd vdd FILL
X_15615_ _15615_/A _15615_/B gnd _15618_/C vdd NOR2X1
XFILL_1__12971_ gnd vdd FILL
XFILL_5__15140_ gnd vdd FILL
XFILL_5__12352_ gnd vdd FILL
XFILL_5__8893_ gnd vdd FILL
XFILL_4__10013_ gnd vdd FILL
XFILL_1_BUFX2_insert430 gnd vdd FILL
X_12827_ vdd _15127_/Y gnd _12827_/Y vdd NAND2X1
XFILL_1_BUFX2_insert441 gnd vdd FILL
XFILL_3__13531_ gnd vdd FILL
XFILL_3__10743_ gnd vdd FILL
XFILL_2__12172_ gnd vdd FILL
XFILL_1__14710_ gnd vdd FILL
XFILL_1_BUFX2_insert452 gnd vdd FILL
XFILL_4__15870_ gnd vdd FILL
XFILL_0__13351_ gnd vdd FILL
XFILL_1__11922_ gnd vdd FILL
XFILL_5__7844_ gnd vdd FILL
XFILL_1__15690_ gnd vdd FILL
XFILL_1_BUFX2_insert463 gnd vdd FILL
XFILL_5__11303_ gnd vdd FILL
XFILL_0__10563_ gnd vdd FILL
XFILL_5__15071_ gnd vdd FILL
X_15546_ _8418_/Q _15978_/B _16014_/C _8290_/Q gnd _15546_/Y vdd AOI22X1
XSFILL114440x29050 gnd vdd FILL
XFILL_1_BUFX2_insert474 gnd vdd FILL
X_12758_ _12812_/Q gnd _12758_/Y vdd INVX1
XFILL_4__14821_ gnd vdd FILL
XFILL_2__11123_ gnd vdd FILL
XFILL_1_BUFX2_insert485 gnd vdd FILL
XFILL_3__16250_ gnd vdd FILL
XFILL_5__12283_ gnd vdd FILL
XFILL_1_BUFX2_insert496 gnd vdd FILL
XFILL_3__13462_ gnd vdd FILL
XFILL_0__12302_ gnd vdd FILL
XFILL_1__14641_ gnd vdd FILL
XFILL_0__16070_ gnd vdd FILL
XFILL_3__10674_ gnd vdd FILL
XFILL_1__11853_ gnd vdd FILL
XFILL_0__13282_ gnd vdd FILL
XFILL_5__14022_ gnd vdd FILL
XFILL_3__15201_ gnd vdd FILL
X_11709_ _11709_/A _11681_/B _11764_/A _11054_/A gnd _11710_/B vdd AOI22X1
XFILL_0__10494_ gnd vdd FILL
XFILL_5__11234_ gnd vdd FILL
XFILL_2__9805_ gnd vdd FILL
XFILL_3__12413_ gnd vdd FILL
XFILL_4__14752_ gnd vdd FILL
X_15477_ _13972_/A _15175_/B _15477_/C gnd _15477_/Y vdd AOI21X1
X_12689_ _12645_/A _12667_/CLK _12689_/R vdd _12689_/D gnd vdd DFFSR
XFILL_3__16181_ gnd vdd FILL
XFILL_0__15021_ gnd vdd FILL
XFILL_2__15931_ gnd vdd FILL
XFILL_4__11964_ gnd vdd FILL
XFILL_2__11054_ gnd vdd FILL
XSFILL43880x20050 gnd vdd FILL
XFILL_3__13393_ gnd vdd FILL
XFILL_0__12233_ gnd vdd FILL
XBUFX2_insert1009 _10928_/Y gnd _12248_/A vdd BUFX2
XFILL_5__9514_ gnd vdd FILL
XFILL_1__10804_ gnd vdd FILL
XFILL_1__14572_ gnd vdd FILL
XFILL_2__7997_ gnd vdd FILL
XFILL_1__11784_ gnd vdd FILL
X_14428_ _8042_/Q gnd _15879_/D vdd INVX1
XFILL_4__10915_ gnd vdd FILL
XFILL_5__11165_ gnd vdd FILL
XFILL_4__13703_ gnd vdd FILL
XFILL_2__10005_ gnd vdd FILL
XFILL_3__15132_ gnd vdd FILL
XFILL_3__12344_ gnd vdd FILL
XFILL_2__9736_ gnd vdd FILL
XFILL_1__16311_ gnd vdd FILL
XFILL_4__14683_ gnd vdd FILL
XFILL_2__6948_ gnd vdd FILL
XFILL_4__11895_ gnd vdd FILL
XFILL_1__13523_ gnd vdd FILL
XFILL_2__15862_ gnd vdd FILL
XFILL_0__12164_ gnd vdd FILL
XSFILL84200x75050 gnd vdd FILL
XFILL_5__10116_ gnd vdd FILL
XFILL_4__13634_ gnd vdd FILL
X_14359_ _15826_/A _14344_/B _13621_/B _14359_/D gnd _14367_/B vdd AOI22X1
XFILL_0__8751_ gnd vdd FILL
XFILL_5__15973_ gnd vdd FILL
XFILL_2__14813_ gnd vdd FILL
XFILL_3__15063_ gnd vdd FILL
XFILL_5__11096_ gnd vdd FILL
X_7290_ _7323_/A _9082_/B gnd _7290_/Y vdd NAND2X1
XFILL_1__16242_ gnd vdd FILL
XFILL_3__8460_ gnd vdd FILL
XFILL_1__13454_ gnd vdd FILL
XFILL_3__12275_ gnd vdd FILL
XFILL_2__9667_ gnd vdd FILL
XSFILL49560x8050 gnd vdd FILL
XFILL_0__11115_ gnd vdd FILL
XFILL_2__15793_ gnd vdd FILL
XFILL_1__10666_ gnd vdd FILL
XFILL_2__6879_ gnd vdd FILL
XFILL_5__9376_ gnd vdd FILL
XSFILL59000x51050 gnd vdd FILL
XFILL_0__12095_ gnd vdd FILL
XFILL_0__7702_ gnd vdd FILL
XFILL_5__10047_ gnd vdd FILL
XFILL_3__14014_ gnd vdd FILL
XFILL_5__14924_ gnd vdd FILL
XFILL_4__16353_ gnd vdd FILL
XFILL_4__13565_ gnd vdd FILL
XFILL_2__8618_ gnd vdd FILL
XFILL_3__11226_ gnd vdd FILL
XFILL_1__12405_ gnd vdd FILL
XFILL_4__10777_ gnd vdd FILL
XSFILL109400x18050 gnd vdd FILL
XFILL_2__14744_ gnd vdd FILL
XFILL_0__15923_ gnd vdd FILL
XFILL_1__16173_ gnd vdd FILL
XFILL_2__11956_ gnd vdd FILL
XFILL_1__13385_ gnd vdd FILL
XFILL_2__9598_ gnd vdd FILL
XFILL_5__8327_ gnd vdd FILL
XFILL_0__11046_ gnd vdd FILL
XFILL_6__7120_ gnd vdd FILL
XFILL_3__8391_ gnd vdd FILL
X_16029_ _9454_/Q _15202_/B _16037_/C gnd _16029_/Y vdd NAND3X1
XFILL_4__15304_ gnd vdd FILL
XFILL_4__12516_ gnd vdd FILL
XFILL_0__7633_ gnd vdd FILL
XFILL_5__14855_ gnd vdd FILL
XFILL_4__16284_ gnd vdd FILL
XFILL_2__10907_ gnd vdd FILL
XFILL112200x57050 gnd vdd FILL
XFILL_3__7342_ gnd vdd FILL
XFILL_1__12336_ gnd vdd FILL
XFILL_4__13496_ gnd vdd FILL
XFILL_3__11157_ gnd vdd FILL
XFILL_1__15124_ gnd vdd FILL
XFILL_2__14675_ gnd vdd FILL
XFILL_2__11887_ gnd vdd FILL
XFILL_0__15854_ gnd vdd FILL
XSFILL89480x44050 gnd vdd FILL
XFILL_5__8258_ gnd vdd FILL
XFILL_5__13806_ gnd vdd FILL
XFILL_4__15235_ gnd vdd FILL
XFILL_0__7564_ gnd vdd FILL
XFILL_4__12447_ gnd vdd FILL
XSFILL64120x42050 gnd vdd FILL
XFILL_2__16414_ gnd vdd FILL
XFILL_3__10108_ gnd vdd FILL
XFILL_2__13626_ gnd vdd FILL
XFILL_5__14786_ gnd vdd FILL
XFILL_0__14805_ gnd vdd FILL
XFILL_5__11998_ gnd vdd FILL
XFILL_1__15055_ gnd vdd FILL
XFILL_3__15965_ gnd vdd FILL
XFILL_1__12267_ gnd vdd FILL
XFILL_3__11088_ gnd vdd FILL
XFILL_5__7209_ gnd vdd FILL
XFILL_0__12997_ gnd vdd FILL
XFILL_0__15785_ gnd vdd FILL
XFILL_5__8189_ gnd vdd FILL
X_9931_ _9865_/A _9803_/B gnd _9932_/C vdd NAND2X1
XFILL_4__15166_ gnd vdd FILL
XFILL_3__9012_ gnd vdd FILL
XFILL_5__13737_ gnd vdd FILL
XFILL_5__10949_ gnd vdd FILL
XFILL_3__10039_ gnd vdd FILL
XFILL_2__16345_ gnd vdd FILL
XFILL_1__14006_ gnd vdd FILL
XFILL_4__12378_ gnd vdd FILL
XFILL_0__7495_ gnd vdd FILL
XFILL_3__14916_ gnd vdd FILL
XFILL_1__11218_ gnd vdd FILL
XFILL_3__15896_ gnd vdd FILL
XFILL_2__13557_ gnd vdd FILL
XFILL_0__11948_ gnd vdd FILL
XFILL_0__14736_ gnd vdd FILL
XFILL_1__12198_ gnd vdd FILL
XFILL_2__10769_ gnd vdd FILL
XFILL_4__14117_ gnd vdd FILL
XFILL_0__9234_ gnd vdd FILL
XFILL_4__11329_ gnd vdd FILL
XFILL_3__14847_ gnd vdd FILL
XFILL_5__13668_ gnd vdd FILL
XFILL_2__12508_ gnd vdd FILL
XFILL_4__15097_ gnd vdd FILL
X_9862_ _9902_/B _8582_/B gnd _9862_/Y vdd NAND2X1
XFILL_1__11149_ gnd vdd FILL
XFILL_2__16276_ gnd vdd FILL
XFILL_2__13488_ gnd vdd FILL
XFILL_0__11879_ gnd vdd FILL
XFILL_5__15407_ gnd vdd FILL
XFILL_0__14667_ gnd vdd FILL
XFILL_6__7953_ gnd vdd FILL
XFILL_5__12619_ gnd vdd FILL
XFILL_0__9165_ gnd vdd FILL
X_8813_ _8813_/Q _7661_/CLK _7533_/R vdd _8765_/Y gnd vdd DFFSR
XFILL_4__14048_ gnd vdd FILL
XFILL_6__14958_ gnd vdd FILL
XFILL_5__16387_ gnd vdd FILL
XFILL_2__15227_ gnd vdd FILL
XSFILL114360x3050 gnd vdd FILL
XFILL_5__13599_ gnd vdd FILL
XFILL_2__12439_ gnd vdd FILL
XFILL_0__16406_ gnd vdd FILL
X_9793_ _9839_/Q gnd _9793_/Y vdd INVX1
XFILL_3__14778_ gnd vdd FILL
XFILL_0__13618_ gnd vdd FILL
XFILL_6__6904_ gnd vdd FILL
XFILL_1__15957_ gnd vdd FILL
XFILL_0__14598_ gnd vdd FILL
XFILL_0__8116_ gnd vdd FILL
XFILL_6_BUFX2_insert602 gnd vdd FILL
XFILL_6__13909_ gnd vdd FILL
XFILL_5__15338_ gnd vdd FILL
XFILL_6_BUFX2_insert613 gnd vdd FILL
X_8744_ _8742_/Y _8714_/B _8744_/C gnd _8744_/Y vdd OAI21X1
XFILL_0__9096_ gnd vdd FILL
XFILL_3__9914_ gnd vdd FILL
XFILL_3__13729_ gnd vdd FILL
XSFILL8680x59050 gnd vdd FILL
XFILL_2__15158_ gnd vdd FILL
XFILL_1__14908_ gnd vdd FILL
XFILL_0__13549_ gnd vdd FILL
XFILL_0__16337_ gnd vdd FILL
XFILL_1__15888_ gnd vdd FILL
XSFILL33880x52050 gnd vdd FILL
X_8675_ _8675_/Q _7530_/CLK _7523_/R vdd _8675_/D gnd vdd DFFSR
XFILL_2__14109_ gnd vdd FILL
XFILL_5__15269_ gnd vdd FILL
XFILL_1__14839_ gnd vdd FILL
XFILL_4__15999_ gnd vdd FILL
XFILL_6_BUFX2_insert679 gnd vdd FILL
XFILL_2__15089_ gnd vdd FILL
XFILL_0__16268_ gnd vdd FILL
XFILL_6__9554_ gnd vdd FILL
X_7626_ _7626_/A gnd _7626_/Y vdd INVX1
XFILL_1__8860_ gnd vdd FILL
XFILL_3__16379_ gnd vdd FILL
XFILL_6__8505_ gnd vdd FILL
XFILL_0__15219_ gnd vdd FILL
XFILL_3__9776_ gnd vdd FILL
XFILL_3__6988_ gnd vdd FILL
XFILL_0__16199_ gnd vdd FILL
XFILL_1__7811_ gnd vdd FILL
X_7557_ _7643_/Q gnd _7557_/Y vdd INVX1
XSFILL108680x66050 gnd vdd FILL
XFILL_3__8727_ gnd vdd FILL
XFILL_0__9998_ gnd vdd FILL
XFILL_1_CLKBUF1_insert117 gnd vdd FILL
XFILL_1_CLKBUF1_insert128 gnd vdd FILL
XSFILL49000x83050 gnd vdd FILL
XFILL_1_CLKBUF1_insert139 gnd vdd FILL
XFILL_1__7742_ gnd vdd FILL
X_7488_ _7486_/Y _7460_/A _7488_/C gnd _7534_/D vdd OAI21X1
XFILL_4__7451_ gnd vdd FILL
XFILL_3__8658_ gnd vdd FILL
XSFILL38680x9050 gnd vdd FILL
X_9227_ _9309_/Q gnd _9227_/Y vdd INVX1
XFILL_3__7609_ gnd vdd FILL
XFILL_1__7673_ gnd vdd FILL
XFILL_3__8589_ gnd vdd FILL
XSFILL28840x41050 gnd vdd FILL
XFILL_1__9412_ gnd vdd FILL
XFILL_3_BUFX2_insert503 gnd vdd FILL
X_9158_ _9158_/A _9112_/A _9158_/C gnd _9200_/D vdd OAI21X1
XFILL_4__9121_ gnd vdd FILL
XFILL_3_BUFX2_insert514 gnd vdd FILL
X_10040_ _15962_/A gnd _10042_/A vdd INVX1
XFILL_3_BUFX2_insert525 gnd vdd FILL
XFILL_3_BUFX2_insert536 gnd vdd FILL
X_8109_ _8100_/A _9517_/B gnd _8110_/C vdd NAND2X1
XFILL_6__7249_ gnd vdd FILL
XFILL_1__9343_ gnd vdd FILL
XFILL_3_BUFX2_insert547 gnd vdd FILL
XFILL_3_BUFX2_insert558 gnd vdd FILL
X_9089_ _9089_/A _9163_/A _9088_/Y gnd _9089_/Y vdd OAI21X1
XSFILL53880x3050 gnd vdd FILL
XFILL_3_BUFX2_insert569 gnd vdd FILL
XSFILL33960x32050 gnd vdd FILL
XFILL_1__9274_ gnd vdd FILL
XFILL_4__8003_ gnd vdd FILL
XSFILL73800x80050 gnd vdd FILL
XFILL_1__8225_ gnd vdd FILL
X_11991_ _12111_/A _11991_/B _12111_/C gnd _11991_/Y vdd NAND3X1
X_13730_ _13728_/Y _14317_/C _14744_/B _13730_/D gnd _13730_/Y vdd OAI22X1
X_10942_ _10941_/Y _10940_/Y gnd _10943_/B vdd NOR2X1
XFILL_6_BUFX2_insert29 gnd vdd FILL
X_13661_ _13659_/Y _13813_/B _13467_/A _15255_/B gnd _13661_/Y vdd OAI22X1
XFILL_1__7107_ gnd vdd FILL
X_10873_ _12701_/A _10873_/B gnd _10874_/B vdd NAND2X1
XFILL_1__8087_ gnd vdd FILL
X_15400_ _7054_/A gnd _15401_/D vdd INVX1
XFILL_4__8905_ gnd vdd FILL
X_12612_ _12612_/A gnd _12614_/A vdd INVX1
XFILL_4__9885_ gnd vdd FILL
X_16380_ _16378_/Y gnd _16379_/Y gnd _16380_/Y vdd OAI21X1
X_13592_ _13592_/A _8191_/A _7039_/A _13592_/D gnd _13595_/A vdd AOI22X1
XFILL_1__7038_ gnd vdd FILL
XSFILL28920x21050 gnd vdd FILL
XFILL_0_BUFX2_insert404 gnd vdd FILL
XFILL_4__8836_ gnd vdd FILL
X_15331_ _15330_/Y _15407_/B _15407_/C _15331_/D gnd _15335_/A vdd OAI22X1
XFILL_0_BUFX2_insert415 gnd vdd FILL
X_12543_ _11912_/B _9050_/CLK _9050_/R vdd _12465_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert426 gnd vdd FILL
XFILL_0_BUFX2_insert437 gnd vdd FILL
XFILL_2__7851_ gnd vdd FILL
XFILL_0_BUFX2_insert448 gnd vdd FILL
XFILL_4__8767_ gnd vdd FILL
XFILL_5__7560_ gnd vdd FILL
XFILL_0_BUFX2_insert459 gnd vdd FILL
XSFILL13640x6050 gnd vdd FILL
X_15262_ _15563_/A _13710_/Y _15563_/C _13704_/D gnd _15264_/B vdd OAI22X1
X_12474_ _12474_/A vdd _12473_/Y gnd _12474_/Y vdd OAI21X1
XFILL_3__10390_ gnd vdd FILL
XFILL_4__7718_ gnd vdd FILL
XFILL_1__8989_ gnd vdd FILL
XSFILL104200x23050 gnd vdd FILL
X_14213_ _14213_/A _9829_/Q _10341_/Q _13621_/B gnd _14215_/A vdd AOI22X1
XFILL_4__10700_ gnd vdd FILL
XFILL_5__7491_ gnd vdd FILL
XFILL_4__8698_ gnd vdd FILL
X_11425_ _11013_/Y _11015_/A gnd _11809_/C vdd NAND2X1
X_15193_ _13597_/Y _15386_/B _15384_/D _13603_/Y gnd _15195_/B vdd OAI22X1
XFILL_2__9521_ gnd vdd FILL
XFILL_1__10520_ gnd vdd FILL
XFILL_4__11680_ gnd vdd FILL
XFILL_5__9230_ gnd vdd FILL
XSFILL18840x73050 gnd vdd FILL
X_14144_ _14144_/A _14144_/B gnd _14171_/B vdd NOR2X1
X_11356_ _11356_/A gnd _12109_/A vdd INVX1
XFILL_4__10631_ gnd vdd FILL
XFILL_3__12060_ gnd vdd FILL
XFILL_5__12970_ gnd vdd FILL
XFILL_2__11810_ gnd vdd FILL
XFILL_1__10451_ gnd vdd FILL
XFILL_2__12790_ gnd vdd FILL
XSFILL108840x26050 gnd vdd FILL
XFILL_5__9161_ gnd vdd FILL
XFILL_4_BUFX2_insert370 gnd vdd FILL
X_10307_ _10305_/Y _10271_/B _10307_/C gnd _10307_/Y vdd OAI21X1
XFILL_4__13350_ gnd vdd FILL
XSFILL99320x71050 gnd vdd FILL
XFILL_4_BUFX2_insert381 gnd vdd FILL
XFILL_5__11921_ gnd vdd FILL
X_14075_ _14074_/Y _14075_/B _15338_/C gnd _12988_/B vdd AOI21X1
XCLKBUF1_insert116 CLKBUF1_insert169/A gnd _9328_/CLK vdd CLKBUF1
XFILL_2__8403_ gnd vdd FILL
XFILL_3__11011_ gnd vdd FILL
XCLKBUF1_insert127 CLKBUF1_insert150/A gnd _7916_/CLK vdd CLKBUF1
X_11287_ _11258_/Y _11281_/Y _11286_/Y gnd _11288_/C vdd OAI21X1
XFILL_4__10562_ gnd vdd FILL
XFILL_2__9383_ gnd vdd FILL
XFILL_4_BUFX2_insert392 gnd vdd FILL
XFILL_1__13170_ gnd vdd FILL
XFILL_5__8112_ gnd vdd FILL
XFILL_2__11741_ gnd vdd FILL
XFILL_1__10382_ gnd vdd FILL
XCLKBUF1_insert138 CLKBUF1_insert220/A gnd _9447_/CLK vdd CLKBUF1
XFILL_5__9092_ gnd vdd FILL
XCLKBUF1_insert149 CLKBUF1_insert216/A gnd _7269_/CLK vdd CLKBUF1
XFILL_4__12301_ gnd vdd FILL
X_13026_ _6895_/A gnd _13026_/Y vdd INVX1
XFILL_5__14640_ gnd vdd FILL
X_10238_ _10236_/Y _10285_/A _10238_/C gnd _10238_/Y vdd OAI21X1
XFILL_4__13281_ gnd vdd FILL
XFILL_2__8334_ gnd vdd FILL
XFILL_1__12121_ gnd vdd FILL
XFILL_5__11852_ gnd vdd FILL
XFILL_2__14460_ gnd vdd FILL
XFILL112280x31050 gnd vdd FILL
XFILL_4__10493_ gnd vdd FILL
XSFILL64040x57050 gnd vdd FILL
XFILL_2__11672_ gnd vdd FILL
XFILL_0__12851_ gnd vdd FILL
XFILL_6__15930_ gnd vdd FILL
XFILL_4__15020_ gnd vdd FILL
X_10169_ _10169_/A _9017_/B gnd _10169_/Y vdd NAND2X1
XFILL_4__12232_ gnd vdd FILL
XFILL_5__10803_ gnd vdd FILL
XFILL_5__14571_ gnd vdd FILL
XFILL_2__13411_ gnd vdd FILL
XFILL_5__11783_ gnd vdd FILL
XFILL_3__15750_ gnd vdd FILL
XFILL_2__10623_ gnd vdd FILL
XFILL_3__12962_ gnd vdd FILL
XFILL_1__12052_ gnd vdd FILL
XFILL_0__11802_ gnd vdd FILL
XFILL_2__8265_ gnd vdd FILL
XFILL_0__15570_ gnd vdd FILL
XFILL_2__14391_ gnd vdd FILL
XFILL_0__12782_ gnd vdd FILL
XFILL_5__16310_ gnd vdd FILL
XFILL_3__14701_ gnd vdd FILL
XFILL_5__13522_ gnd vdd FILL
XFILL_3__11913_ gnd vdd FILL
XFILL_4__12163_ gnd vdd FILL
XFILL_2__7216_ gnd vdd FILL
X_14977_ _14976_/Y _14964_/Y gnd _14978_/A vdd NOR2X1
XFILL_2__16130_ gnd vdd FILL
XFILL_1__11003_ gnd vdd FILL
XFILL_2__13342_ gnd vdd FILL
XFILL_3__15681_ gnd vdd FILL
XSFILL43880x15050 gnd vdd FILL
XFILL_3__12893_ gnd vdd FILL
XFILL_2__8196_ gnd vdd FILL
XFILL_0__14521_ gnd vdd FILL
XFILL_2__10554_ gnd vdd FILL
XFILL_0__11733_ gnd vdd FILL
XFILL_5__16241_ gnd vdd FILL
XFILL_5__9994_ gnd vdd FILL
X_13928_ _13928_/A _13928_/B _13925_/Y gnd _13929_/B vdd NAND3X1
XFILL_4__11114_ gnd vdd FILL
XFILL_3__14632_ gnd vdd FILL
XFILL_5__13453_ gnd vdd FILL
XFILL_6__15792_ gnd vdd FILL
XFILL_5__10665_ gnd vdd FILL
XFILL_4__12094_ gnd vdd FILL
XFILL_1__15811_ gnd vdd FILL
XFILL_2__16061_ gnd vdd FILL
XFILL_3__11844_ gnd vdd FILL
XFILL_2__13273_ gnd vdd FILL
XFILL_0__14452_ gnd vdd FILL
XFILL_0__11664_ gnd vdd FILL
XFILL_5__12404_ gnd vdd FILL
XFILL_6__14743_ gnd vdd FILL
X_13859_ _8926_/Q gnd _13859_/Y vdd INVX1
XFILL_4__15922_ gnd vdd FILL
XFILL_5__16172_ gnd vdd FILL
XFILL_2__15012_ gnd vdd FILL
XFILL_5__13384_ gnd vdd FILL
XFILL_4__11045_ gnd vdd FILL
XFILL_3__14563_ gnd vdd FILL
XSFILL18920x53050 gnd vdd FILL
XFILL_0__13403_ gnd vdd FILL
XFILL_2__12224_ gnd vdd FILL
XFILL_2__7078_ gnd vdd FILL
XFILL_3__7960_ gnd vdd FILL
XFILL_0__10615_ gnd vdd FILL
XFILL_1__15742_ gnd vdd FILL
XFILL_3__11775_ gnd vdd FILL
XFILL_0__14383_ gnd vdd FILL
XFILL_1__12954_ gnd vdd FILL
XFILL_3__16302_ gnd vdd FILL
XFILL_5__8876_ gnd vdd FILL
XFILL_5__12335_ gnd vdd FILL
XFILL_0__11595_ gnd vdd FILL
XFILL_1_BUFX2_insert260 gnd vdd FILL
XFILL_5__15123_ gnd vdd FILL
XFILL_1_BUFX2_insert271 gnd vdd FILL
XFILL_3__13514_ gnd vdd FILL
XFILL_3__6911_ gnd vdd FILL
XFILL_6__11886_ gnd vdd FILL
XFILL_4__15853_ gnd vdd FILL
XFILL_0__13334_ gnd vdd FILL
XFILL_3__14494_ gnd vdd FILL
XFILL_1_BUFX2_insert282 gnd vdd FILL
XSFILL99400x51050 gnd vdd FILL
XFILL_1__11905_ gnd vdd FILL
XFILL_0__16122_ gnd vdd FILL
XFILL_2__12155_ gnd vdd FILL
XFILL_1__15673_ gnd vdd FILL
XFILL_3__7891_ gnd vdd FILL
XFILL_1_BUFX2_insert293 gnd vdd FILL
XFILL_5__7827_ gnd vdd FILL
XFILL_0__10546_ gnd vdd FILL
X_15529_ _9185_/Q gnd _15530_/C vdd INVX1
XFILL_0__9921_ gnd vdd FILL
XFILL_1__12885_ gnd vdd FILL
XFILL_4__14804_ gnd vdd FILL
XFILL_3__16233_ gnd vdd FILL
X_8460_ _8460_/A _6924_/B gnd _8461_/C vdd NAND2X1
XFILL_5__15054_ gnd vdd FILL
XFILL_5__12266_ gnd vdd FILL
XFILL_5_BUFX2_insert609 gnd vdd FILL
XFILL_6__10837_ gnd vdd FILL
XFILL_3__13445_ gnd vdd FILL
XFILL_2__11106_ gnd vdd FILL
XFILL_3__9630_ gnd vdd FILL
XFILL_1__14624_ gnd vdd FILL
XFILL_4__12996_ gnd vdd FILL
XFILL_2__12086_ gnd vdd FILL
XFILL_3__10657_ gnd vdd FILL
XFILL_3__6842_ gnd vdd FILL
XFILL_4__15784_ gnd vdd FILL
XFILL_0__16053_ gnd vdd FILL
XFILL_0__13265_ gnd vdd FILL
XFILL_1__11836_ gnd vdd FILL
XFILL_5__7758_ gnd vdd FILL
X_7411_ _7411_/Q _7411_/CLK _7411_/R vdd _7411_/D gnd vdd DFFSR
XFILL_5__14005_ gnd vdd FILL
XFILL_5__11217_ gnd vdd FILL
XFILL_0_BUFX2_insert960 gnd vdd FILL
XFILL_6__13556_ gnd vdd FILL
XFILL_0__9852_ gnd vdd FILL
XFILL112360x11050 gnd vdd FILL
XFILL_2__15914_ gnd vdd FILL
XFILL_0_BUFX2_insert971 gnd vdd FILL
XFILL_4__14735_ gnd vdd FILL
XFILL_4__11947_ gnd vdd FILL
XSFILL64120x37050 gnd vdd FILL
XFILL_5__12197_ gnd vdd FILL
XFILL_2__11037_ gnd vdd FILL
XFILL_0__15004_ gnd vdd FILL
XFILL_3__16164_ gnd vdd FILL
X_8391_ _8433_/Q gnd _8391_/Y vdd INVX1
XFILL_3__13376_ gnd vdd FILL
XFILL_0_BUFX2_insert982 gnd vdd FILL
XFILL_0__12216_ gnd vdd FILL
XFILL_0_BUFX2_insert993 gnd vdd FILL
XFILL_1__14555_ gnd vdd FILL
XSFILL74280x81050 gnd vdd FILL
XFILL_6__9270_ gnd vdd FILL
XFILL_1__11767_ gnd vdd FILL
XFILL_5__7689_ gnd vdd FILL
X_7342_ _7340_/Y _7323_/A _7342_/C gnd _7400_/D vdd OAI21X1
XFILL_5__11148_ gnd vdd FILL
XFILL_3__15115_ gnd vdd FILL
XFILL_0__9783_ gnd vdd FILL
XFILL_3__8512_ gnd vdd FILL
XFILL_2__9719_ gnd vdd FILL
XFILL_3__12327_ gnd vdd FILL
XFILL_4__11878_ gnd vdd FILL
XFILL_0__6995_ gnd vdd FILL
XFILL_3__16095_ gnd vdd FILL
XFILL_2__15845_ gnd vdd FILL
XFILL_4__14666_ gnd vdd FILL
XFILL_1__13506_ gnd vdd FILL
XFILL_5__9428_ gnd vdd FILL
XFILL_3__9492_ gnd vdd FILL
XFILL_6__8221_ gnd vdd FILL
XFILL_0__12147_ gnd vdd FILL
XFILL_1__14486_ gnd vdd FILL
XFILL_1__11698_ gnd vdd FILL
XFILL_4__16405_ gnd vdd FILL
XFILL_6__12438_ gnd vdd FILL
XFILL_0__8734_ gnd vdd FILL
XFILL_4__10829_ gnd vdd FILL
XFILL_4__13617_ gnd vdd FILL
XFILL_5__15956_ gnd vdd FILL
XFILL_3__15046_ gnd vdd FILL
X_7273_ _7273_/Q _7916_/CLK _7276_/R vdd _7217_/Y gnd vdd DFFSR
XFILL_5__11079_ gnd vdd FILL
XFILL_4__14597_ gnd vdd FILL
XFILL_1__16225_ gnd vdd FILL
XFILL_3__12258_ gnd vdd FILL
XFILL_3__8443_ gnd vdd FILL
XFILL_1__13437_ gnd vdd FILL
XFILL_1__10649_ gnd vdd FILL
XFILL_2__15776_ gnd vdd FILL
XFILL_5__9359_ gnd vdd FILL
XFILL_0__12078_ gnd vdd FILL
XFILL_2__12988_ gnd vdd FILL
X_9012_ _9012_/A _9011_/A _9012_/C gnd _9066_/D vdd OAI21X1
XFILL_5__14907_ gnd vdd FILL
XFILL_4__13548_ gnd vdd FILL
XFILL_4__16336_ gnd vdd FILL
XFILL_3__11209_ gnd vdd FILL
XFILL_2__14727_ gnd vdd FILL
XFILL_5__15887_ gnd vdd FILL
XFILL_3__8374_ gnd vdd FILL
XFILL_0__15906_ gnd vdd FILL
XFILL_3__12189_ gnd vdd FILL
XFILL_2__11939_ gnd vdd FILL
XSFILL115000x34050 gnd vdd FILL
XFILL_0__11029_ gnd vdd FILL
XFILL_1__16156_ gnd vdd FILL
XFILL_1__13368_ gnd vdd FILL
XSFILL69640x68050 gnd vdd FILL
XFILL_0__7616_ gnd vdd FILL
XFILL_5__14838_ gnd vdd FILL
XFILL_0__8596_ gnd vdd FILL
XFILL_3__7325_ gnd vdd FILL
XFILL_1__15107_ gnd vdd FILL
XFILL_4__13479_ gnd vdd FILL
XFILL_4__16267_ gnd vdd FILL
XFILL_1__12319_ gnd vdd FILL
XFILL_2__14658_ gnd vdd FILL
XFILL_1__13299_ gnd vdd FILL
XFILL_0__15837_ gnd vdd FILL
XFILL_1__16087_ gnd vdd FILL
XFILL_4__15218_ gnd vdd FILL
XFILL_0__7547_ gnd vdd FILL
XSFILL104840x77050 gnd vdd FILL
XFILL_2__13609_ gnd vdd FILL
XFILL_4__16198_ gnd vdd FILL
XSFILL33880x47050 gnd vdd FILL
XFILL_5__14769_ gnd vdd FILL
XFILL_1__15038_ gnd vdd FILL
XFILL_3__15948_ gnd vdd FILL
XFILL_2__14589_ gnd vdd FILL
XFILL_0__15768_ gnd vdd FILL
X_9914_ _9912_/Y _9896_/B _9914_/C gnd _9964_/D vdd OAI21X1
XFILL_4__15149_ gnd vdd FILL
XFILL_0__7478_ gnd vdd FILL
XFILL_2__16328_ gnd vdd FILL
XSFILL48920x69050 gnd vdd FILL
XFILL_0__14719_ gnd vdd FILL
XFILL_3__7187_ gnd vdd FILL
XFILL_3__15879_ gnd vdd FILL
XFILL_0__9217_ gnd vdd FILL
XFILL_1__8010_ gnd vdd FILL
XSFILL64200x17050 gnd vdd FILL
XFILL_0__15699_ gnd vdd FILL
XFILL_6_BUFX2_insert1007 gnd vdd FILL
X_9845_ _9811_/A _9589_/CLK _7285_/R vdd _9845_/D gnd vdd DFFSR
XFILL_2__16259_ gnd vdd FILL
XSFILL48520x71050 gnd vdd FILL
XFILL_0__9148_ gnd vdd FILL
XSFILL49000x78050 gnd vdd FILL
X_9776_ _9798_/B _8624_/B gnd _9777_/C vdd NAND2X1
XSFILL23640x1050 gnd vdd FILL
XSFILL89400x83050 gnd vdd FILL
XFILL_4__6951_ gnd vdd FILL
X_6988_ _6988_/A _6988_/B _6988_/C gnd _6988_/Y vdd OAI21X1
XSFILL3640x24050 gnd vdd FILL
XSFILL63800x6050 gnd vdd FILL
X_8727_ _8801_/Q gnd _8727_/Y vdd INVX1
XFILL_0__9079_ gnd vdd FILL
XFILL_6_BUFX2_insert454 gnd vdd FILL
XBUFX2_insert509 BUFX2_insert494/A gnd _7921_/R vdd BUFX2
XFILL_4__9670_ gnd vdd FILL
XSFILL28840x36050 gnd vdd FILL
XFILL_4__6882_ gnd vdd FILL
XFILL_1__8912_ gnd vdd FILL
XSFILL54120x69050 gnd vdd FILL
XFILL_6__7798_ gnd vdd FILL
XFILL112120x5050 gnd vdd FILL
XSFILL68440x22050 gnd vdd FILL
XFILL_1__9892_ gnd vdd FILL
XFILL_4__8621_ gnd vdd FILL
X_8658_ _8656_/Y _8657_/A _8658_/C gnd _8658_/Y vdd OAI21X1
XFILL_4_BUFX2_insert1000 gnd vdd FILL
XFILL_4_BUFX2_insert1011 gnd vdd FILL
X_7609_ _7592_/B _8377_/B gnd _7609_/Y vdd NAND2X1
XFILL_1__8843_ gnd vdd FILL
XFILL_4_BUFX2_insert1022 gnd vdd FILL
XFILL_4_BUFX2_insert1033 gnd vdd FILL
X_8589_ _8589_/A _8589_/B _8588_/Y gnd _8589_/Y vdd OAI21X1
XFILL_3__9759_ gnd vdd FILL
XFILL_4_BUFX2_insert1044 gnd vdd FILL
XFILL_4_BUFX2_insert1055 gnd vdd FILL
XSFILL33960x27050 gnd vdd FILL
XFILL_4_BUFX2_insert1066 gnd vdd FILL
XFILL_4__7503_ gnd vdd FILL
XFILL_1__8774_ gnd vdd FILL
XFILL_4__8483_ gnd vdd FILL
XFILL_4_BUFX2_insert1088 gnd vdd FILL
X_11210_ _11200_/Y _11201_/Y _11209_/Y gnd _11210_/Y vdd OAI21X1
X_12190_ _13200_/Q gnd _12192_/A vdd INVX1
XFILL_1__7725_ gnd vdd FILL
XFILL_4__7434_ gnd vdd FILL
XSFILL58360x74050 gnd vdd FILL
X_11141_ _11141_/A _11519_/C gnd _11141_/Y vdd NAND2X1
XFILL_3_BUFX2_insert300 gnd vdd FILL
XFILL_4__7365_ gnd vdd FILL
XFILL_3_BUFX2_insert311 gnd vdd FILL
XFILL_3_BUFX2_insert322 gnd vdd FILL
X_11072_ _11072_/A _11071_/Y gnd _11713_/C vdd NOR2X1
XFILL_3_BUFX2_insert333 gnd vdd FILL
XSFILL23880x79050 gnd vdd FILL
XFILL_4__9104_ gnd vdd FILL
XFILL_1__7587_ gnd vdd FILL
XFILL_3_BUFX2_insert344 gnd vdd FILL
X_10023_ _10024_/B _9895_/B gnd _10023_/Y vdd NAND2X1
XFILL_3_BUFX2_insert355 gnd vdd FILL
X_14900_ _16268_/A _14344_/B gnd _14900_/Y vdd NAND2X1
XFILL_4__7296_ gnd vdd FILL
XFILL_3_BUFX2_insert366 gnd vdd FILL
XFILL_2_BUFX2_insert1070 gnd vdd FILL
XFILL_3_BUFX2_insert377 gnd vdd FILL
X_15880_ _8426_/Q gnd _15881_/D vdd INVX1
XFILL_3_BUFX2_insert388 gnd vdd FILL
XFILL_4__9035_ gnd vdd FILL
XFILL_2_BUFX2_insert1092 gnd vdd FILL
XFILL_3_BUFX2_insert399 gnd vdd FILL
X_14831_ _14831_/A _14830_/Y gnd _14831_/Y vdd NOR2X1
XFILL_1__9257_ gnd vdd FILL
XSFILL79160x53050 gnd vdd FILL
XFILL_1__8208_ gnd vdd FILL
X_14762_ _7281_/Q _14762_/B _13864_/B _8647_/A gnd _14764_/A vdd AOI22X1
X_11974_ _11974_/A gnd _11976_/A vdd INVX1
X_13713_ _13705_/Y _13713_/B gnd _13713_/Y vdd NAND2X1
XFILL_5__6991_ gnd vdd FILL
X_10925_ _10924_/Y _6837_/A gnd _10925_/Y vdd OR2X2
XFILL_5__10450_ gnd vdd FILL
X_14693_ _8688_/Q _13864_/B _13864_/C _8560_/Q gnd _14702_/A vdd AOI22X1
XFILL_1__8139_ gnd vdd FILL
XFILL_2__10270_ gnd vdd FILL
XFILL_5__8730_ gnd vdd FILL
X_16432_ _16432_/Q _7269_/CLK _9061_/R vdd _16368_/Y gnd vdd DFFSR
XFILL_4_CLKBUF1_insert112 gnd vdd FILL
XFILL_4__9937_ gnd vdd FILL
X_13644_ _13644_/A _13644_/B gnd _13648_/C vdd NOR2X1
XSFILL84280x44050 gnd vdd FILL
XFILL_4_CLKBUF1_insert123 gnd vdd FILL
XFILL_5__10381_ gnd vdd FILL
X_10856_ _10796_/A _7912_/CLK _7911_/R vdd _10798_/Y gnd vdd DFFSR
XFILL_4_CLKBUF1_insert134 gnd vdd FILL
XFILL_0__10400_ gnd vdd FILL
XFILL_4_CLKBUF1_insert145 gnd vdd FILL
XFILL_2__8952_ gnd vdd FILL
XFILL_3__11560_ gnd vdd FILL
XFILL_4_CLKBUF1_insert156 gnd vdd FILL
XFILL_0__11380_ gnd vdd FILL
XFILL_5__8661_ gnd vdd FILL
XFILL_5__12120_ gnd vdd FILL
XFILL_4__9868_ gnd vdd FILL
X_16363_ _16363_/A gnd _16363_/Y vdd INVX1
XFILL_4_CLKBUF1_insert167 gnd vdd FILL
XFILL_3__10511_ gnd vdd FILL
XSFILL99320x66050 gnd vdd FILL
XFILL_4_CLKBUF1_insert178 gnd vdd FILL
XFILL_6__11671_ gnd vdd FILL
X_13575_ _9048_/Q gnd _13577_/B vdd INVX1
XFILL_4__12850_ gnd vdd FILL
XSFILL59080x20050 gnd vdd FILL
X_10787_ _10853_/Q gnd _10787_/Y vdd INVX1
XFILL_4_CLKBUF1_insert189 gnd vdd FILL
XFILL_5__7612_ gnd vdd FILL
XFILL_0_BUFX2_insert234 gnd vdd FILL
XFILL_2__8883_ gnd vdd FILL
XFILL_3__11491_ gnd vdd FILL
XFILL_0_BUFX2_insert245 gnd vdd FILL
X_15314_ _9180_/Q gnd _15314_/Y vdd INVX1
XFILL_5__8592_ gnd vdd FILL
X_12526_ _12430_/A gnd _12526_/Y vdd INVX1
XFILL_5__12051_ gnd vdd FILL
XFILL_0_BUFX2_insert256 gnd vdd FILL
XFILL_4__11801_ gnd vdd FILL
XFILL_4__9799_ gnd vdd FILL
XFILL_3__13230_ gnd vdd FILL
XFILL_0_BUFX2_insert267 gnd vdd FILL
XFILL_6__14390_ gnd vdd FILL
X_16294_ _10869_/Q _15357_/B _16294_/C _14956_/B gnd _16294_/Y vdd AOI22X1
XFILL_4__12781_ gnd vdd FILL
XFILL_3__10442_ gnd vdd FILL
XFILL_2__7834_ gnd vdd FILL
XFILL_0_BUFX2_insert278 gnd vdd FILL
XFILL112280x26050 gnd vdd FILL
XFILL_1__11621_ gnd vdd FILL
XFILL_2__13960_ gnd vdd FILL
XFILL_5__7543_ gnd vdd FILL
XFILL_0_BUFX2_insert289 gnd vdd FILL
XFILL_0__10262_ gnd vdd FILL
XFILL_5__11002_ gnd vdd FILL
XFILL_6__13341_ gnd vdd FILL
X_15245_ _15177_/B _15245_/B _15382_/B gnd _15680_/C vdd NOR3X1
X_12457_ _12361_/A gnd _12457_/Y vdd INVX1
XFILL_4__14520_ gnd vdd FILL
XFILL_6__10553_ gnd vdd FILL
XFILL_4__11732_ gnd vdd FILL
XFILL_2__12911_ gnd vdd FILL
XFILL_0__12001_ gnd vdd FILL
XFILL_3__13161_ gnd vdd FILL
XFILL_2__7765_ gnd vdd FILL
XFILL_1__14340_ gnd vdd FILL
XFILL_3__10373_ gnd vdd FILL
XFILL_1__11552_ gnd vdd FILL
XFILL_2__13891_ gnd vdd FILL
XFILL_5__15810_ gnd vdd FILL
X_11408_ _11408_/A gnd _11409_/C vdd INVX1
XFILL_5__7474_ gnd vdd FILL
XFILL_0__10193_ gnd vdd FILL
XFILL_4__14451_ gnd vdd FILL
X_15176_ _15176_/A _15176_/B _15171_/Y gnd _15185_/B vdd NAND3X1
XFILL_2__9504_ gnd vdd FILL
XFILL_3__12112_ gnd vdd FILL
X_12388_ _12388_/A gnd _12390_/A vdd INVX1
XFILL_2__15630_ gnd vdd FILL
XFILL_4__11663_ gnd vdd FILL
XFILL_1__10503_ gnd vdd FILL
XFILL_2__12842_ gnd vdd FILL
XFILL_3__13092_ gnd vdd FILL
XFILL_5__9213_ gnd vdd FILL
XFILL_2__7696_ gnd vdd FILL
XFILL_2_BUFX2_insert16 gnd vdd FILL
XFILL_1__11483_ gnd vdd FILL
XFILL_1__14271_ gnd vdd FILL
X_14127_ _9188_/Q gnd _14127_/Y vdd INVX1
XFILL_4__13402_ gnd vdd FILL
XFILL_2_BUFX2_insert27 gnd vdd FILL
XFILL_4__10614_ gnd vdd FILL
X_11339_ _11224_/Y _11215_/Y gnd _11835_/C vdd NAND2X1
XFILL_2_BUFX2_insert38 gnd vdd FILL
XFILL_5__15741_ gnd vdd FILL
XFILL_1__16010_ gnd vdd FILL
XFILL_3__12043_ gnd vdd FILL
XFILL_5__12953_ gnd vdd FILL
XFILL_4__14382_ gnd vdd FILL
XFILL_1__13222_ gnd vdd FILL
XFILL_2_BUFX2_insert49 gnd vdd FILL
XFILL_2__15561_ gnd vdd FILL
XFILL_1__10434_ gnd vdd FILL
XFILL_4__11594_ gnd vdd FILL
XFILL_2__12773_ gnd vdd FILL
XFILL_5__9144_ gnd vdd FILL
XSFILL114440x42050 gnd vdd FILL
XFILL_0__13952_ gnd vdd FILL
XFILL_4__13333_ gnd vdd FILL
XFILL_0__8450_ gnd vdd FILL
X_14058_ _14058_/A _13601_/B _14237_/B _14056_/Y gnd _14062_/A vdd OAI22X1
XFILL_4__16121_ gnd vdd FILL
XFILL_5__11904_ gnd vdd FILL
XFILL_5__15672_ gnd vdd FILL
XFILL_2__14512_ gnd vdd FILL
XFILL_4__10545_ gnd vdd FILL
XFILL_1__13153_ gnd vdd FILL
XFILL_2__9366_ gnd vdd FILL
XFILL_2__11724_ gnd vdd FILL
XFILL_5__12884_ gnd vdd FILL
XFILL_0__12903_ gnd vdd FILL
XFILL_1__10365_ gnd vdd FILL
XFILL_2__15492_ gnd vdd FILL
X_13009_ vdd _13009_/B gnd _13010_/C vdd NAND2X1
XFILL_5__14623_ gnd vdd FILL
XFILL_0__13883_ gnd vdd FILL
XFILL_6__12085_ gnd vdd FILL
XFILL_4__16052_ gnd vdd FILL
XFILL_4__13264_ gnd vdd FILL
XFILL_0__8381_ gnd vdd FILL
XFILL_1__12104_ gnd vdd FILL
XFILL_3__7110_ gnd vdd FILL
XFILL_3__15802_ gnd vdd FILL
XFILL_2__8317_ gnd vdd FILL
XFILL_5__11835_ gnd vdd FILL
XFILL_2__14443_ gnd vdd FILL
XFILL_3__8090_ gnd vdd FILL
XFILL_0__15622_ gnd vdd FILL
XFILL_3__13994_ gnd vdd FILL
XFILL_1__13084_ gnd vdd FILL
XFILL_2__11655_ gnd vdd FILL
XFILL_2__9297_ gnd vdd FILL
XFILL_0__12834_ gnd vdd FILL
XSFILL99400x46050 gnd vdd FILL
XFILL_4__15003_ gnd vdd FILL
XFILL_1__10296_ gnd vdd FILL
XFILL_0__7332_ gnd vdd FILL
XFILL_4__12215_ gnd vdd FILL
XFILL_5__14554_ gnd vdd FILL
XFILL_3__7041_ gnd vdd FILL
XFILL_2__8248_ gnd vdd FILL
X_7960_ _7970_/B _8088_/B gnd _7961_/C vdd NAND2X1
XFILL_1__12035_ gnd vdd FILL
XFILL_3__15733_ gnd vdd FILL
XFILL_5__11766_ gnd vdd FILL
XFILL_2__14374_ gnd vdd FILL
XFILL_0__12765_ gnd vdd FILL
XFILL_0__15553_ gnd vdd FILL
XFILL_2__11586_ gnd vdd FILL
XFILL_5__13505_ gnd vdd FILL
X_6911_ _6911_/A gnd _6913_/A vdd INVX1
XFILL_2__16113_ gnd vdd FILL
XFILL_4__12146_ gnd vdd FILL
XFILL_5__14485_ gnd vdd FILL
XFILL_2__13325_ gnd vdd FILL
XFILL_3__15664_ gnd vdd FILL
XFILL_5__11697_ gnd vdd FILL
XFILL_0__14504_ gnd vdd FILL
XFILL_3__12876_ gnd vdd FILL
X_7891_ _7925_/Q gnd _7893_/A vdd INVX1
XFILL_0__11716_ gnd vdd FILL
XFILL_2__10537_ gnd vdd FILL
XFILL_0__9002_ gnd vdd FILL
XFILL_0__12696_ gnd vdd FILL
XFILL_5__16224_ gnd vdd FILL
XFILL_0__15484_ gnd vdd FILL
XFILL_3__14615_ gnd vdd FILL
XFILL_5__10648_ gnd vdd FILL
XFILL_0__7194_ gnd vdd FILL
X_9630_ _9597_/A _7838_/B gnd _9631_/C vdd NAND2X1
XFILL_5__9977_ gnd vdd FILL
XFILL_5__13436_ gnd vdd FILL
XFILL_2__16044_ gnd vdd FILL
XSFILL89880x55050 gnd vdd FILL
XFILL_4__12077_ gnd vdd FILL
X_6842_ _6842_/A gnd memoryAddress[4] vdd BUFX2
XFILL_3__11827_ gnd vdd FILL
XFILL_2__13256_ gnd vdd FILL
XFILL_3__15595_ gnd vdd FILL
XFILL_3__8992_ gnd vdd FILL
XFILL_0__14435_ gnd vdd FILL
XFILL_0__11647_ gnd vdd FILL
XFILL_1__13986_ gnd vdd FILL
XFILL_4__15905_ gnd vdd FILL
XSFILL49080x52050 gnd vdd FILL
XFILL_4__11028_ gnd vdd FILL
XFILL_5__16155_ gnd vdd FILL
X_9561_ _9561_/Q _8942_/CLK _9561_/R vdd _9561_/D gnd vdd DFFSR
XFILL_5__13367_ gnd vdd FILL
XFILL_3__14546_ gnd vdd FILL
XFILL_2__12207_ gnd vdd FILL
XFILL_5__10579_ gnd vdd FILL
XFILL_1__15725_ gnd vdd FILL
XFILL_3__7943_ gnd vdd FILL
XFILL_3__11758_ gnd vdd FILL
XFILL_0__14366_ gnd vdd FILL
XFILL_2__10399_ gnd vdd FILL
XFILL_0__11578_ gnd vdd FILL
XFILL_5__15106_ gnd vdd FILL
X_8512_ _8512_/A _8484_/A _8511_/Y gnd _8512_/Y vdd OAI21X1
XFILL_5__8859_ gnd vdd FILL
XFILL_5__12318_ gnd vdd FILL
XFILL_5__13298_ gnd vdd FILL
XFILL_4__15836_ gnd vdd FILL
XFILL_3__10709_ gnd vdd FILL
XFILL_5__16086_ gnd vdd FILL
XFILL_0__13317_ gnd vdd FILL
XFILL_3__14477_ gnd vdd FILL
XFILL_2__12138_ gnd vdd FILL
XFILL_5_BUFX2_insert406 gnd vdd FILL
XFILL_0__16105_ gnd vdd FILL
X_9492_ _9492_/A gnd _9494_/A vdd INVX1
XSFILL114520x22050 gnd vdd FILL
XFILL_1__15656_ gnd vdd FILL
XFILL_0__10529_ gnd vdd FILL
XFILL_3__7874_ gnd vdd FILL
XFILL_3__11689_ gnd vdd FILL
XFILL_5_BUFX2_insert417 gnd vdd FILL
XFILL_6__13608_ gnd vdd FILL
XFILL_1__12868_ gnd vdd FILL
XFILL_5_BUFX2_insert428 gnd vdd FILL
XFILL_0__9904_ gnd vdd FILL
XFILL_0__14297_ gnd vdd FILL
XFILL_3__16216_ gnd vdd FILL
XFILL_5__15037_ gnd vdd FILL
XFILL_5_BUFX2_insert439 gnd vdd FILL
XFILL_3__9613_ gnd vdd FILL
XSFILL43800x54050 gnd vdd FILL
XFILL_3__13428_ gnd vdd FILL
XFILL_5__12249_ gnd vdd FILL
X_8443_ _8443_/A _8496_/A _8443_/C gnd _8535_/D vdd OAI21X1
XFILL_1__14607_ gnd vdd FILL
XFILL_4__15767_ gnd vdd FILL
XFILL_0__13248_ gnd vdd FILL
XFILL_0__16036_ gnd vdd FILL
XFILL_2__12069_ gnd vdd FILL
XFILL_4__12979_ gnd vdd FILL
XFILL_1__11819_ gnd vdd FILL
XFILL_1__15587_ gnd vdd FILL
XFILL_0_BUFX2_insert790 gnd vdd FILL
X_8374_ _8333_/B _7990_/B gnd _8374_/Y vdd NAND2X1
XSFILL103560x46050 gnd vdd FILL
XFILL_4__14718_ gnd vdd FILL
XSFILL3560x8050 gnd vdd FILL
XFILL_3__16147_ gnd vdd FILL
XFILL_3__13359_ gnd vdd FILL
XSFILL69240x65050 gnd vdd FILL
XFILL_3__9544_ gnd vdd FILL
XFILL_4__15698_ gnd vdd FILL
XFILL_1__14538_ gnd vdd FILL
X_7325_ _7325_/A gnd _7327_/A vdd INVX1
XFILL_6__16258_ gnd vdd FILL
XFILL_0__9766_ gnd vdd FILL
XFILL_2__15828_ gnd vdd FILL
XFILL_0__6978_ gnd vdd FILL
XFILL_4__14649_ gnd vdd FILL
XFILL_3__16078_ gnd vdd FILL
XFILL_3__9475_ gnd vdd FILL
XFILL_1__14469_ gnd vdd FILL
XSFILL33480x44050 gnd vdd FILL
XFILL_6__15209_ gnd vdd FILL
XFILL_0__8717_ gnd vdd FILL
XFILL_3__15029_ gnd vdd FILL
XFILL_5__15939_ gnd vdd FILL
X_7256_ _7256_/Q _7143_/CLK _7015_/R vdd _7256_/D gnd vdd DFFSR
XFILL_1__16208_ gnd vdd FILL
XFILL_1__8490_ gnd vdd FILL
XFILL_2__15759_ gnd vdd FILL
XSFILL23720x21050 gnd vdd FILL
XFILL_4__16319_ gnd vdd FILL
XFILL_1__7441_ gnd vdd FILL
XFILL_0__8648_ gnd vdd FILL
X_7187_ _7187_/A _7250_/B _7186_/Y gnd _7187_/Y vdd OAI21X1
XFILL_3__8357_ gnd vdd FILL
XFILL_1__16139_ gnd vdd FILL
XSFILL89400x78050 gnd vdd FILL
XSFILL3640x19050 gnd vdd FILL
XFILL_1__7372_ gnd vdd FILL
XFILL_3__7308_ gnd vdd FILL
XFILL_0__8579_ gnd vdd FILL
XFILL_2_BUFX2_insert307 gnd vdd FILL
XFILL_1_BUFX2_insert2 gnd vdd FILL
XFILL_4__7081_ gnd vdd FILL
XFILL_1__9111_ gnd vdd FILL
XFILL_2_BUFX2_insert318 gnd vdd FILL
XFILL_2_BUFX2_insert329 gnd vdd FILL
XFILL_3__7239_ gnd vdd FILL
XSFILL13640x73050 gnd vdd FILL
XSFILL94520x69050 gnd vdd FILL
XFILL_1__9042_ gnd vdd FILL
XSFILL69320x45050 gnd vdd FILL
X_9828_ _9760_/A _9306_/CLK _8801_/R vdd _9828_/D gnd vdd DFFSR
XSFILL29320x61050 gnd vdd FILL
X_10710_ _15002_/C _8818_/CLK _9430_/R vdd _10616_/Y gnd vdd DFFSR
XFILL_4__7983_ gnd vdd FILL
X_11690_ _11689_/Y gnd _12041_/A vdd INVX1
X_9759_ _9757_/Y _9813_/B _9759_/C gnd _9827_/D vdd OAI21X1
XBUFX2_insert306 _11983_/Y gnd _12059_/C vdd BUFX2
XFILL_4__6934_ gnd vdd FILL
XFILL_4__9722_ gnd vdd FILL
XBUFX2_insert317 _15000_/Y gnd _16235_/A vdd BUFX2
XSFILL8760x52050 gnd vdd FILL
X_10641_ _15439_/A gnd _10643_/A vdd INVX1
XBUFX2_insert328 _13345_/Y gnd _9920_/B vdd BUFX2
XBUFX2_insert339 _12811_/Q gnd _13381_/A vdd BUFX2
XFILL_6_BUFX2_insert295 gnd vdd FILL
XFILL_4__9653_ gnd vdd FILL
XFILL_4__6865_ gnd vdd FILL
X_13360_ _13244_/A _13239_/B _13363_/B gnd _13360_/Y vdd OAI21X1
XFILL_5_CLKBUF1_insert207 gnd vdd FILL
X_10572_ _10572_/A _10557_/B _10572_/C gnd _10610_/D vdd OAI21X1
XFILL_4__8604_ gnd vdd FILL
XFILL_1__9875_ gnd vdd FILL
XFILL_5_CLKBUF1_insert218 gnd vdd FILL
XFILL_5_BUFX2_insert940 gnd vdd FILL
XFILL_5_BUFX2_insert951 gnd vdd FILL
X_12311_ _12216_/A gnd _12311_/C gnd _12311_/Y vdd NAND3X1
XFILL_5_BUFX2_insert962 gnd vdd FILL
X_13291_ _13291_/A _13290_/Y gnd _13292_/B vdd NAND2X1
XFILL_5_BUFX2_insert973 gnd vdd FILL
XFILL_1__8826_ gnd vdd FILL
XFILL_5_BUFX2_insert984 gnd vdd FILL
XFILL_5_BUFX2_insert995 gnd vdd FILL
X_15030_ _12813_/Q _14980_/Y gnd _15031_/B vdd NAND2X1
X_12242_ _12239_/Y _12242_/B _12242_/C gnd _12242_/Y vdd NAND3X1
XFILL_1__8757_ gnd vdd FILL
XFILL_2__7550_ gnd vdd FILL
XSFILL13720x53050 gnd vdd FILL
XFILL_4__8466_ gnd vdd FILL
XFILL_1__7708_ gnd vdd FILL
X_12173_ _12117_/B _12938_/Q gnd _12174_/C vdd NAND2X1
XFILL_2__7481_ gnd vdd FILL
XFILL_4__7417_ gnd vdd FILL
XFILL_4__8397_ gnd vdd FILL
X_11124_ _12294_/Y gnd _11125_/B vdd INVX1
XFILL_5__7190_ gnd vdd FILL
XFILL_2__9220_ gnd vdd FILL
XSFILL28920x3050 gnd vdd FILL
XFILL_4__7348_ gnd vdd FILL
X_15932_ _15931_/Y _16228_/B _15726_/A _14501_/Y gnd _15932_/Y vdd OAI22X1
XSFILL84280x39050 gnd vdd FILL
X_11055_ _11055_/A _11055_/B gnd _11055_/Y vdd NAND2X1
XFILL_2__9151_ gnd vdd FILL
XFILL_1__10150_ gnd vdd FILL
XFILL_0__10880_ gnd vdd FILL
X_10006_ _10006_/A _10066_/B _10006_/C gnd _10080_/D vdd OAI21X1
XFILL_2__8102_ gnd vdd FILL
XFILL_5__11620_ gnd vdd FILL
X_15863_ _15863_/A _15863_/B _10162_/A _15695_/D gnd _15865_/B vdd AOI22X1
XFILL_4__10261_ gnd vdd FILL
XSFILL59080x15050 gnd vdd FILL
XFILL_4__9018_ gnd vdd FILL
XFILL_2_BUFX2_insert830 gnd vdd FILL
XFILL_2__11440_ gnd vdd FILL
XFILL_2__9082_ gnd vdd FILL
XFILL_3__10991_ gnd vdd FILL
XFILL_5__9900_ gnd vdd FILL
XFILL_4__12000_ gnd vdd FILL
X_14814_ _8778_/A gnd _14814_/Y vdd INVX1
XFILL_2_BUFX2_insert841 gnd vdd FILL
XSFILL99480x20050 gnd vdd FILL
XFILL_2_BUFX2_insert852 gnd vdd FILL
XFILL_5__11551_ gnd vdd FILL
XFILL_3__12730_ gnd vdd FILL
XFILL_2_BUFX2_insert863 gnd vdd FILL
X_15794_ _9448_/Q _15794_/B _15071_/C gnd _15795_/C vdd NAND3X1
XFILL_2_BUFX2_insert874 gnd vdd FILL
XFILL_4__10192_ gnd vdd FILL
XFILL_2__11371_ gnd vdd FILL
XFILL_2_BUFX2_insert885 gnd vdd FILL
XFILL_5__10502_ gnd vdd FILL
XFILL_6__12841_ gnd vdd FILL
XFILL_2_BUFX2_insert896 gnd vdd FILL
X_14745_ _8305_/Q _14323_/B _14745_/C gnd _14754_/B vdd AOI21X1
X_11957_ _11909_/A _12508_/A gnd _11958_/C vdd NAND2X1
XFILL_2__13110_ gnd vdd FILL
XFILL_5__11482_ gnd vdd FILL
XFILL_5__14270_ gnd vdd FILL
XFILL_3__12661_ gnd vdd FILL
XSFILL23560x56050 gnd vdd FILL
XFILL_2__10322_ gnd vdd FILL
XFILL_0__11501_ gnd vdd FILL
XFILL_1__13840_ gnd vdd FILL
XFILL_2__14090_ gnd vdd FILL
XFILL_0__12481_ gnd vdd FILL
XFILL_5__13221_ gnd vdd FILL
XFILL_5__6974_ gnd vdd FILL
X_10908_ _10906_/Y _10938_/A gnd _10963_/A vdd NOR2X1
XSFILL63960x61050 gnd vdd FILL
XFILL_5__9762_ gnd vdd FILL
XFILL_3__14400_ gnd vdd FILL
XFILL_5__10433_ gnd vdd FILL
XSFILL13800x33050 gnd vdd FILL
XFILL_3__11612_ gnd vdd FILL
X_14676_ _7791_/Q gnd _16079_/D vdd INVX1
XFILL_2__10253_ gnd vdd FILL
XFILL_3__15380_ gnd vdd FILL
XFILL_0__14220_ gnd vdd FILL
X_11888_ _12343_/A _11975_/A gnd _11889_/C vdd NAND2X1
XFILL_4__13951_ gnd vdd FILL
XFILL_2__13041_ gnd vdd FILL
XFILL_3__12592_ gnd vdd FILL
XFILL_2__9984_ gnd vdd FILL
XSFILL79240x28050 gnd vdd FILL
XFILL_0__11432_ gnd vdd FILL
XFILL_5__8713_ gnd vdd FILL
XFILL_4_BUFX2_insert6 gnd vdd FILL
XFILL_1__13771_ gnd vdd FILL
X_16415_ gnd gnd gnd _16416_/C vdd NAND2X1
XFILL_1__10983_ gnd vdd FILL
X_13627_ _14868_/A _10623_/A _9177_/Q _14868_/D gnd _13635_/B vdd AOI22X1
XFILL_5__13152_ gnd vdd FILL
XFILL_4__12902_ gnd vdd FILL
XFILL_3__14331_ gnd vdd FILL
XFILL_5__10364_ gnd vdd FILL
X_10839_ _13485_/A _7515_/CLK _7515_/R vdd _10839_/D gnd vdd DFFSR
XFILL_1__15510_ gnd vdd FILL
XFILL_3__11543_ gnd vdd FILL
XSFILL64040x70050 gnd vdd FILL
XFILL_4__13882_ gnd vdd FILL
XFILL_1__12722_ gnd vdd FILL
XFILL_0__14151_ gnd vdd FILL
XFILL_2__10184_ gnd vdd FILL
XFILL_5__8644_ gnd vdd FILL
XFILL_0__11363_ gnd vdd FILL
XBUFX2_insert840 _13324_/Y gnd _8607_/B vdd BUFX2
X_16346_ gnd gnd gnd _16347_/C vdd NAND2X1
XFILL_5__12103_ gnd vdd FILL
XBUFX2_insert851 _13269_/Y gnd _7068_/B vdd BUFX2
XSFILL114440x37050 gnd vdd FILL
XFILL_0__7950_ gnd vdd FILL
XBUFX2_insert862 _13314_/Y gnd _8246_/A vdd BUFX2
XFILL_4__15621_ gnd vdd FILL
XFILL_5__13083_ gnd vdd FILL
X_13558_ _13558_/A _13557_/Y gnd _13558_/Y vdd NOR2X1
XFILL_5__10295_ gnd vdd FILL
XFILL_3__14262_ gnd vdd FILL
XFILL_0__13102_ gnd vdd FILL
XFILL_4__12833_ gnd vdd FILL
XFILL_0__10314_ gnd vdd FILL
XFILL_2__8866_ gnd vdd FILL
XBUFX2_insert873 _13435_/Y gnd _14410_/A vdd BUFX2
XFILL_3__11474_ gnd vdd FILL
XFILL_1__15441_ gnd vdd FILL
XFILL_1__12653_ gnd vdd FILL
XFILL_2__14992_ gnd vdd FILL
XBUFX2_insert884 _12216_/Y gnd _12309_/C vdd BUFX2
XFILL_0__14082_ gnd vdd FILL
XSFILL84360x19050 gnd vdd FILL
XFILL_5__8575_ gnd vdd FILL
XFILL_3__16001_ gnd vdd FILL
XBUFX2_insert895 _13470_/Y gnd _13614_/C vdd BUFX2
X_12509_ vdd _12081_/A gnd _12509_/Y vdd NAND2X1
XFILL_5__12034_ gnd vdd FILL
XFILL_0__6901_ gnd vdd FILL
XFILL_0__11294_ gnd vdd FILL
XFILL_3__13213_ gnd vdd FILL
X_16277_ _8656_/A gnd _16277_/Y vdd INVX1
XFILL_4__12764_ gnd vdd FILL
XFILL_2__7817_ gnd vdd FILL
XFILL_4__15552_ gnd vdd FILL
XFILL_3__10425_ gnd vdd FILL
X_13489_ _13489_/A _13488_/Y _13489_/C gnd _13489_/Y vdd NAND3X1
XFILL_0__7881_ gnd vdd FILL
XFILL_3__14193_ gnd vdd FILL
XFILL_1__11604_ gnd vdd FILL
XFILL_2__13943_ gnd vdd FILL
XFILL_0__13033_ gnd vdd FILL
XFILL_3__7590_ gnd vdd FILL
XFILL_1__15372_ gnd vdd FILL
XFILL_0__10245_ gnd vdd FILL
X_15228_ _15228_/A _15226_/Y gnd _15229_/C vdd NOR2X1
XFILL_1__12584_ gnd vdd FILL
XFILL_0__9620_ gnd vdd FILL
XFILL_4__14503_ gnd vdd FILL
XFILL_3__13144_ gnd vdd FILL
XFILL_4__11715_ gnd vdd FILL
XFILL_4__12695_ gnd vdd FILL
XFILL_1__14323_ gnd vdd FILL
XFILL_4__15483_ gnd vdd FILL
XFILL_2__7748_ gnd vdd FILL
XFILL_2__13874_ gnd vdd FILL
XFILL_1__11535_ gnd vdd FILL
XSFILL84200x83050 gnd vdd FILL
XFILL_0__10176_ gnd vdd FILL
XFILL_6__16043_ gnd vdd FILL
XFILL_5__7457_ gnd vdd FILL
X_7110_ _7110_/A _7064_/A _7109_/Y gnd _7152_/D vdd OAI21X1
XFILL_0__9551_ gnd vdd FILL
XFILL_6__13255_ gnd vdd FILL
X_15159_ _15774_/C _13536_/D _15158_/Y _15801_/C gnd _15160_/A vdd OAI22X1
X_8090_ _8090_/A gnd _8092_/A vdd INVX1
XFILL_2__15613_ gnd vdd FILL
XFILL_4__11646_ gnd vdd FILL
XFILL_4__14434_ gnd vdd FILL
XFILL_5__13985_ gnd vdd FILL
XFILL_2__12825_ gnd vdd FILL
XFILL_3__9260_ gnd vdd FILL
XFILL_2__7679_ gnd vdd FILL
XFILL_1__14254_ gnd vdd FILL
XFILL_3__10287_ gnd vdd FILL
XFILL_1__11466_ gnd vdd FILL
XFILL_0__8502_ gnd vdd FILL
X_7041_ _7041_/A _7100_/A _7040_/Y gnd _7129_/D vdd OAI21X1
XFILL_5__15724_ gnd vdd FILL
XFILL_0__14984_ gnd vdd FILL
XFILL_0__9482_ gnd vdd FILL
XFILL_2__9418_ gnd vdd FILL
XFILL_3__12026_ gnd vdd FILL
XFILL_4__14365_ gnd vdd FILL
XFILL_3__8211_ gnd vdd FILL
XFILL_2__15544_ gnd vdd FILL
XFILL_6__10398_ gnd vdd FILL
XFILL_4__11577_ gnd vdd FILL
XFILL_2__12756_ gnd vdd FILL
XFILL_5__9127_ gnd vdd FILL
XFILL_1__10417_ gnd vdd FILL
XFILL_1__14185_ gnd vdd FILL
XFILL_0__13935_ gnd vdd FILL
XFILL_1__11397_ gnd vdd FILL
XFILL_6__12137_ gnd vdd FILL
XFILL_4__16104_ gnd vdd FILL
XFILL_4__13316_ gnd vdd FILL
XFILL_5__15655_ gnd vdd FILL
XFILL_4__10528_ gnd vdd FILL
XSFILL49080x47050 gnd vdd FILL
XFILL_3__8142_ gnd vdd FILL
XFILL112200x65050 gnd vdd FILL
XFILL_5__12867_ gnd vdd FILL
XFILL_2__11707_ gnd vdd FILL
XFILL_2__9349_ gnd vdd FILL
XFILL_4__14296_ gnd vdd FILL
XFILL_1__13136_ gnd vdd FILL
XFILL_2__15475_ gnd vdd FILL
XFILL_0__13866_ gnd vdd FILL
XFILL_5__14606_ gnd vdd FILL
XFILL_4__13247_ gnd vdd FILL
XFILL_4__16035_ gnd vdd FILL
XSFILL64120x50050 gnd vdd FILL
XFILL_0__8364_ gnd vdd FILL
XFILL_5__11818_ gnd vdd FILL
XFILL_5__15586_ gnd vdd FILL
XFILL_2__14426_ gnd vdd FILL
XFILL_3__8073_ gnd vdd FILL
X_8992_ _8992_/A gnd _8994_/A vdd INVX1
XFILL_3__13977_ gnd vdd FILL
XFILL_2__11638_ gnd vdd FILL
XFILL_0__15605_ gnd vdd FILL
XSFILL114520x17050 gnd vdd FILL
XFILL_5__8009_ gnd vdd FILL
XFILL_1__10279_ gnd vdd FILL
XFILL_0__7315_ gnd vdd FILL
XFILL_0__13797_ gnd vdd FILL
XFILL_5__14537_ gnd vdd FILL
XFILL_3__15716_ gnd vdd FILL
X_7943_ _7941_/Y _7931_/B _7943_/C gnd _7943_/Y vdd OAI21X1
XFILL_5__11749_ gnd vdd FILL
XFILL_1__12018_ gnd vdd FILL
XFILL_2__14357_ gnd vdd FILL
XFILL_0__15536_ gnd vdd FILL
XFILL_2__11569_ gnd vdd FILL
XFILL_0__12748_ gnd vdd FILL
XFILL_0__7246_ gnd vdd FILL
XFILL_4__12129_ gnd vdd FILL
XFILL_2__13308_ gnd vdd FILL
XFILL_5__14468_ gnd vdd FILL
XFILL_3__15647_ gnd vdd FILL
XFILL_3__12859_ gnd vdd FILL
X_7874_ _7892_/A _8642_/B gnd _7875_/C vdd NAND2X1
XSFILL18600x25050 gnd vdd FILL
XFILL_2__14288_ gnd vdd FILL
XFILL_5__16207_ gnd vdd FILL
XFILL_0__15467_ gnd vdd FILL
X_9613_ _9613_/A _9613_/B _9613_/C gnd _9693_/D vdd OAI21X1
XFILL_5__13419_ gnd vdd FILL
XFILL_0__7177_ gnd vdd FILL
XFILL_2__16027_ gnd vdd FILL
XFILL_2__13239_ gnd vdd FILL
XFILL_5__14399_ gnd vdd FILL
XFILL_3__8975_ gnd vdd FILL
XFILL_0__14418_ gnd vdd FILL
XFILL_3__15578_ gnd vdd FILL
XFILL_1__13969_ gnd vdd FILL
XSFILL104440x69050 gnd vdd FILL
XFILL_0__15398_ gnd vdd FILL
XFILL_5__16138_ gnd vdd FILL
X_9544_ _9466_/A _7496_/B gnd _9545_/C vdd NAND2X1
XFILL_1__7990_ gnd vdd FILL
XFILL_1__15708_ gnd vdd FILL
XFILL_3__7926_ gnd vdd FILL
XFILL_3__14529_ gnd vdd FILL
XSFILL8680x67050 gnd vdd FILL
XSFILL23720x16050 gnd vdd FILL
XFILL_0__14349_ gnd vdd FILL
XFILL_5_BUFX2_insert225 gnd vdd FILL
XFILL_4__15819_ gnd vdd FILL
XFILL_1__6941_ gnd vdd FILL
XFILL_5__16069_ gnd vdd FILL
X_9475_ _9551_/B _9475_/B gnd _9475_/Y vdd NAND2X1
XFILL_5_BUFX2_insert236 gnd vdd FILL
XFILL_1__15639_ gnd vdd FILL
XFILL_5_BUFX2_insert247 gnd vdd FILL
XFILL_3__7857_ gnd vdd FILL
XFILL_5_BUFX2_insert258 gnd vdd FILL
XFILL_1__9660_ gnd vdd FILL
XFILL_5_BUFX2_insert269 gnd vdd FILL
X_8426_ _8426_/Q _9716_/CLK _9460_/R vdd _8426_/D gnd vdd DFFSR
XFILL_1__6872_ gnd vdd FILL
XFILL_0__16019_ gnd vdd FILL
XFILL_4_BUFX2_insert903 gnd vdd FILL
XSFILL64200x30050 gnd vdd FILL
XFILL_4_BUFX2_insert914 gnd vdd FILL
XFILL_1__8611_ gnd vdd FILL
XSFILL94440x9050 gnd vdd FILL
XSFILL89000x75050 gnd vdd FILL
XFILL_6__7497_ gnd vdd FILL
XFILL_4_BUFX2_insert925 gnd vdd FILL
XFILL_3__9527_ gnd vdd FILL
XFILL_4__8320_ gnd vdd FILL
X_8357_ _8355_/Y _8356_/A _8357_/C gnd _8421_/D vdd OAI21X1
XFILL_4_BUFX2_insert936 gnd vdd FILL
XFILL_1__9591_ gnd vdd FILL
XFILL_4_BUFX2_insert947 gnd vdd FILL
XFILL_4_BUFX2_insert958 gnd vdd FILL
XFILL_4_BUFX2_insert969 gnd vdd FILL
X_7308_ _7308_/A _7180_/B gnd _7309_/C vdd NAND2X1
XFILL_0__9749_ gnd vdd FILL
XFILL_4__8251_ gnd vdd FILL
X_8288_ _8212_/A _9568_/CLK _7648_/R vdd _8214_/Y gnd vdd DFFSR
XFILL_6__9167_ gnd vdd FILL
XSFILL4120x44050 gnd vdd FILL
XFILL_1__8473_ gnd vdd FILL
XFILL_4__7202_ gnd vdd FILL
X_7239_ _7281_/Q gnd _7241_/A vdd INVX1
XFILL_6__8118_ gnd vdd FILL
XFILL_4__8182_ gnd vdd FILL
XFILL_3__9389_ gnd vdd FILL
XSFILL29320x56050 gnd vdd FILL
XSFILL54120x82050 gnd vdd FILL
XFILL_1__7424_ gnd vdd FILL
XSFILL104520x49050 gnd vdd FILL
XFILL_2_BUFX2_insert104 gnd vdd FILL
XFILL_1__7355_ gnd vdd FILL
XSFILL8760x47050 gnd vdd FILL
XFILL_4__7064_ gnd vdd FILL
X_12860_ vdd _12860_/B gnd _12861_/C vdd NAND2X1
XFILL_1__7286_ gnd vdd FILL
X_11811_ _11810_/Y _11005_/Y gnd _11811_/Y vdd AND2X2
XFILL_1__9025_ gnd vdd FILL
XFILL_1_BUFX2_insert804 gnd vdd FILL
X_12791_ _12695_/A _12667_/CLK _12809_/R vdd _12791_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert815 gnd vdd FILL
XFILL_1_BUFX2_insert826 gnd vdd FILL
X_14530_ _9836_/Q gnd _14532_/A vdd INVX1
XFILL_1_BUFX2_insert837 gnd vdd FILL
XSFILL108760x54050 gnd vdd FILL
X_11742_ _11041_/Y _11028_/Y gnd _11744_/A vdd NOR2X1
XFILL_1_BUFX2_insert848 gnd vdd FILL
XFILL_1_BUFX2_insert859 gnd vdd FILL
XSFILL13720x48050 gnd vdd FILL
XSFILL78680x36050 gnd vdd FILL
XFILL_4__7966_ gnd vdd FILL
X_14461_ _10091_/Q gnd _14461_/Y vdd INVX1
XBUFX2_insert103 _10925_/Y gnd _11955_/B vdd BUFX2
X_11673_ _11671_/Y _11672_/Y _11673_/C gnd _11673_/Y vdd OAI21X1
X_16200_ _16200_/A _16200_/B gnd _16201_/B vdd NOR2X1
XFILL_2__6981_ gnd vdd FILL
X_13412_ _13718_/B _13718_/A gnd _13412_/Y vdd NAND2X1
XFILL_4__6917_ gnd vdd FILL
X_10624_ _10661_/B _8576_/B gnd _10625_/C vdd NAND2X1
XFILL_2__8720_ gnd vdd FILL
X_14392_ _7727_/A gnd _14393_/B vdd INVX1
XFILL_1__9927_ gnd vdd FILL
XFILL_4__9636_ gnd vdd FILL
XFILL_4__6848_ gnd vdd FILL
X_16131_ _16131_/A _16130_/Y _16128_/Y gnd _16140_/A vdd NAND3X1
X_13343_ _13341_/Y _13343_/B gnd _13343_/Y vdd NOR2X1
X_10555_ _14584_/A gnd _10557_/A vdd INVX1
XFILL_2__8651_ gnd vdd FILL
XFILL_1__9858_ gnd vdd FILL
XFILL_5_BUFX2_insert770 gnd vdd FILL
XFILL_5__8360_ gnd vdd FILL
XFILL_5_BUFX2_insert781 gnd vdd FILL
XFILL_5_BUFX2_insert792 gnd vdd FILL
X_16062_ _15841_/C _14686_/D _16062_/C _15813_/C gnd _16065_/B vdd OAI22X1
X_13274_ _13274_/A _13273_/Y _13266_/Y gnd _13275_/B vdd NAND3X1
XFILL_2__7602_ gnd vdd FILL
X_10486_ _10486_/A gnd _10486_/Y vdd INVX1
XFILL_1__9789_ gnd vdd FILL
XFILL_2__10940_ gnd vdd FILL
XFILL_5__7311_ gnd vdd FILL
XFILL_0__10030_ gnd vdd FILL
XFILL_3__11190_ gnd vdd FILL
XFILL_2__8582_ gnd vdd FILL
XFILL_4__8518_ gnd vdd FILL
X_15013_ _12767_/A _12764_/A gnd _15014_/C vdd OR2X2
XFILL_4__9498_ gnd vdd FILL
X_12225_ _6872_/A _12237_/B _12269_/C _12695_/A gnd _12226_/C vdd AOI22X1
XFILL_4__11500_ gnd vdd FILL
XSFILL99480x15050 gnd vdd FILL
XFILL_4__12480_ gnd vdd FILL
XFILL_3__10141_ gnd vdd FILL
XSFILL74120x13050 gnd vdd FILL
XFILL_1__11320_ gnd vdd FILL
XSFILL18840x81050 gnd vdd FILL
XFILL_4__8449_ gnd vdd FILL
XFILL_5__7242_ gnd vdd FILL
XSFILL18040x62050 gnd vdd FILL
XFILL_2__10871_ gnd vdd FILL
XFILL_4__11431_ gnd vdd FILL
X_12156_ _12156_/A _12123_/B _12156_/C gnd _12156_/Y vdd OAI21X1
XFILL_2__12610_ gnd vdd FILL
XFILL_5__13770_ gnd vdd FILL
XFILL_5__10982_ gnd vdd FILL
XFILL_2__7464_ gnd vdd FILL
XFILL_1__11251_ gnd vdd FILL
XFILL_2__13590_ gnd vdd FILL
XFILL_0__11981_ gnd vdd FILL
X_11107_ _11542_/A _11107_/B gnd _11143_/A vdd NOR2X1
XFILL_5__7173_ gnd vdd FILL
XFILL_5__12721_ gnd vdd FILL
XFILL_4__14150_ gnd vdd FILL
X_12087_ _12007_/A _12418_/A _12059_/C gnd _12090_/A vdd NAND3X1
XSFILL13800x28050 gnd vdd FILL
XFILL_3__13900_ gnd vdd FILL
XFILL_4__11362_ gnd vdd FILL
XFILL_3__14880_ gnd vdd FILL
XFILL_0__10932_ gnd vdd FILL
XFILL_0__13720_ gnd vdd FILL
XFILL_1__11182_ gnd vdd FILL
XFILL_4__13101_ gnd vdd FILL
X_15915_ _15915_/A _15972_/B _15915_/C _14454_/Y gnd _15915_/Y vdd OAI22X1
XFILL_4__10313_ gnd vdd FILL
XFILL_5__15440_ gnd vdd FILL
X_11038_ _12138_/Y gnd _11038_/Y vdd INVX1
XFILL_5__12652_ gnd vdd FILL
XFILL_3__13831_ gnd vdd FILL
XFILL_2__9134_ gnd vdd FILL
XFILL_4__14081_ gnd vdd FILL
XFILL_4__11293_ gnd vdd FILL
XFILL_1__10133_ gnd vdd FILL
XFILL_2__15260_ gnd vdd FILL
XSFILL64040x65050 gnd vdd FILL
XFILL_2__12472_ gnd vdd FILL
XFILL_1__15990_ gnd vdd FILL
XFILL_0__13651_ gnd vdd FILL
XFILL_4__13032_ gnd vdd FILL
XFILL_5__11603_ gnd vdd FILL
XFILL_5__15371_ gnd vdd FILL
XFILL_2__14211_ gnd vdd FILL
XFILL_4__10244_ gnd vdd FILL
X_15846_ _15846_/A gnd _15848_/D vdd INVX1
XFILL_5__12583_ gnd vdd FILL
XFILL_3__13762_ gnd vdd FILL
XFILL_2__11423_ gnd vdd FILL
XFILL_0__12602_ gnd vdd FILL
XFILL_3__10974_ gnd vdd FILL
XFILL_2__15191_ gnd vdd FILL
XFILL_2_BUFX2_insert660 gnd vdd FILL
XFILL_1__14941_ gnd vdd FILL
XFILL_1__10064_ gnd vdd FILL
XFILL_0__7100_ gnd vdd FILL
XFILL_0__16370_ gnd vdd FILL
XFILL_2_BUFX2_insert671 gnd vdd FILL
XFILL_0__13582_ gnd vdd FILL
XFILL_5__14322_ gnd vdd FILL
XFILL_2_BUFX2_insert682 gnd vdd FILL
XFILL_0__10794_ gnd vdd FILL
XFILL_0__8080_ gnd vdd FILL
XFILL_3__12713_ gnd vdd FILL
XFILL_3__15501_ gnd vdd FILL
XFILL_2_BUFX2_insert693 gnd vdd FILL
XFILL_5__11534_ gnd vdd FILL
XFILL_2__8016_ gnd vdd FILL
XFILL_4__10175_ gnd vdd FILL
XFILL_2__14142_ gnd vdd FILL
X_12989_ _12987_/Y vdd _12989_/C gnd _13059_/D vdd OAI21X1
X_15777_ _15777_/A _15772_/Y _15777_/C gnd _15786_/B vdd NAND3X1
XSFILL43880x23050 gnd vdd FILL
XFILL_0__15321_ gnd vdd FILL
XFILL_3__13693_ gnd vdd FILL
XFILL_2__11354_ gnd vdd FILL
XSFILL3480x72050 gnd vdd FILL
XFILL_1__14872_ gnd vdd FILL
XFILL_0__12533_ gnd vdd FILL
XFILL_0__7031_ gnd vdd FILL
XFILL_5__14253_ gnd vdd FILL
X_14728_ _16113_/D _14200_/C _14555_/C _14726_/Y gnd _14728_/Y vdd OAI22X1
XSFILL84760x35050 gnd vdd FILL
XFILL_3__12644_ gnd vdd FILL
XFILL_2__10305_ gnd vdd FILL
XFILL_3__15432_ gnd vdd FILL
XFILL_5__11465_ gnd vdd FILL
XFILL_1__13823_ gnd vdd FILL
XFILL_4__14983_ gnd vdd FILL
XFILL_2__14073_ gnd vdd FILL
XFILL_0__15252_ gnd vdd FILL
XFILL_0__12464_ gnd vdd FILL
XFILL_5_BUFX2_insert20 gnd vdd FILL
XFILL_2__11285_ gnd vdd FILL
XSFILL84200x78050 gnd vdd FILL
XFILL_5_BUFX2_insert31 gnd vdd FILL
XFILL_5__9745_ gnd vdd FILL
XFILL_5_BUFX2_insert42 gnd vdd FILL
XFILL_5__6957_ gnd vdd FILL
XFILL_5__10416_ gnd vdd FILL
X_14659_ _7279_/Q _14762_/B _14926_/C _7023_/Q gnd _14667_/B vdd AOI22X1
X_7590_ _7590_/A gnd _7592_/A vdd INVX1
XFILL_3__15363_ gnd vdd FILL
XFILL_5__14184_ gnd vdd FILL
XFILL_5_BUFX2_insert53 gnd vdd FILL
XFILL_2__13024_ gnd vdd FILL
XFILL_5__11396_ gnd vdd FILL
XFILL_4__13934_ gnd vdd FILL
XFILL_0__14203_ gnd vdd FILL
XFILL_3__12575_ gnd vdd FILL
XFILL_3__8760_ gnd vdd FILL
XFILL_2__10236_ gnd vdd FILL
XFILL_0__11415_ gnd vdd FILL
XFILL_0__15183_ gnd vdd FILL
XFILL_1__13754_ gnd vdd FILL
XFILL_5_BUFX2_insert64 gnd vdd FILL
XFILL_1__10966_ gnd vdd FILL
XFILL_5_BUFX2_insert75 gnd vdd FILL
XFILL_0__12395_ gnd vdd FILL
XFILL_5__9676_ gnd vdd FILL
XFILL_5__13135_ gnd vdd FILL
XFILL_5_BUFX2_insert86 gnd vdd FILL
XFILL_3__14314_ gnd vdd FILL
XFILL_5__6888_ gnd vdd FILL
XFILL_3__11526_ gnd vdd FILL
XFILL_0__8982_ gnd vdd FILL
XFILL_3__7711_ gnd vdd FILL
XFILL_5_BUFX2_insert97 gnd vdd FILL
XFILL_1__12705_ gnd vdd FILL
XFILL_4__13865_ gnd vdd FILL
XFILL_3__15294_ gnd vdd FILL
XFILL_2__10167_ gnd vdd FILL
XBUFX2_insert670 _12345_/Y gnd _8567_/A vdd BUFX2
XFILL_0__14134_ gnd vdd FILL
XFILL_0__11346_ gnd vdd FILL
XFILL_2__9898_ gnd vdd FILL
XSFILL19000x70050 gnd vdd FILL
XFILL_1__13685_ gnd vdd FILL
XBUFX2_insert681 _15005_/Y gnd _16306_/A vdd BUFX2
XFILL_5__8627_ gnd vdd FILL
XFILL_1__10897_ gnd vdd FILL
XFILL_0__7933_ gnd vdd FILL
X_16329_ _16329_/A gnd _16328_/Y gnd _16329_/Y vdd OAI21X1
XFILL_4__15604_ gnd vdd FILL
XFILL_3__14245_ gnd vdd FILL
XFILL_5__10278_ gnd vdd FILL
X_9260_ _9320_/Q gnd _9262_/A vdd INVX1
XBUFX2_insert692 _13362_/Y gnd _10539_/B vdd BUFX2
XFILL_1__15424_ gnd vdd FILL
XFILL_3__11457_ gnd vdd FILL
XFILL_1__12636_ gnd vdd FILL
XFILL_4__13796_ gnd vdd FILL
XFILL_0__14065_ gnd vdd FILL
XFILL_2__14975_ gnd vdd FILL
XFILL_2__8849_ gnd vdd FILL
XFILL_0__11277_ gnd vdd FILL
XSFILL38840x12050 gnd vdd FILL
XFILL_5__12017_ gnd vdd FILL
X_8211_ _8209_/Y _8244_/B _8211_/C gnd _8287_/D vdd OAI21X1
XFILL_3__10408_ gnd vdd FILL
XSFILL64120x45050 gnd vdd FILL
XFILL_4__15535_ gnd vdd FILL
XFILL_0__7864_ gnd vdd FILL
X_9191_ _9191_/Q _8551_/CLK _9064_/R vdd _9131_/Y gnd vdd DFFSR
XFILL_4__12747_ gnd vdd FILL
XFILL_0__13016_ gnd vdd FILL
XFILL_3__14176_ gnd vdd FILL
XFILL_2__13926_ gnd vdd FILL
XFILL_1__15355_ gnd vdd FILL
XFILL_3__7573_ gnd vdd FILL
XFILL_3__11388_ gnd vdd FILL
XFILL_1__12567_ gnd vdd FILL
XFILL_0__9603_ gnd vdd FILL
XFILL_5__7509_ gnd vdd FILL
XFILL_5__8489_ gnd vdd FILL
X_8142_ _8142_/A _7502_/B gnd _8143_/C vdd NAND2X1
XFILL_3__13127_ gnd vdd FILL
XFILL_4__15466_ gnd vdd FILL
XFILL_1__14306_ gnd vdd FILL
XFILL_2__13857_ gnd vdd FILL
XFILL_1__11518_ gnd vdd FILL
XFILL_0__10159_ gnd vdd FILL
XFILL_1__15286_ gnd vdd FILL
XFILL_0__9534_ gnd vdd FILL
XFILL_1__12498_ gnd vdd FILL
X_8073_ _8142_/A _6921_/B gnd _8074_/C vdd NAND2X1
XSFILL3560x52050 gnd vdd FILL
XFILL_4__14417_ gnd vdd FILL
XFILL_3__9243_ gnd vdd FILL
XFILL_4__11629_ gnd vdd FILL
XFILL_5__13968_ gnd vdd FILL
XFILL_4__15397_ gnd vdd FILL
XFILL_1__14237_ gnd vdd FILL
XFILL_2__13788_ gnd vdd FILL
XFILL_1__11449_ gnd vdd FILL
XFILL_5__15707_ gnd vdd FILL
X_7024_ _6980_/A _9328_/CLK _7152_/R vdd _7024_/D gnd vdd DFFSR
XFILL_0__14967_ gnd vdd FILL
XFILL_3__12009_ gnd vdd FILL
XFILL_0__9465_ gnd vdd FILL
XFILL_2__15527_ gnd vdd FILL
XFILL_4__14348_ gnd vdd FILL
XFILL_2__12739_ gnd vdd FILL
XSFILL44040x12050 gnd vdd FILL
XFILL_5__13899_ gnd vdd FILL
XFILL_1__14168_ gnd vdd FILL
XFILL_0__13918_ gnd vdd FILL
XFILL_5__15638_ gnd vdd FILL
XFILL_0__14898_ gnd vdd FILL
XFILL_3__8125_ gnd vdd FILL
XFILL_0__9396_ gnd vdd FILL
XFILL_1__13119_ gnd vdd FILL
XFILL_2__15458_ gnd vdd FILL
XFILL_4__14279_ gnd vdd FILL
XFILL_0__13849_ gnd vdd FILL
XFILL_1__14099_ gnd vdd FILL
XFILL_4__16018_ gnd vdd FILL
XFILL_0__8347_ gnd vdd FILL
XFILL_5__15569_ gnd vdd FILL
XFILL_2__14409_ gnd vdd FILL
X_8975_ _8969_/A _7439_/B gnd _8975_/Y vdd NAND2X1
XFILL_3__8056_ gnd vdd FILL
XFILL_2__15389_ gnd vdd FILL
X_7926_ _8022_/Q gnd _7928_/A vdd INVX1
XFILL_1__7071_ gnd vdd FILL
XFILL_0__15519_ gnd vdd FILL
XSFILL64200x25050 gnd vdd FILL
XFILL_0__7229_ gnd vdd FILL
XFILL_4__7820_ gnd vdd FILL
X_7857_ _7857_/A _7878_/B _7856_/Y gnd _7913_/D vdd OAI21X1
XFILL_0_CLKBUF1_insert204 gnd vdd FILL
XFILL_0_CLKBUF1_insert215 gnd vdd FILL
X_7788_ _7736_/A _9958_/CLK _7270_/R vdd _7738_/Y gnd vdd DFFSR
XFILL_4__7751_ gnd vdd FILL
XSFILL3640x32050 gnd vdd FILL
XSFILL28760x50 gnd vdd FILL
XFILL_3__8958_ gnd vdd FILL
XFILL_1_BUFX2_insert1008 gnd vdd FILL
X_9527_ _9525_/Y _9551_/B _9527_/C gnd _9579_/D vdd OAI21X1
XFILL_1_BUFX2_insert1019 gnd vdd FILL
XFILL_1__7973_ gnd vdd FILL
XFILL_4__7682_ gnd vdd FILL
XSFILL28040x25050 gnd vdd FILL
XSFILL79480x79050 gnd vdd FILL
XFILL_3__8889_ gnd vdd FILL
XSFILL94280x20050 gnd vdd FILL
XSFILL54120x77050 gnd vdd FILL
XFILL_1__6924_ gnd vdd FILL
XFILL_4__9421_ gnd vdd FILL
X_9458_ _9418_/A _8562_/CLK _9430_/R vdd _9458_/D gnd vdd DFFSR
X_10340_ _14135_/C _8541_/CLK _7258_/R vdd _10340_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert700 gnd vdd FILL
X_8409_ _8409_/Q _9817_/CLK _8942_/R vdd _8409_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert711 gnd vdd FILL
XFILL_1__9643_ gnd vdd FILL
XFILL_1__6855_ gnd vdd FILL
XFILL_4__9352_ gnd vdd FILL
X_9389_ _9372_/B _7853_/B gnd _9389_/Y vdd NAND2X1
XFILL_4_BUFX2_insert722 gnd vdd FILL
XFILL_4_BUFX2_insert733 gnd vdd FILL
XFILL_4_BUFX2_insert744 gnd vdd FILL
XSFILL33960x35050 gnd vdd FILL
XFILL_4_BUFX2_insert755 gnd vdd FILL
X_10271_ _10269_/Y _10271_/B _10271_/C gnd _10271_/Y vdd OAI21X1
XFILL_4_BUFX2_insert766 gnd vdd FILL
XFILL_3_CLKBUF1_insert1076 gnd vdd FILL
XFILL_4_BUFX2_insert777 gnd vdd FILL
X_12010_ _12010_/A _12010_/B _12010_/C gnd _13095_/B vdd NAND3X1
XFILL_4__9283_ gnd vdd FILL
XFILL_6__9219_ gnd vdd FILL
XFILL_4_BUFX2_insert788 gnd vdd FILL
XFILL_4_BUFX2_insert799 gnd vdd FILL
XFILL_1__8525_ gnd vdd FILL
XFILL_4__8234_ gnd vdd FILL
XFILL_1__8456_ gnd vdd FILL
X_13961_ _7316_/A _14738_/A _14909_/C _7060_/A gnd _13963_/A vdd AOI22X1
XFILL_4__7116_ gnd vdd FILL
XFILL_2__7180_ gnd vdd FILL
XFILL_1__8387_ gnd vdd FILL
X_15700_ _14257_/Y _15169_/A gnd _15702_/C vdd NOR2X1
X_12912_ _12910_/Y vdd _12912_/C gnd _12948_/D vdd OAI21X1
XFILL_4__8096_ gnd vdd FILL
XSFILL93720x34050 gnd vdd FILL
XFILL_1__7338_ gnd vdd FILL
X_13892_ _13892_/A gnd _15436_/C vdd INVX1
XSFILL79560x59050 gnd vdd FILL
XFILL_4__7047_ gnd vdd FILL
X_15631_ _7328_/A _15631_/B _15636_/B gnd _15632_/C vdd NAND3X1
X_12843_ _12843_/A vdd _12843_/C gnd _12925_/D vdd OAI21X1
XFILL_1_BUFX2_insert601 gnd vdd FILL
XFILL_1_BUFX2_insert612 gnd vdd FILL
XSFILL79160x61050 gnd vdd FILL
XFILL_1_BUFX2_insert623 gnd vdd FILL
XFILL_5__7860_ gnd vdd FILL
XFILL_1_BUFX2_insert634 gnd vdd FILL
X_15562_ _14025_/Y _15392_/B _15328_/B _15562_/D gnd _15564_/A vdd OAI22X1
XFILL_1__9008_ gnd vdd FILL
XSFILL13640x9050 gnd vdd FILL
X_12774_ _12789_/A memoryOutData[26] gnd _12775_/C vdd NAND2X1
XFILL_1_BUFX2_insert645 gnd vdd FILL
XFILL_1_BUFX2_insert656 gnd vdd FILL
XFILL_3__10690_ gnd vdd FILL
X_14513_ _16439_/Q gnd _14513_/Y vdd INVX1
XFILL_1_BUFX2_insert667 gnd vdd FILL
X_11725_ _11720_/A _11726_/B _11835_/C gnd _11725_/Y vdd AOI21X1
XFILL_5__11250_ gnd vdd FILL
XFILL_1_BUFX2_insert678 gnd vdd FILL
XFILL_4__8998_ gnd vdd FILL
XFILL_1_BUFX2_insert689 gnd vdd FILL
X_15493_ _15842_/A _15493_/B _15491_/Y _16137_/C gnd _15494_/B vdd OAI22X1
XFILL_4__11980_ gnd vdd FILL
XFILL_1__10820_ gnd vdd FILL
XFILL_2__11070_ gnd vdd FILL
XSFILL18840x76050 gnd vdd FILL
XFILL_5__9530_ gnd vdd FILL
XFILL_4__7949_ gnd vdd FILL
X_14444_ _14444_/A _14045_/A _14894_/B _15875_/D gnd _14444_/Y vdd OAI22X1
X_11656_ _11649_/Y _11656_/B gnd _11656_/Y vdd NOR2X1
XFILL_5__11181_ gnd vdd FILL
XFILL_4__10931_ gnd vdd FILL
XFILL_2__10021_ gnd vdd FILL
XFILL_2__9752_ gnd vdd FILL
XFILL_3__12360_ gnd vdd FILL
XFILL_0__11200_ gnd vdd FILL
XFILL_2__6964_ gnd vdd FILL
XFILL_1__10751_ gnd vdd FILL
XFILL_0__12180_ gnd vdd FILL
XFILL_5__10132_ gnd vdd FILL
X_10607_ _16072_/A _7156_/CLK _7775_/R vdd _10607_/D gnd vdd DFFSR
X_14375_ _9321_/Q _13854_/B _14481_/C _6959_/A gnd _14379_/A vdd AOI22X1
XFILL_3__11311_ gnd vdd FILL
XFILL_2__8703_ gnd vdd FILL
XFILL_4__13650_ gnd vdd FILL
X_11587_ _11587_/A _11150_/Y _11587_/C gnd _11587_/Y vdd OAI21X1
XFILL_2__9683_ gnd vdd FILL
XFILL_3__12291_ gnd vdd FILL
XSFILL59000x8050 gnd vdd FILL
XFILL_0__11131_ gnd vdd FILL
XFILL_1__13470_ gnd vdd FILL
XFILL_1__10682_ gnd vdd FILL
X_16114_ _7876_/A gnd _16114_/Y vdd INVX1
XFILL_2__6895_ gnd vdd FILL
XFILL_4__9619_ gnd vdd FILL
X_13326_ _13326_/A _13326_/B gnd _13326_/Y vdd NOR2X1
XFILL_5__9392_ gnd vdd FILL
XFILL_4__12601_ gnd vdd FILL
XFILL_5__10063_ gnd vdd FILL
XFILL_3__14030_ gnd vdd FILL
XFILL_5__14940_ gnd vdd FILL
X_10538_ _10539_/B _9770_/B gnd _10538_/Y vdd NAND2X1
XFILL_2__8634_ gnd vdd FILL
XSFILL38760x27050 gnd vdd FILL
XFILL_3__11242_ gnd vdd FILL
XFILL_1__12421_ gnd vdd FILL
XFILL112280x34050 gnd vdd FILL
XFILL_4__10793_ gnd vdd FILL
XFILL_4__13581_ gnd vdd FILL
XFILL_2__14760_ gnd vdd FILL
XFILL_2__11972_ gnd vdd FILL
XFILL_5__8343_ gnd vdd FILL
XFILL_0__11062_ gnd vdd FILL
X_16045_ _16044_/Y _16022_/Y _16045_/C gnd _16046_/B vdd NOR3X1
X_13257_ _13231_/A _13288_/B gnd _13270_/A vdd NAND2X1
XFILL_4__15320_ gnd vdd FILL
XFILL_5__14871_ gnd vdd FILL
X_10469_ _10469_/Q _7406_/CLK _9692_/R vdd _10405_/Y gnd vdd DFFSR
XFILL_4__12532_ gnd vdd FILL
XFILL_2__13711_ gnd vdd FILL
XFILL_2__10923_ gnd vdd FILL
XFILL_0__10013_ gnd vdd FILL
XFILL_1__15140_ gnd vdd FILL
XFILL_3__11173_ gnd vdd FILL
XFILL_1__12352_ gnd vdd FILL
XFILL_2__14691_ gnd vdd FILL
X_12208_ _13172_/A gnd _12210_/A vdd INVX1
XSFILL74200x2050 gnd vdd FILL
XFILL_5__8274_ gnd vdd FILL
XFILL_0__15870_ gnd vdd FILL
XFILL_5__13822_ gnd vdd FILL
XSFILL113800x2050 gnd vdd FILL
XFILL_3__10124_ gnd vdd FILL
XFILL_4__15251_ gnd vdd FILL
XFILL_4__12463_ gnd vdd FILL
XFILL_0__7580_ gnd vdd FILL
X_13188_ _13188_/Q _13180_/CLK _13180_/R vdd _13188_/D gnd vdd DFFSR
XFILL_2__13642_ gnd vdd FILL
XSFILL79240x41050 gnd vdd FILL
XFILL_1__11303_ gnd vdd FILL
XSFILL43880x18050 gnd vdd FILL
XFILL_3__15981_ gnd vdd FILL
XFILL_0__14821_ gnd vdd FILL
XFILL_1__15071_ gnd vdd FILL
XFILL_5__7225_ gnd vdd FILL
XFILL_2__8496_ gnd vdd FILL
XSFILL3480x67050 gnd vdd FILL
XFILL_1__12283_ gnd vdd FILL
XFILL_4__14202_ gnd vdd FILL
X_12139_ _13103_/A gnd _12139_/Y vdd INVX1
XFILL_4__11414_ gnd vdd FILL
XFILL_5__13753_ gnd vdd FILL
XFILL_5__10965_ gnd vdd FILL
XFILL_4__15182_ gnd vdd FILL
XFILL_1__14022_ gnd vdd FILL
XFILL_2__7447_ gnd vdd FILL
XFILL_4__12394_ gnd vdd FILL
XFILL_3__14932_ gnd vdd FILL
XFILL_2__16361_ gnd vdd FILL
XFILL_3__10055_ gnd vdd FILL
XSFILL28680x79050 gnd vdd FILL
XFILL_2_CLKBUF1_insert170 gnd vdd FILL
XFILL_2__13573_ gnd vdd FILL
XFILL_1__11234_ gnd vdd FILL
XSFILL114440x50050 gnd vdd FILL
XFILL_2__10785_ gnd vdd FILL
XFILL_0__14752_ gnd vdd FILL
XFILL_2_CLKBUF1_insert181 gnd vdd FILL
XFILL_5__12704_ gnd vdd FILL
XFILL_0__9250_ gnd vdd FILL
XFILL_0__11964_ gnd vdd FILL
XFILL_2_CLKBUF1_insert192 gnd vdd FILL
XFILL_2__15312_ gnd vdd FILL
XFILL_4__14133_ gnd vdd FILL
XFILL_4__11345_ gnd vdd FILL
XFILL_5__13684_ gnd vdd FILL
XFILL_2__12524_ gnd vdd FILL
XFILL_3__14863_ gnd vdd FILL
XFILL_5__10896_ gnd vdd FILL
XFILL_2__16292_ gnd vdd FILL
XFILL_1__11165_ gnd vdd FILL
XFILL_0__13703_ gnd vdd FILL
XFILL_2__7378_ gnd vdd FILL
XFILL_0__10915_ gnd vdd FILL
XFILL_0__8201_ gnd vdd FILL
XFILL_5__7087_ gnd vdd FILL
XFILL_0__14683_ gnd vdd FILL
XFILL_5__15423_ gnd vdd FILL
XFILL_5__12635_ gnd vdd FILL
XSFILL59000x49050 gnd vdd FILL
XFILL_0__11895_ gnd vdd FILL
XFILL_4__14064_ gnd vdd FILL
XFILL_2__9117_ gnd vdd FILL
XFILL_3__13814_ gnd vdd FILL
XFILL_1__10116_ gnd vdd FILL
XFILL_2__15243_ gnd vdd FILL
XFILL_4__11276_ gnd vdd FILL
XFILL_2__12455_ gnd vdd FILL
XFILL_0__13634_ gnd vdd FILL
XFILL_1__15973_ gnd vdd FILL
XSFILL99400x54050 gnd vdd FILL
XFILL_3__14794_ gnd vdd FILL
XFILL_1__11096_ gnd vdd FILL
XFILL_4__13015_ gnd vdd FILL
XBUFX2_insert3 _12381_/Y gnd _9371_/B vdd BUFX2
XFILL_0__8132_ gnd vdd FILL
XFILL_6__13925_ gnd vdd FILL
XFILL_5__15354_ gnd vdd FILL
X_15829_ _15632_/A _15829_/B _15829_/C gnd _15829_/Y vdd OAI21X1
X_8760_ _8760_/A gnd _8760_/Y vdd INVX1
XFILL_2__11406_ gnd vdd FILL
XFILL_3__10957_ gnd vdd FILL
XFILL_2__15174_ gnd vdd FILL
XFILL_1__10047_ gnd vdd FILL
XFILL_3__13745_ gnd vdd FILL
XFILL_3__9930_ gnd vdd FILL
XFILL_2_BUFX2_insert490 gnd vdd FILL
XFILL_1__14924_ gnd vdd FILL
XFILL_2__12386_ gnd vdd FILL
XFILL_0__16353_ gnd vdd FILL
XFILL_0__10777_ gnd vdd FILL
XFILL_5__14305_ gnd vdd FILL
XFILL_0__13565_ gnd vdd FILL
XFILL_0__8063_ gnd vdd FILL
XFILL_5__11517_ gnd vdd FILL
XFILL_6_BUFX2_insert817 gnd vdd FILL
X_7711_ _7711_/A _7753_/B _7711_/C gnd _7711_/Y vdd OAI21X1
XFILL112360x14050 gnd vdd FILL
XFILL_2__14125_ gnd vdd FILL
XFILL_4__10158_ gnd vdd FILL
XFILL_5__15285_ gnd vdd FILL
X_8691_ _8653_/A _8429_/CLK _9062_/R vdd _8691_/D gnd vdd DFFSR
XFILL_0__15304_ gnd vdd FILL
XFILL_3__13676_ gnd vdd FILL
XFILL_5__12497_ gnd vdd FILL
XFILL_2__11337_ gnd vdd FILL
XFILL_1__14855_ gnd vdd FILL
XFILL_0__12516_ gnd vdd FILL
XFILL_3__10888_ gnd vdd FILL
XFILL_3__9861_ gnd vdd FILL
XSFILL79720x19050 gnd vdd FILL
XFILL_0__16284_ gnd vdd FILL
XFILL_5__14236_ gnd vdd FILL
XFILL_0__13496_ gnd vdd FILL
XFILL_5__7989_ gnd vdd FILL
XFILL_3__12627_ gnd vdd FILL
XFILL_6__13787_ gnd vdd FILL
X_7642_ _7554_/A _7642_/CLK _9306_/R vdd _7642_/D gnd vdd DFFSR
XFILL_5__11448_ gnd vdd FILL
XFILL_3__15415_ gnd vdd FILL
XFILL_1__13806_ gnd vdd FILL
XFILL_2__14056_ gnd vdd FILL
XFILL_4__14966_ gnd vdd FILL
XFILL_3__16395_ gnd vdd FILL
XFILL_3__9792_ gnd vdd FILL
XFILL_0__15235_ gnd vdd FILL
XFILL_2__11268_ gnd vdd FILL
XFILL_5__9728_ gnd vdd FILL
XFILL_0__12447_ gnd vdd FILL
XFILL_6__15526_ gnd vdd FILL
XFILL_6__8521_ gnd vdd FILL
XFILL_1__14786_ gnd vdd FILL
XFILL_6__12738_ gnd vdd FILL
XSFILL49080x60050 gnd vdd FILL
XFILL_1__11998_ gnd vdd FILL
XFILL_5__14167_ gnd vdd FILL
XFILL_2__13007_ gnd vdd FILL
XFILL_4__13917_ gnd vdd FILL
XFILL_3__15346_ gnd vdd FILL
X_7573_ _7570_/A _6933_/B gnd _7574_/C vdd NAND2X1
XFILL_5__11379_ gnd vdd FILL
XFILL_3__8743_ gnd vdd FILL
XFILL_1__13737_ gnd vdd FILL
XFILL_4__14897_ gnd vdd FILL
XFILL_1__10949_ gnd vdd FILL
XFILL_0__12378_ gnd vdd FILL
XFILL_0__15166_ gnd vdd FILL
XFILL_2__11199_ gnd vdd FILL
XFILL_5__9659_ gnd vdd FILL
XFILL_5__13118_ gnd vdd FILL
X_9312_ _9312_/Q _8433_/CLK _7921_/R vdd _9312_/D gnd vdd DFFSR
XSFILL28760x59050 gnd vdd FILL
XFILL_0__8965_ gnd vdd FILL
XFILL_3__11509_ gnd vdd FILL
XFILL_4__13848_ gnd vdd FILL
XSFILL114520x30050 gnd vdd FILL
XFILL_5__14098_ gnd vdd FILL
XFILL_3__15277_ gnd vdd FILL
XFILL_3__12489_ gnd vdd FILL
XFILL_0__14117_ gnd vdd FILL
XFILL_0__11329_ gnd vdd FILL
XFILL_1__13668_ gnd vdd FILL
XFILL_0__15097_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1082 gnd vdd FILL
XFILL_6__15388_ gnd vdd FILL
XFILL_3__14228_ gnd vdd FILL
X_9243_ _9208_/B _9371_/B gnd _9243_/Y vdd NAND2X1
XFILL_0__8896_ gnd vdd FILL
XFILL_1__15407_ gnd vdd FILL
XFILL_3__7625_ gnd vdd FILL
XFILL_1__12619_ gnd vdd FILL
XFILL_4__13779_ gnd vdd FILL
XFILL_1__16387_ gnd vdd FILL
XFILL_0__14048_ gnd vdd FILL
XFILL_2__14958_ gnd vdd FILL
XFILL_1__13599_ gnd vdd FILL
XFILL_6__14339_ gnd vdd FILL
XFILL_0__7847_ gnd vdd FILL
XSFILL103560x54050 gnd vdd FILL
XFILL_4__15518_ gnd vdd FILL
XSFILL69240x73050 gnd vdd FILL
XFILL_3__14159_ gnd vdd FILL
X_9174_ _9078_/A _8022_/CLK _8674_/R vdd _9174_/D gnd vdd DFFSR
XFILL_3__7556_ gnd vdd FILL
XFILL_1__15338_ gnd vdd FILL
XFILL_2__13909_ gnd vdd FILL
XFILL_2__14889_ gnd vdd FILL
X_8125_ _8123_/Y _8079_/A _8125_/C gnd _8173_/D vdd OAI21X1
XFILL_3_BUFX2_insert707 gnd vdd FILL
XFILL_4__15449_ gnd vdd FILL
XFILL_3_BUFX2_insert718 gnd vdd FILL
XFILL_3__7487_ gnd vdd FILL
XFILL_3_BUFX2_insert729 gnd vdd FILL
XFILL_1__15269_ gnd vdd FILL
XSFILL104440x82050 gnd vdd FILL
XFILL_1__8310_ gnd vdd FILL
XFILL_0__9517_ gnd vdd FILL
XFILL_0__15999_ gnd vdd FILL
XFILL_3__9226_ gnd vdd FILL
X_8056_ _8054_/Y _8100_/A _8055_/Y gnd _8150_/D vdd OAI21X1
XFILL_1__9290_ gnd vdd FILL
XSFILL8680x80050 gnd vdd FILL
XFILL_1_BUFX2_insert40 gnd vdd FILL
XFILL_1_BUFX2_insert51 gnd vdd FILL
X_7007_ _7007_/Q _7007_/CLK _9332_/R vdd _7007_/D gnd vdd DFFSR
XFILL_1__8241_ gnd vdd FILL
XFILL_1_BUFX2_insert62 gnd vdd FILL
XFILL_1_BUFX2_insert73 gnd vdd FILL
XFILL_3__9157_ gnd vdd FILL
XFILL_1_BUFX2_insert84 gnd vdd FILL
XFILL_1_BUFX2_insert95 gnd vdd FILL
XSFILL3640x27050 gnd vdd FILL
XFILL_0__9379_ gnd vdd FILL
XFILL_3__8108_ gnd vdd FILL
XFILL_3__9088_ gnd vdd FILL
XSFILL28840x39050 gnd vdd FILL
XFILL_6__9906_ gnd vdd FILL
XFILL_1__7123_ gnd vdd FILL
XSFILL114600x10050 gnd vdd FILL
XSFILL94280x15050 gnd vdd FILL
X_8958_ _8956_/Y _9005_/A _8958_/C gnd _9048_/D vdd OAI21X1
XSFILL13640x81050 gnd vdd FILL
XFILL_1__7054_ gnd vdd FILL
X_7909_ _7909_/Q _7781_/CLK _8670_/R vdd _7909_/D gnd vdd DFFSR
X_8889_ _8893_/B _8889_/B gnd _8889_/Y vdd NAND2X1
XFILL_4__8852_ gnd vdd FILL
XSFILL69000x3050 gnd vdd FILL
XFILL_0_BUFX2_insert608 gnd vdd FILL
XFILL_4__7803_ gnd vdd FILL
XFILL_0_BUFX2_insert619 gnd vdd FILL
X_11510_ _11513_/B _11574_/B _11510_/C gnd _11510_/Y vdd OAI21X1
XFILL_4__8783_ gnd vdd FILL
X_12490_ _12055_/B gnd _12492_/A vdd INVX1
XSFILL34040x39050 gnd vdd FILL
XFILL_4__7734_ gnd vdd FILL
XSFILL8760x60050 gnd vdd FILL
X_11441_ _11439_/Y _11440_/Y _11204_/Y gnd _11441_/Y vdd OAI21X1
XFILL_1__7956_ gnd vdd FILL
X_14160_ _14160_/A _14160_/B _14849_/B _15642_/D gnd _14161_/B vdd OAI22X1
XFILL_1__6907_ gnd vdd FILL
X_11372_ _11008_/Y gnd _11377_/B vdd INVX1
XFILL_1__7887_ gnd vdd FILL
XFILL_4__9404_ gnd vdd FILL
X_13111_ _13111_/A _13108_/B _13110_/Y gnd _13111_/Y vdd OAI21X1
XFILL_4_BUFX2_insert530 gnd vdd FILL
XFILL_4__7596_ gnd vdd FILL
X_10323_ _14956_/B gnd _10323_/Y vdd INVX1
X_14091_ _14091_/A _13868_/B _14456_/C _14089_/Y gnd _14092_/B vdd OAI22X1
XFILL_1__6838_ gnd vdd FILL
XFILL_1__9626_ gnd vdd FILL
XFILL_4_BUFX2_insert541 gnd vdd FILL
XFILL_4_BUFX2_insert552 gnd vdd FILL
XFILL_4_BUFX2_insert563 gnd vdd FILL
XFILL_4__9335_ gnd vdd FILL
XFILL_4_BUFX2_insert574 gnd vdd FILL
X_13042_ vdd _13042_/B gnd _13042_/Y vdd NAND2X1
X_10254_ _10334_/Q gnd _10254_/Y vdd INVX1
XFILL_1__9557_ gnd vdd FILL
XFILL_4_BUFX2_insert585 gnd vdd FILL
XFILL_2__8350_ gnd vdd FILL
XSFILL13720x61050 gnd vdd FILL
XSFILL94600x57050 gnd vdd FILL
XFILL_4_BUFX2_insert596 gnd vdd FILL
XFILL_4__9266_ gnd vdd FILL
XSFILL79160x56050 gnd vdd FILL
XFILL_1__8508_ gnd vdd FILL
XFILL_2__7301_ gnd vdd FILL
X_10185_ _10185_/A _10160_/A _10185_/C gnd _10225_/D vdd OAI21X1
XFILL_1__9488_ gnd vdd FILL
XFILL_4__8217_ gnd vdd FILL
XFILL_2__7232_ gnd vdd FILL
XFILL_1__8439_ gnd vdd FILL
XFILL_5__10750_ gnd vdd FILL
X_14993_ _14993_/A _15386_/C _15322_/A _13441_/Y gnd _14994_/A vdd OAI22X1
XFILL_2__10570_ gnd vdd FILL
XFILL_4__8148_ gnd vdd FILL
XSFILL84280x47050 gnd vdd FILL
XFILL_3_CLKBUF1_insert210 gnd vdd FILL
XFILL_4__11130_ gnd vdd FILL
XFILL_3_CLKBUF1_insert221 gnd vdd FILL
X_13944_ _7572_/A gnd _13944_/Y vdd INVX1
XFILL_5__10681_ gnd vdd FILL
XFILL_3__11860_ gnd vdd FILL
XFILL_2__7163_ gnd vdd FILL
XFILL_0__10700_ gnd vdd FILL
XFILL_4__8079_ gnd vdd FILL
XFILL_0__11680_ gnd vdd FILL
XFILL_5__8961_ gnd vdd FILL
XFILL_5__12420_ gnd vdd FILL
XFILL_3__10811_ gnd vdd FILL
XSFILL99320x69050 gnd vdd FILL
X_13875_ _9102_/A gnd _13875_/Y vdd INVX1
XFILL_4__11061_ gnd vdd FILL
XSFILL59080x23050 gnd vdd FILL
XFILL_2__12240_ gnd vdd FILL
XFILL_2__7094_ gnd vdd FILL
XFILL_0__10631_ gnd vdd FILL
XFILL_3__11791_ gnd vdd FILL
XFILL_1__12970_ gnd vdd FILL
XFILL_6__13710_ gnd vdd FILL
X_15614_ _16225_/C _15614_/B _15726_/A _15614_/D gnd _15615_/B vdd OAI22X1
XFILL_4__10012_ gnd vdd FILL
XFILL_1_BUFX2_insert420 gnd vdd FILL
X_12826_ _12119_/B gnd _12826_/Y vdd INVX1
XFILL_5__8892_ gnd vdd FILL
XFILL_5__12351_ gnd vdd FILL
XFILL_3__13530_ gnd vdd FILL
XFILL_1_BUFX2_insert431 gnd vdd FILL
XFILL_3__10742_ gnd vdd FILL
XFILL_1_BUFX2_insert442 gnd vdd FILL
XFILL_1__11921_ gnd vdd FILL
XFILL_2__12171_ gnd vdd FILL
XFILL_1_BUFX2_insert453 gnd vdd FILL
XFILL_0__13350_ gnd vdd FILL
XFILL112280x29050 gnd vdd FILL
XFILL_0__10562_ gnd vdd FILL
XFILL_5__7843_ gnd vdd FILL
XFILL_5__11302_ gnd vdd FILL
XFILL_1_BUFX2_insert464 gnd vdd FILL
X_12757_ _12755_/Y _12723_/A _12757_/C gnd _12757_/Y vdd OAI21X1
XFILL_4__14820_ gnd vdd FILL
XFILL_5__15070_ gnd vdd FILL
XFILL_1_BUFX2_insert475 gnd vdd FILL
X_15545_ _15545_/A _15356_/C _15545_/C gnd _15548_/C vdd AOI21X1
XFILL_3__13461_ gnd vdd FILL
XFILL_5__12282_ gnd vdd FILL
XFILL_2__11122_ gnd vdd FILL
XFILL_1__14640_ gnd vdd FILL
XFILL_3__10673_ gnd vdd FILL
XFILL_0__12301_ gnd vdd FILL
XFILL_1_BUFX2_insert486 gnd vdd FILL
XFILL_0__13281_ gnd vdd FILL
XFILL_1_BUFX2_insert497 gnd vdd FILL
XFILL_1__11852_ gnd vdd FILL
XFILL_5__14021_ gnd vdd FILL
XFILL_6__16360_ gnd vdd FILL
X_11708_ _11573_/C _11275_/A _11708_/C gnd _11708_/Y vdd OAI21X1
XFILL_0__10493_ gnd vdd FILL
XFILL_3__12412_ gnd vdd FILL
XFILL_3__15200_ gnd vdd FILL
XFILL_6__13572_ gnd vdd FILL
X_15476_ _16309_/A _15476_/B _15476_/C _16306_/C gnd _15477_/C vdd OAI22X1
XFILL_5__11233_ gnd vdd FILL
X_12688_ _12642_/A _8171_/CLK _8171_/R vdd _12688_/D gnd vdd DFFSR
XFILL_2__9804_ gnd vdd FILL
XFILL_3__16180_ gnd vdd FILL
XFILL_4__14751_ gnd vdd FILL
XFILL_3__13392_ gnd vdd FILL
XFILL_2__15930_ gnd vdd FILL
XFILL_0__15020_ gnd vdd FILL
XFILL_4__11963_ gnd vdd FILL
XFILL_0__12232_ gnd vdd FILL
XFILL_2__11053_ gnd vdd FILL
XFILL_1__10803_ gnd vdd FILL
XFILL_1__14571_ gnd vdd FILL
XFILL_6__15311_ gnd vdd FILL
XFILL_2__7996_ gnd vdd FILL
XFILL_5__9513_ gnd vdd FILL
X_14427_ _9066_/Q gnd _15884_/B vdd INVX1
XFILL_1__11783_ gnd vdd FILL
XFILL_5__11164_ gnd vdd FILL
X_11639_ _11385_/Y _11379_/Y _11055_/Y gnd _11639_/Y vdd AOI21X1
XFILL_4__13702_ gnd vdd FILL
XFILL_3__15131_ gnd vdd FILL
XFILL_4__10914_ gnd vdd FILL
XFILL_3__12343_ gnd vdd FILL
XFILL_1__16310_ gnd vdd FILL
XFILL_2__10004_ gnd vdd FILL
XFILL_2__6947_ gnd vdd FILL
XFILL_4__14682_ gnd vdd FILL
XFILL_2__9735_ gnd vdd FILL
XFILL_1__13522_ gnd vdd FILL
XFILL_4__11894_ gnd vdd FILL
XFILL_0__12163_ gnd vdd FILL
XSFILL69160x9050 gnd vdd FILL
XFILL_2__15861_ gnd vdd FILL
XFILL_5__10115_ gnd vdd FILL
XSFILL114440x45050 gnd vdd FILL
XFILL_6__12454_ gnd vdd FILL
XFILL_0__8750_ gnd vdd FILL
X_14358_ _14358_/A _14358_/B _14739_/C _15837_/A gnd _14358_/Y vdd AOI22X1
XFILL_5__15972_ gnd vdd FILL
XFILL_4__13633_ gnd vdd FILL
XFILL_3__15062_ gnd vdd FILL
XFILL_5__11095_ gnd vdd FILL
XFILL_1__16241_ gnd vdd FILL
XFILL_2__14812_ gnd vdd FILL
XFILL_3__12274_ gnd vdd FILL
XFILL_0__11114_ gnd vdd FILL
XFILL_1__13453_ gnd vdd FILL
XFILL_2__15792_ gnd vdd FILL
XSFILL84360x27050 gnd vdd FILL
XFILL_2__9666_ gnd vdd FILL
XFILL_2__6878_ gnd vdd FILL
X_13309_ _13297_/C _13308_/Y gnd _13309_/Y vdd NOR2X1
XFILL_0__12094_ gnd vdd FILL
XFILL_1__10665_ gnd vdd FILL
XFILL_0__7701_ gnd vdd FILL
XFILL_6__11405_ gnd vdd FILL
XFILL_5__10046_ gnd vdd FILL
XFILL_6__15173_ gnd vdd FILL
XFILL_3__14013_ gnd vdd FILL
XFILL_5__9375_ gnd vdd FILL
XFILL_5__14923_ gnd vdd FILL
X_14289_ _15747_/A _14344_/B _13884_/C _14289_/D gnd _14298_/A vdd AOI22X1
XFILL_4__16352_ gnd vdd FILL
XFILL_3__11225_ gnd vdd FILL
XFILL_2__8617_ gnd vdd FILL
XFILL_1__12404_ gnd vdd FILL
XFILL_4__10776_ gnd vdd FILL
XFILL_2__14743_ gnd vdd FILL
XFILL_4__13564_ gnd vdd FILL
XFILL_0__15922_ gnd vdd FILL
XFILL_1__16172_ gnd vdd FILL
XFILL_2__11955_ gnd vdd FILL
XFILL_3__8390_ gnd vdd FILL
XFILL_2__9597_ gnd vdd FILL
XFILL_0__11045_ gnd vdd FILL
XFILL_6__14124_ gnd vdd FILL
XSFILL99400x49050 gnd vdd FILL
XFILL_1__13384_ gnd vdd FILL
XFILL_5__8326_ gnd vdd FILL
X_16028_ _9326_/Q gnd _16030_/A vdd INVX1
XFILL_4__15303_ gnd vdd FILL
XFILL_0__7632_ gnd vdd FILL
XFILL_5__14854_ gnd vdd FILL
XFILL_4__12515_ gnd vdd FILL
XFILL_2__10906_ gnd vdd FILL
XFILL_3__7341_ gnd vdd FILL
XFILL_3__11156_ gnd vdd FILL
XFILL_1__15123_ gnd vdd FILL
XFILL_4__16283_ gnd vdd FILL
XFILL_1__12335_ gnd vdd FILL
XFILL_2__14674_ gnd vdd FILL
XFILL_4__13495_ gnd vdd FILL
XFILL_2__11886_ gnd vdd FILL
XFILL_0__15853_ gnd vdd FILL
XFILL_5__8257_ gnd vdd FILL
XFILL_5__13805_ gnd vdd FILL
XFILL_0__7563_ gnd vdd FILL
XFILL_4__15234_ gnd vdd FILL
XFILL_3__10107_ gnd vdd FILL
XFILL_6__11267_ gnd vdd FILL
XFILL_2__13625_ gnd vdd FILL
XFILL_4__12446_ gnd vdd FILL
XFILL_2__16413_ gnd vdd FILL
XFILL_5__14785_ gnd vdd FILL
XFILL_0__14804_ gnd vdd FILL
XFILL_5__11997_ gnd vdd FILL
XFILL_1__15054_ gnd vdd FILL
XFILL_3__15964_ gnd vdd FILL
XFILL_2__8479_ gnd vdd FILL
XFILL_3__11087_ gnd vdd FILL
XFILL_2__10837_ gnd vdd FILL
XFILL_5__7208_ gnd vdd FILL
XFILL_1__12266_ gnd vdd FILL
XFILL_6__13006_ gnd vdd FILL
XFILL_0__15784_ gnd vdd FILL
XFILL_5__8188_ gnd vdd FILL
XSFILL74280x79050 gnd vdd FILL
XFILL_0__12996_ gnd vdd FILL
X_9930_ _9970_/Q gnd _9932_/A vdd INVX1
XSFILL109480x50 gnd vdd FILL
XFILL_5__13736_ gnd vdd FILL
XFILL_3__9011_ gnd vdd FILL
XFILL_5__10948_ gnd vdd FILL
XFILL_3__10038_ gnd vdd FILL
XFILL_2__16344_ gnd vdd FILL
XFILL_4__12377_ gnd vdd FILL
XFILL_1__14005_ gnd vdd FILL
XFILL_0__7494_ gnd vdd FILL
XSFILL89080x39050 gnd vdd FILL
XSFILL109400x34050 gnd vdd FILL
XFILL_4__15165_ gnd vdd FILL
XFILL_3__14915_ gnd vdd FILL
XFILL_2__13556_ gnd vdd FILL
XFILL_1__11217_ gnd vdd FILL
XFILL_2__10768_ gnd vdd FILL
XFILL_3__15895_ gnd vdd FILL
XFILL_0__14735_ gnd vdd FILL
XFILL_0__11947_ gnd vdd FILL
XFILL_1__12197_ gnd vdd FILL
XFILL_0__9233_ gnd vdd FILL
XSFILL49080x55050 gnd vdd FILL
XFILL_4__14116_ gnd vdd FILL
XFILL112200x73050 gnd vdd FILL
XFILL_5__13667_ gnd vdd FILL
XFILL_2__12507_ gnd vdd FILL
X_9861_ _9947_/Q gnd _9863_/A vdd INVX1
XFILL_4__11328_ gnd vdd FILL
XFILL_3__14846_ gnd vdd FILL
XFILL_5__10879_ gnd vdd FILL
XFILL_4__15096_ gnd vdd FILL
XFILL_2__16275_ gnd vdd FILL
XFILL_2__13487_ gnd vdd FILL
XFILL_1__11148_ gnd vdd FILL
XFILL_5__15406_ gnd vdd FILL
XFILL_2__10699_ gnd vdd FILL
XFILL_0__14666_ gnd vdd FILL
XFILL_5__12618_ gnd vdd FILL
XFILL_0__11878_ gnd vdd FILL
XFILL_0__9164_ gnd vdd FILL
X_8812_ _8760_/A _9958_/CLK _8929_/R vdd _8812_/D gnd vdd DFFSR
XFILL_5__16386_ gnd vdd FILL
XFILL_2__15226_ gnd vdd FILL
XFILL_4__14047_ gnd vdd FILL
XFILL_4__11259_ gnd vdd FILL
X_9792_ _9790_/Y _9764_/A _9792_/C gnd _9838_/D vdd OAI21X1
XFILL_5__13598_ gnd vdd FILL
XFILL_0__16405_ gnd vdd FILL
XFILL_2__12438_ gnd vdd FILL
XSFILL114520x25050 gnd vdd FILL
XFILL_0__13617_ gnd vdd FILL
XFILL_3__11989_ gnd vdd FILL
XFILL_1__15956_ gnd vdd FILL
XFILL_1__11079_ gnd vdd FILL
XFILL_3__14777_ gnd vdd FILL
XFILL_0__10829_ gnd vdd FILL
XFILL_0__8115_ gnd vdd FILL
XFILL_0__14597_ gnd vdd FILL
XFILL_5__15337_ gnd vdd FILL
X_8743_ _8714_/B _7079_/B gnd _8744_/C vdd NAND2X1
XSFILL43800x57050 gnd vdd FILL
XFILL_0__9095_ gnd vdd FILL
XFILL_3__9913_ gnd vdd FILL
XFILL_2__15157_ gnd vdd FILL
XFILL_3__13728_ gnd vdd FILL
XFILL_2__12369_ gnd vdd FILL
XFILL_0__16336_ gnd vdd FILL
XFILL_1__14907_ gnd vdd FILL
XFILL_0__13548_ gnd vdd FILL
XFILL_6__9622_ gnd vdd FILL
XFILL_1__15887_ gnd vdd FILL
XFILL_2__14108_ gnd vdd FILL
XFILL_5__15268_ gnd vdd FILL
X_8674_ _8602_/A _7382_/CLK _8674_/R vdd _8604_/Y gnd vdd DFFSR
XFILL_4__15998_ gnd vdd FILL
XFILL_1__14838_ gnd vdd FILL
XFILL_3__13659_ gnd vdd FILL
XFILL_2__15088_ gnd vdd FILL
XFILL_6_BUFX2_insert669 gnd vdd FILL
XFILL_0__16267_ gnd vdd FILL
XFILL_5__14219_ gnd vdd FILL
XFILL_0__13479_ gnd vdd FILL
X_7625_ _7623_/Y _7624_/A _7625_/C gnd _7665_/D vdd OAI21X1
XFILL_5__15199_ gnd vdd FILL
XFILL_2__14039_ gnd vdd FILL
XFILL_4__14949_ gnd vdd FILL
XFILL_0__15218_ gnd vdd FILL
XFILL_3__16378_ gnd vdd FILL
XFILL_3__6987_ gnd vdd FILL
XFILL_3__9775_ gnd vdd FILL
XFILL_1__14769_ gnd vdd FILL
XFILL_1__7810_ gnd vdd FILL
XFILL_0__16198_ gnd vdd FILL
XFILL_3__15329_ gnd vdd FILL
X_7556_ _7556_/A _7606_/A _7556_/C gnd _7642_/D vdd OAI21X1
XFILL_0__9997_ gnd vdd FILL
XSFILL8680x75050 gnd vdd FILL
XFILL_3__8726_ gnd vdd FILL
XSFILL23720x24050 gnd vdd FILL
XFILL_1_CLKBUF1_insert118 gnd vdd FILL
XFILL_0__15149_ gnd vdd FILL
XSFILL89160x19050 gnd vdd FILL
XFILL_1_CLKBUF1_insert129 gnd vdd FILL
XFILL_1__7741_ gnd vdd FILL
X_7487_ _7460_/A _7359_/B gnd _7488_/C vdd NAND2X1
XFILL_4__7450_ gnd vdd FILL
XFILL_3__8657_ gnd vdd FILL
X_9226_ _9226_/A _9277_/B _9226_/C gnd _9226_/Y vdd OAI21X1
XFILL_6__8366_ gnd vdd FILL
XFILL_1__7672_ gnd vdd FILL
XFILL_0__8879_ gnd vdd FILL
XFILL_3__7608_ gnd vdd FILL
XFILL_3__8588_ gnd vdd FILL
XFILL_4__7381_ gnd vdd FILL
XFILL_1__9411_ gnd vdd FILL
XFILL_6__7317_ gnd vdd FILL
XFILL_4__9120_ gnd vdd FILL
X_9157_ _9112_/A _6981_/B gnd _9158_/C vdd NAND2X1
XFILL_3_BUFX2_insert504 gnd vdd FILL
XFILL_3_BUFX2_insert515 gnd vdd FILL
XFILL_3_BUFX2_insert526 gnd vdd FILL
XSFILL54280x26050 gnd vdd FILL
XFILL_1__9342_ gnd vdd FILL
X_8108_ _8168_/Q gnd _8108_/Y vdd INVX1
XFILL_3_BUFX2_insert537 gnd vdd FILL
X_9088_ _9163_/A _9600_/B gnd _9088_/Y vdd NAND2X1
XFILL_3_BUFX2_insert548 gnd vdd FILL
XSFILL94680x31050 gnd vdd FILL
XFILL_3_BUFX2_insert559 gnd vdd FILL
XSFILL69320x48050 gnd vdd FILL
XSFILL103640x29050 gnd vdd FILL
XFILL_1__9273_ gnd vdd FILL
XFILL_4__8002_ gnd vdd FILL
X_8039_ _8039_/Q _7527_/CLK _9959_/R vdd _7979_/Y gnd vdd DFFSR
XFILL_3__9209_ gnd vdd FILL
XFILL_1__8224_ gnd vdd FILL
X_11990_ _11990_/A _11986_/Y _11990_/C gnd _13080_/A vdd NAND3X1
XSFILL104520x57050 gnd vdd FILL
X_10941_ _12773_/A _12818_/Q gnd _10941_/Y vdd NAND2X1
XSFILL74440x39050 gnd vdd FILL
XFILL_6_BUFX2_insert19 gnd vdd FILL
X_13660_ _8450_/A gnd _15255_/B vdd INVX1
XFILL_1__7106_ gnd vdd FILL
X_10872_ _12704_/A gnd _10873_/B vdd INVX1
XFILL_1__8086_ gnd vdd FILL
XSFILL74040x41050 gnd vdd FILL
XFILL_4__8904_ gnd vdd FILL
X_12611_ _12611_/A vdd _12611_/C gnd _12677_/D vdd OAI21X1
XFILL_4__9884_ gnd vdd FILL
X_13591_ _13591_/A _13590_/Y gnd _13595_/C vdd NOR2X1
XFILL_1__7037_ gnd vdd FILL
XFILL_4__8835_ gnd vdd FILL
X_15330_ _8328_/A gnd _15330_/Y vdd INVX1
XFILL_0_BUFX2_insert405 gnd vdd FILL
X_12542_ _12364_/A _12538_/CLK _13199_/R vdd _12542_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert416 gnd vdd FILL
XFILL_0_BUFX2_insert427 gnd vdd FILL
XFILL_2__7850_ gnd vdd FILL
XSFILL13720x56050 gnd vdd FILL
XFILL_0_BUFX2_insert438 gnd vdd FILL
XFILL_0_BUFX2_insert449 gnd vdd FILL
XFILL_4__8766_ gnd vdd FILL
X_15261_ _15261_/A _15175_/B _15087_/B _7643_/Q gnd _15261_/Y vdd AOI22X1
XSFILL28520x16050 gnd vdd FILL
X_12473_ vdd _12473_/B gnd _12473_/Y vdd NAND2X1
XFILL_4__7717_ gnd vdd FILL
X_14212_ _14208_/Y _14212_/B gnd _14212_/Y vdd NOR2X1
XFILL_1__8988_ gnd vdd FILL
XSFILL39160x67050 gnd vdd FILL
XFILL_5__7490_ gnd vdd FILL
X_11424_ _11421_/Y _11424_/B gnd _11457_/A vdd NOR2X1
X_15192_ _15192_/A _15192_/B gnd _15196_/A vdd NOR2X1
XFILL_4__8697_ gnd vdd FILL
XFILL_2__9520_ gnd vdd FILL
XFILL_1__7939_ gnd vdd FILL
X_14143_ _14143_/A _14143_/B _14142_/Y gnd _14144_/A vdd NAND3X1
XFILL_4__10630_ gnd vdd FILL
X_11355_ _11354_/Y _11346_/Y gnd _11356_/A vdd NOR2X1
XFILL_1__10450_ gnd vdd FILL
XFILL_5__9160_ gnd vdd FILL
XFILL_4__7579_ gnd vdd FILL
X_10306_ _10271_/B _9282_/B gnd _10307_/C vdd NAND2X1
XFILL_5__11920_ gnd vdd FILL
X_14074_ _14074_/A _14074_/B gnd _14074_/Y vdd NOR2X1
XFILL_2__8402_ gnd vdd FILL
XFILL_4_BUFX2_insert360 gnd vdd FILL
XFILL_3__11010_ gnd vdd FILL
XFILL_1__9609_ gnd vdd FILL
X_11286_ _11059_/Y _11646_/A _11658_/A gnd _11286_/Y vdd AOI21X1
XFILL_4__10561_ gnd vdd FILL
XSFILL59080x18050 gnd vdd FILL
XFILL_4_BUFX2_insert371 gnd vdd FILL
XFILL_2__9382_ gnd vdd FILL
XFILL_5__8111_ gnd vdd FILL
XCLKBUF1_insert117 CLKBUF1_insert193/A gnd _8551_/CLK vdd CLKBUF1
XFILL_2__11740_ gnd vdd FILL
XFILL_4_BUFX2_insert382 gnd vdd FILL
XFILL_1__10381_ gnd vdd FILL
XFILL_4_BUFX2_insert393 gnd vdd FILL
XCLKBUF1_insert128 CLKBUF1_insert193/A gnd _7400_/CLK vdd CLKBUF1
XFILL_5__9091_ gnd vdd FILL
X_13025_ _13023_/Y vdd _13025_/C gnd _13071_/D vdd OAI21X1
XSFILL99480x23050 gnd vdd FILL
XCLKBUF1_insert139 CLKBUF1_insert150/A gnd _9194_/CLK vdd CLKBUF1
XFILL_4__12300_ gnd vdd FILL
X_10237_ _10285_/A _9981_/B gnd _10238_/C vdd NAND2X1
XFILL_2__8333_ gnd vdd FILL
XFILL_4__13280_ gnd vdd FILL
XSFILL74120x21050 gnd vdd FILL
XFILL_5__11851_ gnd vdd FILL
XFILL_4__10492_ gnd vdd FILL
XFILL_1__12120_ gnd vdd FILL
XFILL_2__11671_ gnd vdd FILL
XFILL_4__9249_ gnd vdd FILL
XFILL_0__12850_ gnd vdd FILL
XFILL_4__12231_ gnd vdd FILL
XFILL_6__11052_ gnd vdd FILL
XFILL_5__10802_ gnd vdd FILL
XFILL_5__14570_ gnd vdd FILL
XFILL_2__13410_ gnd vdd FILL
X_10168_ _10220_/Q gnd _10170_/A vdd INVX1
XFILL_2__10622_ gnd vdd FILL
XFILL_2__8264_ gnd vdd FILL
XFILL_5__11782_ gnd vdd FILL
XFILL_3__12961_ gnd vdd FILL
XFILL_1__12051_ gnd vdd FILL
XFILL_2__14390_ gnd vdd FILL
XFILL_0__11801_ gnd vdd FILL
XFILL_0__12781_ gnd vdd FILL
XFILL_5__13521_ gnd vdd FILL
XFILL_4__12162_ gnd vdd FILL
XFILL_2__7215_ gnd vdd FILL
XFILL_3__14700_ gnd vdd FILL
XFILL_2__13341_ gnd vdd FILL
X_10099_ _10061_/A _7661_/CLK _8819_/R vdd _10099_/D gnd vdd DFFSR
XFILL_3__11912_ gnd vdd FILL
X_14976_ _14976_/A _14976_/B _14975_/Y gnd _14976_/Y vdd NAND3X1
XFILL_1__11002_ gnd vdd FILL
XFILL_3__15680_ gnd vdd FILL
XFILL_2__8195_ gnd vdd FILL
XFILL_3__12892_ gnd vdd FILL
XFILL_0__14520_ gnd vdd FILL
XFILL_2__10553_ gnd vdd FILL
XFILL_0__11732_ gnd vdd FILL
XFILL_5__16240_ gnd vdd FILL
XFILL_4__11113_ gnd vdd FILL
XFILL_5__9993_ gnd vdd FILL
XFILL_5__13452_ gnd vdd FILL
X_13927_ _8415_/Q _14414_/B _14926_/C _7007_/Q gnd _13928_/B vdd AOI22X1
XFILL_3__14631_ gnd vdd FILL
XFILL_5__10664_ gnd vdd FILL
XFILL_4__12093_ gnd vdd FILL
XFILL_1__15810_ gnd vdd FILL
XFILL_2__16060_ gnd vdd FILL
XFILL_3__11843_ gnd vdd FILL
XFILL_2__13272_ gnd vdd FILL
XSFILL64040x73050 gnd vdd FILL
XFILL_0__14451_ gnd vdd FILL
XFILL_5__12403_ gnd vdd FILL
XFILL_0__11663_ gnd vdd FILL
XFILL_4__15921_ gnd vdd FILL
XFILL_5__16171_ gnd vdd FILL
XFILL_2__15011_ gnd vdd FILL
XFILL_4__11044_ gnd vdd FILL
X_13858_ _9566_/Q gnd _13860_/D vdd INVX1
XFILL_5__13383_ gnd vdd FILL
XFILL_2__12223_ gnd vdd FILL
XFILL_2__7077_ gnd vdd FILL
XFILL_3__14562_ gnd vdd FILL
XFILL_0__13402_ gnd vdd FILL
XFILL_3__11774_ gnd vdd FILL
XFILL_1__15741_ gnd vdd FILL
XFILL_0__10614_ gnd vdd FILL
XFILL_1__12953_ gnd vdd FILL
XFILL_6__10905_ gnd vdd FILL
XFILL_0__14382_ gnd vdd FILL
XFILL_0__11594_ gnd vdd FILL
XFILL_5__15122_ gnd vdd FILL
X_12809_ _12809_/Q _12809_/CLK _12809_/R vdd _12751_/Y gnd vdd DFFSR
XFILL_3__16301_ gnd vdd FILL
XFILL_5__8875_ gnd vdd FILL
XFILL_5__12334_ gnd vdd FILL
XFILL_1_BUFX2_insert250 gnd vdd FILL
XFILL_4__15852_ gnd vdd FILL
XSFILL43880x31050 gnd vdd FILL
XFILL_1_BUFX2_insert261 gnd vdd FILL
XFILL_3__13513_ gnd vdd FILL
XFILL_3__14493_ gnd vdd FILL
X_13789_ _13789_/A _13789_/B _15338_/C gnd _12970_/B vdd AOI21X1
XFILL_0__16121_ gnd vdd FILL
XFILL_1__11904_ gnd vdd FILL
XFILL_2__12154_ gnd vdd FILL
XFILL_3__6910_ gnd vdd FILL
XFILL_1_BUFX2_insert272 gnd vdd FILL
XSFILL3480x80050 gnd vdd FILL
XFILL_0__13333_ gnd vdd FILL
XFILL_1__15672_ gnd vdd FILL
XFILL_1_BUFX2_insert283 gnd vdd FILL
XFILL_0__10545_ gnd vdd FILL
XFILL_3__7890_ gnd vdd FILL
XSFILL18520x48050 gnd vdd FILL
XFILL_1_BUFX2_insert294 gnd vdd FILL
XFILL_5__7826_ gnd vdd FILL
XFILL_1__12884_ gnd vdd FILL
XFILL_0__9920_ gnd vdd FILL
XFILL_4__14803_ gnd vdd FILL
XFILL_5__15053_ gnd vdd FILL
X_15528_ _15527_/Y _15528_/B gnd _15528_/Y vdd NOR2X1
XFILL_3__16232_ gnd vdd FILL
XFILL_5__12265_ gnd vdd FILL
XFILL_2__11105_ gnd vdd FILL
XFILL_1__14623_ gnd vdd FILL
XFILL_3__6841_ gnd vdd FILL
XFILL_3__10656_ gnd vdd FILL
XFILL_3__13444_ gnd vdd FILL
XFILL_4__15783_ gnd vdd FILL
XFILL_2__12085_ gnd vdd FILL
XFILL_4__12995_ gnd vdd FILL
XFILL_0__16052_ gnd vdd FILL
XFILL_1__11835_ gnd vdd FILL
XFILL_0__13264_ gnd vdd FILL
XFILL_5__14004_ gnd vdd FILL
XFILL_5__7757_ gnd vdd FILL
X_7410_ _7370_/A _8046_/CLK _9692_/R vdd _7372_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert950 gnd vdd FILL
XFILL_5__11216_ gnd vdd FILL
XFILL_4__14734_ gnd vdd FILL
XFILL_0_BUFX2_insert961 gnd vdd FILL
XFILL_0__9851_ gnd vdd FILL
X_15459_ _9440_/Q gnd _15459_/Y vdd INVX1
XFILL_2__15913_ gnd vdd FILL
XFILL_3__13375_ gnd vdd FILL
XFILL_4__11946_ gnd vdd FILL
XFILL_0__15003_ gnd vdd FILL
X_8390_ _8390_/A _8345_/B _8389_/Y gnd _8432_/D vdd OAI21X1
XFILL_5__12196_ gnd vdd FILL
XFILL_2__11036_ gnd vdd FILL
XFILL_3__16163_ gnd vdd FILL
XFILL_1__14554_ gnd vdd FILL
XFILL_0_BUFX2_insert972 gnd vdd FILL
XFILL_0__12215_ gnd vdd FILL
XFILL_0_BUFX2_insert983 gnd vdd FILL
XFILL_2__7979_ gnd vdd FILL
XFILL_1__11766_ gnd vdd FILL
XFILL_0_BUFX2_insert994 gnd vdd FILL
XSFILL59000x62050 gnd vdd FILL
XSFILL23640x39050 gnd vdd FILL
XFILL_0__9782_ gnd vdd FILL
XFILL_5__7688_ gnd vdd FILL
X_7341_ _7323_/A _9901_/B gnd _7342_/C vdd NAND2X1
XFILL_5__11147_ gnd vdd FILL
XFILL_3__15114_ gnd vdd FILL
XSFILL108920x22050 gnd vdd FILL
XFILL_3__12326_ gnd vdd FILL
XFILL_3__8511_ gnd vdd FILL
XFILL_2__9718_ gnd vdd FILL
XFILL_3__16094_ gnd vdd FILL
XFILL_4__14665_ gnd vdd FILL
XFILL_1__13505_ gnd vdd FILL
XFILL_0__6994_ gnd vdd FILL
XFILL_4__11877_ gnd vdd FILL
XFILL_2__15844_ gnd vdd FILL
XSFILL109400x29050 gnd vdd FILL
XFILL_3__9491_ gnd vdd FILL
XFILL_1__14485_ gnd vdd FILL
XFILL_5__9427_ gnd vdd FILL
XFILL_0__12146_ gnd vdd FILL
XFILL_1__11697_ gnd vdd FILL
XFILL_4__16404_ gnd vdd FILL
XFILL_0__8733_ gnd vdd FILL
XFILL_4__13616_ gnd vdd FILL
XFILL112200x68050 gnd vdd FILL
XFILL_1__16224_ gnd vdd FILL
XFILL_4__10828_ gnd vdd FILL
XFILL_3__15045_ gnd vdd FILL
XFILL_5__15955_ gnd vdd FILL
X_7272_ _7212_/A _7016_/CLK _8424_/R vdd _7272_/D gnd vdd DFFSR
XFILL_3__12257_ gnd vdd FILL
XFILL_5__11078_ gnd vdd FILL
XFILL_3__8442_ gnd vdd FILL
XFILL_4__14596_ gnd vdd FILL
XFILL_2__9649_ gnd vdd FILL
XFILL_1__13436_ gnd vdd FILL
XFILL_0__12077_ gnd vdd FILL
XFILL_1__10648_ gnd vdd FILL
XFILL_2__12987_ gnd vdd FILL
XFILL_2__15775_ gnd vdd FILL
XSFILL38840x20050 gnd vdd FILL
XFILL_5__9358_ gnd vdd FILL
X_9011_ _9011_/A _9011_/B gnd _9012_/C vdd NAND2X1
XFILL_4__16335_ gnd vdd FILL
XSFILL64120x53050 gnd vdd FILL
XFILL_5__10029_ gnd vdd FILL
XFILL_5__14906_ gnd vdd FILL
XFILL_3__11208_ gnd vdd FILL
XFILL_4__13547_ gnd vdd FILL
XFILL_5__15886_ gnd vdd FILL
XFILL_3__8373_ gnd vdd FILL
XFILL_0__15905_ gnd vdd FILL
XFILL_3__12188_ gnd vdd FILL
XFILL_2__14726_ gnd vdd FILL
XFILL_2__11938_ gnd vdd FILL
XFILL_4__10759_ gnd vdd FILL
XFILL_0__11028_ gnd vdd FILL
XFILL_1__16155_ gnd vdd FILL
XFILL_1__13367_ gnd vdd FILL
XFILL_0__7615_ gnd vdd FILL
XFILL_6__8082_ gnd vdd FILL
XSFILL79240x50 gnd vdd FILL
XFILL_1__10579_ gnd vdd FILL
XFILL_5__14837_ gnd vdd FILL
XFILL_5__9289_ gnd vdd FILL
XFILL_3__7324_ gnd vdd FILL
XFILL_3__11139_ gnd vdd FILL
XFILL_0__8595_ gnd vdd FILL
XFILL_1__15106_ gnd vdd FILL
XFILL_4__16266_ gnd vdd FILL
XFILL_4__13478_ gnd vdd FILL
XFILL_1__12318_ gnd vdd FILL
XFILL_2__11869_ gnd vdd FILL
XFILL_0__15836_ gnd vdd FILL
XFILL_6__7033_ gnd vdd FILL
XFILL_2__14657_ gnd vdd FILL
XFILL_1__16086_ gnd vdd FILL
XFILL_1__13298_ gnd vdd FILL
XSFILL43960x11050 gnd vdd FILL
XFILL_4__15217_ gnd vdd FILL
XFILL_0__7546_ gnd vdd FILL
XFILL_4__12429_ gnd vdd FILL
XSFILL3560x60050 gnd vdd FILL
XFILL_5__14768_ gnd vdd FILL
XFILL_2__13608_ gnd vdd FILL
XFILL_4__16197_ gnd vdd FILL
XFILL_1__15037_ gnd vdd FILL
XFILL_3__15947_ gnd vdd FILL
XFILL_2__14588_ gnd vdd FILL
XFILL_1__12249_ gnd vdd FILL
XFILL_0__15767_ gnd vdd FILL
XSFILL28760x72050 gnd vdd FILL
X_9913_ _9896_/B _9657_/B gnd _9914_/C vdd NAND2X1
XFILL_0__12979_ gnd vdd FILL
XFILL_5__13719_ gnd vdd FILL
XFILL_0__7477_ gnd vdd FILL
XFILL_4__15148_ gnd vdd FILL
XFILL_5__14699_ gnd vdd FILL
XFILL_2__16327_ gnd vdd FILL
XFILL_2__13539_ gnd vdd FILL
XSFILL44040x20050 gnd vdd FILL
XFILL_0__14718_ gnd vdd FILL
XFILL_3__7186_ gnd vdd FILL
XFILL_3__15878_ gnd vdd FILL
XFILL_0__9216_ gnd vdd FILL
XFILL_0__15698_ gnd vdd FILL
X_9844_ _9844_/Q _9834_/CLK _7793_/R vdd _9810_/Y gnd vdd DFFSR
XFILL_3__14829_ gnd vdd FILL
XFILL_4__15079_ gnd vdd FILL
XSFILL23720x19050 gnd vdd FILL
XFILL_2__16258_ gnd vdd FILL
XFILL_0__14649_ gnd vdd FILL
XFILL_0__9147_ gnd vdd FILL
XFILL_5__16369_ gnd vdd FILL
X_9775_ _9833_/Q gnd _9775_/Y vdd INVX1
XFILL_2__15209_ gnd vdd FILL
X_6987_ _6988_/B _7883_/B gnd _6988_/C vdd NAND2X1
XFILL_2__16189_ gnd vdd FILL
XFILL_4__6950_ gnd vdd FILL
XFILL_1__15939_ gnd vdd FILL
XFILL_0__9078_ gnd vdd FILL
X_8726_ _8724_/Y _8788_/A _8726_/C gnd _8726_/Y vdd OAI21X1
XFILL_6_BUFX2_insert444 gnd vdd FILL
XFILL_0__16319_ gnd vdd FILL
XFILL_4__6881_ gnd vdd FILL
XSFILL64200x33050 gnd vdd FILL
XSFILL89640x5050 gnd vdd FILL
XFILL_1__8911_ gnd vdd FILL
XSFILL49560x51050 gnd vdd FILL
X_8657_ _8657_/A _8529_/B gnd _8658_/C vdd NAND2X1
XFILL_1__9891_ gnd vdd FILL
XFILL_4__8620_ gnd vdd FILL
X_7608_ _7608_/A gnd _7610_/A vdd INVX1
XFILL_4_BUFX2_insert1001 gnd vdd FILL
XFILL_1__8842_ gnd vdd FILL
XFILL_4_BUFX2_insert1012 gnd vdd FILL
X_8588_ _8589_/B _7948_/B gnd _8588_/Y vdd NAND2X1
XFILL_4_BUFX2_insert1023 gnd vdd FILL
XFILL_4_BUFX2_insert1034 gnd vdd FILL
XFILL_3__9758_ gnd vdd FILL
XSFILL3640x40050 gnd vdd FILL
XFILL_6__9467_ gnd vdd FILL
XFILL_4_BUFX2_insert1045 gnd vdd FILL
X_7539_ _7539_/Q _8051_/CLK _7789_/R vdd _7503_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert1056 gnd vdd FILL
XFILL_1__8773_ gnd vdd FILL
XFILL_4__7502_ gnd vdd FILL
XFILL_3__8709_ gnd vdd FILL
XFILL_4_BUFX2_insert1067 gnd vdd FILL
XSFILL28840x52050 gnd vdd FILL
XFILL_4__8482_ gnd vdd FILL
XFILL_4_BUFX2_insert1089 gnd vdd FILL
XFILL_1__7724_ gnd vdd FILL
XFILL_4__7433_ gnd vdd FILL
X_11140_ _11139_/Y _11140_/B gnd _11519_/C vdd NOR2X1
X_9209_ _9303_/Q gnd _9211_/A vdd INVX1
XFILL_3_BUFX2_insert301 gnd vdd FILL
XFILL_4__7364_ gnd vdd FILL
XSFILL33960x43050 gnd vdd FILL
X_11071_ _12147_/Y gnd _11071_/Y vdd INVX2
XFILL_3_BUFX2_insert312 gnd vdd FILL
XFILL_3_BUFX2_insert323 gnd vdd FILL
XFILL_4__9103_ gnd vdd FILL
XFILL_1__7586_ gnd vdd FILL
XFILL_3_BUFX2_insert334 gnd vdd FILL
XFILL_3_BUFX2_insert345 gnd vdd FILL
XFILL_4__7295_ gnd vdd FILL
X_10022_ _14245_/A gnd _10024_/A vdd INVX1
XFILL_3_BUFX2_insert356 gnd vdd FILL
XFILL_2_BUFX2_insert1060 gnd vdd FILL
XFILL_2_BUFX2_insert1071 gnd vdd FILL
XFILL_3_BUFX2_insert367 gnd vdd FILL
XSFILL49400x8050 gnd vdd FILL
XSFILL34040x52050 gnd vdd FILL
XFILL_3_BUFX2_insert378 gnd vdd FILL
XFILL_4__9034_ gnd vdd FILL
XFILL_3_BUFX2_insert389 gnd vdd FILL
XFILL_2_BUFX2_insert1093 gnd vdd FILL
X_14830_ _14830_/A _14830_/B _13882_/B _14830_/D gnd _14830_/Y vdd OAI22X1
XFILL_1__9256_ gnd vdd FILL
XFILL_1__8207_ gnd vdd FILL
X_11973_ _11973_/A _11909_/A _11973_/C gnd _6866_/A vdd OAI21X1
XSFILL13880x10050 gnd vdd FILL
X_14761_ _14757_/Y _14761_/B gnd _14764_/C vdd NOR2X1
XSFILL3720x20050 gnd vdd FILL
X_10924_ _10924_/A _10938_/B gnd _10924_/Y vdd NOR2X1
X_13712_ _13711_/Y _13712_/B gnd _13713_/B vdd NOR2X1
XFILL_5__6990_ gnd vdd FILL
XFILL_1__8138_ gnd vdd FILL
X_14692_ _14692_/A _14692_/B _14402_/C gnd _13027_/B vdd AOI21X1
XSFILL28920x32050 gnd vdd FILL
XFILL_4__9936_ gnd vdd FILL
X_16431_ _16363_/A _6998_/CLK _7644_/R vdd _16431_/D gnd vdd DFFSR
XFILL_4_CLKBUF1_insert113 gnd vdd FILL
XFILL_5__10380_ gnd vdd FILL
X_13643_ _13643_/A _13803_/A _14567_/D _13643_/D gnd _13644_/A vdd OAI22X1
X_10855_ _14289_/D _7016_/CLK _9064_/R vdd _10855_/D gnd vdd DFFSR
XFILL_4_CLKBUF1_insert124 gnd vdd FILL
XFILL_1__8069_ gnd vdd FILL
XFILL_2__8951_ gnd vdd FILL
XFILL_4_CLKBUF1_insert135 gnd vdd FILL
XFILL_4_CLKBUF1_insert146 gnd vdd FILL
XFILL_4_CLKBUF1_insert157 gnd vdd FILL
XFILL_4__9867_ gnd vdd FILL
XFILL_5__8660_ gnd vdd FILL
XFILL_3__10510_ gnd vdd FILL
XFILL_4_CLKBUF1_insert168 gnd vdd FILL
X_16362_ _16362_/A gnd _16362_/C gnd _16430_/D vdd OAI21X1
X_13574_ _13574_/A _14934_/B _13574_/C _15139_/D gnd _13578_/A vdd OAI22X1
X_10786_ _10786_/A _10792_/B _10785_/Y gnd _10852_/D vdd OAI21X1
XFILL_4_CLKBUF1_insert179 gnd vdd FILL
XFILL_3__11490_ gnd vdd FILL
XFILL_5__7611_ gnd vdd FILL
XFILL_0_BUFX2_insert235 gnd vdd FILL
XFILL_2__8882_ gnd vdd FILL
XFILL_0_BUFX2_insert246 gnd vdd FILL
X_12525_ _12523_/Y vdd _12525_/C gnd _12525_/Y vdd OAI21X1
X_15313_ _13755_/D _15313_/B _15715_/C gnd _15318_/A vdd NOR3X1
XFILL_6__10621_ gnd vdd FILL
XFILL_5__8591_ gnd vdd FILL
XFILL_5__12050_ gnd vdd FILL
X_16293_ _16293_/A _7157_/Q _15380_/C _9973_/Q gnd _16295_/C vdd AOI22X1
XFILL_4__9798_ gnd vdd FILL
XFILL_4__11800_ gnd vdd FILL
XFILL_0_BUFX2_insert257 gnd vdd FILL
XFILL_3__10441_ gnd vdd FILL
XSFILL74120x16050 gnd vdd FILL
XFILL_4__12780_ gnd vdd FILL
XFILL_2__7833_ gnd vdd FILL
XFILL_1__11620_ gnd vdd FILL
XFILL_0_BUFX2_insert268 gnd vdd FILL
XFILL_0__10261_ gnd vdd FILL
XFILL_0_BUFX2_insert279 gnd vdd FILL
XSFILL84280x60050 gnd vdd FILL
XFILL_5__7542_ gnd vdd FILL
XFILL_4__8749_ gnd vdd FILL
XFILL_5__11001_ gnd vdd FILL
X_15244_ _15243_/Y _15031_/Y _15244_/C gnd _15680_/B vdd OAI21X1
X_12456_ _12456_/A vdd _12455_/Y gnd _12540_/D vdd OAI21X1
XFILL_2__12910_ gnd vdd FILL
XFILL_3__13160_ gnd vdd FILL
XFILL_4__11731_ gnd vdd FILL
XFILL_0__12000_ gnd vdd FILL
XFILL_3__10372_ gnd vdd FILL
XFILL_2__7764_ gnd vdd FILL
XFILL_1__11551_ gnd vdd FILL
XFILL_2__13890_ gnd vdd FILL
XFILL_5__7473_ gnd vdd FILL
X_11407_ _11406_/Y _11140_/B _11407_/C gnd _11562_/B vdd OAI21X1
XFILL_0__10192_ gnd vdd FILL
XSFILL99320x82050 gnd vdd FILL
X_15175_ _10457_/Q _15175_/B _15383_/A _7641_/Q gnd _15176_/B vdd AOI22X1
XFILL_3__12111_ gnd vdd FILL
X_12387_ _12385_/Y _12371_/A _12387_/C gnd _12387_/Y vdd OAI21X1
XFILL_2__9503_ gnd vdd FILL
XFILL_4__14450_ gnd vdd FILL
XFILL_2__12841_ gnd vdd FILL
XFILL_3__13091_ gnd vdd FILL
XFILL_4__11662_ gnd vdd FILL
XFILL_1__10502_ gnd vdd FILL
XFILL_2__7695_ gnd vdd FILL
XFILL_5__9212_ gnd vdd FILL
XFILL_1__14270_ gnd vdd FILL
X_14126_ _9888_/A gnd _14128_/D vdd INVX1
XFILL_1__11482_ gnd vdd FILL
XFILL_4__13401_ gnd vdd FILL
XFILL_2_BUFX2_insert17 gnd vdd FILL
XFILL_5__15740_ gnd vdd FILL
X_11338_ _11338_/A _10996_/Y _11231_/Y gnd _11341_/B vdd OAI21X1
XFILL_2_BUFX2_insert28 gnd vdd FILL
XFILL_5__12952_ gnd vdd FILL
XFILL_3__12042_ gnd vdd FILL
XSFILL38760x35050 gnd vdd FILL
XFILL_1__13221_ gnd vdd FILL
XFILL_2__15560_ gnd vdd FILL
XFILL_4__14381_ gnd vdd FILL
XFILL_4__11593_ gnd vdd FILL
XFILL_2_BUFX2_insert39 gnd vdd FILL
XFILL_2__12772_ gnd vdd FILL
XFILL112280x42050 gnd vdd FILL
XFILL_1__10433_ gnd vdd FILL
XFILL_5__9143_ gnd vdd FILL
XSFILL64040x68050 gnd vdd FILL
XFILL_0__13951_ gnd vdd FILL
XFILL_4__16120_ gnd vdd FILL
X_14057_ _9314_/Q gnd _14058_/A vdd INVX1
XFILL_5__11903_ gnd vdd FILL
XFILL_4__13332_ gnd vdd FILL
XFILL_5__15671_ gnd vdd FILL
X_11269_ _12141_/Y gnd _11270_/B vdd INVX2
XFILL_2__14511_ gnd vdd FILL
XFILL_4__10544_ gnd vdd FILL
XFILL_2__9365_ gnd vdd FILL
XFILL_2__11723_ gnd vdd FILL
XFILL_5__12883_ gnd vdd FILL
XFILL_1__13152_ gnd vdd FILL
XFILL_0__12902_ gnd vdd FILL
XFILL_2__15491_ gnd vdd FILL
X_13008_ _6889_/A gnd _13008_/Y vdd INVX1
XFILL_1__10364_ gnd vdd FILL
XFILL_0__13882_ gnd vdd FILL
XFILL_5__14622_ gnd vdd FILL
XFILL_0__8380_ gnd vdd FILL
XFILL_3__15801_ gnd vdd FILL
XFILL_4__16051_ gnd vdd FILL
XFILL_5__11834_ gnd vdd FILL
XFILL_4__13263_ gnd vdd FILL
XFILL_1__12103_ gnd vdd FILL
XFILL_2__8316_ gnd vdd FILL
XFILL_2__14442_ gnd vdd FILL
XSFILL43880x26050 gnd vdd FILL
XSFILL114840x56050 gnd vdd FILL
XFILL_0__15621_ gnd vdd FILL
XFILL_2__11654_ gnd vdd FILL
XFILL_2__9296_ gnd vdd FILL
XFILL_0__12833_ gnd vdd FILL
XFILL_3__13993_ gnd vdd FILL
XFILL_1__13083_ gnd vdd FILL
XFILL_3_BUFX2_insert890 gnd vdd FILL
XFILL_1__10295_ gnd vdd FILL
XFILL_0__7331_ gnd vdd FILL
XFILL_4__15002_ gnd vdd FILL
XFILL_5__14553_ gnd vdd FILL
XFILL_4__12214_ gnd vdd FILL
XFILL_3__7040_ gnd vdd FILL
XFILL_2__8247_ gnd vdd FILL
XFILL_3__15732_ gnd vdd FILL
XFILL_5__11765_ gnd vdd FILL
XFILL_1__12034_ gnd vdd FILL
XFILL_2__14373_ gnd vdd FILL
XFILL_0__15552_ gnd vdd FILL
XFILL_2__11585_ gnd vdd FILL
XFILL_0__12764_ gnd vdd FILL
XFILL_5__13504_ gnd vdd FILL
XFILL_6__15843_ gnd vdd FILL
X_6910_ _6910_/A _6955_/B _6909_/Y gnd _6910_/Y vdd OAI21X1
XFILL_2__13324_ gnd vdd FILL
XFILL_5__14484_ gnd vdd FILL
XFILL_2__16112_ gnd vdd FILL
X_14959_ _14211_/A _14959_/B _13587_/C _14959_/D gnd _14963_/A vdd OAI22X1
XFILL_4__12145_ gnd vdd FILL
XFILL_2__10536_ gnd vdd FILL
XFILL_3__15663_ gnd vdd FILL
XFILL_0__14503_ gnd vdd FILL
XSFILL84360x40050 gnd vdd FILL
XFILL_5__11696_ gnd vdd FILL
X_7890_ _7890_/A _7878_/B _7890_/C gnd _7924_/D vdd OAI21X1
XFILL_3__12875_ gnd vdd FILL
XFILL_0__11715_ gnd vdd FILL
XFILL_0__9001_ gnd vdd FILL
XFILL_5__16223_ gnd vdd FILL
XFILL_0__15483_ gnd vdd FILL
XFILL_0__12695_ gnd vdd FILL
XFILL_5__9976_ gnd vdd FILL
XFILL_5__13435_ gnd vdd FILL
XFILL_3__14614_ gnd vdd FILL
X_6841_ _6841_/A gnd memoryAddress[3] vdd BUFX2
XFILL_2__16043_ gnd vdd FILL
XFILL_4__12076_ gnd vdd FILL
XFILL_5__10647_ gnd vdd FILL
XFILL_0__7193_ gnd vdd FILL
XFILL_6__12986_ gnd vdd FILL
XFILL_2__13255_ gnd vdd FILL
XFILL_3__11826_ gnd vdd FILL
XSFILL99400x62050 gnd vdd FILL
XFILL_3__15594_ gnd vdd FILL
XFILL_0__14434_ gnd vdd FILL
XFILL_6__7720_ gnd vdd FILL
XFILL_1__13985_ gnd vdd FILL
XFILL_0__11646_ gnd vdd FILL
XFILL_3__8991_ gnd vdd FILL
XFILL_4__15904_ gnd vdd FILL
XFILL_6__11937_ gnd vdd FILL
XFILL_4__11027_ gnd vdd FILL
XFILL_5__16154_ gnd vdd FILL
XFILL_5__13366_ gnd vdd FILL
XFILL_2__12206_ gnd vdd FILL
X_9560_ _9468_/A _8152_/CLK _9944_/R vdd _9560_/D gnd vdd DFFSR
XFILL_3__14545_ gnd vdd FILL
XFILL_5__10578_ gnd vdd FILL
XFILL_1__15724_ gnd vdd FILL
XFILL_3__7942_ gnd vdd FILL
XFILL_3__11757_ gnd vdd FILL
XFILL_0__14365_ gnd vdd FILL
XFILL_2__10398_ gnd vdd FILL
XFILL_5__15105_ gnd vdd FILL
X_8511_ _8484_/A _8511_/B gnd _8511_/Y vdd NAND2X1
XFILL_5__8858_ gnd vdd FILL
XFILL_0__11577_ gnd vdd FILL
XFILL112360x22050 gnd vdd FILL
XFILL_5__12317_ gnd vdd FILL
XSFILL64120x48050 gnd vdd FILL
XFILL_4__15835_ gnd vdd FILL
XFILL_6__14656_ gnd vdd FILL
XFILL_5__16085_ gnd vdd FILL
XFILL_5__13297_ gnd vdd FILL
XFILL_2__12137_ gnd vdd FILL
XFILL_0__16104_ gnd vdd FILL
XFILL_3__10708_ gnd vdd FILL
X_9491_ _9489_/Y _9554_/B _9490_/Y gnd _9491_/Y vdd OAI21X1
XFILL_0__13316_ gnd vdd FILL
XFILL_5_BUFX2_insert407 gnd vdd FILL
XFILL_3__14476_ gnd vdd FILL
XFILL_1__15655_ gnd vdd FILL
XFILL_3__11688_ gnd vdd FILL
XFILL_5__7809_ gnd vdd FILL
XFILL_0__10528_ gnd vdd FILL
XFILL_1__12867_ gnd vdd FILL
XSFILL100200x5050 gnd vdd FILL
XFILL_3__7873_ gnd vdd FILL
XFILL_5__15036_ gnd vdd FILL
XFILL_0__9903_ gnd vdd FILL
XFILL_5_BUFX2_insert418 gnd vdd FILL
XFILL_0__14296_ gnd vdd FILL
XFILL_3__16215_ gnd vdd FILL
XFILL_5_BUFX2_insert429 gnd vdd FILL
XFILL_5__12248_ gnd vdd FILL
X_8442_ _8496_/A _9466_/B gnd _8443_/C vdd NAND2X1
XFILL_5__8789_ gnd vdd FILL
XFILL_3__10639_ gnd vdd FILL
XFILL_3__9612_ gnd vdd FILL
XFILL_1__14606_ gnd vdd FILL
XFILL_3__13427_ gnd vdd FILL
XFILL_4__15766_ gnd vdd FILL
XFILL_6__11799_ gnd vdd FILL
XFILL_0__16035_ gnd vdd FILL
XFILL_2__12068_ gnd vdd FILL
XFILL_4__12978_ gnd vdd FILL
XFILL_1__11818_ gnd vdd FILL
XFILL_0__13247_ gnd vdd FILL
XFILL_1__15586_ gnd vdd FILL
XFILL_0_BUFX2_insert780 gnd vdd FILL
XFILL_4__14717_ gnd vdd FILL
XFILL_0_BUFX2_insert791 gnd vdd FILL
X_8373_ _8427_/Q gnd _8375_/A vdd INVX1
XFILL_5__12179_ gnd vdd FILL
XSFILL3560x55050 gnd vdd FILL
XFILL_4__11929_ gnd vdd FILL
XFILL_2__11019_ gnd vdd FILL
XFILL_3__16146_ gnd vdd FILL
XFILL_3__13358_ gnd vdd FILL
XFILL_4__15697_ gnd vdd FILL
XFILL_1__14537_ gnd vdd FILL
XFILL_3__9543_ gnd vdd FILL
XFILL_1__11749_ gnd vdd FILL
XFILL_6__13469_ gnd vdd FILL
X_7324_ _7322_/Y _7359_/A _7323_/Y gnd _7324_/Y vdd OAI21X1
XSFILL109560x2050 gnd vdd FILL
XFILL_0__9765_ gnd vdd FILL
XSFILL28760x67050 gnd vdd FILL
XFILL_3__12309_ gnd vdd FILL
XFILL_0__6977_ gnd vdd FILL
XFILL_4__14648_ gnd vdd FILL
XFILL_3__13289_ gnd vdd FILL
XFILL_2__15827_ gnd vdd FILL
XFILL_3__16077_ gnd vdd FILL
XSFILL44040x15050 gnd vdd FILL
XFILL_3__9474_ gnd vdd FILL
XFILL_1__14468_ gnd vdd FILL
XFILL_0__12129_ gnd vdd FILL
XFILL_0__8716_ gnd vdd FILL
XFILL_1__16207_ gnd vdd FILL
XFILL_3__15028_ gnd vdd FILL
XFILL_5__15938_ gnd vdd FILL
X_7255_ _7161_/A _9205_/CLK _8433_/R vdd _7255_/D gnd vdd DFFSR
XFILL_4__14579_ gnd vdd FILL
XFILL_1__13419_ gnd vdd FILL
XFILL_2__15758_ gnd vdd FILL
XFILL_1__14399_ gnd vdd FILL
XFILL_1__7440_ gnd vdd FILL
XFILL_4__16318_ gnd vdd FILL
XFILL_0__8647_ gnd vdd FILL
XSFILL33880x58050 gnd vdd FILL
XFILL_2__14709_ gnd vdd FILL
XFILL_5__15869_ gnd vdd FILL
X_7186_ _7250_/B _7186_/B gnd _7186_/Y vdd NAND2X1
XFILL_1__16138_ gnd vdd FILL
XFILL_3__8356_ gnd vdd FILL
XFILL_2__15689_ gnd vdd FILL
XFILL_1__7371_ gnd vdd FILL
XFILL_0__8578_ gnd vdd FILL
XFILL_4__16249_ gnd vdd FILL
XFILL_3__7307_ gnd vdd FILL
XFILL_4__7080_ gnd vdd FILL
XSFILL33480x60050 gnd vdd FILL
XFILL_0__15819_ gnd vdd FILL
XFILL_1__16069_ gnd vdd FILL
XSFILL64200x28050 gnd vdd FILL
XFILL_1__9110_ gnd vdd FILL
XFILL_2_BUFX2_insert308 gnd vdd FILL
XFILL_1_BUFX2_insert3 gnd vdd FILL
XFILL_2_BUFX2_insert319 gnd vdd FILL
XFILL_3__7238_ gnd vdd FILL
XFILL_1__9041_ gnd vdd FILL
XFILL_3__7169_ gnd vdd FILL
XSFILL3640x35050 gnd vdd FILL
X_9827_ _9757_/A _7530_/CLK _7665_/R vdd _9827_/D gnd vdd DFFSR
XSFILL13240x68050 gnd vdd FILL
XSFILL28840x47050 gnd vdd FILL
XFILL_4__7982_ gnd vdd FILL
XSFILL94280x23050 gnd vdd FILL
X_9758_ _9813_/B _8606_/B gnd _9759_/C vdd NAND2X1
XFILL_6__8898_ gnd vdd FILL
XFILL_4__9721_ gnd vdd FILL
XFILL_4__6933_ gnd vdd FILL
X_10640_ _10638_/Y _10661_/B _10640_/C gnd _10718_/D vdd OAI21X1
XBUFX2_insert307 _11983_/Y gnd _12111_/C vdd BUFX2
XBUFX2_insert318 _15000_/Y gnd _16106_/A vdd BUFX2
XFILL_6__7849_ gnd vdd FILL
X_8709_ _8795_/Q gnd _8711_/A vdd INVX1
XBUFX2_insert329 _12405_/Y gnd _8243_/B vdd BUFX2
X_9689_ _9689_/Q _7129_/CLK _9062_/R vdd _9601_/Y gnd vdd DFFSR
XFILL_6_BUFX2_insert285 gnd vdd FILL
XFILL_4__9652_ gnd vdd FILL
XSFILL69320x61050 gnd vdd FILL
XFILL_4__6864_ gnd vdd FILL
XSFILL103640x42050 gnd vdd FILL
X_10571_ _10557_/B _8011_/B gnd _10572_/C vdd NAND2X1
XSFILL33960x38050 gnd vdd FILL
XFILL_5_CLKBUF1_insert208 gnd vdd FILL
XFILL_4__8603_ gnd vdd FILL
XFILL_1__9874_ gnd vdd FILL
XFILL_5_BUFX2_insert930 gnd vdd FILL
XFILL_5_CLKBUF1_insert219 gnd vdd FILL
X_12310_ _12307_/Y _12310_/B _12310_/C gnd _12310_/Y vdd NAND3X1
XFILL_5_BUFX2_insert941 gnd vdd FILL
XFILL_6__9519_ gnd vdd FILL
XFILL_5_BUFX2_insert952 gnd vdd FILL
X_13290_ _13289_/Y _13285_/B gnd _13290_/Y vdd AND2X2
XFILL_5_BUFX2_insert963 gnd vdd FILL
XFILL_1__8825_ gnd vdd FILL
XSFILL104520x70050 gnd vdd FILL
XFILL_5_BUFX2_insert974 gnd vdd FILL
XFILL_5_BUFX2_insert985 gnd vdd FILL
X_12241_ _6876_/A _12277_/B _12309_/C _12707_/A gnd _12242_/C vdd AOI22X1
XFILL_5_BUFX2_insert996 gnd vdd FILL
XSFILL74440x52050 gnd vdd FILL
XFILL_1__8756_ gnd vdd FILL
XSFILL89240x12050 gnd vdd FILL
XSFILL59080x3050 gnd vdd FILL
XFILL_4__8465_ gnd vdd FILL
X_12172_ _13194_/Q gnd _12174_/A vdd INVX1
XFILL_1__7707_ gnd vdd FILL
XFILL_2__7480_ gnd vdd FILL
XFILL_4__7416_ gnd vdd FILL
XSFILL3720x15050 gnd vdd FILL
X_11123_ _12174_/Y gnd _11125_/A vdd INVX1
XFILL_4__8396_ gnd vdd FILL
XSFILL28920x27050 gnd vdd FILL
XFILL_4__7347_ gnd vdd FILL
X_15931_ _15931_/A gnd _15931_/Y vdd INVX1
X_11054_ _11054_/A _11720_/A gnd _11055_/B vdd NOR2X1
XFILL_2__9150_ gnd vdd FILL
XFILL_1__7569_ gnd vdd FILL
X_10005_ _10066_/B _7317_/B gnd _10006_/C vdd NAND2X1
XSFILL29000x36050 gnd vdd FILL
XFILL_2__8101_ gnd vdd FILL
XFILL_4__10260_ gnd vdd FILL
X_15862_ _9778_/A _15390_/B _15861_/Y gnd _15862_/Y vdd AOI21X1
XFILL_2__9081_ gnd vdd FILL
XFILL_4__9017_ gnd vdd FILL
XFILL_3__10990_ gnd vdd FILL
XFILL_2_BUFX2_insert820 gnd vdd FILL
XFILL_2_BUFX2_insert831 gnd vdd FILL
X_14813_ _9586_/Q gnd _14813_/Y vdd INVX1
XFILL_2_BUFX2_insert842 gnd vdd FILL
XFILL_5__11550_ gnd vdd FILL
XFILL_4__10191_ gnd vdd FILL
XFILL_2_BUFX2_insert853 gnd vdd FILL
XFILL_1__9239_ gnd vdd FILL
X_15793_ _15790_/Y _15793_/B gnd _15793_/Y vdd NOR2X1
XFILL_2_BUFX2_insert864 gnd vdd FILL
XFILL_2__11370_ gnd vdd FILL
XFILL_2_BUFX2_insert875 gnd vdd FILL
XFILL_2_BUFX2_insert886 gnd vdd FILL
XFILL_5__10501_ gnd vdd FILL
XFILL_2_BUFX2_insert897 gnd vdd FILL
XSFILL84280x55050 gnd vdd FILL
X_14744_ _14743_/Y _14744_/B gnd _14745_/C vdd NOR2X1
X_11956_ _12184_/A gnd _11956_/Y vdd INVX1
XFILL_2__10321_ gnd vdd FILL
XFILL_5__11481_ gnd vdd FILL
XFILL_3__12660_ gnd vdd FILL
XFILL_0__11500_ gnd vdd FILL
XFILL_5__13220_ gnd vdd FILL
XFILL_5__9761_ gnd vdd FILL
XFILL_0__12480_ gnd vdd FILL
XFILL_5__6973_ gnd vdd FILL
X_10907_ _10911_/A _10903_/B gnd _10938_/A vdd NAND2X1
XFILL_5__10432_ gnd vdd FILL
XSFILL59080x31050 gnd vdd FILL
X_11887_ _11887_/A gnd _11889_/A vdd INVX1
XFILL_2__13040_ gnd vdd FILL
XFILL_3__11611_ gnd vdd FILL
X_14675_ _14675_/A _14506_/C _14718_/B _14675_/D gnd _14679_/B vdd OAI22X1
XFILL_4__13950_ gnd vdd FILL
XFILL_3__12591_ gnd vdd FILL
XFILL_2__10252_ gnd vdd FILL
XFILL_2__9983_ gnd vdd FILL
XFILL_4__9919_ gnd vdd FILL
XFILL_5__8712_ gnd vdd FILL
XFILL_1__13770_ gnd vdd FILL
XFILL_0__11431_ gnd vdd FILL
XFILL_1__10982_ gnd vdd FILL
X_16414_ _16448_/Q gnd _16414_/Y vdd INVX1
XFILL_6__11722_ gnd vdd FILL
X_13626_ _13876_/B gnd _14868_/D vdd INVX8
XFILL_5__13151_ gnd vdd FILL
X_10838_ _13410_/A _6998_/CLK _7644_/R vdd _10838_/D gnd vdd DFFSR
XFILL_4__12901_ gnd vdd FILL
XFILL_4_BUFX2_insert7 gnd vdd FILL
XFILL_6__15490_ gnd vdd FILL
XFILL_3__14330_ gnd vdd FILL
XFILL_3__11542_ gnd vdd FILL
XFILL_5__10363_ gnd vdd FILL
XFILL_1__12721_ gnd vdd FILL
XFILL_4__13881_ gnd vdd FILL
XFILL_0__14150_ gnd vdd FILL
XFILL112280x37050 gnd vdd FILL
XBUFX2_insert830 _15046_/Y gnd _15802_/D vdd BUFX2
XFILL_2__10183_ gnd vdd FILL
XFILL_5__12102_ gnd vdd FILL
XFILL_5__8643_ gnd vdd FILL
XFILL_0__11362_ gnd vdd FILL
XFILL_6__14441_ gnd vdd FILL
X_16345_ _16425_/Q gnd _16345_/Y vdd INVX1
XFILL_4__15620_ gnd vdd FILL
XBUFX2_insert841 _13324_/Y gnd _8657_/A vdd BUFX2
XBUFX2_insert852 _13269_/Y gnd _7055_/A vdd BUFX2
XFILL_4__12832_ gnd vdd FILL
XFILL_5__13082_ gnd vdd FILL
X_10769_ _13922_/A gnd _10769_/Y vdd INVX1
X_13557_ _15132_/D _14768_/D _14051_/C _13557_/D gnd _13557_/Y vdd OAI22X1
XFILL_5__10294_ gnd vdd FILL
XFILL_3__14261_ gnd vdd FILL
XFILL_0__13101_ gnd vdd FILL
XBUFX2_insert863 _13314_/Y gnd _8232_/B vdd BUFX2
XFILL_1__15440_ gnd vdd FILL
XFILL_3__11473_ gnd vdd FILL
XFILL_1__12652_ gnd vdd FILL
XFILL_2__8865_ gnd vdd FILL
XBUFX2_insert874 _13435_/Y gnd _13587_/A vdd BUFX2
XFILL_0__10313_ gnd vdd FILL
XFILL_2__14991_ gnd vdd FILL
XBUFX2_insert885 _13432_/Y gnd _13574_/C vdd BUFX2
XSFILL74200x5050 gnd vdd FILL
XFILL_0__11293_ gnd vdd FILL
XFILL_0__14081_ gnd vdd FILL
XFILL_0__6900_ gnd vdd FILL
XFILL_3__16000_ gnd vdd FILL
X_12508_ _12508_/A gnd _12508_/Y vdd INVX1
XFILL_5__12033_ gnd vdd FILL
XFILL_5__8574_ gnd vdd FILL
XFILL_3__13212_ gnd vdd FILL
XBUFX2_insert896 _13470_/Y gnd _14030_/A vdd BUFX2
XFILL_4__15551_ gnd vdd FILL
XFILL_3__10424_ gnd vdd FILL
XFILL_6__11584_ gnd vdd FILL
X_13488_ _7127_/Q _14344_/C _14037_/C _6999_/Q gnd _13488_/Y vdd AOI22X1
XFILL_0__7880_ gnd vdd FILL
X_16276_ _16276_/A _15527_/C _15644_/D _16276_/D gnd _16280_/A vdd OAI22X1
XFILL_4__12763_ gnd vdd FILL
XFILL_3__14192_ gnd vdd FILL
XFILL_2__7816_ gnd vdd FILL
XSFILL79240x44050 gnd vdd FILL
XFILL_1__11603_ gnd vdd FILL
XFILL_1__15371_ gnd vdd FILL
XFILL_0__10244_ gnd vdd FILL
XFILL_0__13032_ gnd vdd FILL
XFILL_2__13942_ gnd vdd FILL
XFILL_1__12583_ gnd vdd FILL
X_15227_ _13659_/Y _16213_/B _16208_/B _13657_/Y gnd _15228_/A vdd OAI22X1
X_12439_ _12343_/A gnd _12441_/A vdd INVX1
XFILL_4__14502_ gnd vdd FILL
XFILL_3__13143_ gnd vdd FILL
XFILL_4__11714_ gnd vdd FILL
XFILL_1__14322_ gnd vdd FILL
XFILL_4__15482_ gnd vdd FILL
XFILL_2__7747_ gnd vdd FILL
XFILL_1__11534_ gnd vdd FILL
XFILL_2__13873_ gnd vdd FILL
XFILL_0__10175_ gnd vdd FILL
XFILL_0__9550_ gnd vdd FILL
XSFILL114440x53050 gnd vdd FILL
XFILL_5__7456_ gnd vdd FILL
X_15158_ _9852_/A gnd _15158_/Y vdd INVX1
XFILL_4__14433_ gnd vdd FILL
XFILL_2__15612_ gnd vdd FILL
XFILL_5__13984_ gnd vdd FILL
XFILL_4__11645_ gnd vdd FILL
XFILL_1__14253_ gnd vdd FILL
XFILL_2__12824_ gnd vdd FILL
XFILL_3__10286_ gnd vdd FILL
XFILL_2__7678_ gnd vdd FILL
XFILL_1__11465_ gnd vdd FILL
XFILL_0__8501_ gnd vdd FILL
XFILL_0__14983_ gnd vdd FILL
X_14109_ _8733_/A _13853_/B _14109_/C gnd _14120_/A vdd AOI21X1
X_7040_ _7100_/A _7424_/B gnd _7040_/Y vdd NAND2X1
XFILL_5__15723_ gnd vdd FILL
XFILL_0__9481_ gnd vdd FILL
XFILL_3__12025_ gnd vdd FILL
X_15089_ _13528_/A _15175_/B gnd _15094_/B vdd NAND2X1
XFILL_2__9417_ gnd vdd FILL
XFILL_4__14364_ gnd vdd FILL
XFILL_3__8210_ gnd vdd FILL
XFILL_2__12755_ gnd vdd FILL
XFILL_2__15543_ gnd vdd FILL
XFILL_1__10416_ gnd vdd FILL
XFILL_4__11576_ gnd vdd FILL
XFILL_1__14184_ gnd vdd FILL
XSFILL99400x57050 gnd vdd FILL
XFILL_5__9126_ gnd vdd FILL
XSFILL59160x11050 gnd vdd FILL
XFILL_0__13934_ gnd vdd FILL
XFILL_4__16103_ gnd vdd FILL
XFILL_1__11396_ gnd vdd FILL
XFILL_4__13315_ gnd vdd FILL
XFILL_5__15654_ gnd vdd FILL
XFILL_3__8141_ gnd vdd FILL
XFILL_5__12866_ gnd vdd FILL
XFILL_2__11706_ gnd vdd FILL
XFILL_4__10527_ gnd vdd FILL
XFILL_2__9348_ gnd vdd FILL
XFILL_1__13135_ gnd vdd FILL
XFILL_4__14295_ gnd vdd FILL
XFILL_2__15474_ gnd vdd FILL
XFILL_0__13865_ gnd vdd FILL
XFILL_5__14605_ gnd vdd FILL
XFILL111880x10050 gnd vdd FILL
XFILL_4__16034_ gnd vdd FILL
XFILL_0__8363_ gnd vdd FILL
XFILL_5__11817_ gnd vdd FILL
XFILL_4__13246_ gnd vdd FILL
XFILL_5__15585_ gnd vdd FILL
XFILL_3__8072_ gnd vdd FILL
XFILL_2__11637_ gnd vdd FILL
X_8991_ _8991_/A _9044_/A _8990_/Y gnd _8991_/Y vdd OAI21X1
XFILL_0__15604_ gnd vdd FILL
XFILL_2__14425_ gnd vdd FILL
XFILL_2__9279_ gnd vdd FILL
XFILL_3__13976_ gnd vdd FILL
XFILL_5__8008_ gnd vdd FILL
XFILL_1__10278_ gnd vdd FILL
XFILL_0__7314_ gnd vdd FILL
XFILL_6__9870_ gnd vdd FILL
XFILL_0__13796_ gnd vdd FILL
XFILL_5__14536_ gnd vdd FILL
XFILL_3__15715_ gnd vdd FILL
X_7942_ _7931_/B _9094_/B gnd _7943_/C vdd NAND2X1
XFILL_5__11748_ gnd vdd FILL
XFILL_1__12017_ gnd vdd FILL
XFILL_2__14356_ gnd vdd FILL
XFILL_4__10389_ gnd vdd FILL
XFILL_0__15535_ gnd vdd FILL
XFILL_2__11568_ gnd vdd FILL
XFILL_0__12747_ gnd vdd FILL
XFILL_0__7245_ gnd vdd FILL
XSFILL79320x24050 gnd vdd FILL
XFILL_2__13307_ gnd vdd FILL
XFILL112200x81050 gnd vdd FILL
XFILL_5__14467_ gnd vdd FILL
XSFILL49080x63050 gnd vdd FILL
XFILL_4__12128_ gnd vdd FILL
XFILL_3__15646_ gnd vdd FILL
XFILL_2__10519_ gnd vdd FILL
X_7873_ _7919_/Q gnd _7873_/Y vdd INVX1
XFILL_5__11679_ gnd vdd FILL
XFILL_3__12858_ gnd vdd FILL
XFILL_2__14287_ gnd vdd FILL
XFILL_2__11499_ gnd vdd FILL
XFILL_0__15466_ gnd vdd FILL
X_9612_ _9613_/B _7564_/B gnd _9613_/C vdd NAND2X1
XFILL_5__16206_ gnd vdd FILL
XFILL_5__13418_ gnd vdd FILL
XFILL_0__7176_ gnd vdd FILL
XFILL_2__13238_ gnd vdd FILL
XFILL_2__16026_ gnd vdd FILL
XFILL_4__12059_ gnd vdd FILL
XFILL_5__14398_ gnd vdd FILL
XFILL_3__11809_ gnd vdd FILL
XSFILL114520x33050 gnd vdd FILL
XFILL_3__15577_ gnd vdd FILL
XFILL_0__14417_ gnd vdd FILL
XFILL_3__12789_ gnd vdd FILL
XFILL_3__8974_ gnd vdd FILL
XFILL_0__11629_ gnd vdd FILL
XFILL_1__13968_ gnd vdd FILL
XFILL_0__15397_ gnd vdd FILL
XFILL_5__16137_ gnd vdd FILL
XFILL_5__13349_ gnd vdd FILL
X_9543_ _9543_/A gnd _9543_/Y vdd INVX1
XFILL_3__14528_ gnd vdd FILL
XFILL_1__15707_ gnd vdd FILL
XFILL_2__13169_ gnd vdd FILL
XFILL_0__14348_ gnd vdd FILL
XFILL_1__13899_ gnd vdd FILL
XFILL_1__6940_ gnd vdd FILL
XFILL_5__16068_ gnd vdd FILL
X_9474_ _9562_/Q gnd _9476_/A vdd INVX1
XFILL_5_BUFX2_insert226 gnd vdd FILL
XFILL_4__15818_ gnd vdd FILL
XFILL_3__14459_ gnd vdd FILL
XFILL_1__15638_ gnd vdd FILL
XFILL_3__7856_ gnd vdd FILL
XFILL_5_BUFX2_insert237 gnd vdd FILL
XFILL_5_BUFX2_insert248 gnd vdd FILL
XFILL_5__15019_ gnd vdd FILL
XFILL_0__14279_ gnd vdd FILL
XFILL_6__7565_ gnd vdd FILL
XFILL_5_BUFX2_insert259 gnd vdd FILL
X_8425_ _8367_/A _9705_/CLK _7914_/R vdd _8369_/Y gnd vdd DFFSR
XFILL_1__6871_ gnd vdd FILL
XFILL_4__15749_ gnd vdd FILL
XFILL_0__16018_ gnd vdd FILL
XFILL_1__15569_ gnd vdd FILL
XFILL_4_BUFX2_insert904 gnd vdd FILL
XFILL_6__16309_ gnd vdd FILL
XFILL_1__8610_ gnd vdd FILL
X_8356_ _8356_/A _8356_/B gnd _8357_/C vdd NAND2X1
XFILL_1__9590_ gnd vdd FILL
XFILL_3__16129_ gnd vdd FILL
XFILL_4_BUFX2_insert915 gnd vdd FILL
XSFILL8680x83050 gnd vdd FILL
XFILL_3__9526_ gnd vdd FILL
XFILL_4_BUFX2_insert926 gnd vdd FILL
XFILL_4_BUFX2_insert937 gnd vdd FILL
XFILL_4_BUFX2_insert948 gnd vdd FILL
XFILL_6__9235_ gnd vdd FILL
X_7307_ _7389_/Q gnd _7307_/Y vdd INVX1
XFILL_4_BUFX2_insert959 gnd vdd FILL
XFILL_0__9748_ gnd vdd FILL
X_8287_ _8209_/A _9568_/CLK _8431_/R vdd _8287_/D gnd vdd DFFSR
XFILL_4__8250_ gnd vdd FILL
XFILL_1__8472_ gnd vdd FILL
X_7238_ _7238_/A _7181_/B _7237_/Y gnd _7280_/D vdd OAI21X1
XFILL_0__9679_ gnd vdd FILL
XFILL_4__7201_ gnd vdd FILL
XFILL_3__9388_ gnd vdd FILL
XFILL_1__7423_ gnd vdd FILL
XSFILL114600x13050 gnd vdd FILL
X_7169_ _7169_/A _7168_/A _7169_/C gnd _7257_/D vdd OAI21X1
XFILL_3__8339_ gnd vdd FILL
XSFILL54280x34050 gnd vdd FILL
XFILL_2_BUFX2_insert105 gnd vdd FILL
XSFILL28440x44050 gnd vdd FILL
XFILL_1__7354_ gnd vdd FILL
XFILL_4__7063_ gnd vdd FILL
XSFILL69320x56050 gnd vdd FILL
XFILL_1__9024_ gnd vdd FILL
X_11810_ _12226_/Y _11002_/B _11810_/C gnd _11810_/Y vdd OAI21X1
X_12790_ _12788_/Y _12789_/A _12790_/C gnd _12822_/D vdd OAI21X1
XFILL_1_BUFX2_insert805 gnd vdd FILL
XFILL_6__9999_ gnd vdd FILL
XFILL_1_BUFX2_insert816 gnd vdd FILL
XSFILL104520x65050 gnd vdd FILL
XFILL_1_BUFX2_insert827 gnd vdd FILL
XFILL_1_BUFX2_insert838 gnd vdd FILL
X_11741_ _11741_/A _11741_/B _11741_/C gnd _12467_/B vdd OAI21X1
XSFILL8760x63050 gnd vdd FILL
XSFILL23800x12050 gnd vdd FILL
XFILL_1_BUFX2_insert849 gnd vdd FILL
XFILL_4__7965_ gnd vdd FILL
X_14460_ _14458_/Y _14460_/B _14460_/C gnd _14473_/B vdd NAND3X1
XBUFX2_insert104 _10925_/Y gnd _11895_/B vdd BUFX2
X_11672_ _11656_/B _11649_/Y _11751_/C gnd _11672_/Y vdd OAI21X1
XFILL_2__6980_ gnd vdd FILL
XFILL_4__6916_ gnd vdd FILL
X_10623_ _10623_/A gnd _10623_/Y vdd INVX1
X_13411_ _9334_/A gnd _13411_/Y vdd INVX1
X_14391_ _7599_/A gnd _15815_/D vdd INVX1
XFILL_1__9926_ gnd vdd FILL
XFILL_4__9635_ gnd vdd FILL
X_13342_ _13240_/Y _13342_/B _13339_/Y gnd _13343_/B vdd NAND3X1
XFILL_4__6847_ gnd vdd FILL
X_16130_ _15390_/B _9841_/Q _9543_/A _15652_/A gnd _16130_/Y vdd AOI22X1
X_10554_ _10552_/Y _10557_/B _10554_/C gnd _10604_/D vdd OAI21X1
XSFILL109240x77050 gnd vdd FILL
XFILL_1__9857_ gnd vdd FILL
XFILL_2__8650_ gnd vdd FILL
XFILL_5_BUFX2_insert760 gnd vdd FILL
XFILL_5_BUFX2_insert771 gnd vdd FILL
XSFILL28520x24050 gnd vdd FILL
X_13273_ _13273_/A _13284_/B _13295_/C gnd _13273_/Y vdd OAI21X1
XFILL_5_BUFX2_insert782 gnd vdd FILL
X_16061_ _15087_/B _7663_/Q _7535_/Q _15383_/D gnd _16066_/B vdd AOI22X1
X_10485_ _14942_/A _9589_/CLK _7911_/R vdd _10485_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert793 gnd vdd FILL
XFILL_2__7601_ gnd vdd FILL
XFILL_1__9788_ gnd vdd FILL
XFILL_5__7310_ gnd vdd FILL
XFILL_4__8517_ gnd vdd FILL
XFILL_2__8581_ gnd vdd FILL
X_15012_ _12813_/Q _12812_/Q gnd _15012_/Y vdd NAND2X1
X_12224_ _12224_/A _12701_/A _12224_/C gnd _12226_/B vdd NAND3X1
XFILL_6__10320_ gnd vdd FILL
XFILL_4__9497_ gnd vdd FILL
XFILL_3__10140_ gnd vdd FILL
XFILL_1__8739_ gnd vdd FILL
XFILL_2__10870_ gnd vdd FILL
XFILL_4__8448_ gnd vdd FILL
XFILL_5__7241_ gnd vdd FILL
X_12155_ _12123_/B _12932_/Q gnd _12156_/C vdd NAND2X1
XFILL_4__11430_ gnd vdd FILL
XFILL_5__10981_ gnd vdd FILL
XFILL_2__7463_ gnd vdd FILL
XFILL_1__11250_ gnd vdd FILL
XFILL_5__7172_ gnd vdd FILL
X_11106_ _11105_/Y _11529_/A gnd _11107_/B vdd NOR2X1
XFILL_5__12720_ gnd vdd FILL
XFILL_4__8379_ gnd vdd FILL
XFILL_0__11980_ gnd vdd FILL
X_12086_ _12086_/A _12084_/Y _12085_/Y gnd _13152_/B vdd NAND3X1
XFILL_4__11361_ gnd vdd FILL
XSFILL59080x26050 gnd vdd FILL
XFILL_0__10931_ gnd vdd FILL
XSFILL99480x31050 gnd vdd FILL
XFILL_1__11181_ gnd vdd FILL
X_15914_ _10859_/Q gnd _15915_/A vdd INVX1
XFILL_4__13100_ gnd vdd FILL
X_11037_ _12242_/Y _11037_/B gnd _11037_/Y vdd NOR2X1
XFILL_5__12651_ gnd vdd FILL
XFILL_4__10312_ gnd vdd FILL
XFILL_3__13830_ gnd vdd FILL
XFILL_2__9133_ gnd vdd FILL
XFILL_4__11292_ gnd vdd FILL
XFILL_4__14080_ gnd vdd FILL
XFILL_2__12471_ gnd vdd FILL
XFILL_1__10132_ gnd vdd FILL
XFILL_0__13650_ gnd vdd FILL
XFILL_5__11602_ gnd vdd FILL
XFILL_2__14210_ gnd vdd FILL
XFILL_5__15370_ gnd vdd FILL
XFILL_4__10243_ gnd vdd FILL
X_15845_ _16089_/B _15845_/B _15899_/C _15845_/D gnd _15849_/B vdd OAI22X1
XFILL_4__13031_ gnd vdd FILL
XFILL_5__12582_ gnd vdd FILL
XFILL_2__11422_ gnd vdd FILL
XFILL_0__12601_ gnd vdd FILL
XFILL_2__15190_ gnd vdd FILL
XFILL_3__13761_ gnd vdd FILL
XFILL_2_BUFX2_insert650 gnd vdd FILL
XFILL_3__10973_ gnd vdd FILL
XFILL_1__10063_ gnd vdd FILL
XFILL_2_BUFX2_insert661 gnd vdd FILL
XFILL_1__14940_ gnd vdd FILL
XFILL_2_BUFX2_insert672 gnd vdd FILL
XFILL_5__14321_ gnd vdd FILL
XFILL_0__13581_ gnd vdd FILL
XFILL_2__8015_ gnd vdd FILL
XSFILL63960x72050 gnd vdd FILL
XFILL_3__15500_ gnd vdd FILL
XFILL_0__10793_ gnd vdd FILL
XFILL_5__11533_ gnd vdd FILL
XFILL_4__10174_ gnd vdd FILL
XFILL_3__12712_ gnd vdd FILL
XFILL_2__14141_ gnd vdd FILL
X_15776_ _15774_/Y _15776_/B gnd _15777_/C vdd NOR2X1
XFILL_2_BUFX2_insert683 gnd vdd FILL
XFILL_0__15320_ gnd vdd FILL
XFILL_2_BUFX2_insert694 gnd vdd FILL
X_12988_ vdd _12988_/B gnd _12989_/C vdd NAND2X1
XFILL_2__11353_ gnd vdd FILL
XFILL_1__14871_ gnd vdd FILL
XFILL_0__12532_ gnd vdd FILL
XFILL_5__9813_ gnd vdd FILL
XFILL_3__13692_ gnd vdd FILL
XFILL_0__7030_ gnd vdd FILL
XFILL_5__14252_ gnd vdd FILL
X_14727_ _7108_/A gnd _16113_/D vdd INVX1
XFILL_2__10304_ gnd vdd FILL
X_11939_ _11969_/A _12055_/B gnd _11940_/C vdd NAND2X1
XFILL_3__15431_ gnd vdd FILL
XFILL_5__11464_ gnd vdd FILL
XFILL_1__13822_ gnd vdd FILL
XFILL_3__12643_ gnd vdd FILL
XFILL_4__14982_ gnd vdd FILL
XFILL_2__14072_ gnd vdd FILL
XSFILL64040x81050 gnd vdd FILL
XFILL_5_BUFX2_insert10 gnd vdd FILL
XFILL_0__15251_ gnd vdd FILL
XFILL_2__11284_ gnd vdd FILL
XFILL_5__9744_ gnd vdd FILL
XFILL_5_BUFX2_insert21 gnd vdd FILL
XFILL_0__12463_ gnd vdd FILL
XSFILL114440x48050 gnd vdd FILL
XFILL_5__6956_ gnd vdd FILL
XFILL_5__10415_ gnd vdd FILL
XFILL_5__14183_ gnd vdd FILL
XFILL_2__13023_ gnd vdd FILL
X_14658_ _8385_/A _14414_/B _13883_/B _9455_/Q gnd _14667_/A vdd AOI22X1
XFILL_4__13933_ gnd vdd FILL
XFILL_5_BUFX2_insert32 gnd vdd FILL
XFILL_0__14202_ gnd vdd FILL
XFILL_3__15362_ gnd vdd FILL
XFILL_5_BUFX2_insert43 gnd vdd FILL
XFILL_5__11395_ gnd vdd FILL
XFILL_2__10235_ gnd vdd FILL
XFILL_3__12574_ gnd vdd FILL
XFILL_1__13753_ gnd vdd FILL
XFILL_0__11414_ gnd vdd FILL
XFILL_5_BUFX2_insert54 gnd vdd FILL
XFILL_1__10965_ gnd vdd FILL
XFILL_0__15182_ gnd vdd FILL
XFILL_5_BUFX2_insert65 gnd vdd FILL
XFILL_5_BUFX2_insert76 gnd vdd FILL
X_13609_ _8793_/Q _13853_/B _13609_/C gnd _13610_/B vdd AOI21X1
XFILL_5__13134_ gnd vdd FILL
XFILL_5__9675_ gnd vdd FILL
XFILL_0__12394_ gnd vdd FILL
XFILL_3__14313_ gnd vdd FILL
XFILL_5__6887_ gnd vdd FILL
XFILL_1__12704_ gnd vdd FILL
XFILL_4__13864_ gnd vdd FILL
X_14589_ _7533_/Q gnd _14589_/Y vdd INVX1
XFILL_5_BUFX2_insert87 gnd vdd FILL
XFILL_3__11525_ gnd vdd FILL
XFILL_0__8981_ gnd vdd FILL
XFILL_3__7710_ gnd vdd FILL
XFILL_2__8917_ gnd vdd FILL
XFILL_2__10166_ gnd vdd FILL
XFILL_5_BUFX2_insert98 gnd vdd FILL
XFILL_0__14133_ gnd vdd FILL
XSFILL98920x45050 gnd vdd FILL
XFILL_3__15293_ gnd vdd FILL
XFILL_1__13684_ gnd vdd FILL
XBUFX2_insert660 _11988_/Y gnd _12001_/C vdd BUFX2
XFILL_5__8626_ gnd vdd FILL
XFILL_0__11345_ gnd vdd FILL
XFILL_2__9897_ gnd vdd FILL
XBUFX2_insert671 _15064_/Y gnd _16228_/B vdd BUFX2
XFILL_1__10896_ gnd vdd FILL
XSFILL84360x6050 gnd vdd FILL
X_16328_ gnd gnd gnd _16328_/Y vdd NAND2X1
XFILL_4__15603_ gnd vdd FILL
XBUFX2_insert682 _15005_/Y gnd _15953_/A vdd BUFX2
XFILL_0__7932_ gnd vdd FILL
XFILL_5__10277_ gnd vdd FILL
XFILL_3__14244_ gnd vdd FILL
XBUFX2_insert693 _13362_/Y gnd _10500_/B vdd BUFX2
XFILL_3__11456_ gnd vdd FILL
XFILL_1__15423_ gnd vdd FILL
XFILL_1__12635_ gnd vdd FILL
XFILL_2__8848_ gnd vdd FILL
XFILL_4__13795_ gnd vdd FILL
XFILL_0__14064_ gnd vdd FILL
XFILL_2__14974_ gnd vdd FILL
XFILL_5__12016_ gnd vdd FILL
XFILL_0__11276_ gnd vdd FILL
X_8210_ _8244_/B _9362_/B gnd _8211_/C vdd NAND2X1
XFILL_4__15534_ gnd vdd FILL
X_16259_ _16259_/A _16258_/Y gnd _16283_/A vdd NOR2X1
XFILL_0__7863_ gnd vdd FILL
XFILL_3__10407_ gnd vdd FILL
XFILL_4__12746_ gnd vdd FILL
X_9190_ _9190_/Q _8562_/CLK _7270_/R vdd _9190_/D gnd vdd DFFSR
XFILL_3__14175_ gnd vdd FILL
XFILL_1__15354_ gnd vdd FILL
XFILL_0__13015_ gnd vdd FILL
XFILL_3__11387_ gnd vdd FILL
XFILL_2__13925_ gnd vdd FILL
XFILL_2__8779_ gnd vdd FILL
XFILL_5__7508_ gnd vdd FILL
XFILL_3__7572_ gnd vdd FILL
XFILL_6__13306_ gnd vdd FILL
XSFILL59000x70050 gnd vdd FILL
XFILL_0__9602_ gnd vdd FILL
X_8141_ _8141_/A gnd _8143_/A vdd INVX1
XFILL_5__8488_ gnd vdd FILL
XFILL_3__13126_ gnd vdd FILL
XFILL_1__14305_ gnd vdd FILL
XFILL_4__15465_ gnd vdd FILL
XSFILL109400x37050 gnd vdd FILL
XFILL_1__11517_ gnd vdd FILL
XFILL_2__13856_ gnd vdd FILL
XFILL_0__10158_ gnd vdd FILL
XFILL_1__15285_ gnd vdd FILL
XFILL_5__7439_ gnd vdd FILL
XFILL_1__12497_ gnd vdd FILL
XFILL_0__9533_ gnd vdd FILL
XFILL_6__10449_ gnd vdd FILL
XFILL_4__14416_ gnd vdd FILL
X_8072_ _8156_/Q gnd _8074_/A vdd INVX1
XSFILL49080x58050 gnd vdd FILL
XFILL_4__11628_ gnd vdd FILL
XFILL_5__13967_ gnd vdd FILL
XFILL112200x76050 gnd vdd FILL
XFILL_4__15396_ gnd vdd FILL
XFILL_1__14236_ gnd vdd FILL
XFILL_3__9242_ gnd vdd FILL
XFILL_3__10269_ gnd vdd FILL
XFILL_1__11448_ gnd vdd FILL
XFILL_2__13787_ gnd vdd FILL
XFILL_0__14966_ gnd vdd FILL
XFILL_2__10999_ gnd vdd FILL
XFILL_5__15706_ gnd vdd FILL
X_7023_ _7023_/Q _7647_/CLK _8047_/R vdd _7023_/D gnd vdd DFFSR
XFILL_0__9464_ gnd vdd FILL
XFILL_3__12008_ gnd vdd FILL
XFILL_4__14347_ gnd vdd FILL
XFILL_5__12918_ gnd vdd FILL
XFILL_2__15526_ gnd vdd FILL
XFILL_5__13898_ gnd vdd FILL
XFILL_4__11559_ gnd vdd FILL
XFILL_2__12738_ gnd vdd FILL
XFILL_1__14167_ gnd vdd FILL
XSFILL114520x28050 gnd vdd FILL
XFILL_5__9109_ gnd vdd FILL
XFILL_0__13917_ gnd vdd FILL
XFILL_3__9173_ gnd vdd FILL
XFILL_1__11379_ gnd vdd FILL
XFILL_0__14897_ gnd vdd FILL
XFILL_5__12849_ gnd vdd FILL
XFILL_5__15637_ gnd vdd FILL
XFILL_0__9395_ gnd vdd FILL
XFILL_3__8124_ gnd vdd FILL
XFILL_1__13118_ gnd vdd FILL
XFILL_4__14278_ gnd vdd FILL
XFILL_2__15457_ gnd vdd FILL
XFILL_0__13848_ gnd vdd FILL
XFILL_1__14098_ gnd vdd FILL
XFILL_4__16017_ gnd vdd FILL
XFILL_0__8346_ gnd vdd FILL
XFILL_4__13229_ gnd vdd FILL
X_8974_ _8974_/A gnd _8976_/A vdd INVX1
XFILL_3__8055_ gnd vdd FILL
XFILL_5__15568_ gnd vdd FILL
XFILL_2__14408_ gnd vdd FILL
XSFILL44120x9050 gnd vdd FILL
XFILL_3__13959_ gnd vdd FILL
XFILL_2__15388_ gnd vdd FILL
XFILL_0__13779_ gnd vdd FILL
XSFILL28760x80050 gnd vdd FILL
XFILL_5__14519_ gnd vdd FILL
XFILL_0__8277_ gnd vdd FILL
X_7925_ _7925_/Q _9589_/CLK _7285_/R vdd _7925_/D gnd vdd DFFSR
XFILL_1__7070_ gnd vdd FILL
XFILL_5__15499_ gnd vdd FILL
XFILL_0__15518_ gnd vdd FILL
XFILL_2__14339_ gnd vdd FILL
XFILL_0__7228_ gnd vdd FILL
XFILL_3__15629_ gnd vdd FILL
XFILL_6__6996_ gnd vdd FILL
X_7856_ _7878_/B _7856_/B gnd _7856_/Y vdd NAND2X1
XSFILL8680x78050 gnd vdd FILL
XFILL_0_CLKBUF1_insert205 gnd vdd FILL
XSFILL23720x27050 gnd vdd FILL
XFILL_0__15449_ gnd vdd FILL
XFILL_0_CLKBUF1_insert216 gnd vdd FILL
XFILL_0__7159_ gnd vdd FILL
XSFILL33880x71050 gnd vdd FILL
XFILL_2__16009_ gnd vdd FILL
X_7787_ _7787_/Q _7915_/CLK _7915_/R vdd _7735_/Y gnd vdd DFFSR
XFILL_3__8957_ gnd vdd FILL
XFILL_4__7750_ gnd vdd FILL
X_9526_ _9551_/B _9782_/B gnd _9527_/C vdd NAND2X1
XFILL_1_BUFX2_insert1009 gnd vdd FILL
XFILL_1__7972_ gnd vdd FILL
XFILL_4__7681_ gnd vdd FILL
XFILL_3__8888_ gnd vdd FILL
XFILL_1__6923_ gnd vdd FILL
X_9457_ _9457_/Q _7786_/CLK _8053_/R vdd _9457_/D gnd vdd DFFSR
XFILL_4__9420_ gnd vdd FILL
XFILL_3__7839_ gnd vdd FILL
X_8408_ _8408_/Q _8151_/CLK _9048_/R vdd _8408_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert701 gnd vdd FILL
XFILL_1__9642_ gnd vdd FILL
XFILL_1__6854_ gnd vdd FILL
XFILL_4_BUFX2_insert712 gnd vdd FILL
X_9388_ _9448_/Q gnd _9388_/Y vdd INVX1
XFILL_4_BUFX2_insert723 gnd vdd FILL
XFILL_4__9351_ gnd vdd FILL
XFILL_4_BUFX2_insert734 gnd vdd FILL
X_10270_ _10271_/B _8606_/B gnd _10271_/C vdd NAND2X1
XFILL_4_BUFX2_insert745 gnd vdd FILL
X_8339_ _8337_/Y _8372_/B _8339_/C gnd _8415_/D vdd OAI21X1
XFILL_3__9509_ gnd vdd FILL
XFILL_4_BUFX2_insert756 gnd vdd FILL
XFILL_3_CLKBUF1_insert1077 gnd vdd FILL
XSFILL28840x60050 gnd vdd FILL
XFILL_4_BUFX2_insert767 gnd vdd FILL
XFILL_4_BUFX2_insert778 gnd vdd FILL
XFILL_4__9282_ gnd vdd FILL
XFILL_1__8524_ gnd vdd FILL
XFILL_4_BUFX2_insert789 gnd vdd FILL
XFILL_4__8233_ gnd vdd FILL
XSFILL8760x58050 gnd vdd FILL
XFILL_1__8455_ gnd vdd FILL
X_13960_ _13959_/Y _13960_/B gnd _13960_/Y vdd NOR2X1
XFILL_1__8386_ gnd vdd FILL
XFILL_4__7115_ gnd vdd FILL
XFILL_4__8095_ gnd vdd FILL
X_12911_ vdd _12911_/B gnd _12912_/C vdd NAND2X1
XFILL_1__7337_ gnd vdd FILL
XSFILL79160x7050 gnd vdd FILL
X_13891_ _15437_/A gnd _13891_/Y vdd INVX1
XFILL_4__7046_ gnd vdd FILL
X_15630_ _15708_/A _14160_/A _15708_/C gnd _15650_/B vdd NOR3X1
XSFILL108760x65050 gnd vdd FILL
X_12842_ vdd _12842_/B gnd _12843_/C vdd NAND2X1
XFILL_1_BUFX2_insert602 gnd vdd FILL
XFILL_1_BUFX2_insert613 gnd vdd FILL
XFILL_1_BUFX2_insert624 gnd vdd FILL
X_15561_ _7906_/Q gnd _15562_/D vdd INVX1
XFILL_1__9007_ gnd vdd FILL
X_12773_ _12773_/A gnd _12773_/Y vdd INVX1
XFILL_1_BUFX2_insert635 gnd vdd FILL
XFILL_1_BUFX2_insert646 gnd vdd FILL
XFILL_1__7199_ gnd vdd FILL
XFILL_1_BUFX2_insert657 gnd vdd FILL
XFILL_1_BUFX2_insert668 gnd vdd FILL
X_14512_ _14510_/Y _14511_/Y _14512_/C gnd _14512_/Y vdd NAND3X1
XFILL_4__8997_ gnd vdd FILL
X_11724_ _11713_/A _11846_/C _11723_/Y gnd _11724_/Y vdd AOI21X1
XFILL_1_BUFX2_insert679 gnd vdd FILL
XSFILL28920x40050 gnd vdd FILL
X_15492_ _8544_/Q gnd _15493_/B vdd INVX1
XSFILL28920x9050 gnd vdd FILL
XFILL_4__7948_ gnd vdd FILL
XSFILL69000x33050 gnd vdd FILL
X_11655_ _11650_/Y _11676_/B _11651_/Y gnd _11656_/B vdd AOI21X1
X_14443_ _7274_/Q gnd _14444_/A vdd INVX1
XFILL_4__10930_ gnd vdd FILL
XFILL_2__10020_ gnd vdd FILL
XFILL_5__11180_ gnd vdd FILL
XFILL_2__9751_ gnd vdd FILL
XFILL_1__10750_ gnd vdd FILL
XFILL_2__6963_ gnd vdd FILL
X_10606_ _10606_/Q _7269_/CLK _9061_/R vdd _10606_/D gnd vdd DFFSR
XFILL_5__10131_ gnd vdd FILL
XFILL_3__11310_ gnd vdd FILL
XFILL_4__7879_ gnd vdd FILL
XFILL_1__9909_ gnd vdd FILL
X_14374_ _14374_/A _14373_/Y gnd _14374_/Y vdd NOR2X1
X_11586_ _11142_/A _11057_/Y _11139_/Y gnd _11587_/A vdd AOI21X1
XFILL_2__8702_ gnd vdd FILL
XFILL_3__12290_ gnd vdd FILL
XFILL_0__11130_ gnd vdd FILL
XFILL_4__9618_ gnd vdd FILL
XFILL_2__9682_ gnd vdd FILL
X_16113_ _14735_/Y _15527_/A _15920_/C _16113_/D gnd _16116_/B vdd OAI22X1
XFILL_1__10681_ gnd vdd FILL
XFILL_2__6894_ gnd vdd FILL
XFILL_4__12600_ gnd vdd FILL
XSFILL58840x76050 gnd vdd FILL
X_13325_ _13295_/C _13242_/B gnd _13326_/B vdd NAND2X1
XFILL_5__9391_ gnd vdd FILL
XSFILL99480x26050 gnd vdd FILL
X_10537_ _14295_/A gnd _10537_/Y vdd INVX1
XFILL_5__10062_ gnd vdd FILL
XFILL_3__11241_ gnd vdd FILL
XSFILL74120x24050 gnd vdd FILL
XFILL_2__8633_ gnd vdd FILL
XFILL_1__12420_ gnd vdd FILL
XFILL_4__13580_ gnd vdd FILL
XFILL_5_BUFX2_insert590 gnd vdd FILL
XFILL_4__10792_ gnd vdd FILL
XFILL_2__11971_ gnd vdd FILL
XFILL_0__11061_ gnd vdd FILL
XFILL_4__9549_ gnd vdd FILL
XFILL_6__14140_ gnd vdd FILL
XFILL_5__8342_ gnd vdd FILL
X_16044_ _16044_/A _16044_/B gnd _16044_/Y vdd NAND2X1
X_13256_ _13235_/C gnd _13337_/A vdd INVX2
XFILL_5__14870_ gnd vdd FILL
X_10468_ _14146_/B _7642_/CLK _8676_/R vdd _10402_/Y gnd vdd DFFSR
XFILL_4__12531_ gnd vdd FILL
XFILL_2__10922_ gnd vdd FILL
XFILL_0__10012_ gnd vdd FILL
XFILL_2__13710_ gnd vdd FILL
XFILL_3__11172_ gnd vdd FILL
XFILL_1__12351_ gnd vdd FILL
XFILL_2__14690_ gnd vdd FILL
X_12207_ _12207_/A _12201_/B _12207_/C gnd _12207_/Y vdd OAI21X1
XFILL_5__8273_ gnd vdd FILL
XFILL_5__13821_ gnd vdd FILL
XFILL_3__10123_ gnd vdd FILL
XFILL_4__15250_ gnd vdd FILL
X_13187_ _12151_/A _12537_/CLK _12536_/R vdd _13187_/D gnd vdd DFFSR
XFILL_4__12462_ gnd vdd FILL
XSFILL13800x39050 gnd vdd FILL
X_10399_ _10399_/A _10363_/B _10398_/Y gnd _10467_/D vdd OAI21X1
XFILL_1__11302_ gnd vdd FILL
XFILL_3__15980_ gnd vdd FILL
XFILL_2__13641_ gnd vdd FILL
XFILL_0__14820_ gnd vdd FILL
XFILL_1__15070_ gnd vdd FILL
XSFILL109480x11050 gnd vdd FILL
XFILL_6__13022_ gnd vdd FILL
XFILL_5__7224_ gnd vdd FILL
XFILL_1__12282_ gnd vdd FILL
XFILL_2__8495_ gnd vdd FILL
XFILL_4__14201_ gnd vdd FILL
X_12138_ _12138_/A _12137_/A _12138_/C gnd _12138_/Y vdd OAI21X1
XSFILL8760x2050 gnd vdd FILL
XFILL_5__13752_ gnd vdd FILL
XFILL_4__11413_ gnd vdd FILL
XFILL_5__10964_ gnd vdd FILL
XFILL_4__15181_ gnd vdd FILL
XFILL_1__14021_ gnd vdd FILL
XFILL_3__10054_ gnd vdd FILL
XFILL_3__14931_ gnd vdd FILL
XFILL_4__12393_ gnd vdd FILL
XFILL112280x50050 gnd vdd FILL
XFILL_2__16360_ gnd vdd FILL
XFILL_2__13572_ gnd vdd FILL
XFILL_2__7446_ gnd vdd FILL
XFILL_1__11233_ gnd vdd FILL
XSFILL64040x76050 gnd vdd FILL
XFILL_2_CLKBUF1_insert160 gnd vdd FILL
XFILL_2__10784_ gnd vdd FILL
XFILL_0__14751_ gnd vdd FILL
XFILL_5__12703_ gnd vdd FILL
XFILL_0__11963_ gnd vdd FILL
XFILL_2_CLKBUF1_insert171 gnd vdd FILL
XFILL_6__10165_ gnd vdd FILL
XFILL_4__14132_ gnd vdd FILL
X_12069_ _12069_/A _12093_/B _12061_/C gnd gnd _12069_/Y vdd AOI22X1
XFILL_2_CLKBUF1_insert182 gnd vdd FILL
XFILL_2_CLKBUF1_insert193 gnd vdd FILL
XFILL_2__15311_ gnd vdd FILL
XFILL_5__13683_ gnd vdd FILL
XFILL_4__11344_ gnd vdd FILL
XFILL_3__14862_ gnd vdd FILL
XFILL_2__12523_ gnd vdd FILL
XFILL_5__10895_ gnd vdd FILL
XFILL_0__13702_ gnd vdd FILL
XFILL_2__7377_ gnd vdd FILL
XFILL_0__10914_ gnd vdd FILL
XFILL_0__8200_ gnd vdd FILL
XFILL_2__16291_ gnd vdd FILL
XFILL_1__11164_ gnd vdd FILL
XFILL_5__7086_ gnd vdd FILL
XFILL_0__14682_ gnd vdd FILL
XFILL_5__12634_ gnd vdd FILL
XFILL_0__11894_ gnd vdd FILL
XFILL_5__15422_ gnd vdd FILL
XFILL_3__13813_ gnd vdd FILL
XFILL_2__9116_ gnd vdd FILL
XFILL_4__14063_ gnd vdd FILL
XFILL_6__14973_ gnd vdd FILL
XFILL_1__10115_ gnd vdd FILL
XFILL_2__15242_ gnd vdd FILL
XFILL_2__12454_ gnd vdd FILL
XSFILL43880x34050 gnd vdd FILL
XFILL_4__11275_ gnd vdd FILL
XFILL_0__13633_ gnd vdd FILL
XFILL_3__14793_ gnd vdd FILL
XFILL_1__15972_ gnd vdd FILL
XFILL_1__11095_ gnd vdd FILL
XFILL_0__8131_ gnd vdd FILL
XFILL_4__13014_ gnd vdd FILL
XFILL_5__15353_ gnd vdd FILL
XBUFX2_insert4 _12381_/Y gnd _8987_/B vdd BUFX2
X_15828_ _7401_/Q _15631_/B _15945_/C gnd _15829_/C vdd NAND3X1
XFILL_2__11405_ gnd vdd FILL
XFILL_3__13744_ gnd vdd FILL
XFILL_2__15173_ gnd vdd FILL
XFILL_2_BUFX2_insert480 gnd vdd FILL
XSFILL18680x10050 gnd vdd FILL
XFILL_3__10956_ gnd vdd FILL
XFILL_1__10046_ gnd vdd FILL
XFILL_2__12385_ gnd vdd FILL
XFILL_0__16352_ gnd vdd FILL
XFILL_2_BUFX2_insert491 gnd vdd FILL
XFILL_1__14923_ gnd vdd FILL
XFILL_5__14304_ gnd vdd FILL
XFILL_0__13564_ gnd vdd FILL
XFILL_5__11516_ gnd vdd FILL
XFILL_0__10776_ gnd vdd FILL
XFILL_0__8062_ gnd vdd FILL
X_7710_ _7753_/B _7326_/B gnd _7711_/C vdd NAND2X1
XSFILL68280x81050 gnd vdd FILL
XFILL_6_BUFX2_insert807 gnd vdd FILL
X_15759_ _7337_/A _15789_/B _15794_/B gnd _15760_/C vdd NAND3X1
XFILL_5__15284_ gnd vdd FILL
XSFILL18920x72050 gnd vdd FILL
X_8690_ _8690_/Q _8537_/CLK _8166_/R vdd _8652_/Y gnd vdd DFFSR
XFILL_0__15303_ gnd vdd FILL
XFILL_2__14124_ gnd vdd FILL
XFILL_5__12496_ gnd vdd FILL
XFILL_4__10157_ gnd vdd FILL
XFILL_2__11336_ gnd vdd FILL
XFILL_3__13675_ gnd vdd FILL
XFILL_3__9860_ gnd vdd FILL
XFILL_0__12515_ gnd vdd FILL
XFILL_1__14854_ gnd vdd FILL
XFILL_3__10887_ gnd vdd FILL
XFILL_0__16283_ gnd vdd FILL
XFILL_5__14235_ gnd vdd FILL
XFILL_0__13495_ gnd vdd FILL
X_7641_ _7641_/Q _8537_/CLK _9054_/R vdd _7553_/Y gnd vdd DFFSR
XFILL_3__15414_ gnd vdd FILL
XSFILL59000x65050 gnd vdd FILL
XFILL_5__11447_ gnd vdd FILL
XFILL_5__7988_ gnd vdd FILL
XFILL_3__12626_ gnd vdd FILL
XFILL_2__14055_ gnd vdd FILL
XFILL_4__14965_ gnd vdd FILL
XSFILL108920x25050 gnd vdd FILL
XSFILL99400x70050 gnd vdd FILL
XFILL_1__13805_ gnd vdd FILL
XFILL_0__15234_ gnd vdd FILL
XFILL_2__11267_ gnd vdd FILL
XFILL_3__16394_ gnd vdd FILL
XFILL_3__9791_ gnd vdd FILL
XFILL_5__9727_ gnd vdd FILL
XFILL_0__12446_ gnd vdd FILL
XFILL_1__14785_ gnd vdd FILL
XFILL_1__11997_ gnd vdd FILL
XFILL_5__6939_ gnd vdd FILL
XFILL_5__14166_ gnd vdd FILL
XFILL_2__13006_ gnd vdd FILL
XFILL_4__13916_ gnd vdd FILL
XFILL_3__15345_ gnd vdd FILL
X_7572_ _7572_/A gnd _7572_/Y vdd INVX1
XFILL_5__11378_ gnd vdd FILL
XFILL_3__8742_ gnd vdd FILL
XSFILL23240x44050 gnd vdd FILL
XFILL_4__14896_ gnd vdd FILL
XFILL_1__10948_ gnd vdd FILL
XFILL_0__15165_ gnd vdd FILL
XFILL_1__13736_ gnd vdd FILL
XFILL_2__11198_ gnd vdd FILL
XFILL_0__12377_ gnd vdd FILL
XSFILL109800x53050 gnd vdd FILL
XFILL_5__13117_ gnd vdd FILL
XFILL_5__9658_ gnd vdd FILL
X_9311_ _9311_/Q _7007_/CLK _9332_/R vdd _9311_/D gnd vdd DFFSR
XFILL112360x30050 gnd vdd FILL
XSFILL64920x75050 gnd vdd FILL
XFILL_4__13847_ gnd vdd FILL
XFILL_0__8964_ gnd vdd FILL
XSFILL64120x56050 gnd vdd FILL
XFILL_3__11508_ gnd vdd FILL
XFILL_5__14097_ gnd vdd FILL
XFILL_2__10149_ gnd vdd FILL
XFILL_0__14116_ gnd vdd FILL
XFILL_3__15276_ gnd vdd FILL
XFILL_1__13667_ gnd vdd FILL
XFILL_5__8609_ gnd vdd FILL
XFILL_3__12488_ gnd vdd FILL
XBUFX2_insert490 _13471_/Y gnd _14643_/C vdd BUFX2
XFILL_0__11328_ gnd vdd FILL
XFILL_1__10879_ gnd vdd FILL
XFILL_0__15096_ gnd vdd FILL
X_9242_ _9314_/Q gnd _9244_/A vdd INVX1
XFILL_2_CLKBUF1_insert1083 gnd vdd FILL
XFILL_3__14227_ gnd vdd FILL
XFILL_0__8895_ gnd vdd FILL
XFILL_1__12618_ gnd vdd FILL
XFILL_1__15406_ gnd vdd FILL
XFILL_4__13778_ gnd vdd FILL
XFILL_3__11439_ gnd vdd FILL
XFILL_3__7624_ gnd vdd FILL
XFILL_0__14047_ gnd vdd FILL
XFILL_2__14957_ gnd vdd FILL
XFILL_1__16386_ gnd vdd FILL
XFILL_1__13598_ gnd vdd FILL
XFILL_0__11259_ gnd vdd FILL
XFILL_4__15517_ gnd vdd FILL
XFILL_4__12729_ gnd vdd FILL
XFILL_0__7846_ gnd vdd FILL
XSFILL3560x63050 gnd vdd FILL
X_9173_ _9173_/A _9086_/B _9172_/Y gnd _9205_/D vdd OAI21X1
XFILL_3__14158_ gnd vdd FILL
XFILL_2__13908_ gnd vdd FILL
XFILL_3__7555_ gnd vdd FILL
XFILL_1__15337_ gnd vdd FILL
XFILL_2__14888_ gnd vdd FILL
X_8124_ _8079_/A _7868_/B gnd _8125_/C vdd NAND2X1
XSFILL28760x75050 gnd vdd FILL
XFILL_3__13109_ gnd vdd FILL
XFILL_4__15448_ gnd vdd FILL
XFILL_3_BUFX2_insert708 gnd vdd FILL
XFILL_2__13839_ gnd vdd FILL
XFILL_3_BUFX2_insert719 gnd vdd FILL
XFILL_5__14999_ gnd vdd FILL
XFILL_3__14089_ gnd vdd FILL
XFILL_1__15268_ gnd vdd FILL
XSFILL44040x23050 gnd vdd FILL
XFILL_3__7486_ gnd vdd FILL
XFILL_0__9516_ gnd vdd FILL
XFILL_0__15998_ gnd vdd FILL
X_8055_ _8567_/A _8100_/A gnd _8055_/Y vdd NAND2X1
XFILL_4__15379_ gnd vdd FILL
XFILL_1__14219_ gnd vdd FILL
XFILL_3__9225_ gnd vdd FILL
XFILL_1__15199_ gnd vdd FILL
XFILL_1_BUFX2_insert30 gnd vdd FILL
X_7006_ _6926_/A _7902_/CLK _7150_/R vdd _7006_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert41 gnd vdd FILL
XFILL_0__14949_ gnd vdd FILL
XFILL_1__8240_ gnd vdd FILL
XFILL_1_BUFX2_insert52 gnd vdd FILL
XFILL_2__15509_ gnd vdd FILL
XFILL_1_BUFX2_insert63 gnd vdd FILL
XFILL_1_BUFX2_insert74 gnd vdd FILL
XFILL_3__9156_ gnd vdd FILL
XFILL111800x44050 gnd vdd FILL
XFILL_1_BUFX2_insert85 gnd vdd FILL
XFILL_1_BUFX2_insert96 gnd vdd FILL
XFILL_0__9378_ gnd vdd FILL
XFILL_3__8107_ gnd vdd FILL
XFILL_3__9087_ gnd vdd FILL
XFILL112440x10050 gnd vdd FILL
XSFILL64200x36050 gnd vdd FILL
XSFILL89640x8050 gnd vdd FILL
XFILL_1__7122_ gnd vdd FILL
XFILL_0__8329_ gnd vdd FILL
XSFILL38920x4050 gnd vdd FILL
X_8957_ _9005_/A _7293_/B gnd _8958_/C vdd NAND2X1
XSFILL39000x12050 gnd vdd FILL
XFILL_1__7053_ gnd vdd FILL
X_7908_ _7840_/A _7642_/CLK _8676_/R vdd _7842_/Y gnd vdd DFFSR
X_8888_ _8888_/A gnd _8888_/Y vdd INVX1
XFILL_4__8851_ gnd vdd FILL
XSFILL3640x43050 gnd vdd FILL
XFILL_6__9767_ gnd vdd FILL
X_7839_ _7837_/Y _7814_/A _7839_/C gnd _7907_/D vdd OAI21X1
XFILL_4__7802_ gnd vdd FILL
XFILL_0_BUFX2_insert609 gnd vdd FILL
XFILL_6__8718_ gnd vdd FILL
XFILL_4__8782_ gnd vdd FILL
XSFILL28840x55050 gnd vdd FILL
XFILL_3__9989_ gnd vdd FILL
XFILL_4__7733_ gnd vdd FILL
X_11440_ _11440_/A gnd _11440_/Y vdd INVX1
X_9509_ _9509_/A _9548_/B _9508_/Y gnd _9573_/D vdd OAI21X1
XFILL_1__7955_ gnd vdd FILL
XSFILL33960x46050 gnd vdd FILL
X_11371_ _12230_/Y _10999_/Y _11370_/Y gnd _11379_/B vdd OAI21X1
XFILL_1__6906_ gnd vdd FILL
XFILL_4__9403_ gnd vdd FILL
XFILL_1__7886_ gnd vdd FILL
X_13110_ _13108_/B _13110_/B gnd _13110_/Y vdd NAND2X1
X_10322_ _10320_/Y _10271_/B _10322_/C gnd _10356_/D vdd OAI21X1
XFILL_4__7595_ gnd vdd FILL
XFILL_4_BUFX2_insert520 gnd vdd FILL
X_14090_ _8221_/A gnd _14091_/A vdd INVX1
XFILL_1__9625_ gnd vdd FILL
XFILL_4_BUFX2_insert531 gnd vdd FILL
XFILL_1__6837_ gnd vdd FILL
XFILL_4_BUFX2_insert542 gnd vdd FILL
XFILL_4__9334_ gnd vdd FILL
XFILL_4_BUFX2_insert553 gnd vdd FILL
X_13041_ _6900_/A gnd _13041_/Y vdd INVX1
X_10253_ _10253_/A _10294_/A _10252_/Y gnd _10253_/Y vdd OAI21X1
XFILL_4_BUFX2_insert564 gnd vdd FILL
XFILL_4_BUFX2_insert575 gnd vdd FILL
XFILL_1__9556_ gnd vdd FILL
XFILL_4_BUFX2_insert586 gnd vdd FILL
XFILL_4_BUFX2_insert597 gnd vdd FILL
XFILL_4__9265_ gnd vdd FILL
XFILL_1__8507_ gnd vdd FILL
XFILL_2__7300_ gnd vdd FILL
X_10184_ _10160_/A _8136_/B gnd _10185_/C vdd NAND2X1
XFILL_1__9487_ gnd vdd FILL
XFILL_4__8216_ gnd vdd FILL
XSFILL3720x23050 gnd vdd FILL
XSFILL38680x58050 gnd vdd FILL
XSFILL93720x45050 gnd vdd FILL
XSFILL64600x5050 gnd vdd FILL
XFILL_2__7231_ gnd vdd FILL
XFILL_1__8438_ gnd vdd FILL
X_14992_ _15064_/A _14981_/Y _15044_/C gnd _14992_/Y vdd NAND3X1
XSFILL28920x35050 gnd vdd FILL
XFILL_4__8147_ gnd vdd FILL
XSFILL94360x11050 gnd vdd FILL
XFILL_3_CLKBUF1_insert200 gnd vdd FILL
X_13943_ _10592_/Q gnd _15479_/D vdd INVX1
XFILL_3_CLKBUF1_insert211 gnd vdd FILL
XFILL_5__10680_ gnd vdd FILL
XFILL_2__7162_ gnd vdd FILL
XFILL_3_CLKBUF1_insert222 gnd vdd FILL
XFILL_1__8369_ gnd vdd FILL
XFILL_5__8960_ gnd vdd FILL
XFILL_4__8078_ gnd vdd FILL
XSFILL79160x72050 gnd vdd FILL
X_13874_ _9870_/A gnd _13874_/Y vdd INVX1
XFILL_3__10810_ gnd vdd FILL
XFILL_4__11060_ gnd vdd FILL
XFILL_2__7093_ gnd vdd FILL
XFILL_0__10630_ gnd vdd FILL
XFILL_3__11790_ gnd vdd FILL
X_15613_ _7584_/A gnd _15614_/D vdd INVX1
XFILL_5__12350_ gnd vdd FILL
XFILL_5__8891_ gnd vdd FILL
XFILL_4__10011_ gnd vdd FILL
X_12825_ _12823_/Y vdd _12825_/C gnd _12919_/D vdd OAI21X1
XFILL_1_BUFX2_insert410 gnd vdd FILL
XFILL_1_BUFX2_insert421 gnd vdd FILL
XFILL_1__11920_ gnd vdd FILL
XFILL_2__12170_ gnd vdd FILL
XFILL_1_BUFX2_insert432 gnd vdd FILL
XSFILL74120x19050 gnd vdd FILL
XFILL_1_BUFX2_insert443 gnd vdd FILL
XFILL_5__7842_ gnd vdd FILL
XFILL_5__11301_ gnd vdd FILL
XFILL_0__10561_ gnd vdd FILL
XFILL_1_BUFX2_insert454 gnd vdd FILL
X_15544_ _15544_/A _15544_/B _15384_/D _14053_/Y gnd _15545_/C vdd OAI22X1
X_12756_ _12718_/B memoryOutData[20] gnd _12757_/C vdd NAND2X1
XFILL_5__12281_ gnd vdd FILL
XFILL_2__11121_ gnd vdd FILL
XFILL_1_BUFX2_insert465 gnd vdd FILL
XFILL_3__13460_ gnd vdd FILL
XFILL_1_BUFX2_insert476 gnd vdd FILL
XFILL_0__12300_ gnd vdd FILL
XFILL_3__10672_ gnd vdd FILL
XFILL_1_BUFX2_insert487 gnd vdd FILL
XFILL_1__11851_ gnd vdd FILL
XFILL_0__13280_ gnd vdd FILL
XFILL_5__14020_ gnd vdd FILL
XFILL_1_BUFX2_insert498 gnd vdd FILL
X_11707_ _12262_/Y _12150_/Y _11682_/B gnd _11708_/C vdd OAI21X1
XFILL_0__10492_ gnd vdd FILL
XFILL_5__11232_ gnd vdd FILL
XFILL_3__12411_ gnd vdd FILL
XFILL_2__9803_ gnd vdd FILL
XFILL_4__14750_ gnd vdd FILL
X_15475_ _15475_/A gnd _15476_/B vdd INVX1
X_12687_ _12639_/A _7005_/CLK _7133_/R vdd _12687_/D gnd vdd DFFSR
XFILL_4__11962_ gnd vdd FILL
XFILL_2__11052_ gnd vdd FILL
XFILL_1__10802_ gnd vdd FILL
XFILL_1__14570_ gnd vdd FILL
XFILL_5__9512_ gnd vdd FILL
XFILL_3__13391_ gnd vdd FILL
XFILL_0__12231_ gnd vdd FILL
XFILL_2__7995_ gnd vdd FILL
XFILL_1__11782_ gnd vdd FILL
XSFILL23160x59050 gnd vdd FILL
XFILL_4__13701_ gnd vdd FILL
X_14426_ _14426_/A _14506_/C _14718_/C _14425_/Y gnd _14430_/B vdd OAI22X1
XFILL_4__10913_ gnd vdd FILL
XFILL_5__11163_ gnd vdd FILL
XFILL_2__10003_ gnd vdd FILL
X_11638_ _11638_/A _11637_/Y _11631_/Y gnd _12053_/A vdd NAND3X1
XFILL_3__15130_ gnd vdd FILL
XSFILL109720x68050 gnd vdd FILL
XFILL_3__12342_ gnd vdd FILL
XFILL_4__14681_ gnd vdd FILL
XFILL_2__9734_ gnd vdd FILL
XFILL_1__13521_ gnd vdd FILL
XFILL_2__6946_ gnd vdd FILL
XFILL_4__11893_ gnd vdd FILL
XFILL_2__15860_ gnd vdd FILL
XFILL_0__12162_ gnd vdd FILL
XFILL_5__10114_ gnd vdd FILL
XFILL_4__13632_ gnd vdd FILL
X_14357_ _14357_/A _14357_/B _15812_/C gnd _13006_/B vdd AOI21X1
XFILL_5__15971_ gnd vdd FILL
XFILL_2__14811_ gnd vdd FILL
XFILL_3__15061_ gnd vdd FILL
XFILL_5__11094_ gnd vdd FILL
X_11569_ _11630_/B _11569_/B _11569_/C gnd _11570_/A vdd OAI21X1
XFILL_1__16240_ gnd vdd FILL
XFILL_1__13452_ gnd vdd FILL
XSFILL38360x40050 gnd vdd FILL
XFILL_3__12273_ gnd vdd FILL
XFILL_2__9665_ gnd vdd FILL
XFILL_0__11113_ gnd vdd FILL
XFILL_1__10664_ gnd vdd FILL
XFILL_2__6877_ gnd vdd FILL
XFILL_2__15791_ gnd vdd FILL
X_13308_ _13308_/A _13308_/B gnd _13308_/Y vdd NAND2X1
XFILL_0__12093_ gnd vdd FILL
XFILL_0__7700_ gnd vdd FILL
XFILL_5__9374_ gnd vdd FILL
XFILL_5__10045_ gnd vdd FILL
XFILL_3__14012_ gnd vdd FILL
XFILL_4__16351_ gnd vdd FILL
XFILL_5__14922_ gnd vdd FILL
XFILL_2__8616_ gnd vdd FILL
XFILL_1__12403_ gnd vdd FILL
XFILL_4__13563_ gnd vdd FILL
XFILL_3__11224_ gnd vdd FILL
X_14288_ _14288_/A _14287_/Y gnd _14288_/Y vdd NOR2X1
XFILL_1__16171_ gnd vdd FILL
XSFILL79240x52050 gnd vdd FILL
XFILL_4__10775_ gnd vdd FILL
XFILL_2__14742_ gnd vdd FILL
XFILL_0__15921_ gnd vdd FILL
XFILL_2__11954_ gnd vdd FILL
XFILL_1__13383_ gnd vdd FILL
XFILL_2__9596_ gnd vdd FILL
XFILL_0__11044_ gnd vdd FILL
XFILL_5__8325_ gnd vdd FILL
X_16027_ _16027_/A _16024_/Y gnd _16033_/B vdd NOR2X1
XFILL_4__15302_ gnd vdd FILL
X_13239_ _13281_/B _13239_/B gnd _13242_/B vdd NOR2X1
XFILL_0__7631_ gnd vdd FILL
XFILL_4__12514_ gnd vdd FILL
XFILL_5__14853_ gnd vdd FILL
XFILL_3__11155_ gnd vdd FILL
XFILL_1__15122_ gnd vdd FILL
XFILL_4__16282_ gnd vdd FILL
XFILL_2__10905_ gnd vdd FILL
XFILL_4__13494_ gnd vdd FILL
XFILL_3__7340_ gnd vdd FILL
XFILL_1__12334_ gnd vdd FILL
XFILL_2__14673_ gnd vdd FILL
XFILL_5__8256_ gnd vdd FILL
XSFILL83720x77050 gnd vdd FILL
XFILL_2__11885_ gnd vdd FILL
XSFILL114440x61050 gnd vdd FILL
XFILL_0__15852_ gnd vdd FILL
XFILL_5__13804_ gnd vdd FILL
XFILL_4__15233_ gnd vdd FILL
XFILL_0__7562_ gnd vdd FILL
XFILL_3__10106_ gnd vdd FILL
XFILL_4__12445_ gnd vdd FILL
XFILL_2__16412_ gnd vdd FILL
XFILL_2__13624_ gnd vdd FILL
XSFILL18920x67050 gnd vdd FILL
XFILL_1__15053_ gnd vdd FILL
XFILL_5__11996_ gnd vdd FILL
XFILL_3__15963_ gnd vdd FILL
XFILL_3__11086_ gnd vdd FILL
XFILL_5__14784_ gnd vdd FILL
XFILL_0__14803_ gnd vdd FILL
XFILL_5__7207_ gnd vdd FILL
XSFILL84360x43050 gnd vdd FILL
XFILL_1__12265_ gnd vdd FILL
XFILL_2__8478_ gnd vdd FILL
XFILL_2__10836_ gnd vdd FILL
XFILL_0__15783_ gnd vdd FILL
XFILL_0__9301_ gnd vdd FILL
XFILL_0__12995_ gnd vdd FILL
XFILL_5__8187_ gnd vdd FILL
XFILL_5__10947_ gnd vdd FILL
XFILL_3__10037_ gnd vdd FILL
XFILL_1__14004_ gnd vdd FILL
XFILL_0__7493_ gnd vdd FILL
XFILL_4__15164_ gnd vdd FILL
XFILL_3__9010_ gnd vdd FILL
XFILL_5__13735_ gnd vdd FILL
XFILL_3__14914_ gnd vdd FILL
XFILL_2__16343_ gnd vdd FILL
XFILL_4__12376_ gnd vdd FILL
XFILL_2__7429_ gnd vdd FILL
XFILL_1__11216_ gnd vdd FILL
XFILL_2__10767_ gnd vdd FILL
XFILL_3__15894_ gnd vdd FILL
XFILL_0__14734_ gnd vdd FILL
XFILL_2__13555_ gnd vdd FILL
XSFILL99400x65050 gnd vdd FILL
XFILL_0__11946_ gnd vdd FILL
XFILL_1__12196_ gnd vdd FILL
XFILL_0__9232_ gnd vdd FILL
XFILL_4__14115_ gnd vdd FILL
X_9860_ _9858_/Y _9868_/A _9859_/Y gnd _9946_/D vdd OAI21X1
XFILL_5__13666_ gnd vdd FILL
XFILL_4__11327_ gnd vdd FILL
XFILL_3__14845_ gnd vdd FILL
XFILL_2__12506_ gnd vdd FILL
XFILL_5__10878_ gnd vdd FILL
XFILL_4__15095_ gnd vdd FILL
XFILL_1__11147_ gnd vdd FILL
XFILL_2__16274_ gnd vdd FILL
XFILL_2__10698_ gnd vdd FILL
XFILL_2__13486_ gnd vdd FILL
XFILL_0__14665_ gnd vdd FILL
XFILL_5__12617_ gnd vdd FILL
XFILL_0__11877_ gnd vdd FILL
XFILL_5__15405_ gnd vdd FILL
XFILL_0__9163_ gnd vdd FILL
XFILL_5__7069_ gnd vdd FILL
XSFILL38840x18050 gnd vdd FILL
X_8811_ _8811_/Q _7147_/CLK _7133_/R vdd _8811_/D gnd vdd DFFSR
XFILL_4__14046_ gnd vdd FILL
XFILL112360x25050 gnd vdd FILL
XFILL_5__13597_ gnd vdd FILL
X_9791_ _9764_/A _7743_/B gnd _9792_/C vdd NAND2X1
XFILL_5__16385_ gnd vdd FILL
XFILL_2__15225_ gnd vdd FILL
XFILL_4__11258_ gnd vdd FILL
XFILL_2__12437_ gnd vdd FILL
XFILL_0__13616_ gnd vdd FILL
XFILL_0__16404_ gnd vdd FILL
XFILL_3__14776_ gnd vdd FILL
XFILL_0__10828_ gnd vdd FILL
XFILL_3__11988_ gnd vdd FILL
XFILL_1__15955_ gnd vdd FILL
XFILL_1__11078_ gnd vdd FILL
XFILL_0__14596_ gnd vdd FILL
XFILL_0__8114_ gnd vdd FILL
XSFILL24120x67050 gnd vdd FILL
X_8742_ _8806_/Q gnd _8742_/Y vdd INVX1
XFILL_5__15336_ gnd vdd FILL
XFILL_0__9094_ gnd vdd FILL
XSFILL109400x50050 gnd vdd FILL
XFILL_3__9912_ gnd vdd FILL
XFILL_3__13727_ gnd vdd FILL
XFILL_3__10939_ gnd vdd FILL
XFILL_2__12368_ gnd vdd FILL
XFILL_0__16335_ gnd vdd FILL
XFILL_1__10029_ gnd vdd FILL
XFILL_2__15156_ gnd vdd FILL
XFILL_4__11189_ gnd vdd FILL
XFILL_1__14906_ gnd vdd FILL
XFILL_0__13547_ gnd vdd FILL
XSFILL79320x32050 gnd vdd FILL
XFILL_0__10759_ gnd vdd FILL
XFILL_1__15886_ gnd vdd FILL
XFILL_6__13838_ gnd vdd FILL
XFILL_5__15267_ gnd vdd FILL
XSFILL3560x58050 gnd vdd FILL
XFILL_6_BUFX2_insert648 gnd vdd FILL
X_8673_ _8599_/A _9818_/CLK _9441_/R vdd _8673_/D gnd vdd DFFSR
XFILL_5__12479_ gnd vdd FILL
XFILL_2__14107_ gnd vdd FILL
XFILL_2__11319_ gnd vdd FILL
XFILL_3__13658_ gnd vdd FILL
XFILL_6_BUFX2_insert659 gnd vdd FILL
XFILL_1__14837_ gnd vdd FILL
XFILL_4__15997_ gnd vdd FILL
XFILL_2__12299_ gnd vdd FILL
XFILL_2__15087_ gnd vdd FILL
XFILL_0__16266_ gnd vdd FILL
XFILL_5__14218_ gnd vdd FILL
XFILL_0__13478_ gnd vdd FILL
X_7624_ _7624_/A _7240_/B gnd _7625_/C vdd NAND2X1
XFILL_5__15198_ gnd vdd FILL
XFILL_3__12609_ gnd vdd FILL
XSFILL109560x5050 gnd vdd FILL
XFILL_0__15217_ gnd vdd FILL
XSFILL114520x41050 gnd vdd FILL
XFILL_2__14038_ gnd vdd FILL
XFILL_4__14948_ gnd vdd FILL
XFILL_3__16377_ gnd vdd FILL
XFILL_3__13589_ gnd vdd FILL
XFILL_0__12429_ gnd vdd FILL
XFILL_3__9774_ gnd vdd FILL
XSFILL44040x18050 gnd vdd FILL
XFILL_3__6986_ gnd vdd FILL
XFILL_0__16197_ gnd vdd FILL
XFILL_1__14768_ gnd vdd FILL
XFILL_6__9483_ gnd vdd FILL
XFILL_5__14149_ gnd vdd FILL
XFILL_3__15328_ gnd vdd FILL
X_7555_ _7606_/A _7555_/B gnd _7556_/C vdd NAND2X1
XSFILL84440x23050 gnd vdd FILL
XFILL_0__9996_ gnd vdd FILL
XFILL_4__14879_ gnd vdd FILL
XFILL_3__8725_ gnd vdd FILL
XFILL_0__15148_ gnd vdd FILL
XFILL_1__13719_ gnd vdd FILL
XFILL_1_CLKBUF1_insert119 gnd vdd FILL
XFILL_1__14699_ gnd vdd FILL
XFILL_6__15439_ gnd vdd FILL
XFILL_1__7740_ gnd vdd FILL
X_7486_ _7534_/Q gnd _7486_/Y vdd INVX1
XFILL_3__15259_ gnd vdd FILL
XFILL_3__8656_ gnd vdd FILL
XFILL_2__15989_ gnd vdd FILL
XFILL_0__15079_ gnd vdd FILL
X_9225_ _9277_/B _9353_/B gnd _9226_/C vdd NAND2X1
XFILL_3__7607_ gnd vdd FILL
XFILL_1__7671_ gnd vdd FILL
XFILL_0__8878_ gnd vdd FILL
XFILL_3__8587_ gnd vdd FILL
XSFILL33480x63050 gnd vdd FILL
XFILL_1__16369_ gnd vdd FILL
XFILL_4__7380_ gnd vdd FILL
XFILL_1__9410_ gnd vdd FILL
X_9156_ _9200_/Q gnd _9158_/A vdd INVX1
XFILL_0__7829_ gnd vdd FILL
XFILL_3_BUFX2_insert505 gnd vdd FILL
XFILL_3_BUFX2_insert516 gnd vdd FILL
X_8107_ _8107_/A _8107_/B _8107_/C gnd _8167_/D vdd OAI21X1
XFILL_1__9341_ gnd vdd FILL
XFILL_3_BUFX2_insert527 gnd vdd FILL
X_9087_ _9177_/Q gnd _9089_/A vdd INVX1
XFILL_3_BUFX2_insert538 gnd vdd FILL
XFILL_3_BUFX2_insert549 gnd vdd FILL
XFILL_3__7469_ gnd vdd FILL
XSFILL3640x38050 gnd vdd FILL
X_8038_ _8038_/Q _8038_/CLK _8038_/R vdd _7976_/Y gnd vdd DFFSR
XFILL_6__7178_ gnd vdd FILL
XSFILL88760x4050 gnd vdd FILL
XSFILL12760x64050 gnd vdd FILL
XFILL_3__9208_ gnd vdd FILL
XFILL_1__9272_ gnd vdd FILL
XFILL_4__8001_ gnd vdd FILL
XSFILL94280x26050 gnd vdd FILL
XFILL_1__8223_ gnd vdd FILL
XFILL_3__9139_ gnd vdd FILL
XSFILL54280x42050 gnd vdd FILL
X_10940_ _12788_/A _10939_/Y gnd _10940_/Y vdd NAND2X1
X_9989_ _9989_/A gnd _9989_/Y vdd INVX1
XFILL_1__7105_ gnd vdd FILL
X_10871_ _12710_/A _10871_/B gnd _10871_/Y vdd NAND2X1
XFILL_1__8085_ gnd vdd FILL
XFILL_4__8903_ gnd vdd FILL
X_12610_ vdd memoryOutData[14] gnd _12611_/C vdd NAND2X1
XFILL_4__9883_ gnd vdd FILL
XFILL_1__7036_ gnd vdd FILL
X_13590_ _13846_/A _13588_/Y _13590_/C _14203_/B gnd _13590_/Y vdd OAI22X1
XSFILL104520x73050 gnd vdd FILL
XFILL_4__8834_ gnd vdd FILL
XSFILL8760x71050 gnd vdd FILL
XFILL_0_BUFX2_insert406 gnd vdd FILL
X_12541_ _12361_/A _9060_/CLK _9060_/R vdd _12459_/Y gnd vdd DFFSR
XSFILL23800x20050 gnd vdd FILL
XFILL_0_BUFX2_insert417 gnd vdd FILL
XFILL_0_BUFX2_insert428 gnd vdd FILL
XFILL_0_BUFX2_insert439 gnd vdd FILL
XSFILL89240x15050 gnd vdd FILL
XFILL_4__8765_ gnd vdd FILL
X_15260_ _8795_/Q _15821_/B _15978_/C _8453_/A gnd _15265_/A vdd AOI22X1
X_12472_ _12031_/B gnd _12474_/A vdd INVX1
XFILL_4__7716_ gnd vdd FILL
XFILL_1__8987_ gnd vdd FILL
XSFILL3720x18050 gnd vdd FILL
X_14211_ _14211_/A _14210_/Y _13882_/B _15663_/B gnd _14212_/B vdd OAI22X1
XFILL_4__8696_ gnd vdd FILL
X_11423_ _11203_/Y _11423_/B _11423_/C gnd _11424_/B vdd OAI21X1
X_15191_ _15681_/C _15190_/Y _15191_/C _15394_/C gnd _15192_/B vdd OAI22X1
XFILL_1__7938_ gnd vdd FILL
X_14142_ _14142_/A _14138_/Y gnd _14142_/Y vdd NOR2X1
X_11354_ _11351_/Y _11353_/Y _11354_/C gnd _11354_/Y vdd OAI21X1
XFILL_1__7869_ gnd vdd FILL
XSFILL13720x72050 gnd vdd FILL
XSFILL94600x68050 gnd vdd FILL
XSFILL78680x60050 gnd vdd FILL
X_10305_ _10305_/A gnd _10305_/Y vdd INVX1
XSFILL79160x67050 gnd vdd FILL
XFILL_4__7578_ gnd vdd FILL
XFILL_4_BUFX2_insert350 gnd vdd FILL
XFILL_1__9608_ gnd vdd FILL
X_14073_ _14073_/A _14065_/Y _14073_/C gnd _14074_/B vdd NAND3X1
X_11285_ _11285_/A gnd _11646_/A vdd INVX2
XFILL_4_BUFX2_insert361 gnd vdd FILL
XFILL_2__8401_ gnd vdd FILL
XFILL_4_BUFX2_insert372 gnd vdd FILL
XFILL_4__10560_ gnd vdd FILL
XFILL_2__9381_ gnd vdd FILL
XFILL_5__8110_ gnd vdd FILL
XCLKBUF1_insert118 CLKBUF1_insert169/A gnd _7156_/CLK vdd CLKBUF1
XFILL_1__10380_ gnd vdd FILL
XFILL_4_BUFX2_insert383 gnd vdd FILL
XFILL_5__9090_ gnd vdd FILL
X_13024_ vdd _13024_/B gnd _13025_/C vdd NAND2X1
XFILL_4_BUFX2_insert394 gnd vdd FILL
X_10236_ _13537_/A gnd _10236_/Y vdd INVX1
XCLKBUF1_insert129 CLKBUF1_insert193/A gnd _7527_/CLK vdd CLKBUF1
XFILL_5__11850_ gnd vdd FILL
XFILL_2__8332_ gnd vdd FILL
XFILL_1__9539_ gnd vdd FILL
XFILL_2__11670_ gnd vdd FILL
XFILL_4__10491_ gnd vdd FILL
XFILL_4__9248_ gnd vdd FILL
XFILL_5__10801_ gnd vdd FILL
X_10167_ _10165_/Y _10166_/A _10167_/C gnd _10219_/D vdd OAI21X1
XSFILL84280x58050 gnd vdd FILL
XFILL_4__12230_ gnd vdd FILL
XFILL_2__10621_ gnd vdd FILL
XFILL_5__11781_ gnd vdd FILL
XFILL_3__12960_ gnd vdd FILL
XFILL_1__12050_ gnd vdd FILL
XFILL_0__11800_ gnd vdd FILL
XFILL_2__8263_ gnd vdd FILL
XFILL_0__12780_ gnd vdd FILL
XFILL_5__13520_ gnd vdd FILL
X_10098_ _10098_/Q _7282_/CLK _7411_/R vdd _10098_/D gnd vdd DFFSR
XFILL_3__11911_ gnd vdd FILL
XFILL_4__12161_ gnd vdd FILL
XFILL_2__7214_ gnd vdd FILL
X_14975_ _14974_/Y _14975_/B gnd _14975_/Y vdd NOR2X1
XFILL_1__11001_ gnd vdd FILL
XFILL_2__13340_ gnd vdd FILL
XFILL_2__10552_ gnd vdd FILL
XFILL_2__8194_ gnd vdd FILL
XSFILL34520x51050 gnd vdd FILL
XFILL_3__12891_ gnd vdd FILL
XFILL_0__11731_ gnd vdd FILL
XFILL_6__14810_ gnd vdd FILL
XFILL_5__9992_ gnd vdd FILL
XFILL_5__13451_ gnd vdd FILL
XFILL_4__11112_ gnd vdd FILL
X_13926_ _8671_/Q _13864_/B _14403_/C _8465_/A gnd _13928_/A vdd AOI22X1
XFILL_3__14630_ gnd vdd FILL
XFILL_5__10663_ gnd vdd FILL
XFILL_2__13271_ gnd vdd FILL
XFILL_4__12092_ gnd vdd FILL
XFILL_3__11842_ gnd vdd FILL
XFILL_0__14450_ gnd vdd FILL
XFILL_5__12402_ gnd vdd FILL
XFILL_0__11662_ gnd vdd FILL
XFILL_5__16170_ gnd vdd FILL
XFILL_4__15920_ gnd vdd FILL
X_13857_ _13856_/Y _13857_/B _13857_/C _13855_/Y gnd _13857_/Y vdd OAI22X1
XFILL_5__13382_ gnd vdd FILL
XFILL_2__15010_ gnd vdd FILL
XFILL_4__11043_ gnd vdd FILL
XFILL_2__12222_ gnd vdd FILL
XFILL_2__7076_ gnd vdd FILL
XFILL_3__14561_ gnd vdd FILL
XFILL_0__13401_ gnd vdd FILL
XFILL_1__15740_ gnd vdd FILL
XFILL_3__11773_ gnd vdd FILL
XFILL_1__12952_ gnd vdd FILL
XFILL_0__14381_ gnd vdd FILL
XFILL_5__15121_ gnd vdd FILL
X_12808_ _12808_/Q _12685_/CLK _12685_/R vdd _12808_/D gnd vdd DFFSR
XSFILL63960x80050 gnd vdd FILL
XFILL_1_BUFX2_insert240 gnd vdd FILL
XFILL_3__16300_ gnd vdd FILL
XFILL_5__12333_ gnd vdd FILL
XFILL_0__11593_ gnd vdd FILL
XFILL_5__8874_ gnd vdd FILL
XSFILL74200x8050 gnd vdd FILL
XSFILL13800x52050 gnd vdd FILL
XSFILL113800x8050 gnd vdd FILL
XFILL_6__14672_ gnd vdd FILL
XFILL_3__13512_ gnd vdd FILL
XFILL_1_BUFX2_insert251 gnd vdd FILL
X_13788_ _13788_/A _13788_/B gnd _13789_/B vdd NOR2X1
XFILL_0__16120_ gnd vdd FILL
XFILL_2__12153_ gnd vdd FILL
XFILL_4__15851_ gnd vdd FILL
XFILL_1_BUFX2_insert262 gnd vdd FILL
XFILL_3__14492_ gnd vdd FILL
XFILL_0__13332_ gnd vdd FILL
XSFILL79240x47050 gnd vdd FILL
XFILL_1__11903_ gnd vdd FILL
XFILL_1_BUFX2_insert273 gnd vdd FILL
XFILL_1__15671_ gnd vdd FILL
XFILL_0__10544_ gnd vdd FILL
XFILL_6__16411_ gnd vdd FILL
XFILL_5__7825_ gnd vdd FILL
XFILL_1__12883_ gnd vdd FILL
XFILL_6__13623_ gnd vdd FILL
X_15527_ _15527_/A _15527_/B _15527_/C _15527_/D gnd _15527_/Y vdd OAI22X1
XFILL_1_BUFX2_insert284 gnd vdd FILL
XFILL_5__15052_ gnd vdd FILL
XFILL_1_BUFX2_insert295 gnd vdd FILL
X_12739_ _12737_/Y _12768_/A _12739_/C gnd _12739_/Y vdd OAI21X1
XFILL_3__16231_ gnd vdd FILL
XFILL_4__14802_ gnd vdd FILL
XFILL_5__12264_ gnd vdd FILL
XFILL_2__11104_ gnd vdd FILL
XFILL_3__13443_ gnd vdd FILL
XFILL_4__15782_ gnd vdd FILL
XFILL_1__14622_ gnd vdd FILL
XFILL_2__12084_ gnd vdd FILL
XFILL_4__12994_ gnd vdd FILL
XFILL_3__6840_ gnd vdd FILL
XFILL_3__10655_ gnd vdd FILL
XFILL_0__16051_ gnd vdd FILL
XFILL_1__11834_ gnd vdd FILL
XFILL_0__13263_ gnd vdd FILL
XFILL_5__14003_ gnd vdd FILL
XFILL_5__7756_ gnd vdd FILL
XFILL_0_BUFX2_insert940 gnd vdd FILL
XFILL_5__11215_ gnd vdd FILL
XFILL_4__14733_ gnd vdd FILL
XFILL_0__9850_ gnd vdd FILL
X_15458_ _15458_/A _16089_/B gnd _15458_/Y vdd NOR2X1
XFILL_2__15912_ gnd vdd FILL
XFILL_0__15002_ gnd vdd FILL
XFILL_0_BUFX2_insert951 gnd vdd FILL
XFILL_4__11945_ gnd vdd FILL
XFILL_5__12195_ gnd vdd FILL
XFILL_3__16162_ gnd vdd FILL
XFILL_2__11035_ gnd vdd FILL
XFILL_0_BUFX2_insert962 gnd vdd FILL
XFILL_3__13374_ gnd vdd FILL
XFILL_0__12214_ gnd vdd FILL
XFILL_1__14553_ gnd vdd FILL
XFILL_0_BUFX2_insert973 gnd vdd FILL
XSFILL84360x38050 gnd vdd FILL
XFILL_2__7978_ gnd vdd FILL
XFILL_1__11765_ gnd vdd FILL
XFILL_6__12505_ gnd vdd FILL
X_14409_ _7786_/Q gnd _14410_/B vdd INVX1
XFILL_0_BUFX2_insert984 gnd vdd FILL
X_7340_ _7400_/Q gnd _7340_/Y vdd INVX1
XFILL_5__11146_ gnd vdd FILL
XFILL_5__7687_ gnd vdd FILL
XFILL_3__15113_ gnd vdd FILL
XFILL_6__16273_ gnd vdd FILL
XFILL_0__9781_ gnd vdd FILL
XFILL_0_BUFX2_insert995 gnd vdd FILL
X_15389_ _15389_/A _15381_/Y gnd _15414_/B vdd NOR2X1
XFILL_3__8510_ gnd vdd FILL
XFILL_4__14664_ gnd vdd FILL
XFILL_6__13485_ gnd vdd FILL
XFILL_6__10697_ gnd vdd FILL
XFILL_3__12325_ gnd vdd FILL
XFILL_4__11876_ gnd vdd FILL
XFILL_3__16093_ gnd vdd FILL
XFILL_2__15843_ gnd vdd FILL
XFILL_2__6929_ gnd vdd FILL
XFILL_1__13504_ gnd vdd FILL
XFILL_0__6993_ gnd vdd FILL
XFILL_1__14484_ gnd vdd FILL
XFILL_0__12145_ gnd vdd FILL
XFILL_3__9490_ gnd vdd FILL
XFILL_5__9426_ gnd vdd FILL
XFILL_6__15224_ gnd vdd FILL
XFILL_1__11696_ gnd vdd FILL
XSFILL59160x14050 gnd vdd FILL
XFILL_4__13615_ gnd vdd FILL
XFILL_0__8732_ gnd vdd FILL
XFILL_4__16403_ gnd vdd FILL
XFILL_4__10827_ gnd vdd FILL
XFILL_3__15044_ gnd vdd FILL
XFILL_5__15954_ gnd vdd FILL
XFILL_5__11077_ gnd vdd FILL
X_7271_ _7271_/Q _9447_/CLK _9447_/R vdd _7271_/D gnd vdd DFFSR
XFILL_4__14595_ gnd vdd FILL
XFILL_1__16223_ gnd vdd FILL
XFILL_1__13435_ gnd vdd FILL
XFILL_2__9648_ gnd vdd FILL
XFILL_3__12256_ gnd vdd FILL
XFILL_3__8441_ gnd vdd FILL
XFILL_1__10647_ gnd vdd FILL
XFILL_2__15774_ gnd vdd FILL
XFILL_5__9357_ gnd vdd FILL
XFILL_0__12076_ gnd vdd FILL
XFILL_2__12986_ gnd vdd FILL
X_9010_ _9066_/Q gnd _9012_/A vdd INVX1
XFILL_6__12367_ gnd vdd FILL
XFILL_4__16334_ gnd vdd FILL
XFILL_5__10028_ gnd vdd FILL
XFILL111880x13050 gnd vdd FILL
XFILL_5__14905_ gnd vdd FILL
XFILL_4__13546_ gnd vdd FILL
XFILL_3__11207_ gnd vdd FILL
XFILL_2__14725_ gnd vdd FILL
XFILL_4__10758_ gnd vdd FILL
XFILL_5__15885_ gnd vdd FILL
XFILL_0__15904_ gnd vdd FILL
XFILL_3__12187_ gnd vdd FILL
XFILL_1__13366_ gnd vdd FILL
XFILL_2__11937_ gnd vdd FILL
XFILL_3__8372_ gnd vdd FILL
XFILL_0__11027_ gnd vdd FILL
XFILL_1__16154_ gnd vdd FILL
XFILL_1__10578_ gnd vdd FILL
XFILL_0__7614_ gnd vdd FILL
XFILL_5__9288_ gnd vdd FILL
XFILL_6__11318_ gnd vdd FILL
XFILL_5__14836_ gnd vdd FILL
XFILL_6__15086_ gnd vdd FILL
XFILL_4__16265_ gnd vdd FILL
XSFILL109400x45050 gnd vdd FILL
XFILL_3__7323_ gnd vdd FILL
XFILL_3__11138_ gnd vdd FILL
XSFILL38440x15050 gnd vdd FILL
XFILL_0__8594_ gnd vdd FILL
XFILL_1__15105_ gnd vdd FILL
XFILL_4__13477_ gnd vdd FILL
XFILL_1__12317_ gnd vdd FILL
XFILL_2__14656_ gnd vdd FILL
XFILL_1__16085_ gnd vdd FILL
XFILL_4__10689_ gnd vdd FILL
XFILL_1__13297_ gnd vdd FILL
XFILL_0__15835_ gnd vdd FILL
XFILL_2__11868_ gnd vdd FILL
XFILL_5__8239_ gnd vdd FILL
XFILL_4__15216_ gnd vdd FILL
XFILL_6__14037_ gnd vdd FILL
XFILL_4__12428_ gnd vdd FILL
XSFILL49080x66050 gnd vdd FILL
XSFILL79320x27050 gnd vdd FILL
XFILL_0__7545_ gnd vdd FILL
XFILL_2__13607_ gnd vdd FILL
XFILL_4__16196_ gnd vdd FILL
XFILL_1__15036_ gnd vdd FILL
XFILL_3__15946_ gnd vdd FILL
XFILL_5__11979_ gnd vdd FILL
XFILL_5__14767_ gnd vdd FILL
XFILL_1__12248_ gnd vdd FILL
XFILL_2__10819_ gnd vdd FILL
XFILL_3__11069_ gnd vdd FILL
XFILL_2__14587_ gnd vdd FILL
XSFILL39320x43050 gnd vdd FILL
XFILL_0__15766_ gnd vdd FILL
XFILL_0__12978_ gnd vdd FILL
XFILL_2__11799_ gnd vdd FILL
XFILL_5__13718_ gnd vdd FILL
X_9912_ _9964_/Q gnd _9912_/Y vdd INVX1
XFILL_4__15147_ gnd vdd FILL
XFILL_4__12359_ gnd vdd FILL
XFILL_2__16326_ gnd vdd FILL
XFILL_0__7476_ gnd vdd FILL
XSFILL114520x36050 gnd vdd FILL
XFILL_5__14698_ gnd vdd FILL
XFILL_2__13538_ gnd vdd FILL
XFILL_3__15877_ gnd vdd FILL
XFILL_1__12179_ gnd vdd FILL
XFILL_0__11929_ gnd vdd FILL
XFILL_0__14717_ gnd vdd FILL
XFILL_3__7185_ gnd vdd FILL
XFILL_0__9215_ gnd vdd FILL
XFILL_0__15697_ gnd vdd FILL
X_9843_ _9843_/Q _8051_/CLK _8051_/R vdd _9843_/D gnd vdd DFFSR
XFILL_5__13649_ gnd vdd FILL
XFILL_3__14828_ gnd vdd FILL
XFILL_4__15078_ gnd vdd FILL
XFILL_2__16257_ gnd vdd FILL
XFILL_2__13469_ gnd vdd FILL
XFILL_0__14648_ gnd vdd FILL
XSFILL83400x54050 gnd vdd FILL
XFILL_4__14029_ gnd vdd FILL
XFILL_0__9146_ gnd vdd FILL
XFILL_2__15208_ gnd vdd FILL
XSFILL69080x1050 gnd vdd FILL
XFILL_5__16368_ gnd vdd FILL
X_6986_ _6986_/A gnd _6988_/A vdd INVX1
XSFILL18600x44050 gnd vdd FILL
X_9774_ _9774_/A _9770_/A _9773_/Y gnd _9832_/D vdd OAI21X1
XFILL_3__14759_ gnd vdd FILL
XFILL_2__16188_ gnd vdd FILL
XFILL_1__15938_ gnd vdd FILL
XFILL_0__14579_ gnd vdd FILL
XFILL_5__15319_ gnd vdd FILL
XFILL_6_BUFX2_insert423 gnd vdd FILL
X_8725_ _8788_/A _6933_/B gnd _8726_/C vdd NAND2X1
XFILL_6_BUFX2_insert434 gnd vdd FILL
XFILL_5__16299_ gnd vdd FILL
XFILL_2__15139_ gnd vdd FILL
XFILL_0__16318_ gnd vdd FILL
XFILL_1__15869_ gnd vdd FILL
XFILL_4__6880_ gnd vdd FILL
XFILL_1__8910_ gnd vdd FILL
X_8656_ _8656_/A gnd _8656_/Y vdd INVX1
XFILL_1__9890_ gnd vdd FILL
XSFILL23720x35050 gnd vdd FILL
XFILL_0__16249_ gnd vdd FILL
XSFILL88680x23050 gnd vdd FILL
X_7607_ _7607_/A _7606_/A _7607_/C gnd _7659_/D vdd OAI21X1
XFILL_1__8841_ gnd vdd FILL
XFILL_4_BUFX2_insert1002 gnd vdd FILL
X_8587_ _8669_/Q gnd _8589_/A vdd INVX1
XSFILL18840x3050 gnd vdd FILL
XFILL_4_BUFX2_insert1013 gnd vdd FILL
XFILL_3__9757_ gnd vdd FILL
XFILL_4_BUFX2_insert1024 gnd vdd FILL
XFILL_3__6969_ gnd vdd FILL
XSFILL105000x4050 gnd vdd FILL
XFILL_4_BUFX2_insert1035 gnd vdd FILL
X_7538_ _7538_/Q _7406_/CLK _8430_/R vdd _7500_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert1046 gnd vdd FILL
XFILL_4__7501_ gnd vdd FILL
XFILL_3__8708_ gnd vdd FILL
XFILL_4_BUFX2_insert1057 gnd vdd FILL
XFILL_1__8772_ gnd vdd FILL
XFILL_0__9979_ gnd vdd FILL
XFILL_4__8481_ gnd vdd FILL
XFILL_4_BUFX2_insert1068 gnd vdd FILL
XSFILL114600x16050 gnd vdd FILL
XFILL_1__7723_ gnd vdd FILL
X_7469_ _7470_/B _9901_/B gnd _7469_/Y vdd NAND2X1
XFILL_3__8639_ gnd vdd FILL
XFILL_4__7432_ gnd vdd FILL
X_9208_ _9208_/A _9208_/B _9207_/Y gnd _9302_/D vdd OAI21X1
XFILL_4__7363_ gnd vdd FILL
XFILL_3_BUFX2_insert302 gnd vdd FILL
X_11070_ _12258_/Y gnd _11072_/A vdd INVX1
XSFILL69320x59050 gnd vdd FILL
XFILL_3_BUFX2_insert313 gnd vdd FILL
X_9139_ _9112_/A _9267_/B gnd _9139_/Y vdd NAND2X1
XFILL_4__9102_ gnd vdd FILL
XFILL_3_BUFX2_insert324 gnd vdd FILL
XFILL_1__7585_ gnd vdd FILL
X_10021_ _10019_/Y _9975_/B _10021_/C gnd _10085_/D vdd OAI21X1
XFILL_3_BUFX2_insert335 gnd vdd FILL
XFILL_2_BUFX2_insert1050 gnd vdd FILL
XFILL_4__7294_ gnd vdd FILL
XFILL_3_BUFX2_insert346 gnd vdd FILL
XFILL_3_BUFX2_insert357 gnd vdd FILL
XFILL_2_BUFX2_insert1061 gnd vdd FILL
XFILL_3_BUFX2_insert368 gnd vdd FILL
XFILL_2_BUFX2_insert1072 gnd vdd FILL
XFILL_4__9033_ gnd vdd FILL
XFILL_3_BUFX2_insert379 gnd vdd FILL
XSFILL73960x43050 gnd vdd FILL
XSFILL3480x3050 gnd vdd FILL
XFILL_1__9255_ gnd vdd FILL
XSFILL23800x15050 gnd vdd FILL
XSFILL84200x3050 gnd vdd FILL
XFILL_1__8206_ gnd vdd FILL
X_14760_ _14760_/A _14897_/D _13876_/C _16155_/C gnd _14761_/B vdd OAI22X1
X_11972_ _11909_/A _12427_/A gnd _11973_/C vdd NAND2X1
X_13711_ _13710_/Y _14200_/C _13479_/C _13711_/D gnd _13711_/Y vdd OAI22X1
X_10923_ _10929_/A _10906_/Y gnd _6837_/A vdd NOR2X1
XFILL_1__8137_ gnd vdd FILL
X_14691_ _14691_/A _14691_/B gnd _14692_/B vdd NOR2X1
XFILL_4__9935_ gnd vdd FILL
X_16430_ _14099_/A _8152_/CLK _8664_/R vdd _16430_/D gnd vdd DFFSR
X_13642_ _8066_/A gnd _13643_/D vdd INVX1
XFILL_4_CLKBUF1_insert114 gnd vdd FILL
X_10854_ _14252_/D _7411_/CLK _7411_/R vdd _10854_/D gnd vdd DFFSR
XFILL_2__8950_ gnd vdd FILL
XFILL_1__8068_ gnd vdd FILL
XFILL_4_CLKBUF1_insert125 gnd vdd FILL
XSFILL13720x67050 gnd vdd FILL
XFILL_4_CLKBUF1_insert136 gnd vdd FILL
XFILL_4__9866_ gnd vdd FILL
X_16361_ gnd gnd gnd _16362_/C vdd NAND2X1
XFILL_4_CLKBUF1_insert147 gnd vdd FILL
XFILL_4_CLKBUF1_insert158 gnd vdd FILL
X_13573_ _8828_/A gnd _13574_/A vdd INVX1
X_10785_ _10792_/B _7713_/B gnd _10785_/Y vdd NAND2X1
XFILL_4_CLKBUF1_insert169 gnd vdd FILL
XFILL_5__7610_ gnd vdd FILL
XFILL_2__8881_ gnd vdd FILL
XFILL_0_BUFX2_insert225 gnd vdd FILL
XSFILL39160x78050 gnd vdd FILL
X_15312_ _9352_/A _15380_/B gnd _15324_/A vdd NAND2X1
XFILL_5__8590_ gnd vdd FILL
X_12524_ vdd _12101_/A gnd _12525_/C vdd NAND2X1
XFILL_4__9797_ gnd vdd FILL
XFILL_0_BUFX2_insert236 gnd vdd FILL
XFILL_0_BUFX2_insert247 gnd vdd FILL
X_16292_ _9811_/A _15390_/B _16291_/Y gnd _16292_/Y vdd AOI21X1
XSFILL79560x83050 gnd vdd FILL
XFILL_2__7832_ gnd vdd FILL
XFILL_0_BUFX2_insert258 gnd vdd FILL
XFILL_3__10440_ gnd vdd FILL
XFILL_4__8748_ gnd vdd FILL
XFILL_0__10260_ gnd vdd FILL
XFILL_0_BUFX2_insert269 gnd vdd FILL
XFILL_5__11000_ gnd vdd FILL
X_15243_ _15220_/Y _15243_/B _15656_/B gnd _15243_/Y vdd AOI21X1
XSFILL69000x41050 gnd vdd FILL
X_12455_ vdd _12009_/A gnd _12455_/Y vdd NAND2X1
XSFILL3640x50 gnd vdd FILL
XFILL_4__11730_ gnd vdd FILL
XFILL_3__10371_ gnd vdd FILL
XFILL_2__7763_ gnd vdd FILL
XFILL_1__11550_ gnd vdd FILL
XFILL_0__10191_ gnd vdd FILL
XFILL_6__13270_ gnd vdd FILL
XFILL_5__7472_ gnd vdd FILL
X_11406_ _11150_/Y gnd _11406_/Y vdd INVX2
X_15174_ _15390_/B _9817_/Q _9689_/Q _15652_/D gnd _15176_/A vdd AOI22X1
XFILL_3__12110_ gnd vdd FILL
XFILL_2__9502_ gnd vdd FILL
X_12386_ _12371_/A _12609_/A gnd _12387_/C vdd NAND2X1
XSFILL59080x29050 gnd vdd FILL
XFILL_1__10501_ gnd vdd FILL
XFILL_4__11661_ gnd vdd FILL
XFILL_3__13090_ gnd vdd FILL
XFILL_2__12840_ gnd vdd FILL
XFILL_5__9211_ gnd vdd FILL
XFILL_2__7694_ gnd vdd FILL
XFILL_1__11481_ gnd vdd FILL
X_14125_ _14125_/A _14466_/C _14872_/C _14125_/D gnd _14129_/A vdd OAI22X1
XFILL_4__13400_ gnd vdd FILL
XSFILL99480x34050 gnd vdd FILL
XFILL_2_BUFX2_insert18 gnd vdd FILL
X_11337_ _11337_/A _11358_/B _11337_/C gnd _11338_/A vdd AOI21X1
XFILL_1__13220_ gnd vdd FILL
XFILL_2_BUFX2_insert29 gnd vdd FILL
XFILL_3__12041_ gnd vdd FILL
XFILL_5__12951_ gnd vdd FILL
XSFILL74120x32050 gnd vdd FILL
XFILL_4__14380_ gnd vdd FILL
XFILL_1__10432_ gnd vdd FILL
XFILL_4__11592_ gnd vdd FILL
XFILL_5__9142_ gnd vdd FILL
XFILL_2__12771_ gnd vdd FILL
XFILL_0__13950_ gnd vdd FILL
XFILL_6__12152_ gnd vdd FILL
XFILL_4__13331_ gnd vdd FILL
X_14056_ _9186_/Q gnd _14056_/Y vdd INVX1
XFILL_5__11902_ gnd vdd FILL
XFILL_5__15670_ gnd vdd FILL
XFILL_2__14510_ gnd vdd FILL
XFILL_5__12882_ gnd vdd FILL
XFILL_4__10543_ gnd vdd FILL
X_11268_ _11267_/Y gnd _11268_/Y vdd INVX1
XFILL_1__13151_ gnd vdd FILL
XFILL_0__12901_ gnd vdd FILL
XFILL_2__9364_ gnd vdd FILL
XFILL_2__11722_ gnd vdd FILL
XFILL_6__11103_ gnd vdd FILL
XFILL_1__10363_ gnd vdd FILL
XFILL_2__15490_ gnd vdd FILL
XFILL_0__13881_ gnd vdd FILL
X_13007_ _13005_/Y vdd _13007_/C gnd _13007_/Y vdd OAI21X1
X_10219_ _10219_/Q _9963_/CLK _9963_/R vdd _10219_/D gnd vdd DFFSR
XFILL_5__14621_ gnd vdd FILL
XFILL_3__15800_ gnd vdd FILL
XFILL_4__16050_ gnd vdd FILL
XFILL_5__11833_ gnd vdd FILL
XFILL_4__13262_ gnd vdd FILL
XFILL_1__12102_ gnd vdd FILL
XSFILL13800x47050 gnd vdd FILL
XFILL_2__8315_ gnd vdd FILL
X_11199_ _12334_/Y gnd _11199_/Y vdd INVX1
XSFILL78760x35050 gnd vdd FILL
XFILL_2__14441_ gnd vdd FILL
XFILL_2__9295_ gnd vdd FILL
XFILL_0__15620_ gnd vdd FILL
XFILL_0__12832_ gnd vdd FILL
XFILL_3__13992_ gnd vdd FILL
XFILL_1__13082_ gnd vdd FILL
XFILL_2__11653_ gnd vdd FILL
XFILL_1__10294_ gnd vdd FILL
XFILL_4__15001_ gnd vdd FILL
XFILL_0__7330_ gnd vdd FILL
XFILL_3_BUFX2_insert880 gnd vdd FILL
XFILL_4__12213_ gnd vdd FILL
XSFILL109720x81050 gnd vdd FILL
XFILL_3_BUFX2_insert891 gnd vdd FILL
XFILL_5__14552_ gnd vdd FILL
XFILL_3__15731_ gnd vdd FILL
XSFILL38760x51050 gnd vdd FILL
XFILL_5__11764_ gnd vdd FILL
XFILL_2__8246_ gnd vdd FILL
XFILL_1__12033_ gnd vdd FILL
XFILL_0__15551_ gnd vdd FILL
XFILL_2__14372_ gnd vdd FILL
XFILL_2__11584_ gnd vdd FILL
XFILL_0__12763_ gnd vdd FILL
XSFILL113960x44050 gnd vdd FILL
XFILL_5__13503_ gnd vdd FILL
XFILL_5__14483_ gnd vdd FILL
XFILL_2__16111_ gnd vdd FILL
X_14958_ _7763_/A gnd _14959_/B vdd INVX1
XFILL_4__12144_ gnd vdd FILL
XFILL_2__10535_ gnd vdd FILL
XFILL_2__13323_ gnd vdd FILL
XFILL_3__15662_ gnd vdd FILL
XFILL_0__14502_ gnd vdd FILL
XFILL_5__11695_ gnd vdd FILL
XFILL_3__12874_ gnd vdd FILL
XFILL_0__11714_ gnd vdd FILL
XFILL_0__9000_ gnd vdd FILL
XFILL_0__15482_ gnd vdd FILL
XFILL_5__16222_ gnd vdd FILL
XFILL_5__9975_ gnd vdd FILL
X_13909_ _13909_/A _14344_/B _14145_/D _7647_/Q gnd _13909_/Y vdd AOI22X1
XFILL_3__14613_ gnd vdd FILL
X_6840_ _6840_/A gnd memoryAddress[2] vdd BUFX2
XFILL_5__13434_ gnd vdd FILL
XFILL_0__7192_ gnd vdd FILL
XFILL_5__10646_ gnd vdd FILL
XFILL_2__16042_ gnd vdd FILL
XFILL_4__12075_ gnd vdd FILL
XSFILL43880x42050 gnd vdd FILL
XFILL_3__11825_ gnd vdd FILL
X_14889_ _9332_/Q _13854_/B _13853_/B _8820_/Q gnd _14889_/Y vdd AOI22X1
XSFILL8920x26050 gnd vdd FILL
XFILL_2__13254_ gnd vdd FILL
XFILL_3__15593_ gnd vdd FILL
XFILL_0__14433_ gnd vdd FILL
XFILL_0__11645_ gnd vdd FILL
XFILL_3__8990_ gnd vdd FILL
XFILL_1__13984_ gnd vdd FILL
XFILL_5__13365_ gnd vdd FILL
XFILL_4__15903_ gnd vdd FILL
XFILL_4__11026_ gnd vdd FILL
XFILL_5__16153_ gnd vdd FILL
XFILL_3__14544_ gnd vdd FILL
XFILL_2__12205_ gnd vdd FILL
XFILL_5__10577_ gnd vdd FILL
XFILL_1__15723_ gnd vdd FILL
XSFILL33640x5050 gnd vdd FILL
XFILL_3__7941_ gnd vdd FILL
XFILL_2__7059_ gnd vdd FILL
XFILL_3__11756_ gnd vdd FILL
XFILL_0__14364_ gnd vdd FILL
XFILL_2__10397_ gnd vdd FILL
X_8510_ _8558_/Q gnd _8512_/A vdd INVX1
XFILL_5__8857_ gnd vdd FILL
XFILL_5__12316_ gnd vdd FILL
XFILL_0__11576_ gnd vdd FILL
XSFILL74200x12050 gnd vdd FILL
XFILL_5__15104_ gnd vdd FILL
XFILL_5__16084_ gnd vdd FILL
XFILL_5__13296_ gnd vdd FILL
XFILL_4__15834_ gnd vdd FILL
XFILL_3__10707_ gnd vdd FILL
X_9490_ _9554_/B _8466_/B gnd _9490_/Y vdd NAND2X1
XFILL_0__13315_ gnd vdd FILL
XFILL_3__14475_ gnd vdd FILL
XFILL_2__12136_ gnd vdd FILL
XFILL_0__16103_ gnd vdd FILL
XFILL_3__7872_ gnd vdd FILL
XFILL_5__7808_ gnd vdd FILL
XFILL_1__15654_ gnd vdd FILL
XFILL_3__11687_ gnd vdd FILL
XFILL_0__10527_ gnd vdd FILL
XFILL_5_BUFX2_insert408 gnd vdd FILL
XFILL_1__12866_ gnd vdd FILL
XFILL_0__14295_ gnd vdd FILL
XFILL_0__9902_ gnd vdd FILL
XSFILL59000x73050 gnd vdd FILL
XFILL_3__16214_ gnd vdd FILL
XFILL_5__15035_ gnd vdd FILL
XFILL_5_BUFX2_insert419 gnd vdd FILL
XFILL_5__12247_ gnd vdd FILL
X_8441_ _8441_/A gnd _8443_/A vdd INVX1
XFILL_5__8788_ gnd vdd FILL
XFILL_3__9611_ gnd vdd FILL
XFILL_3__13426_ gnd vdd FILL
XSFILL108920x33050 gnd vdd FILL
XFILL_3__10638_ gnd vdd FILL
XFILL_1__14605_ gnd vdd FILL
XFILL_4__12977_ gnd vdd FILL
XFILL_0__16034_ gnd vdd FILL
XFILL_2__12067_ gnd vdd FILL
XFILL_4__15765_ gnd vdd FILL
XFILL_0__13246_ gnd vdd FILL
XFILL_1__11817_ gnd vdd FILL
XFILL_5__7739_ gnd vdd FILL
XFILL_1__15585_ gnd vdd FILL
XFILL_0_BUFX2_insert770 gnd vdd FILL
XFILL_5__12178_ gnd vdd FILL
XFILL_4__14716_ gnd vdd FILL
XFILL_4__11928_ gnd vdd FILL
XFILL_0_BUFX2_insert781 gnd vdd FILL
X_8372_ _8370_/Y _8372_/B _8372_/C gnd _8426_/D vdd OAI21X1
XFILL_2__11018_ gnd vdd FILL
XFILL_3__16145_ gnd vdd FILL
XFILL_3__13357_ gnd vdd FILL
XFILL_4__15696_ gnd vdd FILL
XFILL_0_BUFX2_insert792 gnd vdd FILL
XFILL_3__9542_ gnd vdd FILL
XFILL_1__14536_ gnd vdd FILL
XFILL_3__10569_ gnd vdd FILL
XFILL_1__11748_ gnd vdd FILL
X_7323_ _7323_/A _7451_/B gnd _7323_/Y vdd NAND2X1
XFILL_0__10389_ gnd vdd FILL
XFILL_5__11129_ gnd vdd FILL
XFILL_0__9764_ gnd vdd FILL
XSFILL64120x64050 gnd vdd FILL
XFILL_3__12308_ gnd vdd FILL
XFILL_0__6976_ gnd vdd FILL
XFILL_4__14647_ gnd vdd FILL
XFILL_2__15826_ gnd vdd FILL
XFILL_4__11859_ gnd vdd FILL
XFILL_3__16076_ gnd vdd FILL
XFILL_3__9473_ gnd vdd FILL
XFILL_3__13288_ gnd vdd FILL
XFILL_0__12128_ gnd vdd FILL
XFILL_5__9409_ gnd vdd FILL
XFILL_1__14467_ gnd vdd FILL
XFILL_1__11679_ gnd vdd FILL
XFILL_0__8715_ gnd vdd FILL
XFILL_3__15027_ gnd vdd FILL
X_7254_ _7158_/A _6998_/CLK _7644_/R vdd _7254_/D gnd vdd DFFSR
XFILL_5__15937_ gnd vdd FILL
XFILL_4__14578_ gnd vdd FILL
XFILL_1__16206_ gnd vdd FILL
XFILL_3__12239_ gnd vdd FILL
XFILL_1__13418_ gnd vdd FILL
XFILL_2__15757_ gnd vdd FILL
XFILL_0__12059_ gnd vdd FILL
XFILL_2__12969_ gnd vdd FILL
XFILL_6__8133_ gnd vdd FILL
XFILL_1__14398_ gnd vdd FILL
XSFILL43960x22050 gnd vdd FILL
XSFILL3560x71050 gnd vdd FILL
XFILL_0__8646_ gnd vdd FILL
XFILL_4__16317_ gnd vdd FILL
XFILL_4__13529_ gnd vdd FILL
XFILL_2__14708_ gnd vdd FILL
XFILL_5__15868_ gnd vdd FILL
X_7185_ _7185_/A gnd _7187_/A vdd INVX1
XFILL_3__8355_ gnd vdd FILL
XSFILL18600x39050 gnd vdd FILL
XSFILL59080x50 gnd vdd FILL
XFILL_1__16137_ gnd vdd FILL
XFILL_1__13349_ gnd vdd FILL
XFILL_2__15688_ gnd vdd FILL
XFILL_5__14819_ gnd vdd FILL
XFILL_0__8577_ gnd vdd FILL
XFILL_1__7370_ gnd vdd FILL
XFILL_3__7306_ gnd vdd FILL
XFILL_4__16248_ gnd vdd FILL
XFILL_2__14639_ gnd vdd FILL
XFILL_5__15799_ gnd vdd FILL
XFILL_0__15818_ gnd vdd FILL
XFILL_1__16068_ gnd vdd FILL
XFILL_1_BUFX2_insert4 gnd vdd FILL
XFILL_2_BUFX2_insert309 gnd vdd FILL
XFILL_4__16179_ gnd vdd FILL
XFILL_3__15929_ gnd vdd FILL
XFILL_3__7237_ gnd vdd FILL
XFILL_1__15019_ gnd vdd FILL
XFILL_0__15749_ gnd vdd FILL
XFILL_1__9040_ gnd vdd FILL
XSFILL33880x74050 gnd vdd FILL
XFILL_0__7459_ gnd vdd FILL
XFILL_2__16309_ gnd vdd FILL
XFILL_3__7168_ gnd vdd FILL
XSFILL23320x32050 gnd vdd FILL
XFILL_6__8966_ gnd vdd FILL
X_9826_ _9826_/Q _8022_/CLK _8674_/R vdd _9826_/D gnd vdd DFFSR
XSFILL38920x11050 gnd vdd FILL
XFILL_3__7099_ gnd vdd FILL
XSFILL64200x44050 gnd vdd FILL
XFILL_4__7981_ gnd vdd FILL
XFILL_0__9129_ gnd vdd FILL
XFILL_4__9720_ gnd vdd FILL
X_9757_ _9757_/A gnd _9757_/Y vdd INVX1
X_6969_ _6937_/B _9657_/B gnd _6969_/Y vdd NAND2X1
XFILL_4__6932_ gnd vdd FILL
XBUFX2_insert308 _11983_/Y gnd _11999_/C vdd BUFX2
X_8708_ _8706_/Y _8765_/B _8708_/C gnd _8794_/D vdd OAI21X1
XBUFX2_insert319 _15000_/Y gnd _16301_/A vdd BUFX2
XFILL_6_BUFX2_insert275 gnd vdd FILL
X_9688_ _9596_/A _8151_/CLK _9048_/R vdd _9598_/Y gnd vdd DFFSR
XFILL_4__9651_ gnd vdd FILL
XSFILL3640x51050 gnd vdd FILL
XFILL_4__6863_ gnd vdd FILL
X_10570_ _16187_/A gnd _10572_/A vdd INVX1
X_8639_ _8577_/B _7231_/B gnd _8640_/C vdd NAND2X1
XFILL_4__8602_ gnd vdd FILL
XFILL_5_BUFX2_insert920 gnd vdd FILL
XFILL_1__9873_ gnd vdd FILL
XFILL_3__9809_ gnd vdd FILL
XSFILL28840x63050 gnd vdd FILL
XFILL_5_CLKBUF1_insert209 gnd vdd FILL
XFILL_5_BUFX2_insert931 gnd vdd FILL
XFILL_5_BUFX2_insert942 gnd vdd FILL
XSFILL115160x5050 gnd vdd FILL
XFILL_1__8824_ gnd vdd FILL
XFILL_5_BUFX2_insert953 gnd vdd FILL
XFILL_5_BUFX2_insert964 gnd vdd FILL
XFILL_5_BUFX2_insert975 gnd vdd FILL
XFILL_4__8533_ gnd vdd FILL
XSFILL104600x6050 gnd vdd FILL
XFILL_5_BUFX2_insert986 gnd vdd FILL
X_12240_ _12272_/A _12713_/A _12272_/C gnd _12242_/B vdd NAND3X1
XFILL_5_BUFX2_insert997 gnd vdd FILL
XFILL_1__8755_ gnd vdd FILL
XFILL_4__8464_ gnd vdd FILL
XSFILL33960x54050 gnd vdd FILL
X_12171_ _12171_/A _12117_/B _12171_/C gnd _12171_/Y vdd OAI21X1
XFILL_1__7706_ gnd vdd FILL
XFILL_4__7415_ gnd vdd FILL
XFILL_4__8395_ gnd vdd FILL
X_11122_ _11121_/Y gnd _11130_/B vdd INVX2
XSFILL89640x26050 gnd vdd FILL
XFILL_1__7637_ gnd vdd FILL
XFILL_3_BUFX2_insert110 gnd vdd FILL
XFILL_4__7346_ gnd vdd FILL
X_15930_ _15369_/D _14540_/Y _15972_/C _14520_/Y gnd _15930_/Y vdd OAI22X1
X_11053_ _12258_/Y _12147_/Y gnd _11720_/A vdd XOR2X1
XFILL_1__7568_ gnd vdd FILL
X_10004_ _15475_/A gnd _10006_/A vdd INVX1
XFILL_2__8100_ gnd vdd FILL
X_15861_ _14407_/A _15940_/B _16099_/C _14433_/A gnd _15861_/Y vdd OAI22X1
XFILL_2__9080_ gnd vdd FILL
XFILL_4__9016_ gnd vdd FILL
XSFILL3720x31050 gnd vdd FILL
XFILL_2_BUFX2_insert810 gnd vdd FILL
XFILL_1__7499_ gnd vdd FILL
XFILL_2_BUFX2_insert821 gnd vdd FILL
X_14812_ _14812_/A _14812_/B gnd _14834_/A vdd NOR2X1
XSFILL94360x4050 gnd vdd FILL
XFILL_2_BUFX2_insert832 gnd vdd FILL
X_15792_ _15791_/Y _15792_/B _15633_/D _14348_/D gnd _15793_/B vdd OAI22X1
XFILL_2_BUFX2_insert843 gnd vdd FILL
XFILL_1__9238_ gnd vdd FILL
XFILL_4__10190_ gnd vdd FILL
XFILL_2_BUFX2_insert854 gnd vdd FILL
XFILL_2_BUFX2_insert865 gnd vdd FILL
XFILL_5__10500_ gnd vdd FILL
XFILL_2_BUFX2_insert876 gnd vdd FILL
X_14743_ _7495_/A gnd _14743_/Y vdd INVX1
XFILL_2_BUFX2_insert887 gnd vdd FILL
X_11955_ _11955_/A _11955_/B _11954_/Y gnd _6860_/A vdd OAI21X1
XFILL_2__10320_ gnd vdd FILL
XFILL_5__11480_ gnd vdd FILL
XFILL_2_BUFX2_insert898 gnd vdd FILL
XFILL_1__9169_ gnd vdd FILL
XSFILL79160x80050 gnd vdd FILL
XFILL_5__9760_ gnd vdd FILL
XFILL_5__6972_ gnd vdd FILL
X_10906_ _10906_/A _10910_/B gnd _10906_/Y vdd NAND2X1
XFILL_5__10431_ gnd vdd FILL
X_14674_ _9583_/Q gnd _14675_/D vdd INVX1
XFILL_3__11610_ gnd vdd FILL
XFILL_2__10251_ gnd vdd FILL
X_11886_ _11884_/Y _11874_/B _11885_/Y gnd _13289_/B vdd OAI21X1
XFILL_3__12590_ gnd vdd FILL
XFILL_5__8711_ gnd vdd FILL
XFILL_0__11430_ gnd vdd FILL
XFILL_2__9982_ gnd vdd FILL
XFILL_1__10981_ gnd vdd FILL
XFILL_4__9918_ gnd vdd FILL
X_16413_ _16413_/A gnd _16412_/Y gnd _16413_/Y vdd OAI21X1
X_13625_ _9817_/Q _14213_/A _13625_/C gnd _13635_/A vdd AOI21X1
XFILL_5__13150_ gnd vdd FILL
XSFILL99480x29050 gnd vdd FILL
XFILL_4_BUFX2_insert8 gnd vdd FILL
XFILL_5__10362_ gnd vdd FILL
XFILL_4__12900_ gnd vdd FILL
X_10837_ _10837_/A _10797_/A _10837_/C gnd _10869_/D vdd OAI21X1
XFILL_4__13880_ gnd vdd FILL
XSFILL74120x27050 gnd vdd FILL
XFILL_3__11541_ gnd vdd FILL
XFILL_1__12720_ gnd vdd FILL
XFILL_2__10182_ gnd vdd FILL
XFILL_5__12101_ gnd vdd FILL
XFILL_5__8642_ gnd vdd FILL
XBUFX2_insert820 _12384_/Y gnd _7326_/B vdd BUFX2
XFILL_0__11361_ gnd vdd FILL
X_16344_ _16344_/A gnd _16343_/Y gnd _16424_/D vdd OAI21X1
XBUFX2_insert831 _15046_/Y gnd _15384_/A vdd BUFX2
XFILL_4__9849_ gnd vdd FILL
XFILL_5__13081_ gnd vdd FILL
XBUFX2_insert842 _13324_/Y gnd _8609_/A vdd BUFX2
X_13556_ _9340_/A gnd _13557_/D vdd INVX1
XFILL_4__12831_ gnd vdd FILL
X_10768_ _10766_/Y _10789_/B _10768_/C gnd _10846_/D vdd OAI21X1
XFILL_5__10293_ gnd vdd FILL
XBUFX2_insert853 _13269_/Y gnd _7100_/A vdd BUFX2
XFILL_3__14260_ gnd vdd FILL
XFILL_0__13100_ gnd vdd FILL
XFILL_1__12651_ gnd vdd FILL
XFILL_2__8864_ gnd vdd FILL
XFILL_0__10312_ gnd vdd FILL
XFILL_3__11472_ gnd vdd FILL
XFILL_2__14990_ gnd vdd FILL
XBUFX2_insert864 _13438_/Y gnd _13592_/A vdd BUFX2
XFILL_0__14080_ gnd vdd FILL
X_12507_ _12505_/Y vdd _12506_/Y gnd _12557_/D vdd OAI21X1
XFILL_5__12032_ gnd vdd FILL
XBUFX2_insert875 _13435_/Y gnd _14700_/A vdd BUFX2
XFILL_0__11292_ gnd vdd FILL
XFILL_5__8573_ gnd vdd FILL
XFILL_3__13211_ gnd vdd FILL
XBUFX2_insert886 _13432_/Y gnd _14466_/C vdd BUFX2
XFILL_4__15550_ gnd vdd FILL
X_16275_ _8272_/A gnd _16276_/D vdd INVX1
XFILL_3__10423_ gnd vdd FILL
XFILL_4__12762_ gnd vdd FILL
XBUFX2_insert897 _13470_/Y gnd _13836_/B vdd BUFX2
X_13487_ _14200_/C gnd _13487_/Y vdd INVX8
XFILL_2__7815_ gnd vdd FILL
XFILL_3__14191_ gnd vdd FILL
X_10699_ _10700_/B _7883_/B gnd _10699_/Y vdd NAND2X1
XFILL_0__13031_ gnd vdd FILL
XFILL_1__11602_ gnd vdd FILL
XFILL_2__13941_ gnd vdd FILL
XFILL_1__15370_ gnd vdd FILL
XFILL_1__12582_ gnd vdd FILL
XFILL_0__10243_ gnd vdd FILL
X_15226_ _15351_/A _15226_/B _13643_/D _15351_/D gnd _15226_/Y vdd OAI22X1
XSFILL8760x5050 gnd vdd FILL
XFILL_4__14501_ gnd vdd FILL
X_12438_ _12436_/Y _12359_/A _12438_/C gnd _12438_/Y vdd OAI21X1
XFILL_4__11713_ gnd vdd FILL
XFILL_3__13142_ gnd vdd FILL
XSFILL38760x46050 gnd vdd FILL
XFILL_4__15481_ gnd vdd FILL
XFILL112280x53050 gnd vdd FILL
XFILL_1__14321_ gnd vdd FILL
XFILL_2__7746_ gnd vdd FILL
XFILL_1__11533_ gnd vdd FILL
XSFILL64040x79050 gnd vdd FILL
XFILL_2__13872_ gnd vdd FILL
XFILL_0__10174_ gnd vdd FILL
XSFILL113960x39050 gnd vdd FILL
XFILL_5__7455_ gnd vdd FILL
X_15157_ _15802_/A _15157_/B _15157_/C _15802_/D gnd _15157_/Y vdd OAI22X1
XFILL_4__14432_ gnd vdd FILL
X_12369_ _12367_/Y _12368_/A _12369_/C gnd _12369_/Y vdd OAI21X1
XFILL_2__15611_ gnd vdd FILL
XFILL_4__11644_ gnd vdd FILL
XFILL_5__13983_ gnd vdd FILL
XFILL_2__12823_ gnd vdd FILL
XFILL_1__14252_ gnd vdd FILL
XFILL_3__10285_ gnd vdd FILL
XFILL_2__7677_ gnd vdd FILL
XFILL_1__11464_ gnd vdd FILL
X_14108_ _15599_/D _14949_/C gnd _14109_/C vdd NOR2X1
XFILL_0__8500_ gnd vdd FILL
XFILL_5__15722_ gnd vdd FILL
XFILL_0__14982_ gnd vdd FILL
X_15088_ _16228_/B gnd _15175_/B vdd INVX8
XFILL_0__9480_ gnd vdd FILL
XFILL_3__12024_ gnd vdd FILL
XFILL_2__9416_ gnd vdd FILL
XFILL_4__14363_ gnd vdd FILL
XFILL_2__15542_ gnd vdd FILL
XFILL_1__10415_ gnd vdd FILL
XFILL_4__11575_ gnd vdd FILL
XFILL_5__9125_ gnd vdd FILL
XFILL_2__12754_ gnd vdd FILL
XFILL_1__14183_ gnd vdd FILL
XFILL_1__11395_ gnd vdd FILL
XFILL_0__13933_ gnd vdd FILL
XFILL_4__13314_ gnd vdd FILL
X_14039_ _7138_/Q gnd _14039_/Y vdd INVX1
XFILL_4__16102_ gnd vdd FILL
XFILL_5__15653_ gnd vdd FILL
XFILL_4__10526_ gnd vdd FILL
XFILL_2__9347_ gnd vdd FILL
XFILL_1__13134_ gnd vdd FILL
XFILL_5__12865_ gnd vdd FILL
XFILL_3__8140_ gnd vdd FILL
XFILL_4__14294_ gnd vdd FILL
XFILL_2__11705_ gnd vdd FILL
XSFILL18680x13050 gnd vdd FILL
XFILL_2__15473_ gnd vdd FILL
XFILL_0__13864_ gnd vdd FILL
XFILL_5__14604_ gnd vdd FILL
XFILL_4__16033_ gnd vdd FILL
XFILL_4__13245_ gnd vdd FILL
XFILL_0__8362_ gnd vdd FILL
XFILL_5__11816_ gnd vdd FILL
XFILL_5__15584_ gnd vdd FILL
XFILL_2__14424_ gnd vdd FILL
XFILL_2__9278_ gnd vdd FILL
XSFILL84360x51050 gnd vdd FILL
XFILL_2__11636_ gnd vdd FILL
X_8990_ _9044_/A _7838_/B gnd _8990_/Y vdd NAND2X1
XFILL_3__8071_ gnd vdd FILL
XFILL_0__15603_ gnd vdd FILL
XFILL_3__13975_ gnd vdd FILL
XFILL_5__8007_ gnd vdd FILL
XFILL_1__10277_ gnd vdd FILL
XFILL_0__13795_ gnd vdd FILL
XSFILL58520x61050 gnd vdd FILL
XFILL_0__7313_ gnd vdd FILL
XSFILL59000x68050 gnd vdd FILL
XFILL_5__14535_ gnd vdd FILL
XFILL_2__8229_ gnd vdd FILL
XFILL_3__15714_ gnd vdd FILL
XFILL_1__12016_ gnd vdd FILL
X_7941_ _7941_/A gnd _7941_/Y vdd INVX1
XFILL_5__11747_ gnd vdd FILL
XFILL_2__14355_ gnd vdd FILL
XFILL_4__10388_ gnd vdd FILL
XFILL_0__12746_ gnd vdd FILL
XSFILL99400x73050 gnd vdd FILL
XFILL_0__15534_ gnd vdd FILL
XFILL_2__11567_ gnd vdd FILL
XFILL_0__7244_ gnd vdd FILL
XFILL_4__12127_ gnd vdd FILL
XFILL_2__13306_ gnd vdd FILL
X_7872_ _7872_/A _7872_/B _7871_/Y gnd _7872_/Y vdd OAI21X1
XFILL_5__14466_ gnd vdd FILL
XFILL_3__15645_ gnd vdd FILL
XFILL_5__11678_ gnd vdd FILL
XFILL_3__12857_ gnd vdd FILL
XFILL_2__10518_ gnd vdd FILL
XFILL_2__14286_ gnd vdd FILL
XFILL_5__16205_ gnd vdd FILL
XFILL_2__11498_ gnd vdd FILL
XFILL_0__15465_ gnd vdd FILL
XSFILL38840x26050 gnd vdd FILL
X_9611_ _9611_/A gnd _9613_/A vdd INVX1
XFILL_5__13417_ gnd vdd FILL
XFILL112360x33050 gnd vdd FILL
XFILL_5__10629_ gnd vdd FILL
XFILL_0__7175_ gnd vdd FILL
XFILL_6__15756_ gnd vdd FILL
XFILL_2__16025_ gnd vdd FILL
XFILL_4__12058_ gnd vdd FILL
XFILL_3__11808_ gnd vdd FILL
XFILL_2__13237_ gnd vdd FILL
XFILL_5__14397_ gnd vdd FILL
XFILL_3__15576_ gnd vdd FILL
XFILL_3__12788_ gnd vdd FILL
XSFILL49480x77050 gnd vdd FILL
XFILL_3__8973_ gnd vdd FILL
XFILL_2__10449_ gnd vdd FILL
XFILL_0__11628_ gnd vdd FILL
XFILL_0__14416_ gnd vdd FILL
XFILL_5__8909_ gnd vdd FILL
XFILL_0__15396_ gnd vdd FILL
XFILL_6__14707_ gnd vdd FILL
XFILL_1__13967_ gnd vdd FILL
XFILL_5__16136_ gnd vdd FILL
XFILL_4__11009_ gnd vdd FILL
XFILL_5__13348_ gnd vdd FILL
XFILL_5__9889_ gnd vdd FILL
XFILL_3__14527_ gnd vdd FILL
X_9542_ _9540_/Y _9529_/A _9542_/C gnd _9584_/D vdd OAI21X1
XFILL_1__15706_ gnd vdd FILL
XSFILL114600x1050 gnd vdd FILL
XFILL_3__11739_ gnd vdd FILL
XFILL_2__13168_ gnd vdd FILL
XFILL_0__14347_ gnd vdd FILL
XFILL_1__12918_ gnd vdd FILL
XFILL_0__11559_ gnd vdd FILL
XSFILL79320x40050 gnd vdd FILL
XFILL_1__13898_ gnd vdd FILL
XSFILL43960x17050 gnd vdd FILL
XFILL_5__13279_ gnd vdd FILL
XFILL_4__15817_ gnd vdd FILL
XFILL_5__16067_ gnd vdd FILL
X_9473_ _9471_/Y _9548_/B _9472_/Y gnd _9561_/D vdd OAI21X1
XFILL_3__14458_ gnd vdd FILL
XFILL_2__12119_ gnd vdd FILL
XFILL_5_BUFX2_insert227 gnd vdd FILL
XFILL_1__15637_ gnd vdd FILL
XFILL_3__7855_ gnd vdd FILL
XFILL_1__12849_ gnd vdd FILL
XFILL_2__13099_ gnd vdd FILL
XFILL_0__14278_ gnd vdd FILL
XFILL_5_BUFX2_insert238 gnd vdd FILL
XFILL_5__15018_ gnd vdd FILL
XFILL_5_BUFX2_insert249 gnd vdd FILL
XSFILL28760x78050 gnd vdd FILL
XFILL_6__14569_ gnd vdd FILL
XFILL_3__13409_ gnd vdd FILL
X_8424_ _8424_/Q _7016_/CLK _8424_/R vdd _8366_/Y gnd vdd DFFSR
XFILL_1__6870_ gnd vdd FILL
XFILL_4__15748_ gnd vdd FILL
XFILL_0__13229_ gnd vdd FILL
XFILL_0__16017_ gnd vdd FILL
XFILL_3__14389_ gnd vdd FILL
XFILL_1__15568_ gnd vdd FILL
XFILL_4_BUFX2_insert905 gnd vdd FILL
X_8355_ _8421_/Q gnd _8355_/Y vdd INVX1
XFILL_3__16128_ gnd vdd FILL
XFILL_3__9525_ gnd vdd FILL
XFILL_4_BUFX2_insert916 gnd vdd FILL
XFILL_4__15679_ gnd vdd FILL
XFILL_1__14519_ gnd vdd FILL
XFILL_4_BUFX2_insert927 gnd vdd FILL
X_7306_ _7304_/Y _7359_/A _7305_/Y gnd _7388_/D vdd OAI21X1
XFILL_1__15499_ gnd vdd FILL
XFILL_4_BUFX2_insert938 gnd vdd FILL
XFILL_4_BUFX2_insert949 gnd vdd FILL
XFILL_0__9747_ gnd vdd FILL
X_8286_ _8206_/A _8025_/CLK _8025_/R vdd _8286_/D gnd vdd DFFSR
XSFILL33880x69050 gnd vdd FILL
XFILL_0__6959_ gnd vdd FILL
XFILL_2__15809_ gnd vdd FILL
XFILL_3__16059_ gnd vdd FILL
X_7237_ _7181_/B _9413_/B gnd _7237_/Y vdd NAND2X1
XFILL_0__9678_ gnd vdd FILL
XFILL_1__8471_ gnd vdd FILL
XFILL_4__7200_ gnd vdd FILL
XFILL_3__9387_ gnd vdd FILL
XFILL112440x13050 gnd vdd FILL
XSFILL64200x39050 gnd vdd FILL
XFILL_0__8629_ gnd vdd FILL
XFILL_1__7422_ gnd vdd FILL
X_7168_ _7168_/A _9600_/B gnd _7169_/C vdd NAND2X1
XSFILL38920x7050 gnd vdd FILL
XFILL_3__8338_ gnd vdd FILL
XSFILL89160x43050 gnd vdd FILL
XFILL_1__7353_ gnd vdd FILL
X_7099_ _7149_/Q gnd _7099_/Y vdd INVX1
XFILL_2_BUFX2_insert106 gnd vdd FILL
XFILL_3__8269_ gnd vdd FILL
XFILL_4__7062_ gnd vdd FILL
XSFILL79400x20050 gnd vdd FILL
XSFILL3640x46050 gnd vdd FILL
XSFILL13240x79050 gnd vdd FILL
XFILL_1__9023_ gnd vdd FILL
XSFILL68440x44050 gnd vdd FILL
XFILL_1_BUFX2_insert806 gnd vdd FILL
XFILL_1_BUFX2_insert817 gnd vdd FILL
XFILL_1_BUFX2_insert828 gnd vdd FILL
X_11740_ _11739_/Y _11740_/B _11735_/Y gnd _11741_/C vdd AOI21X1
XFILL_1_BUFX2_insert839 gnd vdd FILL
XSFILL69080x10050 gnd vdd FILL
X_9809_ _9785_/A _8529_/B gnd _9809_/Y vdd NAND2X1
XSFILL104680x17050 gnd vdd FILL
XFILL_4__7964_ gnd vdd FILL
XSFILL33960x49050 gnd vdd FILL
X_11671_ _11656_/B _11649_/Y gnd _11671_/Y vdd AND2X2
XBUFX2_insert105 _10925_/Y gnd _11909_/A vdd BUFX2
XFILL_4__6915_ gnd vdd FILL
X_13410_ _13410_/A gnd _13410_/Y vdd INVX1
X_10622_ _10622_/A _10619_/B _10621_/Y gnd _10622_/Y vdd OAI21X1
XSFILL64120x2050 gnd vdd FILL
XFILL_1__9925_ gnd vdd FILL
X_14390_ _14390_/A _14390_/B _14387_/Y gnd _14390_/Y vdd NAND3X1
XSFILL104520x81050 gnd vdd FILL
XFILL_4__9634_ gnd vdd FILL
XFILL_4__6846_ gnd vdd FILL
X_13341_ _13236_/B _13310_/A _13337_/B gnd _13341_/Y vdd OAI21X1
X_10553_ _10557_/B _8889_/B gnd _10554_/C vdd NAND2X1
XFILL_1__9856_ gnd vdd FILL
XFILL_5_BUFX2_insert750 gnd vdd FILL
XFILL_5_BUFX2_insert761 gnd vdd FILL
XFILL_5_BUFX2_insert772 gnd vdd FILL
X_16060_ _7023_/Q _15382_/B _16096_/C _7361_/A gnd _16066_/A vdd AOI22X1
X_13272_ _13337_/A _13283_/A gnd _13273_/A vdd NOR2X1
XFILL_5_BUFX2_insert783 gnd vdd FILL
XFILL_2__7600_ gnd vdd FILL
XFILL_5_BUFX2_insert794 gnd vdd FILL
X_10484_ _14918_/A _8815_/CLK _8047_/R vdd _10484_/D gnd vdd DFFSR
XFILL_1__9787_ gnd vdd FILL
XFILL_2__8580_ gnd vdd FILL
XFILL_4__8516_ gnd vdd FILL
X_15011_ _7766_/Q _15969_/C gnd _15011_/Y vdd NAND2X1
XSFILL64600x8050 gnd vdd FILL
XFILL_4__9496_ gnd vdd FILL
X_12223_ _12227_/A vdd _12307_/C gnd _12226_/A vdd NAND3X1
XFILL_1__8738_ gnd vdd FILL
XFILL_4__8447_ gnd vdd FILL
XSFILL94360x14050 gnd vdd FILL
XFILL_5__7240_ gnd vdd FILL
X_12154_ _13188_/Q gnd _12156_/A vdd INVX1
XFILL_5__10980_ gnd vdd FILL
XFILL_2__7462_ gnd vdd FILL
XSFILL79160x75050 gnd vdd FILL
XFILL_4__8378_ gnd vdd FILL
XFILL_5__7171_ gnd vdd FILL
X_11105_ _12186_/Y _12310_/Y gnd _11105_/Y vdd NOR2X1
XFILL_6__10181_ gnd vdd FILL
X_12085_ _12512_/B _12105_/B _12001_/C gnd gnd _12085_/Y vdd AOI22X1
XFILL_4__11360_ gnd vdd FILL
XFILL_0__10930_ gnd vdd FILL
XFILL_4__7329_ gnd vdd FILL
XFILL_1__11180_ gnd vdd FILL
XSFILL109400x2050 gnd vdd FILL
X_15913_ _10475_/Q _15175_/B _15912_/Y gnd _15917_/C vdd AOI21X1
XFILL_4__10311_ gnd vdd FILL
X_11036_ _12135_/Y gnd _11037_/B vdd INVX1
XFILL_5__12650_ gnd vdd FILL
XSFILL8440x38050 gnd vdd FILL
XFILL_2__9132_ gnd vdd FILL
XFILL_4__11291_ gnd vdd FILL
XFILL_1__10131_ gnd vdd FILL
XFILL_2__12470_ gnd vdd FILL
XSFILL84280x66050 gnd vdd FILL
XFILL_4__13030_ gnd vdd FILL
X_15844_ _9961_/Q gnd _15845_/D vdd INVX1
XFILL_5__11601_ gnd vdd FILL
XFILL_6__13940_ gnd vdd FILL
XFILL_5__12581_ gnd vdd FILL
XFILL_4__10242_ gnd vdd FILL
XFILL_0__12600_ gnd vdd FILL
XFILL_3__13760_ gnd vdd FILL
XFILL_2_BUFX2_insert640 gnd vdd FILL
XFILL_2__11421_ gnd vdd FILL
XFILL_1__10062_ gnd vdd FILL
XFILL_3__10972_ gnd vdd FILL
XFILL_2_BUFX2_insert651 gnd vdd FILL
XFILL_0__13580_ gnd vdd FILL
XFILL_0__10792_ gnd vdd FILL
XFILL_5__14320_ gnd vdd FILL
XFILL_5__11532_ gnd vdd FILL
XFILL_2_BUFX2_insert662 gnd vdd FILL
XFILL_2__8014_ gnd vdd FILL
XFILL_3__12711_ gnd vdd FILL
XSFILL59080x42050 gnd vdd FILL
XFILL_2_BUFX2_insert673 gnd vdd FILL
X_15775_ _14316_/Y _15565_/B _15563_/C _14336_/A gnd _15776_/B vdd OAI22X1
XFILL_4__10173_ gnd vdd FILL
XFILL_2_BUFX2_insert684 gnd vdd FILL
XFILL_2__14140_ gnd vdd FILL
X_12987_ _6882_/A gnd _12987_/Y vdd INVX1
XFILL_0__12531_ gnd vdd FILL
XFILL_2__11352_ gnd vdd FILL
XFILL_3__13691_ gnd vdd FILL
XFILL_2_BUFX2_insert695 gnd vdd FILL
XFILL_1__14870_ gnd vdd FILL
XFILL_5__9812_ gnd vdd FILL
X_14726_ _6980_/A gnd _14726_/Y vdd INVX1
XFILL_5__14251_ gnd vdd FILL
X_11938_ _13192_/Q gnd _11940_/A vdd INVX1
XFILL_3__15430_ gnd vdd FILL
XFILL_5__11463_ gnd vdd FILL
XFILL_2__10303_ gnd vdd FILL
XFILL_3__12642_ gnd vdd FILL
XFILL_1__13821_ gnd vdd FILL
XFILL_0__15250_ gnd vdd FILL
XFILL112280x48050 gnd vdd FILL
XFILL_4__14981_ gnd vdd FILL
XFILL_2__14071_ gnd vdd FILL
XFILL_2__11283_ gnd vdd FILL
XFILL_0__12462_ gnd vdd FILL
XFILL_5__9743_ gnd vdd FILL
XFILL_5_BUFX2_insert11 gnd vdd FILL
XFILL_6__15541_ gnd vdd FILL
XFILL_5__10414_ gnd vdd FILL
XFILL_5__6955_ gnd vdd FILL
XFILL_5__14182_ gnd vdd FILL
XFILL_6__12753_ gnd vdd FILL
X_14657_ _14655_/Y _14657_/B _14654_/Y gnd _14668_/A vdd NAND3X1
XFILL_5_BUFX2_insert22 gnd vdd FILL
XFILL_0__14201_ gnd vdd FILL
XFILL_2__13022_ gnd vdd FILL
XFILL_3__15361_ gnd vdd FILL
X_11869_ _12521_/B _12081_/A gnd _11869_/Y vdd NOR2X1
XFILL_2__10234_ gnd vdd FILL
XFILL_5__11394_ gnd vdd FILL
XFILL_4__13932_ gnd vdd FILL
XFILL_5_BUFX2_insert33 gnd vdd FILL
XFILL_3__12573_ gnd vdd FILL
XFILL_5_BUFX2_insert44 gnd vdd FILL
XFILL_0__11413_ gnd vdd FILL
XFILL_0__15181_ gnd vdd FILL
XFILL_1__13752_ gnd vdd FILL
XFILL_1__10964_ gnd vdd FILL
X_13608_ _13607_/Y _14203_/C gnd _13609_/C vdd NOR2X1
XFILL_5_BUFX2_insert55 gnd vdd FILL
XFILL_0__12393_ gnd vdd FILL
XFILL_5__9674_ gnd vdd FILL
XFILL_5__13133_ gnd vdd FILL
XSFILL13800x60050 gnd vdd FILL
XFILL_5__6886_ gnd vdd FILL
XFILL_5_BUFX2_insert66 gnd vdd FILL
XFILL_3__14312_ gnd vdd FILL
X_14588_ _8507_/A gnd _14588_/Y vdd INVX1
XFILL_5_BUFX2_insert77 gnd vdd FILL
XFILL_3__11524_ gnd vdd FILL
XFILL_0__8980_ gnd vdd FILL
XFILL_2__8916_ gnd vdd FILL
XFILL_2__10165_ gnd vdd FILL
XFILL_1__12703_ gnd vdd FILL
XFILL_4__13863_ gnd vdd FILL
XFILL_0__14132_ gnd vdd FILL
XFILL_5_BUFX2_insert88 gnd vdd FILL
XFILL_3__15292_ gnd vdd FILL
XFILL_2__9896_ gnd vdd FILL
XBUFX2_insert650 _10915_/Y gnd _12028_/A vdd BUFX2
XFILL_5__8625_ gnd vdd FILL
XFILL_0__11344_ gnd vdd FILL
XFILL_1__13683_ gnd vdd FILL
XBUFX2_insert661 _11988_/Y gnd _12113_/C vdd BUFX2
XFILL_5_BUFX2_insert99 gnd vdd FILL
XFILL_1__10895_ gnd vdd FILL
X_16327_ _16419_/Q gnd _16329_/A vdd INVX1
XBUFX2_insert672 _15064_/Y gnd _15394_/B vdd BUFX2
XFILL_6__11635_ gnd vdd FILL
XFILL_4__15602_ gnd vdd FILL
X_13539_ _14887_/B _13537_/Y _13539_/C _14068_/C gnd _13539_/Y vdd OAI22X1
XFILL_0__7931_ gnd vdd FILL
XFILL_5__10276_ gnd vdd FILL
XFILL_3__14243_ gnd vdd FILL
XFILL_4__13794_ gnd vdd FILL
XFILL_2__8847_ gnd vdd FILL
XFILL_3__11455_ gnd vdd FILL
XFILL_1__15422_ gnd vdd FILL
XBUFX2_insert683 _15005_/Y gnd _16247_/C vdd BUFX2
XFILL_1__12634_ gnd vdd FILL
XBUFX2_insert694 _13362_/Y gnd _10557_/B vdd BUFX2
XFILL_0__14063_ gnd vdd FILL
XFILL_2__14973_ gnd vdd FILL
XSFILL114440x64050 gnd vdd FILL
XFILL_5__12015_ gnd vdd FILL
XFILL_0__11275_ gnd vdd FILL
XSFILL8520x18050 gnd vdd FILL
XFILL_6__14354_ gnd vdd FILL
X_16258_ _16252_/Y _16253_/Y _16258_/C gnd _16258_/Y vdd NAND3X1
XFILL_0__7862_ gnd vdd FILL
XFILL_3__10406_ gnd vdd FILL
XFILL_4__12745_ gnd vdd FILL
XFILL_4__15533_ gnd vdd FILL
XFILL_0__13014_ gnd vdd FILL
XFILL_3__14174_ gnd vdd FILL
XFILL_2__13924_ gnd vdd FILL
XFILL_1__15353_ gnd vdd FILL
XFILL_2__8778_ gnd vdd FILL
XFILL_5__7507_ gnd vdd FILL
XFILL_3__7571_ gnd vdd FILL
XFILL_3__11386_ gnd vdd FILL
XFILL_0__9601_ gnd vdd FILL
X_15209_ _15802_/A gnd _15652_/A vdd INVX4
XFILL_5__8487_ gnd vdd FILL
X_8140_ _8140_/A _8098_/B _8139_/Y gnd _8178_/D vdd OAI21X1
XSFILL48920x2050 gnd vdd FILL
XFILL_6__10517_ gnd vdd FILL
XFILL_3__13125_ gnd vdd FILL
X_16189_ _16186_/Y _16189_/B gnd _16190_/A vdd NOR2X1
XFILL_2__7729_ gnd vdd FILL
XFILL_1__14304_ gnd vdd FILL
XFILL_4__15464_ gnd vdd FILL
XFILL_6__11497_ gnd vdd FILL
XFILL_2__13855_ gnd vdd FILL
XFILL_1__11516_ gnd vdd FILL
XFILL_5__7438_ gnd vdd FILL
XSFILL99400x68050 gnd vdd FILL
XFILL_1__12496_ gnd vdd FILL
XFILL_0__10157_ gnd vdd FILL
XFILL_1__15284_ gnd vdd FILL
XSFILL59160x22050 gnd vdd FILL
XFILL_0__9532_ gnd vdd FILL
X_8071_ _8071_/A _8107_/B _8070_/Y gnd _8155_/D vdd OAI21X1
XFILL_4__11627_ gnd vdd FILL
XFILL_4__14415_ gnd vdd FILL
XFILL_4__15395_ gnd vdd FILL
XFILL_3__9241_ gnd vdd FILL
XFILL_5__13966_ gnd vdd FILL
XFILL_1__14235_ gnd vdd FILL
XFILL_3__10268_ gnd vdd FILL
XFILL_1__11447_ gnd vdd FILL
XFILL_2__13786_ gnd vdd FILL
X_7022_ _6974_/A _7902_/CLK _9561_/R vdd _7022_/D gnd vdd DFFSR
XFILL_5__15705_ gnd vdd FILL
XFILL_5__7369_ gnd vdd FILL
XFILL_0__14965_ gnd vdd FILL
XFILL111880x21050 gnd vdd FILL
XFILL_2__10998_ gnd vdd FILL
XFILL_0__9463_ gnd vdd FILL
XFILL_3__12007_ gnd vdd FILL
XFILL_4__14346_ gnd vdd FILL
XFILL_5__12917_ gnd vdd FILL
XFILL112360x28050 gnd vdd FILL
XFILL_2__15525_ gnd vdd FILL
XFILL_4__11558_ gnd vdd FILL
XFILL_2__12737_ gnd vdd FILL
XFILL_5__9108_ gnd vdd FILL
XFILL_5__13897_ gnd vdd FILL
XFILL_3__9172_ gnd vdd FILL
XFILL_1__14166_ gnd vdd FILL
XFILL_0__13916_ gnd vdd FILL
XFILL_1__11378_ gnd vdd FILL
XFILL_4__10509_ gnd vdd FILL
XFILL_5__15636_ gnd vdd FILL
XFILL_0__14896_ gnd vdd FILL
XFILL_3__8123_ gnd vdd FILL
XFILL_5__12848_ gnd vdd FILL
XFILL_0__9394_ gnd vdd FILL
XFILL_4__14277_ gnd vdd FILL
XFILL_1__13117_ gnd vdd FILL
XFILL_4__11489_ gnd vdd FILL
XFILL_2__15456_ gnd vdd FILL
XFILL_5__9039_ gnd vdd FILL
XFILL_1__14097_ gnd vdd FILL
XFILL_0__13847_ gnd vdd FILL
XFILL_6__9921_ gnd vdd FILL
XFILL_4__13228_ gnd vdd FILL
XFILL_4__16016_ gnd vdd FILL
XFILL_0__8345_ gnd vdd FILL
XFILL_5__15567_ gnd vdd FILL
XFILL_2__14407_ gnd vdd FILL
XFILL_5__12779_ gnd vdd FILL
X_8973_ _8971_/Y _9014_/A _8973_/C gnd _8973_/Y vdd OAI21X1
XFILL_3__13958_ gnd vdd FILL
XFILL_2__11619_ gnd vdd FILL
XFILL_3__8054_ gnd vdd FILL
XFILL_2__15387_ gnd vdd FILL
XFILL_2__12599_ gnd vdd FILL
XFILL_0__13778_ gnd vdd FILL
XFILL_5__14518_ gnd vdd FILL
XFILL_4__13159_ gnd vdd FILL
XFILL_3__12909_ gnd vdd FILL
XFILL_0__8276_ gnd vdd FILL
X_7924_ _7888_/A _7156_/CLK _7775_/R vdd _7924_/D gnd vdd DFFSR
XFILL_5__15498_ gnd vdd FILL
XFILL_2__14338_ gnd vdd FILL
XFILL_0__15517_ gnd vdd FILL
XFILL_3__13889_ gnd vdd FILL
XFILL_0__12729_ gnd vdd FILL
XFILL_0__7227_ gnd vdd FILL
XFILL_5__14449_ gnd vdd FILL
XFILL_3__15628_ gnd vdd FILL
X_7855_ _7913_/Q gnd _7857_/A vdd INVX1
XFILL_2__14269_ gnd vdd FILL
XFILL_0__15448_ gnd vdd FILL
XFILL_0_CLKBUF1_insert206 gnd vdd FILL
XFILL_1__14999_ gnd vdd FILL
XFILL_0_CLKBUF1_insert217 gnd vdd FILL
XFILL_2__16008_ gnd vdd FILL
XFILL_0__7158_ gnd vdd FILL
XSFILL18600x52050 gnd vdd FILL
XFILL_3__15559_ gnd vdd FILL
X_7786_ _7786_/Q _7786_/CLK _9964_/R vdd _7786_/D gnd vdd DFFSR
XFILL_3__8956_ gnd vdd FILL
XFILL_0__15379_ gnd vdd FILL
XFILL_5__16119_ gnd vdd FILL
X_9525_ _9579_/Q gnd _9525_/Y vdd INVX1
XFILL_1__7971_ gnd vdd FILL
XFILL_0__7089_ gnd vdd FILL
XFILL_4__7680_ gnd vdd FILL
XFILL_3__8887_ gnd vdd FILL
XFILL_6__7616_ gnd vdd FILL
XFILL_1__6922_ gnd vdd FILL
X_9456_ _9412_/A _7642_/CLK _8676_/R vdd _9456_/D gnd vdd DFFSR
XFILL_3__7838_ gnd vdd FILL
XSFILL105080x62050 gnd vdd FILL
XFILL112040x10050 gnd vdd FILL
X_8407_ _8407_/Q _9077_/CLK _8433_/R vdd _8315_/Y gnd vdd DFFSR
XFILL_1__9641_ gnd vdd FILL
XFILL_1__6853_ gnd vdd FILL
XFILL_4_BUFX2_insert702 gnd vdd FILL
X_9387_ _9387_/A _9372_/B _9387_/C gnd _9447_/D vdd OAI21X1
XFILL_4__9350_ gnd vdd FILL
XFILL_4_BUFX2_insert713 gnd vdd FILL
XFILL_4_BUFX2_insert724 gnd vdd FILL
XFILL_4_BUFX2_insert735 gnd vdd FILL
XFILL_3__9508_ gnd vdd FILL
XFILL_4_BUFX2_insert746 gnd vdd FILL
X_8338_ _8372_/B _9362_/B gnd _8339_/C vdd NAND2X1
XFILL_4_BUFX2_insert757 gnd vdd FILL
XFILL_4__9281_ gnd vdd FILL
XFILL_3_CLKBUF1_insert1078 gnd vdd FILL
XFILL_4_BUFX2_insert768 gnd vdd FILL
XFILL_1__8523_ gnd vdd FILL
XFILL_4_BUFX2_insert779 gnd vdd FILL
XSFILL94280x29050 gnd vdd FILL
XSFILL114600x24050 gnd vdd FILL
X_8269_ _8269_/A gnd _8271_/A vdd INVX1
XFILL_4__8232_ gnd vdd FILL
XFILL_1__8454_ gnd vdd FILL
XSFILL69320x67050 gnd vdd FILL
XFILL_4__7114_ gnd vdd FILL
XFILL_1__8385_ gnd vdd FILL
X_12910_ _12910_/A gnd _12910_/Y vdd INVX1
XFILL_4__8094_ gnd vdd FILL
XFILL_1__7336_ gnd vdd FILL
X_13890_ _15416_/A _14721_/A _13876_/C _15423_/D gnd _13894_/B vdd OAI22X1
XSFILL104520x76050 gnd vdd FILL
XFILL_4__7045_ gnd vdd FILL
X_12841_ _12841_/A gnd _12843_/A vdd INVX1
XSFILL8760x74050 gnd vdd FILL
XSFILL23800x23050 gnd vdd FILL
XSFILL89240x18050 gnd vdd FILL
XFILL_1_BUFX2_insert603 gnd vdd FILL
XSFILL59080x9050 gnd vdd FILL
XFILL_1_BUFX2_insert614 gnd vdd FILL
X_15560_ _15560_/A _15559_/Y gnd _15572_/C vdd NAND2X1
XFILL_1__9006_ gnd vdd FILL
X_12772_ _12770_/Y _12723_/A _12772_/C gnd _12816_/D vdd OAI21X1
XFILL_1_BUFX2_insert625 gnd vdd FILL
XFILL_1_BUFX2_insert636 gnd vdd FILL
XSFILL74040x60050 gnd vdd FILL
XFILL_1__7198_ gnd vdd FILL
X_14511_ _9144_/A _14868_/D _14878_/C _10552_/A gnd _14511_/Y vdd AOI22X1
XFILL_1_BUFX2_insert647 gnd vdd FILL
XFILL_4__8996_ gnd vdd FILL
XFILL_1_BUFX2_insert658 gnd vdd FILL
X_11723_ _11703_/C _11748_/A _11722_/Y gnd _11723_/Y vdd OAI21X1
XFILL_1_BUFX2_insert669 gnd vdd FILL
X_15491_ _8596_/A gnd _15491_/Y vdd INVX1
XFILL_4__7947_ gnd vdd FILL
X_14442_ _14442_/A gnd _15875_/D vdd INVX1
X_11654_ _11257_/Y _11654_/B _11654_/C gnd _11676_/B vdd OAI21X1
XFILL_2__9750_ gnd vdd FILL
XSFILL13720x75050 gnd vdd FILL
XFILL_2__6962_ gnd vdd FILL
X_10605_ _14584_/A _9453_/CLK _9453_/R vdd _10557_/Y gnd vdd DFFSR
XFILL_4__7878_ gnd vdd FILL
XFILL_5__10130_ gnd vdd FILL
X_14373_ _13868_/B _15842_/C _14711_/B _15829_/B gnd _14373_/Y vdd OAI22X1
XFILL_2__8701_ gnd vdd FILL
XFILL_1__9908_ gnd vdd FILL
X_11585_ _11582_/C gnd _11587_/C vdd INVX2
XFILL_2__9681_ gnd vdd FILL
XFILL_2__6893_ gnd vdd FILL
X_16112_ _14713_/A _15680_/B _15680_/C gnd _16112_/Y vdd NAND3X1
XFILL_1__10680_ gnd vdd FILL
XFILL_4__9617_ gnd vdd FILL
X_13324_ _13297_/C _13323_/Y gnd _13324_/Y vdd NOR2X1
XFILL_5__9390_ gnd vdd FILL
XFILL_6__11420_ gnd vdd FILL
X_10536_ _10536_/A _10535_/A _10536_/C gnd _10536_/Y vdd OAI21X1
XFILL_5__10061_ gnd vdd FILL
XFILL112040x3050 gnd vdd FILL
XFILL_2__8632_ gnd vdd FILL
XFILL_3__11240_ gnd vdd FILL
XFILL_4__10791_ gnd vdd FILL
XFILL_5_BUFX2_insert580 gnd vdd FILL
XFILL_4__9548_ gnd vdd FILL
XFILL_5_BUFX2_insert591 gnd vdd FILL
XFILL_2__11970_ gnd vdd FILL
XFILL_5__8341_ gnd vdd FILL
XFILL_0__11060_ gnd vdd FILL
X_16043_ _16041_/Y _16043_/B gnd _16044_/B vdd NOR2X1
X_13255_ _13289_/B _13274_/A gnd _13259_/C vdd NAND2X1
XFILL_4__12530_ gnd vdd FILL
X_10467_ _14078_/A _6999_/CLK _7000_/R vdd _10467_/D gnd vdd DFFSR
XFILL_2__10921_ gnd vdd FILL
XFILL_1__12350_ gnd vdd FILL
XFILL_0__10011_ gnd vdd FILL
XFILL_3__11171_ gnd vdd FILL
X_12206_ _12117_/B _12949_/Q gnd _12207_/C vdd NAND2X1
XFILL_4__9479_ gnd vdd FILL
XFILL_5__8272_ gnd vdd FILL
XSFILL98840x76050 gnd vdd FILL
XFILL_5__13820_ gnd vdd FILL
XFILL_6__11282_ gnd vdd FILL
XFILL_3__10122_ gnd vdd FILL
XFILL_4__12461_ gnd vdd FILL
X_13186_ _13186_/Q _13184_/CLK _8033_/R vdd _13114_/Y gnd vdd DFFSR
XSFILL59080x37050 gnd vdd FILL
XFILL_1__11301_ gnd vdd FILL
XFILL_2__13640_ gnd vdd FILL
X_10398_ _10363_/B _7838_/B gnd _10398_/Y vdd NAND2X1
XFILL_5__7223_ gnd vdd FILL
XFILL_1__12281_ gnd vdd FILL
XFILL_2__8494_ gnd vdd FILL
XFILL_4__14200_ gnd vdd FILL
XSFILL99480x42050 gnd vdd FILL
XFILL_6__10233_ gnd vdd FILL
X_12137_ _12137_/A _12844_/A gnd _12138_/C vdd NAND2X1
XFILL_4__11412_ gnd vdd FILL
XFILL_4__15180_ gnd vdd FILL
XFILL_5__13751_ gnd vdd FILL
XSFILL74120x40050 gnd vdd FILL
XFILL_4__12392_ gnd vdd FILL
XFILL_5__10963_ gnd vdd FILL
XFILL_1__14020_ gnd vdd FILL
XFILL_3__14930_ gnd vdd FILL
XFILL_3__10053_ gnd vdd FILL
XFILL_2__7445_ gnd vdd FILL
XFILL_1__11232_ gnd vdd FILL
XFILL_2_CLKBUF1_insert150 gnd vdd FILL
XFILL_2__13571_ gnd vdd FILL
XFILL_0__11962_ gnd vdd FILL
XFILL_0__14750_ gnd vdd FILL
XFILL_2__10783_ gnd vdd FILL
XFILL_2_CLKBUF1_insert161 gnd vdd FILL
XFILL_5__12702_ gnd vdd FILL
XFILL_4__14131_ gnd vdd FILL
XFILL_2__15310_ gnd vdd FILL
X_12068_ _12012_/A _12809_/Q _11996_/C gnd _12070_/B vdd NAND3X1
XFILL_2_CLKBUF1_insert172 gnd vdd FILL
XFILL_4__11343_ gnd vdd FILL
XFILL_3__14861_ gnd vdd FILL
XFILL_5__13682_ gnd vdd FILL
XFILL_2__12522_ gnd vdd FILL
XSFILL53800x39050 gnd vdd FILL
XFILL_2_CLKBUF1_insert183 gnd vdd FILL
XFILL_5__10894_ gnd vdd FILL
XFILL_2_CLKBUF1_insert194 gnd vdd FILL
XFILL_0__10913_ gnd vdd FILL
XFILL_2__16290_ gnd vdd FILL
XSFILL34040x6050 gnd vdd FILL
XFILL_1__11163_ gnd vdd FILL
XFILL_0__13701_ gnd vdd FILL
XFILL_2__7376_ gnd vdd FILL
XSFILL63960x83050 gnd vdd FILL
XFILL_0__11893_ gnd vdd FILL
XFILL_5__7085_ gnd vdd FILL
XFILL_0__14681_ gnd vdd FILL
XFILL_5__15421_ gnd vdd FILL
X_11019_ _12242_/Y _12135_/Y gnd _11019_/Y vdd AND2X2
XFILL_5__12633_ gnd vdd FILL
XFILL_3__13812_ gnd vdd FILL
XSFILL13800x55050 gnd vdd FILL
XFILL_2__9115_ gnd vdd FILL
XFILL_4__14062_ gnd vdd FILL
XFILL_1__10114_ gnd vdd FILL
XFILL_2__15241_ gnd vdd FILL
XFILL_4__11274_ gnd vdd FILL
XFILL_3__14792_ gnd vdd FILL
XFILL_2__12453_ gnd vdd FILL
XFILL_0__13632_ gnd vdd FILL
XFILL_1__15971_ gnd vdd FILL
XFILL_1__11094_ gnd vdd FILL
XFILL_0__8130_ gnd vdd FILL
XFILL_4__13013_ gnd vdd FILL
XFILL_5__15352_ gnd vdd FILL
X_15827_ _15708_/A _15826_/Y _15708_/C gnd _15851_/B vdd NOR3X1
XFILL_3__13743_ gnd vdd FILL
XBUFX2_insert5 _13280_/Y gnd _7369_/B vdd BUFX2
XFILL_2__11404_ gnd vdd FILL
XFILL_3__10955_ gnd vdd FILL
XFILL_1__10045_ gnd vdd FILL
XFILL_2_BUFX2_insert470 gnd vdd FILL
XFILL_2__15172_ gnd vdd FILL
XFILL_1__14922_ gnd vdd FILL
XFILL_2_BUFX2_insert481 gnd vdd FILL
XFILL_2__12384_ gnd vdd FILL
XFILL_0__16351_ gnd vdd FILL
XFILL_0__13563_ gnd vdd FILL
XFILL_0__10775_ gnd vdd FILL
XFILL_5__14303_ gnd vdd FILL
XFILL_2_BUFX2_insert492 gnd vdd FILL
XFILL_0__8061_ gnd vdd FILL
XFILL_5__11515_ gnd vdd FILL
X_15758_ _15758_/A _15758_/B gnd _15758_/Y vdd NAND2X1
XFILL_2__14123_ gnd vdd FILL
XFILL_5__12495_ gnd vdd FILL
XFILL_4__10156_ gnd vdd FILL
XFILL_5__15283_ gnd vdd FILL
XFILL_0__15302_ gnd vdd FILL
XFILL_3__13674_ gnd vdd FILL
XFILL_0__12514_ gnd vdd FILL
XFILL_2__11335_ gnd vdd FILL
XFILL_1__14853_ gnd vdd FILL
XFILL_3__10886_ gnd vdd FILL
XFILL_0__13494_ gnd vdd FILL
XFILL_0__16282_ gnd vdd FILL
XFILL_3__15413_ gnd vdd FILL
XFILL_5__14234_ gnd vdd FILL
X_14709_ _14709_/A _14705_/Y gnd _14714_/C vdd NOR2X1
XFILL_5__11446_ gnd vdd FILL
XFILL_5__7987_ gnd vdd FILL
X_15689_ _15689_/A _15688_/Y _15689_/C gnd _15690_/B vdd NAND3X1
XFILL_3__12625_ gnd vdd FILL
X_7640_ _7548_/A _7640_/CLK _7515_/R vdd _7640_/D gnd vdd DFFSR
XFILL_1__13804_ gnd vdd FILL
XFILL_3__16393_ gnd vdd FILL
XFILL_2__14054_ gnd vdd FILL
XFILL_4__14964_ gnd vdd FILL
XFILL_3__9790_ gnd vdd FILL
XFILL_0__15233_ gnd vdd FILL
XFILL_0__12445_ gnd vdd FILL
XFILL_2__11266_ gnd vdd FILL
XFILL_5__6938_ gnd vdd FILL
XFILL_5__9726_ gnd vdd FILL
XFILL_1__14784_ gnd vdd FILL
XFILL_1__11996_ gnd vdd FILL
XFILL_3__15344_ gnd vdd FILL
XFILL_5__14165_ gnd vdd FILL
XFILL_2__13005_ gnd vdd FILL
X_7571_ _7569_/Y _7570_/A _7571_/C gnd _7647_/D vdd OAI21X1
XFILL_4__13915_ gnd vdd FILL
XFILL_5__11377_ gnd vdd FILL
XFILL_3__8741_ gnd vdd FILL
XSFILL99560x22050 gnd vdd FILL
XFILL_0__15164_ gnd vdd FILL
XFILL_1__13735_ gnd vdd FILL
XFILL_2__11197_ gnd vdd FILL
XFILL_4__14895_ gnd vdd FILL
XFILL_1__10947_ gnd vdd FILL
XFILL_0__12376_ gnd vdd FILL
XSFILL74200x20050 gnd vdd FILL
X_9310_ _9310_/Q _7790_/CLK _9561_/R vdd _9310_/D gnd vdd DFFSR
XFILL_5__6869_ gnd vdd FILL
XFILL_5__13116_ gnd vdd FILL
XFILL_5__9657_ gnd vdd FILL
XFILL_0__8963_ gnd vdd FILL
XFILL_3__11507_ gnd vdd FILL
XFILL_5__14096_ gnd vdd FILL
XFILL_4__13846_ gnd vdd FILL
XFILL_0__14115_ gnd vdd FILL
XFILL_3__15275_ gnd vdd FILL
XFILL_2__10148_ gnd vdd FILL
XBUFX2_insert480 _14979_/Y gnd _15244_/C vdd BUFX2
XFILL_2__9879_ gnd vdd FILL
XFILL_3__12487_ gnd vdd FILL
XFILL_0__11327_ gnd vdd FILL
XFILL_1__13666_ gnd vdd FILL
XFILL_5__8608_ gnd vdd FILL
XFILL_6__14406_ gnd vdd FILL
XFILL_0__15095_ gnd vdd FILL
XBUFX2_insert491 _13471_/Y gnd _13479_/C vdd BUFX2
XSFILL59000x81050 gnd vdd FILL
XFILL_6__8381_ gnd vdd FILL
XFILL_1__10878_ gnd vdd FILL
XFILL_3__14226_ gnd vdd FILL
X_9241_ _9241_/A _9240_/A _9241_/C gnd _9313_/D vdd OAI21X1
XFILL_5__10259_ gnd vdd FILL
XFILL_0__8894_ gnd vdd FILL
XFILL_1__15405_ gnd vdd FILL
XFILL_6__12598_ gnd vdd FILL
XSFILL109400x48050 gnd vdd FILL
XFILL_3__11438_ gnd vdd FILL
XFILL_3__7623_ gnd vdd FILL
XFILL_1__12617_ gnd vdd FILL
XFILL_4__13777_ gnd vdd FILL
XFILL_0__14046_ gnd vdd FILL
XFILL_4__10989_ gnd vdd FILL
XFILL_2__14956_ gnd vdd FILL
XFILL_1__16385_ gnd vdd FILL
XFILL_6__7332_ gnd vdd FILL
XFILL_0__11258_ gnd vdd FILL
XFILL_1__13597_ gnd vdd FILL
XFILL_0__7845_ gnd vdd FILL
XFILL_4__15516_ gnd vdd FILL
X_9172_ _9086_/B _9172_/B gnd _9172_/Y vdd NAND2X1
XFILL_4__12728_ gnd vdd FILL
XSFILL49080x69050 gnd vdd FILL
XFILL_3__14157_ gnd vdd FILL
XFILL_2__13907_ gnd vdd FILL
XFILL_1__15336_ gnd vdd FILL
XFILL_3__7554_ gnd vdd FILL
XFILL_3__11369_ gnd vdd FILL
XFILL_2__14887_ gnd vdd FILL
X_8123_ _8173_/Q gnd _8123_/Y vdd INVX1
XFILL_0__11189_ gnd vdd FILL
XSFILL64120x72050 gnd vdd FILL
XFILL_3__13108_ gnd vdd FILL
XFILL_4__15447_ gnd vdd FILL
XFILL_4__12659_ gnd vdd FILL
XFILL_2__13838_ gnd vdd FILL
XFILL_5__14998_ gnd vdd FILL
XFILL_3__14088_ gnd vdd FILL
XFILL_6__9002_ gnd vdd FILL
XFILL_3__7485_ gnd vdd FILL
XFILL_6__16007_ gnd vdd FILL
XFILL_3_BUFX2_insert709 gnd vdd FILL
XFILL_1__15267_ gnd vdd FILL
XFILL_6__13219_ gnd vdd FILL
XFILL_1__12479_ gnd vdd FILL
XFILL_0__9515_ gnd vdd FILL
XFILL_0__15997_ gnd vdd FILL
X_8054_ _8150_/Q gnd _8054_/Y vdd INVX1
XFILL_3__9224_ gnd vdd FILL
XFILL_3__13039_ gnd vdd FILL
XFILL_5__13949_ gnd vdd FILL
XFILL_1__14218_ gnd vdd FILL
XFILL_4__15378_ gnd vdd FILL
XFILL_2__13769_ gnd vdd FILL
XFILL_1_BUFX2_insert20 gnd vdd FILL
X_7005_ _7005_/Q _7005_/CLK _7133_/R vdd _6925_/Y gnd vdd DFFSR
XFILL_1__15198_ gnd vdd FILL
XFILL_1_BUFX2_insert31 gnd vdd FILL
XFILL_0__14948_ gnd vdd FILL
XSFILL43960x30050 gnd vdd FILL
XFILL_1_BUFX2_insert42 gnd vdd FILL
XFILL_2__15508_ gnd vdd FILL
XFILL_4__14329_ gnd vdd FILL
XFILL_1_BUFX2_insert53 gnd vdd FILL
XFILL_3__9155_ gnd vdd FILL
XFILL_1__14149_ gnd vdd FILL
XFILL_1_BUFX2_insert64 gnd vdd FILL
XFILL_1_BUFX2_insert75 gnd vdd FILL
XFILL_0__14879_ gnd vdd FILL
XFILL_5__15619_ gnd vdd FILL
XFILL_1_BUFX2_insert86 gnd vdd FILL
XFILL_0__9377_ gnd vdd FILL
XFILL_3__8106_ gnd vdd FILL
XFILL_1_BUFX2_insert97 gnd vdd FILL
XFILL_2__15439_ gnd vdd FILL
XFILL_3__9086_ gnd vdd FILL
XFILL_0__8328_ gnd vdd FILL
XFILL_1__7121_ gnd vdd FILL
X_8956_ _9048_/Q gnd _8956_/Y vdd INVX1
XSFILL23720x38050 gnd vdd FILL
XSFILL33880x82050 gnd vdd FILL
XFILL_1__7052_ gnd vdd FILL
X_7907_ _7907_/Q _6999_/CLK _7011_/R vdd _7907_/D gnd vdd DFFSR
XFILL_0__8259_ gnd vdd FILL
X_8887_ _8887_/A _8845_/B _8887_/C gnd _8887_/Y vdd OAI21X1
XSFILL18840x6050 gnd vdd FILL
XFILL_4__8850_ gnd vdd FILL
XFILL_4__7801_ gnd vdd FILL
X_7838_ _7814_/A _7838_/B gnd _7839_/C vdd NAND2X1
XFILL_4__8781_ gnd vdd FILL
XSFILL64200x52050 gnd vdd FILL
XFILL_3__9988_ gnd vdd FILL
XSFILL49560x70050 gnd vdd FILL
X_7769_ _7769_/Q _8921_/CLK _9049_/R vdd _7769_/D gnd vdd DFFSR
XFILL_4__7732_ gnd vdd FILL
X_9508_ _9548_/B _8228_/B gnd _9508_/Y vdd NAND2X1
XFILL_1__7954_ gnd vdd FILL
XFILL_1__6905_ gnd vdd FILL
X_11370_ _11235_/Y _11236_/Y _11006_/A gnd _11370_/Y vdd OAI21X1
XFILL_4__9402_ gnd vdd FILL
X_9439_ _9361_/A _7274_/CLK _7274_/R vdd _9439_/D gnd vdd DFFSR
XSFILL84920x22050 gnd vdd FILL
XFILL_1__7885_ gnd vdd FILL
XSFILL28840x71050 gnd vdd FILL
XSFILL69480x21050 gnd vdd FILL
XFILL_4_BUFX2_insert510 gnd vdd FILL
XFILL_4__7594_ gnd vdd FILL
X_10321_ _10271_/B _7889_/B gnd _10322_/C vdd NAND2X1
XFILL_4_BUFX2_insert521 gnd vdd FILL
XFILL_1__9624_ gnd vdd FILL
XFILL_1__6836_ gnd vdd FILL
XFILL_4_BUFX2_insert532 gnd vdd FILL
XFILL_4_BUFX2_insert543 gnd vdd FILL
X_13040_ _13038_/Y vdd _13040_/C gnd _13076_/D vdd OAI21X1
XFILL_4_BUFX2_insert554 gnd vdd FILL
X_10252_ _10294_/A _7180_/B gnd _10252_/Y vdd NAND2X1
XFILL_4_BUFX2_insert565 gnd vdd FILL
XSFILL8760x69050 gnd vdd FILL
XFILL_1__9555_ gnd vdd FILL
XSFILL44040x1050 gnd vdd FILL
XSFILL23800x18050 gnd vdd FILL
XFILL_4_BUFX2_insert576 gnd vdd FILL
XFILL_4__9264_ gnd vdd FILL
XSFILL84200x6050 gnd vdd FILL
XFILL_4_BUFX2_insert587 gnd vdd FILL
XFILL_4_BUFX2_insert598 gnd vdd FILL
XFILL_1__8506_ gnd vdd FILL
X_10183_ _10225_/Q gnd _10185_/A vdd INVX1
XFILL_1__9486_ gnd vdd FILL
XFILL_4__8215_ gnd vdd FILL
XFILL_2__7230_ gnd vdd FILL
X_14991_ _12767_/A _16216_/B gnd _14991_/Y vdd NOR2X1
XFILL_4__8146_ gnd vdd FILL
X_13942_ _13931_/Y _13934_/Y _13941_/Y gnd _13942_/Y vdd NAND3X1
XFILL_3_CLKBUF1_insert201 gnd vdd FILL
XFILL_3_CLKBUF1_insert212 gnd vdd FILL
XFILL_1__8368_ gnd vdd FILL
XFILL_2__7161_ gnd vdd FILL
XFILL_3_CLKBUF1_insert223 gnd vdd FILL
XFILL_4__8077_ gnd vdd FILL
X_13873_ _13864_/Y _13873_/B _13872_/Y gnd _13873_/Y vdd NAND3X1
XFILL_1__7319_ gnd vdd FILL
XFILL_2__7092_ gnd vdd FILL
X_15612_ _14135_/C gnd _15614_/B vdd INVX1
XFILL_6__10920_ gnd vdd FILL
XFILL_5__8890_ gnd vdd FILL
X_12824_ _12824_/A vdd gnd _12825_/C vdd NAND2X1
XFILL_4__10010_ gnd vdd FILL
XFILL_1_BUFX2_insert400 gnd vdd FILL
XFILL_1_BUFX2_insert411 gnd vdd FILL
XSFILL28920x51050 gnd vdd FILL
XFILL_1_BUFX2_insert422 gnd vdd FILL
XFILL_1_BUFX2_insert433 gnd vdd FILL
XFILL_0__10560_ gnd vdd FILL
XFILL_5__7841_ gnd vdd FILL
XFILL_5__11300_ gnd vdd FILL
XFILL_1_BUFX2_insert444 gnd vdd FILL
X_15543_ _7706_/A gnd _15544_/B vdd INVX1
X_12755_ _11884_/A gnd _12755_/Y vdd INVX1
XFILL_1_BUFX2_insert455 gnd vdd FILL
XFILL_5__12280_ gnd vdd FILL
XFILL_2__11120_ gnd vdd FILL
XFILL_1_BUFX2_insert466 gnd vdd FILL
XFILL_3__10671_ gnd vdd FILL
XFILL_1_BUFX2_insert477 gnd vdd FILL
XFILL_1__11850_ gnd vdd FILL
XFILL_1_BUFX2_insert488 gnd vdd FILL
X_11706_ _11074_/C _11704_/Y _11706_/C gnd _11717_/B vdd AOI21X1
XFILL_0__10491_ gnd vdd FILL
XFILL_5__11231_ gnd vdd FILL
XFILL_3__12410_ gnd vdd FILL
XFILL_4__8979_ gnd vdd FILL
X_15474_ _15474_/A _16294_/C gnd _15481_/A vdd NAND2X1
XFILL_1_BUFX2_insert499 gnd vdd FILL
X_12686_ _12413_/B _12809_/CLK _12809_/R vdd _12686_/D gnd vdd DFFSR
XFILL_4__11961_ gnd vdd FILL
XFILL_2__9802_ gnd vdd FILL
XFILL_2__11051_ gnd vdd FILL
XFILL_3__13390_ gnd vdd FILL
XFILL_0__12230_ gnd vdd FILL
XFILL_1__10801_ gnd vdd FILL
XFILL_5__9511_ gnd vdd FILL
XFILL_2__7994_ gnd vdd FILL
XSFILL99480x37050 gnd vdd FILL
XFILL_1__11781_ gnd vdd FILL
X_14425_ _9394_/A gnd _14425_/Y vdd INVX1
XFILL_4__10912_ gnd vdd FILL
X_11637_ _11615_/Y _11637_/B _11636_/Y gnd _11637_/Y vdd OAI21X1
XFILL_5__11162_ gnd vdd FILL
XFILL_4__13700_ gnd vdd FILL
XSFILL74120x35050 gnd vdd FILL
XFILL_3__12341_ gnd vdd FILL
XFILL_2__10002_ gnd vdd FILL
XFILL_2__9733_ gnd vdd FILL
XFILL_2__6945_ gnd vdd FILL
XFILL_4__11892_ gnd vdd FILL
XFILL_4__14680_ gnd vdd FILL
XFILL_1__13520_ gnd vdd FILL
XFILL_0__12161_ gnd vdd FILL
XFILL_5__10113_ gnd vdd FILL
X_14356_ _14356_/A _14345_/Y gnd _14357_/B vdd NOR2X1
XFILL_5__15970_ gnd vdd FILL
XFILL_4__13631_ gnd vdd FILL
XFILL_2__14810_ gnd vdd FILL
XFILL_3__15060_ gnd vdd FILL
XFILL_5__11093_ gnd vdd FILL
X_11568_ _11623_/B _11623_/A gnd _11630_/B vdd NOR2X1
XFILL_2__9664_ gnd vdd FILL
XFILL_3__12272_ gnd vdd FILL
XFILL_0__11112_ gnd vdd FILL
XFILL_1__10663_ gnd vdd FILL
XFILL_1__13451_ gnd vdd FILL
XFILL_2__6876_ gnd vdd FILL
XFILL_2__15790_ gnd vdd FILL
X_13307_ _13266_/A _13248_/A _13300_/B gnd _13308_/A vdd AOI21X1
XFILL_0__12092_ gnd vdd FILL
XFILL_5__9373_ gnd vdd FILL
XFILL_5__10044_ gnd vdd FILL
XFILL_3__14011_ gnd vdd FILL
X_10519_ _13983_/A gnd _10521_/A vdd INVX1
XFILL_5__14921_ gnd vdd FILL
XFILL_2__8615_ gnd vdd FILL
XFILL_4__13562_ gnd vdd FILL
XFILL_4__16350_ gnd vdd FILL
X_14287_ _14287_/A _14286_/Y _14287_/C gnd _14287_/Y vdd NAND3X1
XFILL_3__11223_ gnd vdd FILL
XFILL_1__12402_ gnd vdd FILL
XFILL_2__14741_ gnd vdd FILL
X_11499_ _11185_/A _11185_/B _11513_/B gnd _11500_/C vdd OAI21X1
XFILL_4__10774_ gnd vdd FILL
XFILL_0__15920_ gnd vdd FILL
XFILL_5__8324_ gnd vdd FILL
XFILL_1__16170_ gnd vdd FILL
XFILL_2__11953_ gnd vdd FILL
XFILL_0__11043_ gnd vdd FILL
XFILL_2__9595_ gnd vdd FILL
X_16026_ _15394_/C _14598_/Y _16026_/C _16026_/D gnd _16027_/A vdd OAI22X1
XFILL_1__13382_ gnd vdd FILL
X_13238_ _13237_/Y _13335_/A gnd _13297_/C vdd NAND2X1
XFILL_0__7630_ gnd vdd FILL
XFILL_4__15301_ gnd vdd FILL
XFILL_5__14852_ gnd vdd FILL
XFILL_4__12513_ gnd vdd FILL
XFILL_2__10904_ gnd vdd FILL
XFILL112280x61050 gnd vdd FILL
XFILL_3__11154_ gnd vdd FILL
XFILL_4__13493_ gnd vdd FILL
XFILL_1__15121_ gnd vdd FILL
XFILL_4__16281_ gnd vdd FILL
XFILL_1__12333_ gnd vdd FILL
XFILL_2__14672_ gnd vdd FILL
XFILL_5__8255_ gnd vdd FILL
XFILL_2__11884_ gnd vdd FILL
XFILL_0__15851_ gnd vdd FILL
XFILL_5__13803_ gnd vdd FILL
XSFILL113960x47050 gnd vdd FILL
XFILL_6__14053_ gnd vdd FILL
XFILL_4__15232_ gnd vdd FILL
XFILL_0__7561_ gnd vdd FILL
X_13169_ _12108_/B gnd _13169_/Y vdd INVX1
XFILL_4__12444_ gnd vdd FILL
XFILL_2__16411_ gnd vdd FILL
XFILL_3__10105_ gnd vdd FILL
XFILL_2__13623_ gnd vdd FILL
XFILL_5__14783_ gnd vdd FILL
XFILL_0__14802_ gnd vdd FILL
XFILL_5__7206_ gnd vdd FILL
XFILL_5__11995_ gnd vdd FILL
XFILL_3__15962_ gnd vdd FILL
XFILL_1__15052_ gnd vdd FILL
XFILL_1__12264_ gnd vdd FILL
XFILL_2__8477_ gnd vdd FILL
XFILL_3__11085_ gnd vdd FILL
XFILL_2__10835_ gnd vdd FILL
XFILL_0__9300_ gnd vdd FILL
XFILL_0__15782_ gnd vdd FILL
XFILL_5__8186_ gnd vdd FILL
XFILL_0__12994_ gnd vdd FILL
XFILL_5__13734_ gnd vdd FILL
XFILL_5__10946_ gnd vdd FILL
XFILL_2__16342_ gnd vdd FILL
XFILL_2__7428_ gnd vdd FILL
XFILL_1__14003_ gnd vdd FILL
XFILL_0__7492_ gnd vdd FILL
XFILL_4__12375_ gnd vdd FILL
XFILL_3__10036_ gnd vdd FILL
XFILL_4__15163_ gnd vdd FILL
XFILL_3__14913_ gnd vdd FILL
XFILL_2__13554_ gnd vdd FILL
XFILL_1__11215_ gnd vdd FILL
XFILL_2__10766_ gnd vdd FILL
XFILL_3__15893_ gnd vdd FILL
XFILL_0__14733_ gnd vdd FILL
XFILL_1__12195_ gnd vdd FILL
XFILL_0__9231_ gnd vdd FILL
XFILL_0__11945_ gnd vdd FILL
XFILL_4__14114_ gnd vdd FILL
XFILL_4__11326_ gnd vdd FILL
XFILL_5__13665_ gnd vdd FILL
XFILL_2__12505_ gnd vdd FILL
XSFILL28840x1050 gnd vdd FILL
XFILL_4__15094_ gnd vdd FILL
XFILL_3__14844_ gnd vdd FILL
XFILL_2__7359_ gnd vdd FILL
XFILL_5__10877_ gnd vdd FILL
XFILL_1__11146_ gnd vdd FILL
XFILL_2__16273_ gnd vdd FILL
XSFILL18680x21050 gnd vdd FILL
XFILL_2__13485_ gnd vdd FILL
XFILL_0__11876_ gnd vdd FILL
XFILL_5__15404_ gnd vdd FILL
XFILL_5__7068_ gnd vdd FILL
XFILL_0__14664_ gnd vdd FILL
XSFILL74200x15050 gnd vdd FILL
XFILL_2__10697_ gnd vdd FILL
XFILL_5__12616_ gnd vdd FILL
XFILL_0__9162_ gnd vdd FILL
XFILL_4__14045_ gnd vdd FILL
X_8810_ _8810_/Q _7535_/CLK _7523_/R vdd _8810_/D gnd vdd DFFSR
XFILL_5__16384_ gnd vdd FILL
XFILL_2__15224_ gnd vdd FILL
XFILL_4__11257_ gnd vdd FILL
X_9790_ _9838_/Q gnd _9790_/Y vdd INVX1
XFILL_5__13596_ gnd vdd FILL
XFILL_2__12436_ gnd vdd FILL
XFILL_0__16403_ gnd vdd FILL
XFILL_0__13615_ gnd vdd FILL
XFILL_3__11987_ gnd vdd FILL
XFILL_1__15954_ gnd vdd FILL
XFILL_1__11077_ gnd vdd FILL
XFILL_3__14775_ gnd vdd FILL
XFILL_0__10827_ gnd vdd FILL
XFILL_0__8113_ gnd vdd FILL
XSFILL59000x76050 gnd vdd FILL
XFILL_0__14595_ gnd vdd FILL
XFILL_5__15335_ gnd vdd FILL
X_8741_ _8741_/A _8740_/A _8741_/C gnd _8741_/Y vdd OAI21X1
XFILL_2__9029_ gnd vdd FILL
XFILL_0__9093_ gnd vdd FILL
XFILL_6__14886_ gnd vdd FILL
XFILL_3__9911_ gnd vdd FILL
XFILL_3__10938_ gnd vdd FILL
XFILL_1__10028_ gnd vdd FILL
XFILL_2__15155_ gnd vdd FILL
XFILL_4__11188_ gnd vdd FILL
XFILL_3__13726_ gnd vdd FILL
XFILL_1__14905_ gnd vdd FILL
XSFILL99400x81050 gnd vdd FILL
XFILL_2__12367_ gnd vdd FILL
XFILL_0__16334_ gnd vdd FILL
XFILL_0__13546_ gnd vdd FILL
XFILL_0__10758_ gnd vdd FILL
XFILL_1__15885_ gnd vdd FILL
XFILL_4__10139_ gnd vdd FILL
XFILL_2__14106_ gnd vdd FILL
XFILL_5__15266_ gnd vdd FILL
XFILL_3__13657_ gnd vdd FILL
XFILL_6_BUFX2_insert638 gnd vdd FILL
XFILL_5__12478_ gnd vdd FILL
XFILL_2__11318_ gnd vdd FILL
X_8672_ _8596_/A _7535_/CLK _8682_/R vdd _8598_/Y gnd vdd DFFSR
XFILL_1__14836_ gnd vdd FILL
XFILL_4__15996_ gnd vdd FILL
XFILL_2__15086_ gnd vdd FILL
XSFILL38840x34050 gnd vdd FILL
XFILL_0__16265_ gnd vdd FILL
XFILL_2__12298_ gnd vdd FILL
XFILL_5__14217_ gnd vdd FILL
XFILL112360x41050 gnd vdd FILL
XFILL_0__10689_ gnd vdd FILL
XFILL_0__13477_ gnd vdd FILL
XSFILL64120x67050 gnd vdd FILL
XFILL_3__12608_ gnd vdd FILL
X_7623_ _7623_/A gnd _7623_/Y vdd INVX1
XFILL_5__11429_ gnd vdd FILL
XFILL_5__15197_ gnd vdd FILL
XFILL_2__14037_ gnd vdd FILL
XFILL_4__14947_ gnd vdd FILL
XFILL_3__13588_ gnd vdd FILL
XFILL_0__15216_ gnd vdd FILL
XFILL_3__16376_ gnd vdd FILL
XFILL_3__9773_ gnd vdd FILL
XFILL_2__11249_ gnd vdd FILL
XFILL_0__12428_ gnd vdd FILL
XFILL_3__6985_ gnd vdd FILL
XFILL_1__14767_ gnd vdd FILL
XFILL_0__16196_ gnd vdd FILL
XFILL_1__11979_ gnd vdd FILL
XFILL_5__14148_ gnd vdd FILL
XFILL_0__9995_ gnd vdd FILL
XFILL_3__15327_ gnd vdd FILL
X_7554_ _7554_/A gnd _7556_/A vdd INVX1
XFILL_3__8724_ gnd vdd FILL
XFILL_4__14878_ gnd vdd FILL
XFILL_1__13718_ gnd vdd FILL
XFILL_0__12359_ gnd vdd FILL
XFILL_0__15147_ gnd vdd FILL
XFILL_1__14698_ gnd vdd FILL
XSFILL3560x74050 gnd vdd FILL
X_7485_ _7483_/Y _7425_/B _7485_/C gnd _7485_/Y vdd OAI21X1
XFILL_4__13829_ gnd vdd FILL
XFILL_3__15258_ gnd vdd FILL
XFILL_5__14079_ gnd vdd FILL
XFILL_3__8655_ gnd vdd FILL
XFILL_1__13649_ gnd vdd FILL
XFILL_2__15988_ gnd vdd FILL
XFILL_0__15078_ gnd vdd FILL
XFILL_3__14209_ gnd vdd FILL
X_9224_ _9224_/A gnd _9226_/A vdd INVX1
XFILL_3__7606_ gnd vdd FILL
XFILL_1__7670_ gnd vdd FILL
XFILL_0__8877_ gnd vdd FILL
XSFILL99160x50 gnd vdd FILL
XSFILL8600x11050 gnd vdd FILL
XFILL_3__15189_ gnd vdd FILL
XFILL_3__8586_ gnd vdd FILL
XFILL_0__14029_ gnd vdd FILL
XFILL_2__14939_ gnd vdd FILL
XFILL_1__16368_ gnd vdd FILL
XFILL_0__7828_ gnd vdd FILL
X_9155_ _9155_/A _9170_/B _9154_/Y gnd _9155_/Y vdd OAI21X1
XFILL_1__15319_ gnd vdd FILL
XFILL_3_BUFX2_insert506 gnd vdd FILL
XFILL_1__16299_ gnd vdd FILL
XFILL_1__9340_ gnd vdd FILL
XFILL_3_BUFX2_insert517 gnd vdd FILL
X_8106_ _8107_/B _9770_/B gnd _8107_/C vdd NAND2X1
XFILL_0__7759_ gnd vdd FILL
XSFILL33880x77050 gnd vdd FILL
XFILL_3_BUFX2_insert528 gnd vdd FILL
X_9086_ _9084_/Y _9086_/B _9086_/C gnd _9176_/D vdd OAI21X1
XFILL_3_BUFX2_insert539 gnd vdd FILL
XFILL_3__7468_ gnd vdd FILL
XFILL_4__8000_ gnd vdd FILL
XFILL_1__9271_ gnd vdd FILL
X_8037_ _7971_/A _8165_/CLK _8165_/R vdd _8037_/D gnd vdd DFFSR
XFILL_3__9207_ gnd vdd FILL
XFILL112440x21050 gnd vdd FILL
XSFILL64200x47050 gnd vdd FILL
XFILL_0__9429_ gnd vdd FILL
XFILL_1__8222_ gnd vdd FILL
XFILL_3__9138_ gnd vdd FILL
XSFILL68680x6050 gnd vdd FILL
XSFILL24200x63050 gnd vdd FILL
XSFILL104120x3050 gnd vdd FILL
X_9988_ _9988_/A _9996_/A _9988_/C gnd _9988_/Y vdd OAI21X1
XSFILL8600x2050 gnd vdd FILL
XFILL_1__7104_ gnd vdd FILL
XSFILL3640x54050 gnd vdd FILL
X_10870_ _12707_/A gnd _10871_/B vdd INVX1
X_8939_ _8939_/Q _7389_/CLK _8285_/R vdd _8887_/Y gnd vdd DFFSR
XFILL_1__8084_ gnd vdd FILL
XFILL_4__8902_ gnd vdd FILL
XSFILL28840x66050 gnd vdd FILL
XFILL_4__9882_ gnd vdd FILL
XFILL_1__7035_ gnd vdd FILL
XFILL_4__8833_ gnd vdd FILL
X_12540_ _12454_/A _12537_/CLK _12536_/R vdd _12540_/D gnd vdd DFFSR
XSFILL104600x9050 gnd vdd FILL
XFILL_0_BUFX2_insert407 gnd vdd FILL
XFILL_0_BUFX2_insert418 gnd vdd FILL
XFILL_4__8764_ gnd vdd FILL
XFILL_0_BUFX2_insert429 gnd vdd FILL
X_12471_ _12469_/Y vdd _12470_/Y gnd _12471_/Y vdd OAI21X1
XFILL_1__8986_ gnd vdd FILL
X_14210_ _7781_/Q gnd _14210_/Y vdd INVX1
XFILL_4__7715_ gnd vdd FILL
XFILL_4__8695_ gnd vdd FILL
X_11422_ _11202_/Y _11848_/A gnd _11423_/C vdd NAND2X1
X_15190_ _7039_/A gnd _15190_/Y vdd INVX1
XSFILL89640x29050 gnd vdd FILL
XFILL_1__7937_ gnd vdd FILL
X_14141_ _14567_/A _14141_/B _14141_/C _13978_/B gnd _14142_/A vdd OAI22X1
X_11353_ _11338_/A _11348_/A _11360_/C gnd _11353_/Y vdd OAI21X1
XFILL_1__7868_ gnd vdd FILL
XSFILL89240x31050 gnd vdd FILL
X_10304_ _10302_/Y _10304_/B _10303_/Y gnd _10350_/D vdd OAI21X1
XFILL_4_BUFX2_insert340 gnd vdd FILL
XFILL_4__7577_ gnd vdd FILL
X_14072_ _14068_/Y _14072_/B gnd _14073_/C vdd NOR2X1
XFILL_2__8400_ gnd vdd FILL
XFILL_4_BUFX2_insert351 gnd vdd FILL
XFILL_1__9607_ gnd vdd FILL
X_11284_ _12278_/Y _12162_/Y gnd _11285_/A vdd NOR2X1
XSFILL13880x24050 gnd vdd FILL
XFILL_2__9380_ gnd vdd FILL
XFILL_4_BUFX2_insert362 gnd vdd FILL
XFILL_4_BUFX2_insert373 gnd vdd FILL
XFILL_1__7799_ gnd vdd FILL
XSFILL3720x34050 gnd vdd FILL
XCLKBUF1_insert119 CLKBUF1_insert187/A gnd _7005_/CLK vdd CLKBUF1
X_13023_ _6894_/A gnd _13023_/Y vdd INVX1
XFILL_4_BUFX2_insert384 gnd vdd FILL
X_10235_ _10235_/A _10325_/B _10235_/C gnd _10327_/D vdd OAI21X1
XFILL_2__8331_ gnd vdd FILL
XFILL_1__9538_ gnd vdd FILL
XFILL_4_BUFX2_insert395 gnd vdd FILL
XSFILL28920x46050 gnd vdd FILL
XFILL_4__10490_ gnd vdd FILL
XSFILL53720x72050 gnd vdd FILL
XFILL_4__9247_ gnd vdd FILL
XSFILL94360x22050 gnd vdd FILL
XFILL_5__10800_ gnd vdd FILL
X_10166_ _10166_/A _8630_/B gnd _10167_/C vdd NAND2X1
XSFILL69000x39050 gnd vdd FILL
XFILL_2__8262_ gnd vdd FILL
XFILL_1__9469_ gnd vdd FILL
XFILL_2__10620_ gnd vdd FILL
XFILL_5__11780_ gnd vdd FILL
XFILL_3__11910_ gnd vdd FILL
XFILL_4__12160_ gnd vdd FILL
XFILL_2__7213_ gnd vdd FILL
XFILL_1__11000_ gnd vdd FILL
X_14974_ _14045_/A _14973_/Y _14068_/C _14974_/D gnd _14974_/Y vdd OAI22X1
X_10097_ _14777_/A _9834_/CLK _7921_/R vdd _10057_/Y gnd vdd DFFSR
XFILL_2__8193_ gnd vdd FILL
XFILL_2__10551_ gnd vdd FILL
XFILL_3__12890_ gnd vdd FILL
XFILL_4__8129_ gnd vdd FILL
XFILL_0__11730_ gnd vdd FILL
XFILL_4__11111_ gnd vdd FILL
XFILL_5__13450_ gnd vdd FILL
XFILL_5__9991_ gnd vdd FILL
X_13925_ _13921_/Y _13925_/B gnd _13925_/Y vdd NOR2X1
XFILL_5__10662_ gnd vdd FILL
XFILL_4__12091_ gnd vdd FILL
XFILL_3__11841_ gnd vdd FILL
XFILL_2__13270_ gnd vdd FILL
XFILL_0__11661_ gnd vdd FILL
XFILL_5__12401_ gnd vdd FILL
X_13856_ _8158_/Q gnd _13856_/Y vdd INVX1
XFILL_6__11952_ gnd vdd FILL
XFILL_4__11042_ gnd vdd FILL
XFILL_3__14560_ gnd vdd FILL
XFILL_5__13381_ gnd vdd FILL
XFILL_2__12221_ gnd vdd FILL
XFILL_2__7075_ gnd vdd FILL
XFILL_0__13400_ gnd vdd FILL
XFILL_3__11772_ gnd vdd FILL
XFILL_1__12951_ gnd vdd FILL
XFILL_0__14380_ gnd vdd FILL
X_12807_ _12807_/Q _12685_/CLK _12685_/R vdd _12745_/Y gnd vdd DFFSR
XFILL_0__11592_ gnd vdd FILL
XFILL_1_BUFX2_insert230 gnd vdd FILL
XFILL_5__15120_ gnd vdd FILL
XSFILL59080x50050 gnd vdd FILL
XFILL_5__8873_ gnd vdd FILL
XFILL_5__12332_ gnd vdd FILL
XSFILL89320x11050 gnd vdd FILL
XFILL_3__13511_ gnd vdd FILL
X_13787_ _13787_/A _13787_/B gnd _13788_/A vdd NAND2X1
XFILL_1_BUFX2_insert241 gnd vdd FILL
XFILL_4__15850_ gnd vdd FILL
XFILL_3__14491_ gnd vdd FILL
XFILL_1_BUFX2_insert252 gnd vdd FILL
XFILL_1__11902_ gnd vdd FILL
XFILL_2__12152_ gnd vdd FILL
X_10999_ _12126_/Y gnd _10999_/Y vdd INVX1
XFILL_0__13331_ gnd vdd FILL
XFILL_1__15670_ gnd vdd FILL
XFILL_0__10543_ gnd vdd FILL
XSFILL109480x17050 gnd vdd FILL
XFILL_1_BUFX2_insert263 gnd vdd FILL
XFILL_5__7824_ gnd vdd FILL
XFILL_1_BUFX2_insert274 gnd vdd FILL
XFILL_1__12882_ gnd vdd FILL
X_12738_ _12768_/A memoryOutData[14] gnd _12739_/C vdd NAND2X1
XFILL_4__14801_ gnd vdd FILL
XFILL_5__15051_ gnd vdd FILL
X_15526_ _7191_/A gnd _15527_/B vdd INVX1
XFILL_1_BUFX2_insert285 gnd vdd FILL
XSFILL8760x8050 gnd vdd FILL
XFILL_3__16230_ gnd vdd FILL
XFILL_3__13442_ gnd vdd FILL
XFILL_5__12263_ gnd vdd FILL
XFILL_2__11103_ gnd vdd FILL
XFILL_1_BUFX2_insert296 gnd vdd FILL
XSFILL110200x67050 gnd vdd FILL
XFILL_1__14621_ gnd vdd FILL
XFILL_4__15781_ gnd vdd FILL
XFILL_3__10654_ gnd vdd FILL
XFILL_0__13262_ gnd vdd FILL
XFILL_2__12083_ gnd vdd FILL
XFILL112280x56050 gnd vdd FILL
XFILL_4__12993_ gnd vdd FILL
XFILL_0__16050_ gnd vdd FILL
XFILL_1__11833_ gnd vdd FILL
XFILL_5__14002_ gnd vdd FILL
XFILL_5__7755_ gnd vdd FILL
X_15457_ _9312_/Q _15892_/B gnd _15466_/A vdd NAND2X1
XFILL_0_BUFX2_insert930 gnd vdd FILL
XFILL_5__11214_ gnd vdd FILL
XFILL_6__10765_ gnd vdd FILL
X_12669_ _12362_/B _12669_/CLK _12799_/R vdd _12669_/D gnd vdd DFFSR
XFILL_4__14732_ gnd vdd FILL
XFILL_5__12194_ gnd vdd FILL
XFILL_3__16161_ gnd vdd FILL
XFILL_0_BUFX2_insert941 gnd vdd FILL
XFILL_2__15911_ gnd vdd FILL
XFILL_0__15001_ gnd vdd FILL
XFILL_4__11944_ gnd vdd FILL
XFILL_0__12213_ gnd vdd FILL
XFILL_3__13373_ gnd vdd FILL
XFILL_2__11034_ gnd vdd FILL
XFILL_0_BUFX2_insert952 gnd vdd FILL
XFILL_1__14552_ gnd vdd FILL
XFILL_2__7977_ gnd vdd FILL
XFILL_0_BUFX2_insert963 gnd vdd FILL
X_14408_ _8170_/Q gnd _14408_/Y vdd INVX1
XFILL_1__11764_ gnd vdd FILL
XFILL_0_BUFX2_insert974 gnd vdd FILL
XFILL_5__11145_ gnd vdd FILL
XFILL_5__7686_ gnd vdd FILL
XFILL_3__15112_ gnd vdd FILL
X_15388_ _15388_/A _15388_/B _15388_/C gnd _15389_/A vdd NAND3X1
XFILL_3__12324_ gnd vdd FILL
XFILL_0__9780_ gnd vdd FILL
XFILL_0_BUFX2_insert985 gnd vdd FILL
XFILL_2__6928_ gnd vdd FILL
XSFILL79240x63050 gnd vdd FILL
XFILL_3__16092_ gnd vdd FILL
XFILL_0_BUFX2_insert996 gnd vdd FILL
XFILL_4__14663_ gnd vdd FILL
XFILL_1__13503_ gnd vdd FILL
XFILL_0__6992_ gnd vdd FILL
XFILL_4__11875_ gnd vdd FILL
XFILL_2__15842_ gnd vdd FILL
XFILL_0__12144_ gnd vdd FILL
XFILL_1__14483_ gnd vdd FILL
XSFILL49800x9050 gnd vdd FILL
XFILL_5__9425_ gnd vdd FILL
XFILL_0__8731_ gnd vdd FILL
X_14339_ _14643_/C _15805_/D _13461_/C _14338_/Y gnd _14340_/A vdd OAI22X1
XFILL_1__11695_ gnd vdd FILL
XFILL_4__16402_ gnd vdd FILL
XFILL_4__13614_ gnd vdd FILL
X_7270_ _7206_/A _8562_/CLK _7270_/R vdd _7208_/Y gnd vdd DFFSR
XFILL_3__15043_ gnd vdd FILL
XFILL_5__15953_ gnd vdd FILL
XFILL_5__11076_ gnd vdd FILL
XFILL_1__16222_ gnd vdd FILL
XFILL_4__10826_ gnd vdd FILL
XFILL_3__8440_ gnd vdd FILL
XFILL_3__12255_ gnd vdd FILL
XFILL_4__14594_ gnd vdd FILL
XFILL_2__6859_ gnd vdd FILL
XFILL_1__13434_ gnd vdd FILL
XFILL_2__9647_ gnd vdd FILL
XFILL_2__15773_ gnd vdd FILL
XSFILL18680x16050 gnd vdd FILL
XFILL_0__12075_ gnd vdd FILL
XFILL_2__12985_ gnd vdd FILL
XFILL_1__10646_ gnd vdd FILL
XSFILL114440x72050 gnd vdd FILL
XFILL_5__9356_ gnd vdd FILL
XFILL_5__14904_ gnd vdd FILL
XFILL_5__10027_ gnd vdd FILL
XFILL_4__16333_ gnd vdd FILL
XFILL_3__11206_ gnd vdd FILL
XFILL_2__14724_ gnd vdd FILL
XFILL_4__10757_ gnd vdd FILL
XFILL_4__13545_ gnd vdd FILL
XFILL_5__15884_ gnd vdd FILL
XFILL_0__15903_ gnd vdd FILL
XFILL_3__12186_ gnd vdd FILL
XFILL_2__11936_ gnd vdd FILL
XFILL_0__11026_ gnd vdd FILL
XFILL_3__8371_ gnd vdd FILL
XFILL_1__16153_ gnd vdd FILL
XFILL_1__13365_ gnd vdd FILL
X_16009_ _16007_/Y _16009_/B gnd _16009_/Y vdd NOR2X1
XFILL_0__7613_ gnd vdd FILL
XFILL_5__9287_ gnd vdd FILL
XFILL_1__10577_ gnd vdd FILL
XFILL_5__14835_ gnd vdd FILL
XFILL_3__7322_ gnd vdd FILL
XFILL_3__11137_ gnd vdd FILL
XFILL_1__15104_ gnd vdd FILL
XFILL_0__8593_ gnd vdd FILL
XFILL_2__8529_ gnd vdd FILL
XFILL_4__16264_ gnd vdd FILL
XFILL_4__10688_ gnd vdd FILL
XFILL_4__13476_ gnd vdd FILL
XFILL_1__12316_ gnd vdd FILL
XFILL_2__14655_ gnd vdd FILL
XFILL_0__15834_ gnd vdd FILL
XFILL_2__11867_ gnd vdd FILL
XSFILL59160x30050 gnd vdd FILL
XFILL_5__8238_ gnd vdd FILL
XFILL_1__16084_ gnd vdd FILL
XFILL_1__13296_ gnd vdd FILL
XFILL_4__15215_ gnd vdd FILL
XFILL_0__7544_ gnd vdd FILL
XFILL_4__12427_ gnd vdd FILL
XFILL_2__13606_ gnd vdd FILL
XFILL_5__14766_ gnd vdd FILL
XFILL_4__16195_ gnd vdd FILL
XFILL_1__15035_ gnd vdd FILL
XFILL_3__15945_ gnd vdd FILL
XFILL_5__11978_ gnd vdd FILL
XFILL_2__10818_ gnd vdd FILL
XFILL_3__11068_ gnd vdd FILL
XFILL_3__7253_ gnd vdd FILL
XFILL_2__14586_ gnd vdd FILL
XFILL_1__12247_ gnd vdd FILL
XSFILL38840x29050 gnd vdd FILL
XFILL_0__15765_ gnd vdd FILL
XFILL_2__11798_ gnd vdd FILL
X_9911_ _9909_/Y _9917_/B _9911_/C gnd _9911_/Y vdd OAI21X1
XFILL_0__12977_ gnd vdd FILL
XFILL_5__13717_ gnd vdd FILL
XFILL_3__10019_ gnd vdd FILL
XFILL_5__10929_ gnd vdd FILL
XFILL_4__12358_ gnd vdd FILL
XFILL112360x36050 gnd vdd FILL
XFILL_2__16325_ gnd vdd FILL
XFILL_0__7475_ gnd vdd FILL
XFILL_4__15146_ gnd vdd FILL
XFILL_5__14697_ gnd vdd FILL
XFILL_2__13537_ gnd vdd FILL
XFILL_3__7184_ gnd vdd FILL
XFILL_0__14716_ gnd vdd FILL
XFILL_2__10749_ gnd vdd FILL
XFILL_3__15876_ gnd vdd FILL
XFILL_1__12178_ gnd vdd FILL
XFILL_0__11928_ gnd vdd FILL
XFILL_0__9214_ gnd vdd FILL
XFILL_0__15696_ gnd vdd FILL
XFILL_4__11309_ gnd vdd FILL
XFILL_5__13648_ gnd vdd FILL
X_9842_ _9802_/A _9436_/CLK _9430_/R vdd _9842_/D gnd vdd DFFSR
XFILL_3__14827_ gnd vdd FILL
XFILL_4__15077_ gnd vdd FILL
XFILL_4__12289_ gnd vdd FILL
XFILL_2__16256_ gnd vdd FILL
XFILL_2__13468_ gnd vdd FILL
XFILL_1__11129_ gnd vdd FILL
XFILL_0__14647_ gnd vdd FILL
XSFILL49080x82050 gnd vdd FILL
XFILL_0__9145_ gnd vdd FILL
XSFILL79320x43050 gnd vdd FILL
XFILL_0__11859_ gnd vdd FILL
XFILL_5__16367_ gnd vdd FILL
XFILL_2__15207_ gnd vdd FILL
XFILL_4__14028_ gnd vdd FILL
XFILL_6__14938_ gnd vdd FILL
XSFILL3560x69050 gnd vdd FILL
XFILL_2__12419_ gnd vdd FILL
X_9773_ _9770_/A _9901_/B gnd _9773_/Y vdd NAND2X1
XFILL_5__13579_ gnd vdd FILL
XFILL_2__16187_ gnd vdd FILL
XFILL_1__15937_ gnd vdd FILL
X_6985_ _6985_/A _6985_/B _6984_/Y gnd _7025_/D vdd OAI21X1
XFILL_3__14758_ gnd vdd FILL
XFILL_2__13399_ gnd vdd FILL
XFILL_0__14578_ gnd vdd FILL
XFILL_5__15318_ gnd vdd FILL
XFILL_6_BUFX2_insert413 gnd vdd FILL
XFILL_6__7864_ gnd vdd FILL
X_8724_ _8724_/A gnd _8724_/Y vdd INVX1
XFILL_5__16298_ gnd vdd FILL
XFILL_3__13709_ gnd vdd FILL
XFILL_2__15138_ gnd vdd FILL
XSFILL114520x52050 gnd vdd FILL
XFILL_0__16317_ gnd vdd FILL
XSFILL44040x29050 gnd vdd FILL
XFILL_1__15868_ gnd vdd FILL
XFILL_3__14689_ gnd vdd FILL
XFILL_0__13529_ gnd vdd FILL
XFILL_5__15249_ gnd vdd FILL
X_8655_ _8655_/A _8655_/B _8655_/C gnd _8691_/D vdd OAI21X1
XFILL_4__15979_ gnd vdd FILL
XFILL_1__14819_ gnd vdd FILL
XFILL_2__15069_ gnd vdd FILL
XFILL_0__16248_ gnd vdd FILL
XFILL_6__9534_ gnd vdd FILL
XFILL_1__15799_ gnd vdd FILL
XFILL_1__8840_ gnd vdd FILL
X_7606_ _7606_/A _8630_/B gnd _7607_/C vdd NAND2X1
XFILL_3__16359_ gnd vdd FILL
XFILL_4_BUFX2_insert1003 gnd vdd FILL
X_8586_ _8584_/Y _8577_/B _8586_/C gnd _8668_/D vdd OAI21X1
XFILL_4_BUFX2_insert1014 gnd vdd FILL
XFILL_3__9756_ gnd vdd FILL
XFILL_3__6968_ gnd vdd FILL
XFILL_4_BUFX2_insert1025 gnd vdd FILL
XFILL_0__16179_ gnd vdd FILL
XFILL_4_BUFX2_insert1036 gnd vdd FILL
XFILL_4__7500_ gnd vdd FILL
X_7537_ _7495_/A _7537_/CLK _7537_/R vdd _7537_/D gnd vdd DFFSR
XFILL_1__8771_ gnd vdd FILL
XFILL_3__8707_ gnd vdd FILL
XFILL_4_BUFX2_insert1047 gnd vdd FILL
XFILL_0__9978_ gnd vdd FILL
XFILL_4__8480_ gnd vdd FILL
XFILL_4_BUFX2_insert1058 gnd vdd FILL
XFILL112440x16050 gnd vdd FILL
XFILL_3__6899_ gnd vdd FILL
XFILL_4_BUFX2_insert1069 gnd vdd FILL
XFILL_4_BUFX2_insert90 gnd vdd FILL
XFILL_1__7722_ gnd vdd FILL
XSFILL23720x51050 gnd vdd FILL
X_7468_ _7468_/A gnd _7470_/A vdd INVX1
XFILL_4__7431_ gnd vdd FILL
XFILL_3__8638_ gnd vdd FILL
X_9207_ _8183_/A _9208_/B gnd _9207_/Y vdd NAND2X1
XSFILL39000x18050 gnd vdd FILL
X_7399_ _7337_/A _7527_/CLK _8935_/R vdd _7399_/D gnd vdd DFFSR
XFILL_4__7362_ gnd vdd FILL
XFILL_3__8569_ gnd vdd FILL
XSFILL79400x23050 gnd vdd FILL
XSFILL3640x49050 gnd vdd FILL
XFILL_4__9101_ gnd vdd FILL
XFILL_3_BUFX2_insert303 gnd vdd FILL
X_9138_ _9194_/Q gnd _9140_/A vdd INVX1
XFILL_1__7584_ gnd vdd FILL
XFILL_3_BUFX2_insert314 gnd vdd FILL
XFILL_3_BUFX2_insert325 gnd vdd FILL
X_10020_ _9975_/B _8868_/B gnd _10021_/C vdd NAND2X1
XFILL_6__7229_ gnd vdd FILL
XFILL_3_BUFX2_insert336 gnd vdd FILL
XFILL_2_BUFX2_insert1040 gnd vdd FILL
XFILL_4__7293_ gnd vdd FILL
XSFILL114600x32050 gnd vdd FILL
XSFILL94280x37050 gnd vdd FILL
XFILL_2_BUFX2_insert1051 gnd vdd FILL
XFILL_3_BUFX2_insert347 gnd vdd FILL
X_9069_ _9069_/Q _8947_/CLK _9069_/R vdd _9069_/D gnd vdd DFFSR
XFILL_2_BUFX2_insert1062 gnd vdd FILL
XFILL_3_BUFX2_insert358 gnd vdd FILL
XFILL_4__9032_ gnd vdd FILL
XFILL_2_BUFX2_insert1073 gnd vdd FILL
XFILL_3_BUFX2_insert369 gnd vdd FILL
XFILL_2_BUFX2_insert1084 gnd vdd FILL
XSFILL54280x53050 gnd vdd FILL
XFILL_1__9254_ gnd vdd FILL
XFILL_1__8205_ gnd vdd FILL
X_11971_ _11971_/A gnd _11973_/A vdd INVX1
X_13710_ _7045_/A gnd _13710_/Y vdd INVX1
XSFILL104280x22050 gnd vdd FILL
X_10922_ _10922_/A _10944_/B gnd _10922_/Y vdd AND2X2
XFILL_1__8136_ gnd vdd FILL
X_14690_ _14690_/A _14690_/B _14687_/Y gnd _14691_/A vdd NAND3X1
XFILL_4__9934_ gnd vdd FILL
X_13641_ _9306_/Q gnd _13643_/A vdd INVX1
XSFILL8760x82050 gnd vdd FILL
X_10853_ _10853_/Q _7781_/CLK _8025_/R vdd _10789_/Y gnd vdd DFFSR
XFILL_1__8067_ gnd vdd FILL
XFILL_4_CLKBUF1_insert115 gnd vdd FILL
XFILL_4_CLKBUF1_insert126 gnd vdd FILL
XFILL_4__9865_ gnd vdd FILL
X_16360_ _14099_/A gnd _16362_/A vdd INVX1
XFILL_4_CLKBUF1_insert137 gnd vdd FILL
XFILL_4_CLKBUF1_insert148 gnd vdd FILL
X_13572_ _13572_/A gnd _15139_/D vdd INVX1
X_10784_ _14156_/A gnd _10786_/A vdd INVX1
XSFILL49240x42050 gnd vdd FILL
XFILL_2__8880_ gnd vdd FILL
XFILL_4_CLKBUF1_insert159 gnd vdd FILL
X_15311_ _15656_/B _15656_/C gnd _15380_/B vdd NOR2X1
XSFILL3720x29050 gnd vdd FILL
XFILL_0_BUFX2_insert226 gnd vdd FILL
X_12523_ _12427_/A gnd _12523_/Y vdd INVX1
XFILL_6_BUFX2_insert991 gnd vdd FILL
XFILL_4__9796_ gnd vdd FILL
X_16291_ _14934_/A _15940_/B _15569_/C _14974_/D gnd _16291_/Y vdd OAI22X1
XFILL_0_BUFX2_insert237 gnd vdd FILL
XFILL_2__7831_ gnd vdd FILL
XFILL_0_BUFX2_insert248 gnd vdd FILL
XFILL_0_BUFX2_insert259 gnd vdd FILL
XSFILL94360x17050 gnd vdd FILL
X_15242_ _15220_/B _14980_/Y gnd _15243_/B vdd NAND2X1
XFILL_4__8747_ gnd vdd FILL
X_12454_ _12454_/A gnd _12456_/A vdd INVX1
XSFILL13720x83050 gnd vdd FILL
XFILL_3__10370_ gnd vdd FILL
XFILL_2__7762_ gnd vdd FILL
XFILL_1__8969_ gnd vdd FILL
XFILL_0__10190_ gnd vdd FILL
XSFILL28520x43050 gnd vdd FILL
XFILL_5__7471_ gnd vdd FILL
X_11405_ _11623_/A _11623_/B _11404_/Y gnd _11411_/B vdd OAI21X1
XSFILL79160x78050 gnd vdd FILL
X_15173_ _15322_/D gnd _15652_/D vdd INVX8
X_12385_ _12385_/A gnd _12385_/Y vdd INVX1
XFILL_4__11660_ gnd vdd FILL
XFILL_2__9501_ gnd vdd FILL
XFILL_1__10500_ gnd vdd FILL
XFILL_2__7693_ gnd vdd FILL
XFILL_5__9210_ gnd vdd FILL
XFILL_4__7629_ gnd vdd FILL
X_14124_ _10016_/A gnd _14125_/D vdd INVX1
XFILL_1__11480_ gnd vdd FILL
XSFILL109400x5050 gnd vdd FILL
X_11336_ _11198_/Y _11199_/Y _11336_/C gnd _11337_/C vdd OAI21X1
XFILL_3__12040_ gnd vdd FILL
XFILL_2_BUFX2_insert19 gnd vdd FILL
XFILL_4__11591_ gnd vdd FILL
XFILL_5__9141_ gnd vdd FILL
XFILL_2__12770_ gnd vdd FILL
XFILL_1__10431_ gnd vdd FILL
XFILL_5__11901_ gnd vdd FILL
X_14055_ _14055_/A _14051_/Y gnd _14055_/Y vdd NOR2X1
XFILL_4__13330_ gnd vdd FILL
XSFILL84280x69050 gnd vdd FILL
XSFILL104600x64050 gnd vdd FILL
XFILL_4__10542_ gnd vdd FILL
X_11267_ _12254_/Y _12144_/Y gnd _11267_/Y vdd NOR2X1
XFILL_5__12881_ gnd vdd FILL
XFILL_2__9363_ gnd vdd FILL
XFILL_2__11721_ gnd vdd FILL
XFILL_1__13150_ gnd vdd FILL
XFILL_1__10362_ gnd vdd FILL
XFILL_0__12900_ gnd vdd FILL
X_13006_ vdd _13006_/B gnd _13007_/C vdd NAND2X1
XFILL_0__13880_ gnd vdd FILL
XFILL_5__14620_ gnd vdd FILL
X_10218_ _10162_/A _9578_/CLK _7153_/R vdd _10218_/D gnd vdd DFFSR
XFILL_4__13261_ gnd vdd FILL
XFILL_2__8314_ gnd vdd FILL
XFILL_5__11832_ gnd vdd FILL
XFILL_1__12101_ gnd vdd FILL
XSFILL59080x45050 gnd vdd FILL
XFILL_2__14440_ gnd vdd FILL
X_11198_ _12204_/Y gnd _11198_/Y vdd INVX2
XFILL_2__9294_ gnd vdd FILL
XFILL_2__11652_ gnd vdd FILL
XFILL_1__10293_ gnd vdd FILL
XFILL_1__13081_ gnd vdd FILL
XFILL_3__13991_ gnd vdd FILL
XSFILL99480x50050 gnd vdd FILL
XFILL_0__12831_ gnd vdd FILL
XFILL_6__15910_ gnd vdd FILL
XFILL_4__15000_ gnd vdd FILL
XFILL_3_BUFX2_insert870 gnd vdd FILL
XFILL_4__12212_ gnd vdd FILL
XFILL_5__14551_ gnd vdd FILL
X_10149_ _10147_/Y _10127_/A _10148_/Y gnd _10149_/Y vdd OAI21X1
XFILL_3_BUFX2_insert881 gnd vdd FILL
XFILL_2__8245_ gnd vdd FILL
XFILL_3__15730_ gnd vdd FILL
XFILL_5__11763_ gnd vdd FILL
XFILL_3_BUFX2_insert892 gnd vdd FILL
XFILL_1__12032_ gnd vdd FILL
XFILL_2__14371_ gnd vdd FILL
XFILL_0__15550_ gnd vdd FILL
XFILL_2__11583_ gnd vdd FILL
XFILL_0__12762_ gnd vdd FILL
XFILL_5__13502_ gnd vdd FILL
XFILL_2__16110_ gnd vdd FILL
XFILL_4__12143_ gnd vdd FILL
XFILL_2__13322_ gnd vdd FILL
XFILL_5__14482_ gnd vdd FILL
XSFILL53800x47050 gnd vdd FILL
X_14957_ _7669_/Q gnd _14959_/D vdd INVX1
XFILL_2__10534_ gnd vdd FILL
XFILL_3__15661_ gnd vdd FILL
XFILL_0__14501_ gnd vdd FILL
XFILL_3__12873_ gnd vdd FILL
XFILL_5__11694_ gnd vdd FILL
XFILL_0__11713_ gnd vdd FILL
XFILL_5__16221_ gnd vdd FILL
XFILL_0__15481_ gnd vdd FILL
XSFILL13800x63050 gnd vdd FILL
XFILL_5__9974_ gnd vdd FILL
XFILL_5__13433_ gnd vdd FILL
XFILL_6__15772_ gnd vdd FILL
X_13908_ _13908_/A _13908_/B gnd _13930_/B vdd NOR2X1
XFILL_3__14612_ gnd vdd FILL
XFILL_2__16041_ gnd vdd FILL
XFILL_4__12074_ gnd vdd FILL
XFILL_0__7191_ gnd vdd FILL
XFILL_5__10645_ gnd vdd FILL
XFILL_3__11824_ gnd vdd FILL
XFILL_2__13253_ gnd vdd FILL
X_14888_ _14888_/A _14887_/Y gnd _14891_/C vdd NOR2X1
XFILL_3__15592_ gnd vdd FILL
XFILL_0__14432_ gnd vdd FILL
XFILL_1__13983_ gnd vdd FILL
XFILL_6__14723_ gnd vdd FILL
XFILL_0__11644_ gnd vdd FILL
XFILL_4__15902_ gnd vdd FILL
XFILL_4__11025_ gnd vdd FILL
XFILL_5__16152_ gnd vdd FILL
XFILL_5__13364_ gnd vdd FILL
X_13839_ _13839_/A _13839_/B gnd _13840_/B vdd NOR2X1
XFILL_2__12204_ gnd vdd FILL
XFILL_1__15722_ gnd vdd FILL
XFILL_3__7940_ gnd vdd FILL
XFILL_3__14543_ gnd vdd FILL
XFILL_2__7058_ gnd vdd FILL
XFILL_3__11755_ gnd vdd FILL
XFILL_5__10576_ gnd vdd FILL
XFILL_2__10396_ gnd vdd FILL
XFILL_0__14363_ gnd vdd FILL
XFILL_0__11575_ gnd vdd FILL
XFILL_5__15103_ gnd vdd FILL
XSFILL114440x67050 gnd vdd FILL
XFILL_5__8856_ gnd vdd FILL
XFILL_5__12315_ gnd vdd FILL
XFILL_4__15833_ gnd vdd FILL
XFILL_5__16083_ gnd vdd FILL
XFILL_3__10706_ gnd vdd FILL
XFILL_5__13295_ gnd vdd FILL
XFILL_3__14474_ gnd vdd FILL
XFILL_2__12135_ gnd vdd FILL
XFILL_0__16102_ gnd vdd FILL
XFILL_0__13314_ gnd vdd FILL
XFILL_3__7871_ gnd vdd FILL
XFILL_1__15653_ gnd vdd FILL
XFILL_3__11686_ gnd vdd FILL
XFILL_0__10526_ gnd vdd FILL
XFILL_5__7807_ gnd vdd FILL
XFILL_1__12865_ gnd vdd FILL
X_15509_ _15509_/A _15357_/B _16166_/A _15509_/D gnd _15509_/Y vdd AOI22X1
XFILL_5__15034_ gnd vdd FILL
XFILL_6__7580_ gnd vdd FILL
XFILL_0__14294_ gnd vdd FILL
XFILL_0__9901_ gnd vdd FILL
XFILL_3__16213_ gnd vdd FILL
XFILL_6__14585_ gnd vdd FILL
XFILL_3__13425_ gnd vdd FILL
XFILL_5_BUFX2_insert409 gnd vdd FILL
X_8440_ _8438_/Y _8440_/B _8439_/Y gnd _8534_/D vdd OAI21X1
XFILL_5__12246_ gnd vdd FILL
XFILL_5__8787_ gnd vdd FILL
XFILL_3__10637_ gnd vdd FILL
XFILL_3__9610_ gnd vdd FILL
XFILL_1__14604_ gnd vdd FILL
XFILL_4__15764_ gnd vdd FILL
XFILL_4__12976_ gnd vdd FILL
XFILL_0__16033_ gnd vdd FILL
XFILL_2__12066_ gnd vdd FILL
XFILL_1__11816_ gnd vdd FILL
XFILL_0__13245_ gnd vdd FILL
XFILL_6__16324_ gnd vdd FILL
XFILL_1__15584_ gnd vdd FILL
XSFILL59160x25050 gnd vdd FILL
XFILL_0_BUFX2_insert760 gnd vdd FILL
XFILL_5__7738_ gnd vdd FILL
XFILL_6__13536_ gnd vdd FILL
XFILL_0_BUFX2_insert771 gnd vdd FILL
XFILL_4__14715_ gnd vdd FILL
XFILL_3__13356_ gnd vdd FILL
XFILL_0_BUFX2_insert782 gnd vdd FILL
XFILL_4__11927_ gnd vdd FILL
X_8371_ _8372_/B _8243_/B gnd _8372_/C vdd NAND2X1
XFILL_5__12177_ gnd vdd FILL
XFILL_2__11017_ gnd vdd FILL
XFILL_3__16144_ gnd vdd FILL
XFILL_4__15695_ gnd vdd FILL
XFILL_1__14535_ gnd vdd FILL
XFILL_3__9541_ gnd vdd FILL
XFILL_3__10568_ gnd vdd FILL
XFILL_0_BUFX2_insert793 gnd vdd FILL
XFILL_1__11747_ gnd vdd FILL
XFILL_6__9250_ gnd vdd FILL
XFILL_0__10388_ gnd vdd FILL
XFILL_0__9763_ gnd vdd FILL
X_7322_ _7394_/Q gnd _7322_/Y vdd INVX1
XFILL_3__12307_ gnd vdd FILL
XFILL_5__11128_ gnd vdd FILL
XFILL_0__6975_ gnd vdd FILL
XFILL_4__14646_ gnd vdd FILL
XFILL_3__16075_ gnd vdd FILL
XFILL_3__9472_ gnd vdd FILL
XFILL_3__13287_ gnd vdd FILL
XFILL_0__12127_ gnd vdd FILL
XFILL_2__15825_ gnd vdd FILL
XFILL_4__11858_ gnd vdd FILL
XFILL_1__14466_ gnd vdd FILL
XFILL_5__9408_ gnd vdd FILL
XFILL_6__8201_ gnd vdd FILL
XFILL_3__10499_ gnd vdd FILL
XFILL_0__8714_ gnd vdd FILL
XFILL_6__12418_ gnd vdd FILL
XFILL_1__11678_ gnd vdd FILL
XFILL_6__16186_ gnd vdd FILL
XFILL_3__15026_ gnd vdd FILL
XFILL_5__15936_ gnd vdd FILL
XFILL_1__16205_ gnd vdd FILL
XFILL_6__13398_ gnd vdd FILL
XFILL_4__10809_ gnd vdd FILL
XFILL_3__12238_ gnd vdd FILL
XFILL_5__11059_ gnd vdd FILL
X_7253_ _7253_/A _7210_/A _7253_/C gnd _7285_/D vdd OAI21X1
XFILL_4__14577_ gnd vdd FILL
XSFILL109400x56050 gnd vdd FILL
XFILL_1__13417_ gnd vdd FILL
XFILL_0__12058_ gnd vdd FILL
XFILL_1__10629_ gnd vdd FILL
XFILL_4__11789_ gnd vdd FILL
XFILL_2__15756_ gnd vdd FILL
XFILL_2__12968_ gnd vdd FILL
XFILL_1__14397_ gnd vdd FILL
XFILL_6__15137_ gnd vdd FILL
XFILL_5__9339_ gnd vdd FILL
XFILL_0__8645_ gnd vdd FILL
XSFILL79320x38050 gnd vdd FILL
XFILL_4__16316_ gnd vdd FILL
X_7184_ _7182_/Y _7184_/B _7183_/Y gnd _7184_/Y vdd OAI21X1
XFILL_5__15867_ gnd vdd FILL
XFILL_4__13528_ gnd vdd FILL
XFILL_3__8354_ gnd vdd FILL
XFILL_2__14707_ gnd vdd FILL
XFILL_2__11919_ gnd vdd FILL
XFILL_3__12169_ gnd vdd FILL
XFILL_1__16136_ gnd vdd FILL
XFILL_0__11009_ gnd vdd FILL
XFILL_1__13348_ gnd vdd FILL
XFILL_2__15687_ gnd vdd FILL
XFILL_2__12899_ gnd vdd FILL
XFILL_5__14818_ gnd vdd FILL
XFILL_0__8576_ gnd vdd FILL
XFILL_3__7305_ gnd vdd FILL
XFILL_4__16247_ gnd vdd FILL
XFILL_2__14638_ gnd vdd FILL
XFILL_4__13459_ gnd vdd FILL
XFILL_5__15798_ gnd vdd FILL
XFILL_0__15817_ gnd vdd FILL
XFILL_1__16067_ gnd vdd FILL
XFILL_1__13279_ gnd vdd FILL
XFILL_5__14749_ gnd vdd FILL
XFILL_3__15928_ gnd vdd FILL
XFILL_4__16178_ gnd vdd FILL
XFILL_3__7236_ gnd vdd FILL
XFILL_1__15018_ gnd vdd FILL
XFILL_1_BUFX2_insert5 gnd vdd FILL
XFILL_2__14569_ gnd vdd FILL
XFILL_0__15748_ gnd vdd FILL
XFILL_0__7458_ gnd vdd FILL
XFILL_4__15129_ gnd vdd FILL
XFILL_2__16308_ gnd vdd FILL
XFILL_3__7167_ gnd vdd FILL
XFILL_3__15859_ gnd vdd FILL
XFILL_0__15679_ gnd vdd FILL
X_9825_ _9751_/A _9188_/CLK _9441_/R vdd _9825_/D gnd vdd DFFSR
XFILL_2__16239_ gnd vdd FILL
XFILL_3__7098_ gnd vdd FILL
XFILL_0__9128_ gnd vdd FILL
XFILL_4__7980_ gnd vdd FILL
X_9756_ _9756_/A _9737_/A _9755_/Y gnd _9826_/D vdd OAI21X1
XSFILL23720x46050 gnd vdd FILL
X_6968_ _7020_/Q gnd _6968_/Y vdd INVX1
XFILL_4__6931_ gnd vdd FILL
X_8707_ _8765_/B _9475_/B gnd _8708_/C vdd NAND2X1
XFILL112040x13050 gnd vdd FILL
XFILL_6_BUFX2_insert254 gnd vdd FILL
XBUFX2_insert309 _11222_/Y gnd _11764_/D vdd BUFX2
XFILL_1__9941_ gnd vdd FILL
XFILL_6_BUFX2_insert265 gnd vdd FILL
X_9687_ _9593_/A _7143_/CLK _7131_/R vdd _9687_/D gnd vdd DFFSR
XFILL_4__6862_ gnd vdd FILL
X_6899_ _6899_/A gnd memoryWriteData[29] vdd BUFX2
XFILL_4__9650_ gnd vdd FILL
X_8638_ _8638_/A gnd _8638_/Y vdd INVX1
XFILL_1__9872_ gnd vdd FILL
XFILL_5_BUFX2_insert910 gnd vdd FILL
XFILL_4__8601_ gnd vdd FILL
XFILL_3__9808_ gnd vdd FILL
XFILL_5_BUFX2_insert921 gnd vdd FILL
XFILL_5_BUFX2_insert932 gnd vdd FILL
XFILL_5_BUFX2_insert943 gnd vdd FILL
XFILL_1__8823_ gnd vdd FILL
XSFILL114600x27050 gnd vdd FILL
XFILL_5_BUFX2_insert954 gnd vdd FILL
X_8569_ _8663_/Q gnd _8571_/A vdd INVX1
XFILL_5_BUFX2_insert965 gnd vdd FILL
XFILL_3__9739_ gnd vdd FILL
XFILL_4__8532_ gnd vdd FILL
XFILL_5_BUFX2_insert976 gnd vdd FILL
XFILL_5_BUFX2_insert987 gnd vdd FILL
XFILL_5_BUFX2_insert998 gnd vdd FILL
XFILL_1__8754_ gnd vdd FILL
XFILL_4__8463_ gnd vdd FILL
XSFILL94680x53050 gnd vdd FILL
XFILL_1__7705_ gnd vdd FILL
X_12170_ _12150_/B _12170_/B gnd _12171_/C vdd NAND2X1
XFILL_6__9379_ gnd vdd FILL
XFILL_4__7414_ gnd vdd FILL
XFILL_4__8394_ gnd vdd FILL
X_11121_ _12171_/Y _12290_/Y gnd _11121_/Y vdd NAND2X1
XFILL_1__7636_ gnd vdd FILL
XFILL_3_BUFX2_insert100 gnd vdd FILL
XFILL_4__7345_ gnd vdd FILL
X_11052_ _12262_/Y _12150_/Y gnd _11054_/A vdd XOR2X1
XSFILL8760x77050 gnd vdd FILL
XFILL_1__7567_ gnd vdd FILL
XSFILL33960x70050 gnd vdd FILL
X_10003_ _10001_/Y _10054_/B _10002_/Y gnd _10079_/D vdd OAI21X1
X_15860_ _15860_/A _15860_/B _15860_/C gnd _15860_/Y vdd NAND3X1
XFILL_4__9015_ gnd vdd FILL
XFILL_2_BUFX2_insert800 gnd vdd FILL
XFILL_1__7498_ gnd vdd FILL
XFILL_2_BUFX2_insert811 gnd vdd FILL
X_14811_ _14802_/Y _14803_/Y _14811_/C gnd _14812_/B vdd NAND3X1
XSFILL90120x30050 gnd vdd FILL
XFILL_2_BUFX2_insert822 gnd vdd FILL
XFILL_2_BUFX2_insert833 gnd vdd FILL
XFILL_1__9237_ gnd vdd FILL
X_15791_ _10412_/A gnd _15791_/Y vdd INVX1
XFILL_2_BUFX2_insert844 gnd vdd FILL
XFILL_2_BUFX2_insert855 gnd vdd FILL
XFILL_2_BUFX2_insert866 gnd vdd FILL
X_11954_ _11955_/B _12409_/A gnd _11954_/Y vdd NAND2X1
XFILL_2_BUFX2_insert877 gnd vdd FILL
X_14742_ _14742_/A _14741_/Y _15651_/C gnd _13030_/B vdd AOI21X1
XSFILL74280x6050 gnd vdd FILL
XFILL_2_BUFX2_insert888 gnd vdd FILL
XFILL_1__9168_ gnd vdd FILL
XFILL_2_BUFX2_insert899 gnd vdd FILL
XSFILL54360x28050 gnd vdd FILL
X_10905_ _10987_/Q gnd _10910_/B vdd INVX2
XFILL_5__6971_ gnd vdd FILL
XFILL_1__8119_ gnd vdd FILL
XFILL_5__10430_ gnd vdd FILL
X_14673_ _9711_/Q gnd _14675_/A vdd INVX1
X_11885_ _11874_/B _11885_/B gnd _11885_/Y vdd NAND2X1
XFILL_1__9099_ gnd vdd FILL
XFILL_2__10250_ gnd vdd FILL
XFILL_4__9917_ gnd vdd FILL
XFILL_5__8710_ gnd vdd FILL
XFILL_2__9981_ gnd vdd FILL
XFILL_1__10980_ gnd vdd FILL
X_13624_ _13623_/Y _14593_/C gnd _13625_/C vdd NOR2X1
X_16412_ gnd gnd gnd _16412_/Y vdd NAND2X1
XFILL112040x6050 gnd vdd FILL
XFILL_5__10361_ gnd vdd FILL
X_10836_ _10797_/A _7380_/B gnd _10837_/C vdd NAND2X1
XFILL_3__11540_ gnd vdd FILL
XFILL_4_BUFX2_insert9 gnd vdd FILL
XFILL_2__10181_ gnd vdd FILL
XBUFX2_insert810 _13329_/Y gnd _9011_/A vdd BUFX2
XFILL_0__11360_ gnd vdd FILL
XFILL_5__12100_ gnd vdd FILL
XFILL_4__9848_ gnd vdd FILL
XFILL_5__8641_ gnd vdd FILL
XBUFX2_insert821 _12384_/Y gnd _9374_/B vdd BUFX2
X_16343_ gnd gnd gnd _16343_/Y vdd NAND2X1
XFILL_6__11651_ gnd vdd FILL
X_13555_ _9596_/A gnd _15132_/D vdd INVX1
X_10767_ _10789_/B _8207_/B gnd _10768_/C vdd NAND2X1
XFILL_5__13080_ gnd vdd FILL
XBUFX2_insert832 _15046_/Y gnd _15170_/D vdd BUFX2
XFILL_4__12830_ gnd vdd FILL
XFILL_5__10292_ gnd vdd FILL
XFILL_0__10311_ gnd vdd FILL
XBUFX2_insert843 _12375_/Y gnd _6933_/B vdd BUFX2
XFILL_3__11471_ gnd vdd FILL
XFILL_1__12650_ gnd vdd FILL
XBUFX2_insert854 _13269_/Y gnd _7095_/B vdd BUFX2
XFILL_2__8863_ gnd vdd FILL
X_12506_ vdd _12077_/A gnd _12506_/Y vdd NAND2X1
XFILL_0__11291_ gnd vdd FILL
XBUFX2_insert865 _13438_/Y gnd _14323_/B vdd BUFX2
XFILL_3__13210_ gnd vdd FILL
XFILL_5__12031_ gnd vdd FILL
XBUFX2_insert876 _15019_/Y gnd _15948_/D vdd BUFX2
XFILL_6__14370_ gnd vdd FILL
XFILL_5__8572_ gnd vdd FILL
X_16274_ _8436_/Q gnd _16276_/A vdd INVX1
XFILL_4__9779_ gnd vdd FILL
XFILL_3__10422_ gnd vdd FILL
X_13486_ _14555_/C gnd _13486_/Y vdd INVX8
XFILL_4__12761_ gnd vdd FILL
XFILL_3__14190_ gnd vdd FILL
X_10698_ _10738_/Q gnd _10700_/A vdd INVX1
XBUFX2_insert887 _13432_/Y gnd _13846_/A vdd BUFX2
XFILL_0__13030_ gnd vdd FILL
XFILL_1__11601_ gnd vdd FILL
XFILL_2__7814_ gnd vdd FILL
XFILL_2__13940_ gnd vdd FILL
XSFILL104200x61050 gnd vdd FILL
XBUFX2_insert898 _13470_/Y gnd _14643_/B vdd BUFX2
XFILL_0__10242_ gnd vdd FILL
XFILL_6__13321_ gnd vdd FILL
XFILL_1__12581_ gnd vdd FILL
X_15225_ _15225_/A _7554_/A _7514_/Q _15383_/D gnd _15225_/Y vdd AOI22X1
X_12437_ _12407_/A _12694_/Q gnd _12438_/C vdd NAND2X1
XFILL_4__14500_ gnd vdd FILL
XFILL_3__13141_ gnd vdd FILL
XSFILL74120x43050 gnd vdd FILL
XFILL_4__11712_ gnd vdd FILL
XFILL_1__14320_ gnd vdd FILL
XFILL_2__7745_ gnd vdd FILL
XFILL_4__15480_ gnd vdd FILL
XFILL_2__13871_ gnd vdd FILL
XFILL_1__11532_ gnd vdd FILL
XFILL_0__10173_ gnd vdd FILL
XFILL_5__7454_ gnd vdd FILL
X_15156_ _15156_/A _15156_/B gnd _15166_/A vdd NAND2X1
X_12368_ _12368_/A _12591_/A gnd _12369_/C vdd NAND2X1
XSFILL109880x28050 gnd vdd FILL
XFILL_4__14431_ gnd vdd FILL
XFILL_5__13982_ gnd vdd FILL
XFILL_4__11643_ gnd vdd FILL
XFILL_2__15610_ gnd vdd FILL
XFILL_1__14251_ gnd vdd FILL
XFILL_3__10284_ gnd vdd FILL
XFILL_2__7676_ gnd vdd FILL
XFILL_6__12203_ gnd vdd FILL
X_14107_ _8035_/Q gnd _15599_/D vdd INVX1
XFILL_1__11463_ gnd vdd FILL
XFILL_5__15721_ gnd vdd FILL
XFILL_0__14981_ gnd vdd FILL
X_11319_ _11173_/Y _11195_/A gnd _11461_/A vdd NOR2X1
XFILL_3__12023_ gnd vdd FILL
X_15087_ _7639_/Q _15087_/B gnd _15094_/A vdd NAND2X1
XFILL_2__15541_ gnd vdd FILL
XFILL_2__9415_ gnd vdd FILL
XFILL_4__14362_ gnd vdd FILL
X_12299_ _12216_/A gnd _12311_/C gnd _12302_/A vdd NAND3X1
XFILL_4__11574_ gnd vdd FILL
XFILL_2__12753_ gnd vdd FILL
XFILL_1__10414_ gnd vdd FILL
XFILL_5__9124_ gnd vdd FILL
XFILL_1__14182_ gnd vdd FILL
XFILL_0__13932_ gnd vdd FILL
X_14038_ _15566_/A _14868_/A _13771_/D _8474_/A gnd _14047_/B vdd AOI22X1
XFILL_4__16101_ gnd vdd FILL
XFILL_1__11394_ gnd vdd FILL
XFILL_4__13313_ gnd vdd FILL
XFILL_5__15652_ gnd vdd FILL
XFILL_2__9346_ gnd vdd FILL
XFILL_2__11704_ gnd vdd FILL
XFILL_4__10525_ gnd vdd FILL
XFILL_5__12864_ gnd vdd FILL
XFILL_1__13133_ gnd vdd FILL
XSFILL54040x10050 gnd vdd FILL
XFILL_2__15472_ gnd vdd FILL
XFILL_4__14293_ gnd vdd FILL
XFILL_0__13863_ gnd vdd FILL
XFILL_5__14603_ gnd vdd FILL
XFILL_4__16032_ gnd vdd FILL
XFILL_6__12065_ gnd vdd FILL
XFILL_0__8361_ gnd vdd FILL
XFILL_5__11815_ gnd vdd FILL
XFILL_4__13244_ gnd vdd FILL
XFILL_5__15583_ gnd vdd FILL
XFILL_2__14423_ gnd vdd FILL
XFILL_2__9277_ gnd vdd FILL
XFILL_3__8070_ gnd vdd FILL
XFILL_2__11635_ gnd vdd FILL
XFILL_0__15602_ gnd vdd FILL
XFILL_1__10276_ gnd vdd FILL
XFILL_5__8006_ gnd vdd FILL
XFILL_3__13974_ gnd vdd FILL
XFILL_0__7312_ gnd vdd FILL
XFILL_6__11016_ gnd vdd FILL
XFILL_0__13794_ gnd vdd FILL
XFILL_5__14534_ gnd vdd FILL
XFILL_2__8228_ gnd vdd FILL
XFILL_3__15713_ gnd vdd FILL
X_7940_ _7938_/Y _7970_/B _7940_/C gnd _8026_/D vdd OAI21X1
XFILL_5__11746_ gnd vdd FILL
X_15989_ _9325_/Q gnd _15989_/Y vdd INVX1
XFILL_1__12015_ gnd vdd FILL
XSFILL43880x53050 gnd vdd FILL
XFILL_2__14354_ gnd vdd FILL
XFILL_4__10387_ gnd vdd FILL
XFILL_0__15533_ gnd vdd FILL
XFILL_2__11566_ gnd vdd FILL
XFILL_0__12745_ gnd vdd FILL
XFILL_0__7243_ gnd vdd FILL
XFILL_2__13305_ gnd vdd FILL
XFILL_5__14465_ gnd vdd FILL
XFILL_4__12126_ gnd vdd FILL
X_7871_ _7872_/B _7743_/B gnd _7871_/Y vdd NAND2X1
XFILL_3__15644_ gnd vdd FILL
XFILL_5__11677_ gnd vdd FILL
XFILL_2__10517_ gnd vdd FILL
XSFILL99560x25050 gnd vdd FILL
XFILL_3__12856_ gnd vdd FILL
XFILL_2__14285_ gnd vdd FILL
XFILL_5__16204_ gnd vdd FILL
XFILL_0__15464_ gnd vdd FILL
XFILL_2__11497_ gnd vdd FILL
XSFILL74200x23050 gnd vdd FILL
X_9610_ _9608_/Y _9615_/A _9610_/C gnd _9692_/D vdd OAI21X1
XFILL_5__13416_ gnd vdd FILL
XFILL_2__16024_ gnd vdd FILL
XFILL_5__10628_ gnd vdd FILL
XFILL_4__12057_ gnd vdd FILL
XFILL_0__7174_ gnd vdd FILL
XFILL_2__13236_ gnd vdd FILL
XFILL_5__14396_ gnd vdd FILL
XFILL_3__11807_ gnd vdd FILL
XFILL_3__12787_ gnd vdd FILL
XFILL_2__10448_ gnd vdd FILL
XFILL_3__15575_ gnd vdd FILL
XFILL_0__14415_ gnd vdd FILL
XFILL_3__8972_ gnd vdd FILL
XFILL_5__8908_ gnd vdd FILL
XFILL_0__11627_ gnd vdd FILL
XFILL_1__13966_ gnd vdd FILL
XFILL_0__15395_ gnd vdd FILL
XFILL_5__16135_ gnd vdd FILL
XFILL_4__11008_ gnd vdd FILL
XFILL_5__13347_ gnd vdd FILL
XFILL_5__9888_ gnd vdd FILL
X_9541_ _9529_/A _7877_/B gnd _9542_/C vdd NAND2X1
XFILL_5__10559_ gnd vdd FILL
XFILL_3__14526_ gnd vdd FILL
XFILL_6__12898_ gnd vdd FILL
XFILL_1__15705_ gnd vdd FILL
XFILL_2__13167_ gnd vdd FILL
XFILL_1__12917_ gnd vdd FILL
XFILL_3__11738_ gnd vdd FILL
XFILL_2__10379_ gnd vdd FILL
XFILL_0__14346_ gnd vdd FILL
XFILL_5__8839_ gnd vdd FILL
XFILL_1__13897_ gnd vdd FILL
XFILL_0__11558_ gnd vdd FILL
XFILL_6__7632_ gnd vdd FILL
XFILL_4__15816_ gnd vdd FILL
XSFILL109560x10050 gnd vdd FILL
XFILL_5__16066_ gnd vdd FILL
X_9472_ _9548_/B _8576_/B gnd _9472_/Y vdd NAND2X1
XFILL_5__13278_ gnd vdd FILL
XFILL_2__12118_ gnd vdd FILL
XFILL_3__14457_ gnd vdd FILL
XFILL_1__15636_ gnd vdd FILL
XFILL_3__11669_ gnd vdd FILL
XFILL_0__10509_ gnd vdd FILL
XFILL_1__12848_ gnd vdd FILL
XFILL_2__13098_ gnd vdd FILL
XFILL_3__7854_ gnd vdd FILL
XSFILL38040x23050 gnd vdd FILL
XFILL_5_BUFX2_insert228 gnd vdd FILL
XFILL_5__15017_ gnd vdd FILL
XFILL_0__11489_ gnd vdd FILL
XFILL_0__14277_ gnd vdd FILL
XFILL_5_BUFX2_insert239 gnd vdd FILL
XFILL_5__12229_ gnd vdd FILL
X_8423_ _8423_/Q _7016_/CLK _9064_/R vdd _8423_/D gnd vdd DFFSR
XFILL_3__13408_ gnd vdd FILL
XFILL_4__15747_ gnd vdd FILL
XFILL_0__16016_ gnd vdd FILL
XFILL_2__12049_ gnd vdd FILL
XFILL_4__12959_ gnd vdd FILL
XFILL_0__13228_ gnd vdd FILL
XFILL_1__15567_ gnd vdd FILL
XFILL_3__14388_ gnd vdd FILL
XFILL_1__12779_ gnd vdd FILL
XFILL_0_BUFX2_insert590 gnd vdd FILL
X_8354_ _8354_/A _8333_/B _8354_/C gnd _8354_/Y vdd OAI21X1
XFILL_3__16127_ gnd vdd FILL
XFILL_4_BUFX2_insert906 gnd vdd FILL
XFILL_3__13339_ gnd vdd FILL
XFILL_4__15678_ gnd vdd FILL
XFILL_1__14518_ gnd vdd FILL
XFILL_3__9524_ gnd vdd FILL
XFILL_4_BUFX2_insert917 gnd vdd FILL
XFILL_1__15498_ gnd vdd FILL
XFILL_0__13159_ gnd vdd FILL
XFILL_4_BUFX2_insert928 gnd vdd FILL
X_7305_ _7359_/A _6921_/B gnd _7305_/Y vdd NAND2X1
XFILL_4_BUFX2_insert939 gnd vdd FILL
XFILL_4__14629_ gnd vdd FILL
XFILL_0__6958_ gnd vdd FILL
XFILL_0__9746_ gnd vdd FILL
X_8285_ _8203_/A _7389_/CLK _8285_/R vdd _8205_/Y gnd vdd DFFSR
XFILL_2__15808_ gnd vdd FILL
XSFILL69080x7050 gnd vdd FILL
XFILL_3__16058_ gnd vdd FILL
XFILL_1__14449_ gnd vdd FILL
XFILL_0__9677_ gnd vdd FILL
XFILL_5__15919_ gnd vdd FILL
X_7236_ _7236_/A gnd _7238_/A vdd INVX1
XFILL_3__15009_ gnd vdd FILL
XFILL_1__8470_ gnd vdd FILL
XFILL_0__6889_ gnd vdd FILL
XSFILL68360x80050 gnd vdd FILL
XFILL_2__15739_ gnd vdd FILL
XFILL_3__9386_ gnd vdd FILL
XFILL_6__9095_ gnd vdd FILL
XFILL_1__7421_ gnd vdd FILL
XFILL_0__8628_ gnd vdd FILL
X_7167_ _7167_/A gnd _7169_/A vdd INVX1
XFILL_1__16119_ gnd vdd FILL
XFILL_3__8337_ gnd vdd FILL
XSFILL84280x1050 gnd vdd FILL
XFILL_1__7352_ gnd vdd FILL
XSFILL33080x66050 gnd vdd FILL
X_7098_ _7096_/Y _7068_/B _7098_/C gnd _7098_/Y vdd OAI21X1
XFILL_3__8268_ gnd vdd FILL
XFILL_2_BUFX2_insert107 gnd vdd FILL
XSFILL18840x9050 gnd vdd FILL
XFILL_4__7061_ gnd vdd FILL
XFILL_3__7219_ gnd vdd FILL
XSFILL38920x22050 gnd vdd FILL
XFILL_3__8199_ gnd vdd FILL
XFILL_1__9022_ gnd vdd FILL
XSFILL79000x15050 gnd vdd FILL
XSFILL24200x71050 gnd vdd FILL
XFILL_1_BUFX2_insert807 gnd vdd FILL
XSFILL39000x31050 gnd vdd FILL
XFILL_1_BUFX2_insert818 gnd vdd FILL
XFILL_1_BUFX2_insert829 gnd vdd FILL
X_9808_ _9844_/Q gnd _9808_/Y vdd INVX1
XFILL_4__7963_ gnd vdd FILL
X_11670_ _11669_/Y _11670_/B gnd _11673_/C vdd NOR2X1
X_9739_ _9821_/Q gnd _9741_/A vdd INVX1
XFILL_4__6914_ gnd vdd FILL
XBUFX2_insert106 _10925_/Y gnd _11921_/A vdd BUFX2
XSFILL28840x74050 gnd vdd FILL
X_10621_ _10619_/B _7037_/B gnd _10621_/Y vdd NAND2X1
XSFILL94280x50050 gnd vdd FILL
XFILL_1__9924_ gnd vdd FILL
XFILL_4__9633_ gnd vdd FILL
X_13340_ _13326_/A _13339_/Y gnd _13340_/Y vdd NOR2X1
XFILL_4__6845_ gnd vdd FILL
X_10552_ _10552_/A gnd _10552_/Y vdd INVX1
XFILL_1__9855_ gnd vdd FILL
XFILL_5_BUFX2_insert740 gnd vdd FILL
XFILL_5_BUFX2_insert751 gnd vdd FILL
XFILL_5_BUFX2_insert762 gnd vdd FILL
X_13271_ _13222_/B gnd _13283_/A vdd INVX2
XFILL_5_BUFX2_insert773 gnd vdd FILL
X_10483_ _10483_/Q _7021_/CLK _9062_/R vdd _10483_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert784 gnd vdd FILL
XFILL_5_BUFX2_insert795 gnd vdd FILL
XFILL_1__9786_ gnd vdd FILL
X_15010_ _15010_/A gnd _15969_/C vdd INVX8
XFILL_4__8515_ gnd vdd FILL
X_12222_ _12219_/Y _12222_/B _12222_/C gnd _12222_/Y vdd NAND3X1
XFILL_4__9495_ gnd vdd FILL
XFILL_1__8737_ gnd vdd FILL
XFILL_4__8446_ gnd vdd FILL
X_12153_ _12153_/A _12150_/B _12153_/C gnd _12153_/Y vdd OAI21X1
XFILL_2__7461_ gnd vdd FILL
XFILL_4__8377_ gnd vdd FILL
XFILL_5__7170_ gnd vdd FILL
X_11104_ _11102_/Y _11103_/Y gnd _11529_/A vdd NOR2X1
X_12084_ _12084_/A _12813_/Q _12084_/C gnd _12084_/Y vdd NAND3X1
XFILL_1__7619_ gnd vdd FILL
XFILL_1__8599_ gnd vdd FILL
XSFILL3720x42050 gnd vdd FILL
XFILL_4__7328_ gnd vdd FILL
X_15912_ _16002_/C _14461_/Y _14464_/Y _15912_/D gnd _15912_/Y vdd OAI22X1
XFILL_4__10310_ gnd vdd FILL
X_11035_ _11384_/A _12138_/Y gnd _11035_/Y vdd XNOR2X1
XFILL_2__9131_ gnd vdd FILL
XSFILL28920x54050 gnd vdd FILL
XFILL_4__11290_ gnd vdd FILL
XFILL_1__10130_ gnd vdd FILL
XFILL_5__11600_ gnd vdd FILL
XFILL_4__10241_ gnd vdd FILL
X_15843_ _15843_/A _15841_/Y gnd _15843_/Y vdd NOR2X1
XFILL_5__12580_ gnd vdd FILL
XFILL_2__11420_ gnd vdd FILL
XFILL_3__10971_ gnd vdd FILL
XFILL_1__10061_ gnd vdd FILL
XFILL_2_BUFX2_insert630 gnd vdd FILL
XFILL_2_BUFX2_insert641 gnd vdd FILL
XFILL_2_BUFX2_insert652 gnd vdd FILL
XFILL_0__10791_ gnd vdd FILL
XFILL_2__8013_ gnd vdd FILL
XFILL_5__11531_ gnd vdd FILL
XFILL_2_BUFX2_insert663 gnd vdd FILL
XFILL_4__10172_ gnd vdd FILL
XFILL_3__12710_ gnd vdd FILL
X_12986_ _12984_/Y vdd _12986_/C gnd _13058_/D vdd OAI21X1
X_15774_ _15563_/A _15773_/Y _15774_/C _14318_/Y gnd _15774_/Y vdd OAI22X1
XFILL_2_BUFX2_insert674 gnd vdd FILL
XFILL_3__13690_ gnd vdd FILL
XFILL_2__11351_ gnd vdd FILL
XFILL_2_BUFX2_insert685 gnd vdd FILL
XFILL_0__12530_ gnd vdd FILL
XFILL_5__9811_ gnd vdd FILL
XFILL_2_BUFX2_insert696 gnd vdd FILL
XFILL_5__14250_ gnd vdd FILL
X_14725_ _14725_/A _14725_/B _14725_/C _13824_/B gnd _14729_/A vdd OAI22X1
XFILL_2__10302_ gnd vdd FILL
XFILL_3__12641_ gnd vdd FILL
X_11937_ _11937_/A _11934_/B _11937_/C gnd _6854_/A vdd OAI21X1
XFILL_5__11462_ gnd vdd FILL
XFILL_1__13820_ gnd vdd FILL
XFILL_4__14980_ gnd vdd FILL
XFILL_2__14070_ gnd vdd FILL
XSFILL74120x38050 gnd vdd FILL
XFILL_2__11282_ gnd vdd FILL
XFILL_5__9742_ gnd vdd FILL
XFILL_0__12461_ gnd vdd FILL
XSFILL84280x82050 gnd vdd FILL
XFILL_5_BUFX2_insert12 gnd vdd FILL
XFILL_5__10413_ gnd vdd FILL
XFILL_5__6954_ gnd vdd FILL
XFILL_2__13021_ gnd vdd FILL
XFILL_5__14181_ gnd vdd FILL
X_11868_ _11866_/Y _11868_/B gnd _11868_/Y vdd AND2X2
X_14656_ _10305_/A _13621_/B _14283_/C _9967_/Q gnd _14657_/B vdd AOI22X1
XFILL_4__13931_ gnd vdd FILL
XFILL_0__14200_ gnd vdd FILL
XFILL_3__15360_ gnd vdd FILL
XFILL_3__12572_ gnd vdd FILL
XFILL_5__11393_ gnd vdd FILL
XFILL_2__10233_ gnd vdd FILL
XFILL_5_BUFX2_insert23 gnd vdd FILL
XFILL_5_BUFX2_insert34 gnd vdd FILL
XFILL_1__13751_ gnd vdd FILL
XFILL_0__11412_ gnd vdd FILL
XFILL_0__15180_ gnd vdd FILL
XFILL_0__12392_ gnd vdd FILL
XFILL_1__10963_ gnd vdd FILL
XFILL_5_BUFX2_insert45 gnd vdd FILL
X_13607_ _9561_/Q gnd _13607_/Y vdd INVX1
XFILL_5_BUFX2_insert56 gnd vdd FILL
XFILL_5__13132_ gnd vdd FILL
XFILL_5__9673_ gnd vdd FILL
X_10819_ _10819_/A _10773_/A _10818_/Y gnd _10819_/Y vdd OAI21X1
XFILL_5__6885_ gnd vdd FILL
XFILL_5_BUFX2_insert67 gnd vdd FILL
XFILL_3__14311_ gnd vdd FILL
XFILL_3__11523_ gnd vdd FILL
XFILL_1__12702_ gnd vdd FILL
XFILL_4__13862_ gnd vdd FILL
X_14587_ _14583_/Y _14586_/Y gnd _14587_/Y vdd NOR2X1
XFILL_3__15291_ gnd vdd FILL
X_11799_ _11798_/Y _11799_/B gnd _11800_/A vdd NOR2X1
XFILL_2__8915_ gnd vdd FILL
XFILL_0__14131_ gnd vdd FILL
XFILL_5_BUFX2_insert78 gnd vdd FILL
XBUFX2_insert640 _12438_/Y gnd _9940_/B vdd BUFX2
XFILL_2__10164_ gnd vdd FILL
XFILL_0__11343_ gnd vdd FILL
XFILL_2__9895_ gnd vdd FILL
XFILL_5_BUFX2_insert89 gnd vdd FILL
XFILL_1__13682_ gnd vdd FILL
XFILL_5__8624_ gnd vdd FILL
XBUFX2_insert651 _10915_/Y gnd _12084_/A vdd BUFX2
XFILL_1__10894_ gnd vdd FILL
X_16326_ _16326_/A gnd _16325_/Y gnd _16326_/Y vdd OAI21X1
XFILL_4__15601_ gnd vdd FILL
XFILL_0__7930_ gnd vdd FILL
XBUFX2_insert662 _11364_/Y gnd _11681_/B vdd BUFX2
X_13538_ _8700_/A gnd _13539_/C vdd INVX1
XFILL_5__10275_ gnd vdd FILL
XFILL_3__14242_ gnd vdd FILL
XBUFX2_insert673 _15064_/Y gnd _15622_/A vdd BUFX2
XFILL_3__11454_ gnd vdd FILL
XFILL_1__15421_ gnd vdd FILL
XFILL_1__12633_ gnd vdd FILL
XFILL_2__8846_ gnd vdd FILL
XFILL_4__13793_ gnd vdd FILL
XFILL112280x64050 gnd vdd FILL
XBUFX2_insert684 _13459_/Y gnd _13882_/B vdd BUFX2
XBUFX2_insert695 _13362_/Y gnd _10511_/A vdd BUFX2
XFILL_0__14062_ gnd vdd FILL
XFILL_0__11274_ gnd vdd FILL
XFILL_2__14972_ gnd vdd FILL
XFILL_5__12014_ gnd vdd FILL
XFILL_0__7861_ gnd vdd FILL
XFILL_3__10405_ gnd vdd FILL
X_13469_ _8662_/Q gnd _13469_/Y vdd INVX1
XFILL_4__15532_ gnd vdd FILL
XSFILL94440x10050 gnd vdd FILL
X_16257_ _16257_/A _16257_/B gnd _16258_/C vdd NOR2X1
XFILL_4__12744_ gnd vdd FILL
XFILL_3__14173_ gnd vdd FILL
XFILL_1__15352_ gnd vdd FILL
XFILL_2__13923_ gnd vdd FILL
XFILL_3__7570_ gnd vdd FILL
XFILL_3__11385_ gnd vdd FILL
XFILL_0__13013_ gnd vdd FILL
XFILL_5__7506_ gnd vdd FILL
XFILL_2__8777_ gnd vdd FILL
XFILL_0__9600_ gnd vdd FILL
X_15208_ _15208_/A _15208_/B _14265_/C gnd _12833_/B vdd AOI21X1
XFILL_5__8486_ gnd vdd FILL
XFILL_3__13124_ gnd vdd FILL
XSFILL79240x71050 gnd vdd FILL
X_16188_ _15392_/C _16187_/Y _15677_/D _14797_/Y gnd _16189_/B vdd OAI22X1
XFILL_1__14303_ gnd vdd FILL
XFILL_4__15463_ gnd vdd FILL
XFILL_2__7728_ gnd vdd FILL
XFILL_1__11515_ gnd vdd FILL
XFILL_2__13854_ gnd vdd FILL
XFILL_0__10156_ gnd vdd FILL
XFILL_1__15283_ gnd vdd FILL
XFILL_0__9531_ gnd vdd FILL
XFILL_5__7437_ gnd vdd FILL
XFILL_1__12495_ gnd vdd FILL
X_15139_ _16225_/C _13537_/Y _15558_/D _15139_/D gnd _15139_/Y vdd OAI22X1
XFILL_4__14414_ gnd vdd FILL
XFILL_3__9240_ gnd vdd FILL
X_8070_ _8107_/B _9094_/B gnd _8070_/Y vdd NAND2X1
XSFILL28840x4050 gnd vdd FILL
XFILL_4__11626_ gnd vdd FILL
XFILL_5__13965_ gnd vdd FILL
XFILL_4__15394_ gnd vdd FILL
XFILL_1__14234_ gnd vdd FILL
XFILL_3__10267_ gnd vdd FILL
XFILL_2__13785_ gnd vdd FILL
XSFILL115000x5050 gnd vdd FILL
XFILL_1__11446_ gnd vdd FILL
XSFILL18680x24050 gnd vdd FILL
XSFILL114440x80050 gnd vdd FILL
XFILL_0__14964_ gnd vdd FILL
XSFILL74200x18050 gnd vdd FILL
XFILL_2__10997_ gnd vdd FILL
X_7021_ _7021_/Q _7021_/CLK _9069_/R vdd _7021_/D gnd vdd DFFSR
XFILL_6__13166_ gnd vdd FILL
XFILL_5__15704_ gnd vdd FILL
XFILL_0__9462_ gnd vdd FILL
XFILL_3__12006_ gnd vdd FILL
XFILL_5__7368_ gnd vdd FILL
XFILL_5__12916_ gnd vdd FILL
XFILL_6__10378_ gnd vdd FILL
XFILL_4__14345_ gnd vdd FILL
XFILL_2__12736_ gnd vdd FILL
XFILL_2__15524_ gnd vdd FILL
XFILL_3__9171_ gnd vdd FILL
XFILL_5__13896_ gnd vdd FILL
XFILL_4__11557_ gnd vdd FILL
XSFILL84360x62050 gnd vdd FILL
XFILL_1__14165_ gnd vdd FILL
XFILL_5__9107_ gnd vdd FILL
XFILL_0__13915_ gnd vdd FILL
XFILL_1__11377_ gnd vdd FILL
XFILL_5__7299_ gnd vdd FILL
XFILL_5__15635_ gnd vdd FILL
XFILL_0__14895_ gnd vdd FILL
XFILL_4__10508_ gnd vdd FILL
XFILL_3__8122_ gnd vdd FILL
XFILL_5__12847_ gnd vdd FILL
XFILL_0__9393_ gnd vdd FILL
XFILL_1__13116_ gnd vdd FILL
XFILL_4__14276_ gnd vdd FILL
XFILL_2__15455_ gnd vdd FILL
XFILL_4__11488_ gnd vdd FILL
XFILL_5__9038_ gnd vdd FILL
XFILL_0__13846_ gnd vdd FILL
XFILL_1__14096_ gnd vdd FILL
XFILL_4__16015_ gnd vdd FILL
XFILL_0__8344_ gnd vdd FILL
XFILL_4__13227_ gnd vdd FILL
XFILL_5__15566_ gnd vdd FILL
XFILL_5__12778_ gnd vdd FILL
X_8972_ _9014_/A _6924_/B gnd _8973_/C vdd NAND2X1
XFILL_4__10439_ gnd vdd FILL
XFILL_2__14406_ gnd vdd FILL
XFILL_2__11618_ gnd vdd FILL
XFILL_2__15386_ gnd vdd FILL
XFILL_3__13957_ gnd vdd FILL
XFILL_2__12598_ gnd vdd FILL
XFILL_1__10259_ gnd vdd FILL
XFILL_0__13777_ gnd vdd FILL
XFILL_5__14517_ gnd vdd FILL
XSFILL38840x37050 gnd vdd FILL
X_7923_ _7885_/A _8051_/CLK _8051_/R vdd _7923_/D gnd vdd DFFSR
XFILL112360x44050 gnd vdd FILL
XFILL_0__8275_ gnd vdd FILL
XFILL_0__10989_ gnd vdd FILL
XFILL_5__11729_ gnd vdd FILL
XFILL_3__12908_ gnd vdd FILL
XFILL_4__13158_ gnd vdd FILL
XFILL_2__14337_ gnd vdd FILL
XFILL_5__15497_ gnd vdd FILL
XFILL_0__15516_ gnd vdd FILL
XFILL_2__11549_ gnd vdd FILL
XFILL_0__12728_ gnd vdd FILL
XSFILL79720x49050 gnd vdd FILL
XFILL_3__13888_ gnd vdd FILL
XFILL_0__7226_ gnd vdd FILL
XFILL_6__15807_ gnd vdd FILL
XFILL_6__9782_ gnd vdd FILL
XFILL_4__12109_ gnd vdd FILL
XFILL_5__14448_ gnd vdd FILL
XFILL_3__15627_ gnd vdd FILL
X_7854_ _7852_/Y _7800_/B _7854_/C gnd _7912_/D vdd OAI21X1
XFILL_4__13089_ gnd vdd FILL
XFILL_3__12839_ gnd vdd FILL
XFILL_2__14268_ gnd vdd FILL
XFILL_0__15447_ gnd vdd FILL
XFILL_0__12659_ gnd vdd FILL
XSFILL79320x51050 gnd vdd FILL
XFILL_1__14998_ gnd vdd FILL
XFILL_6__8733_ gnd vdd FILL
XFILL_0_CLKBUF1_insert207 gnd vdd FILL
XSFILL43960x28050 gnd vdd FILL
XFILL_2__13219_ gnd vdd FILL
XSFILL3560x77050 gnd vdd FILL
XFILL_2__16007_ gnd vdd FILL
XFILL_5__14379_ gnd vdd FILL
XFILL_0_CLKBUF1_insert218 gnd vdd FILL
XFILL_3__15558_ gnd vdd FILL
X_7785_ _7727_/A _7664_/CLK _7920_/R vdd _7785_/D gnd vdd DFFSR
XSFILL94200x4050 gnd vdd FILL
XFILL_2__14199_ gnd vdd FILL
XFILL_3__8955_ gnd vdd FILL
XFILL_1__13949_ gnd vdd FILL
XFILL_0__15378_ gnd vdd FILL
XFILL_5__16118_ gnd vdd FILL
X_9524_ _9522_/Y _9529_/A _9524_/C gnd _9578_/D vdd OAI21X1
XFILL_6__15669_ gnd vdd FILL
XFILL_1__7970_ gnd vdd FILL
XFILL_3__14509_ gnd vdd FILL
XFILL_0__7088_ gnd vdd FILL
XSFILL114520x60050 gnd vdd FILL
XSFILL8600x14050 gnd vdd FILL
XSFILL44040x37050 gnd vdd FILL
XFILL_3__15489_ gnd vdd FILL
XFILL_0__14329_ gnd vdd FILL
XFILL_3__8886_ gnd vdd FILL
XFILL_1__6921_ gnd vdd FILL
XFILL_5__16049_ gnd vdd FILL
X_9455_ _9455_/Q _9568_/CLK _8431_/R vdd _9411_/Y gnd vdd DFFSR
XFILL_1__15619_ gnd vdd FILL
XFILL_3__7837_ gnd vdd FILL
X_8406_ _8310_/A _7382_/CLK _8674_/R vdd _8406_/D gnd vdd DFFSR
XFILL_1__9640_ gnd vdd FILL
XFILL_1__6852_ gnd vdd FILL
X_9386_ _9372_/B _9258_/B gnd _9387_/C vdd NAND2X1
XFILL_4_BUFX2_insert703 gnd vdd FILL
XFILL_4_BUFX2_insert714 gnd vdd FILL
XFILL_6__7477_ gnd vdd FILL
XFILL_4_BUFX2_insert725 gnd vdd FILL
X_8337_ _8415_/Q gnd _8337_/Y vdd INVX1
XFILL_3__9507_ gnd vdd FILL
XFILL_4_BUFX2_insert736 gnd vdd FILL
XFILL_4__9280_ gnd vdd FILL
XFILL_4_BUFX2_insert747 gnd vdd FILL
XFILL_4_BUFX2_insert758 gnd vdd FILL
XFILL112440x24050 gnd vdd FILL
XFILL_4_BUFX2_insert769 gnd vdd FILL
XFILL_1__8522_ gnd vdd FILL
XFILL_3__7699_ gnd vdd FILL
XFILL_0__9729_ gnd vdd FILL
XFILL_3_CLKBUF1_insert1079 gnd vdd FILL
X_8268_ _8268_/A _8249_/A _8267_/Y gnd _8268_/Y vdd OAI21X1
XSFILL49560x68050 gnd vdd FILL
XFILL_4__8231_ gnd vdd FILL
XSFILL89160x54050 gnd vdd FILL
XSFILL39000x26050 gnd vdd FILL
X_7219_ _7250_/B _8243_/B gnd _7220_/C vdd NAND2X1
XFILL_1__8453_ gnd vdd FILL
XSFILL8600x5050 gnd vdd FILL
X_8199_ _8197_/Y _8237_/A _8199_/C gnd _8199_/Y vdd OAI21X1
XFILL_3__9369_ gnd vdd FILL
XFILL_1__8384_ gnd vdd FILL
XFILL_4__7113_ gnd vdd FILL
XFILL_4__8093_ gnd vdd FILL
XSFILL28840x69050 gnd vdd FILL
XFILL_1__7335_ gnd vdd FILL
XFILL_4__7044_ gnd vdd FILL
X_12840_ _12838_/Y vdd _12840_/C gnd _12924_/D vdd OAI21X1
XFILL_1_BUFX2_insert604 gnd vdd FILL
XFILL_1__9005_ gnd vdd FILL
X_12771_ _12723_/A memoryOutData[25] gnd _12772_/C vdd NAND2X1
XFILL_1_BUFX2_insert615 gnd vdd FILL
XFILL_1_BUFX2_insert626 gnd vdd FILL
XFILL_1__7197_ gnd vdd FILL
XFILL_1_BUFX2_insert637 gnd vdd FILL
XFILL_1_BUFX2_insert648 gnd vdd FILL
X_14510_ _9964_/Q _13645_/C _14510_/C gnd _14510_/Y vdd AOI21X1
X_11722_ _11713_/C _11681_/B _11573_/C _11073_/Y gnd _11722_/Y vdd AOI22X1
XFILL_4__8995_ gnd vdd FILL
XFILL_1_BUFX2_insert659 gnd vdd FILL
X_15490_ _15488_/Y _15527_/C _15449_/C _15490_/D gnd _15490_/Y vdd OAI22X1
XFILL_4__7946_ gnd vdd FILL
X_11653_ _11653_/A gnd _11654_/C vdd INVX1
X_14441_ _15870_/A _14441_/B _14555_/C _15870_/D gnd _14445_/A vdd OAI22X1
XFILL_2__6961_ gnd vdd FILL
XSFILL89240x34050 gnd vdd FILL
X_10604_ _10552_/A _9958_/CLK _8929_/R vdd _10604_/D gnd vdd DFFSR
XFILL_4__7877_ gnd vdd FILL
X_14372_ _7471_/A gnd _15829_/B vdd INVX1
XFILL_1__9907_ gnd vdd FILL
XFILL_2__8700_ gnd vdd FILL
X_11584_ _11153_/Y gnd _11588_/B vdd INVX1
XFILL_4__9616_ gnd vdd FILL
XFILL_2__6892_ gnd vdd FILL
XFILL_2__9680_ gnd vdd FILL
X_13323_ _13289_/B _13322_/Y _13316_/Y gnd _13323_/Y vdd OAI21X1
X_16111_ _16111_/A _16110_/Y _16111_/C gnd _16123_/A vdd NAND3X1
X_10535_ _10535_/A _7975_/B gnd _10536_/C vdd NAND2X1
XFILL_5__10060_ gnd vdd FILL
XFILL_5_BUFX2_insert570 gnd vdd FILL
XFILL_2__8631_ gnd vdd FILL
XFILL_4__10790_ gnd vdd FILL
XFILL_5_BUFX2_insert581 gnd vdd FILL
XFILL_4__9547_ gnd vdd FILL
XFILL_5_BUFX2_insert592 gnd vdd FILL
XFILL_5__8340_ gnd vdd FILL
XSFILL94360x25050 gnd vdd FILL
X_13254_ _13274_/A gnd _13326_/A vdd INVX4
X_16042_ _15169_/D _14635_/Y _15677_/A _14632_/Y gnd _16043_/B vdd OAI22X1
X_10466_ _15547_/A _7778_/CLK _8424_/R vdd _10466_/D gnd vdd DFFSR
XFILL_2__10920_ gnd vdd FILL
XFILL_0__10010_ gnd vdd FILL
XFILL_3__11170_ gnd vdd FILL
XFILL_1__9769_ gnd vdd FILL
XFILL_5__8271_ gnd vdd FILL
X_12205_ _12108_/B gnd _12207_/A vdd INVX1
XFILL_4__9478_ gnd vdd FILL
XFILL_3__10121_ gnd vdd FILL
X_13185_ _13185_/Q _13184_/CLK _8033_/R vdd _13111_/Y gnd vdd DFFSR
XFILL_4__12460_ gnd vdd FILL
X_10397_ _14078_/A gnd _10399_/A vdd INVX1
XFILL_1__11300_ gnd vdd FILL
XFILL_2__8493_ gnd vdd FILL
XFILL_5__7222_ gnd vdd FILL
XFILL_1__12280_ gnd vdd FILL
X_12136_ _13182_/Q gnd _12138_/A vdd INVX1
XFILL_5__13750_ gnd vdd FILL
XFILL_4__11411_ gnd vdd FILL
XFILL_5__10962_ gnd vdd FILL
XFILL_3__10052_ gnd vdd FILL
XFILL_2__7444_ gnd vdd FILL
XSFILL104360x10050 gnd vdd FILL
XFILL_4__12391_ gnd vdd FILL
XFILL_2__13570_ gnd vdd FILL
XFILL_1__11231_ gnd vdd FILL
XFILL_2_CLKBUF1_insert140 gnd vdd FILL
XFILL_2__10782_ gnd vdd FILL
XFILL_5__12701_ gnd vdd FILL
XFILL_0__11961_ gnd vdd FILL
XFILL_2_CLKBUF1_insert151 gnd vdd FILL
XFILL_4__14130_ gnd vdd FILL
XFILL_2_CLKBUF1_insert162 gnd vdd FILL
X_12067_ _11987_/A _12403_/A _12059_/C gnd _12070_/A vdd NAND3X1
XFILL_2_CLKBUF1_insert173 gnd vdd FILL
XFILL_5__13681_ gnd vdd FILL
XFILL_2__12521_ gnd vdd FILL
XFILL_4__11342_ gnd vdd FILL
XFILL_3__14860_ gnd vdd FILL
XFILL_2__7375_ gnd vdd FILL
XFILL_2_CLKBUF1_insert184 gnd vdd FILL
XFILL_5__10893_ gnd vdd FILL
XFILL_0__13700_ gnd vdd FILL
XFILL_0__10912_ gnd vdd FILL
XFILL_1__11162_ gnd vdd FILL
XFILL_2_CLKBUF1_insert195 gnd vdd FILL
XFILL_5__7084_ gnd vdd FILL
XFILL_0__14680_ gnd vdd FILL
XFILL_5__15420_ gnd vdd FILL
X_11018_ _11384_/A _12138_/Y gnd _11018_/Y vdd NOR2X1
XFILL_5__12632_ gnd vdd FILL
XFILL_0__11892_ gnd vdd FILL
XSFILL89320x14050 gnd vdd FILL
XFILL_3__13811_ gnd vdd FILL
XSFILL59080x53050 gnd vdd FILL
XFILL_2__15240_ gnd vdd FILL
XFILL_2__9114_ gnd vdd FILL
XFILL_4__14061_ gnd vdd FILL
XFILL_4__11273_ gnd vdd FILL
XFILL_1__10113_ gnd vdd FILL
XFILL_2__12452_ gnd vdd FILL
XFILL_1__15970_ gnd vdd FILL
XFILL_0__13631_ gnd vdd FILL
XFILL_3__14791_ gnd vdd FILL
XFILL_1__11093_ gnd vdd FILL
XFILL_5__15351_ gnd vdd FILL
X_15826_ _15826_/A gnd _15826_/Y vdd INVX1
XFILL_4__13012_ gnd vdd FILL
XFILL_2__11403_ gnd vdd FILL
XFILL_2__9045_ gnd vdd FILL
XFILL_2__15171_ gnd vdd FILL
XFILL_3__13742_ gnd vdd FILL
XFILL_2_BUFX2_insert460 gnd vdd FILL
XFILL_3__10954_ gnd vdd FILL
XFILL_2_BUFX2_insert471 gnd vdd FILL
XFILL_1__10044_ gnd vdd FILL
XFILL112280x59050 gnd vdd FILL
XFILL_2__12383_ gnd vdd FILL
XBUFX2_insert6 _13280_/Y gnd _7359_/A vdd BUFX2
XFILL_1__14921_ gnd vdd FILL
XFILL_0__16350_ gnd vdd FILL
XFILL_2_BUFX2_insert482 gnd vdd FILL
XFILL_0__13562_ gnd vdd FILL
XFILL_5__14302_ gnd vdd FILL
XFILL_0__8060_ gnd vdd FILL
XFILL_5__11514_ gnd vdd FILL
XFILL_0__10774_ gnd vdd FILL
XFILL_6__13853_ gnd vdd FILL
XFILL_2_BUFX2_insert493 gnd vdd FILL
XFILL_4__10155_ gnd vdd FILL
XFILL_2__14122_ gnd vdd FILL
XFILL_5__15282_ gnd vdd FILL
X_15757_ _15756_/Y _15757_/B gnd _15758_/B vdd NOR2X1
XFILL_0__15301_ gnd vdd FILL
XFILL_5__12494_ gnd vdd FILL
X_12969_ _6876_/A gnd _12969_/Y vdd INVX1
XFILL_2__11334_ gnd vdd FILL
XFILL_1__14852_ gnd vdd FILL
XFILL_0__12513_ gnd vdd FILL
XFILL_3__13673_ gnd vdd FILL
XFILL_3__10885_ gnd vdd FILL
XFILL_0__16281_ gnd vdd FILL
XSFILL13800x71050 gnd vdd FILL
XFILL_5__14233_ gnd vdd FILL
X_14708_ _14708_/A _14865_/B _14555_/B _16106_/B gnd _14709_/A vdd OAI22X1
XFILL_0__13493_ gnd vdd FILL
XFILL_3__15412_ gnd vdd FILL
XFILL_5__11445_ gnd vdd FILL
XFILL_5__7986_ gnd vdd FILL
X_15688_ _15688_/A _15687_/Y gnd _15688_/Y vdd NOR2X1
XFILL_1__13803_ gnd vdd FILL
XFILL_3__12624_ gnd vdd FILL
XFILL_2__14053_ gnd vdd FILL
XFILL_4__14963_ gnd vdd FILL
XFILL_6__10996_ gnd vdd FILL
XSFILL79240x66050 gnd vdd FILL
XFILL_0__15232_ gnd vdd FILL
XFILL_3__16392_ gnd vdd FILL
XFILL_2__11265_ gnd vdd FILL
XFILL_0__12444_ gnd vdd FILL
XFILL_5__9725_ gnd vdd FILL
XFILL_1__14783_ gnd vdd FILL
XFILL_1__11995_ gnd vdd FILL
XFILL_5__6937_ gnd vdd FILL
X_14639_ _7534_/Q gnd _16024_/D vdd INVX1
XFILL_5__14164_ gnd vdd FILL
XFILL_4__13914_ gnd vdd FILL
XFILL_2__13004_ gnd vdd FILL
XFILL_3__15343_ gnd vdd FILL
X_7570_ _7570_/A _8466_/B gnd _7571_/C vdd NAND2X1
XFILL_5__11376_ gnd vdd FILL
XFILL_3__8740_ gnd vdd FILL
XFILL_1__13734_ gnd vdd FILL
XFILL_4__14894_ gnd vdd FILL
XFILL_1__10946_ gnd vdd FILL
XFILL_0__15163_ gnd vdd FILL
XFILL_2__11196_ gnd vdd FILL
XSFILL18680x19050 gnd vdd FILL
XSFILL114440x75050 gnd vdd FILL
XFILL_5__13115_ gnd vdd FILL
XFILL_0__12375_ gnd vdd FILL
XFILL_5__9656_ gnd vdd FILL
XSFILL8520x29050 gnd vdd FILL
XFILL_5__6868_ gnd vdd FILL
XFILL_6__15454_ gnd vdd FILL
XFILL_4__13845_ gnd vdd FILL
XFILL_0__8962_ gnd vdd FILL
XFILL_3__11506_ gnd vdd FILL
XFILL_5__14095_ gnd vdd FILL
XFILL_3__12486_ gnd vdd FILL
XFILL_2__10147_ gnd vdd FILL
XFILL_0__14114_ gnd vdd FILL
XFILL_3__15274_ gnd vdd FILL
XSFILL33720x22050 gnd vdd FILL
XSFILL84360x57050 gnd vdd FILL
XFILL_1__13665_ gnd vdd FILL
XBUFX2_insert470 _13318_/Y gnd _8345_/B vdd BUFX2
XFILL_2__9878_ gnd vdd FILL
XFILL_0__11326_ gnd vdd FILL
XFILL_5__8607_ gnd vdd FILL
XBUFX2_insert481 _14979_/Y gnd _14983_/A vdd BUFX2
XFILL_1__10877_ gnd vdd FILL
X_16309_ _16309_/A _14969_/Y _14949_/D _15802_/D gnd _16312_/B vdd OAI22X1
XFILL_0__15094_ gnd vdd FILL
X_9240_ _9240_/A _8088_/B gnd _9241_/C vdd NAND2X1
XFILL_5__13046_ gnd vdd FILL
XBUFX2_insert492 _13471_/Y gnd _14721_/A vdd BUFX2
XFILL_1__15404_ gnd vdd FILL
XFILL_3__14225_ gnd vdd FILL
XFILL_0__8893_ gnd vdd FILL
XFILL_5__10258_ gnd vdd FILL
XFILL_3__11437_ gnd vdd FILL
XFILL_1__12616_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1074 gnd vdd FILL
XFILL_4__13776_ gnd vdd FILL
XFILL_3__7622_ gnd vdd FILL
XFILL_2__8829_ gnd vdd FILL
XFILL_1__16384_ gnd vdd FILL
XFILL_0__14045_ gnd vdd FILL
XFILL_4__10988_ gnd vdd FILL
XFILL_2__14955_ gnd vdd FILL
XFILL_1__13596_ gnd vdd FILL
XSFILL59160x33050 gnd vdd FILL
XFILL_0__11257_ gnd vdd FILL
XFILL_0__7844_ gnd vdd FILL
XFILL_4__15515_ gnd vdd FILL
XFILL_6__11548_ gnd vdd FILL
XFILL_4__12727_ gnd vdd FILL
X_9171_ _9205_/Q gnd _9173_/A vdd INVX1
XFILL_5__10189_ gnd vdd FILL
XFILL_1__15335_ gnd vdd FILL
XFILL_3__14156_ gnd vdd FILL
XFILL_2__13906_ gnd vdd FILL
XFILL_3__11368_ gnd vdd FILL
XFILL_3__7553_ gnd vdd FILL
XFILL_0__11188_ gnd vdd FILL
XFILL_2__14886_ gnd vdd FILL
X_8122_ _8122_/A _8142_/A _8122_/C gnd _8172_/D vdd OAI21X1
XFILL_5__8469_ gnd vdd FILL
XFILL_6__14267_ gnd vdd FILL
XFILL_3__10319_ gnd vdd FILL
XFILL_3__13107_ gnd vdd FILL
XFILL_4__15446_ gnd vdd FILL
XFILL_4__12658_ gnd vdd FILL
XFILL_5__14997_ gnd vdd FILL
XFILL_3__14087_ gnd vdd FILL
XFILL_3__7484_ gnd vdd FILL
XFILL_2__13837_ gnd vdd FILL
XFILL_0__10139_ gnd vdd FILL
XFILL_3__11299_ gnd vdd FILL
XFILL_1__15266_ gnd vdd FILL
XFILL_1__12478_ gnd vdd FILL
XSFILL23640x74050 gnd vdd FILL
XFILL_0__15996_ gnd vdd FILL
XFILL_6__7193_ gnd vdd FILL
XFILL_0__9514_ gnd vdd FILL
XFILL_3__13038_ gnd vdd FILL
X_8053_ _8019_/A _7537_/CLK _8053_/R vdd _8053_/D gnd vdd DFFSR
XFILL_4__11609_ gnd vdd FILL
XFILL_5__13948_ gnd vdd FILL
XFILL_4__15377_ gnd vdd FILL
XFILL_1__14217_ gnd vdd FILL
XSFILL109400x64050 gnd vdd FILL
XFILL_3__9223_ gnd vdd FILL
XFILL_4__12589_ gnd vdd FILL
XFILL_1_BUFX2_insert10 gnd vdd FILL
XFILL_1__11429_ gnd vdd FILL
XFILL_1__15197_ gnd vdd FILL
XFILL_2__13768_ gnd vdd FILL
XSFILL24280x40050 gnd vdd FILL
XFILL_0__14947_ gnd vdd FILL
X_7004_ _7004_/Q _7406_/CLK _8430_/R vdd _7004_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert21 gnd vdd FILL
XSFILL79320x46050 gnd vdd FILL
XFILL_4__14328_ gnd vdd FILL
XFILL_1_BUFX2_insert32 gnd vdd FILL
XFILL_5__13879_ gnd vdd FILL
XFILL_1_BUFX2_insert43 gnd vdd FILL
XFILL_2__15507_ gnd vdd FILL
XFILL_2__12719_ gnd vdd FILL
XFILL_1__14148_ gnd vdd FILL
XFILL_3__9154_ gnd vdd FILL
XFILL_1_BUFX2_insert54 gnd vdd FILL
XFILL_1_BUFX2_insert65 gnd vdd FILL
XFILL_2__13699_ gnd vdd FILL
XFILL_0__14878_ gnd vdd FILL
XFILL_1_BUFX2_insert76 gnd vdd FILL
XFILL_0__9376_ gnd vdd FILL
XFILL_5__15618_ gnd vdd FILL
XFILL_4__14259_ gnd vdd FILL
XFILL_1_BUFX2_insert87 gnd vdd FILL
XFILL_3__8105_ gnd vdd FILL
XFILL_1_BUFX2_insert98 gnd vdd FILL
XFILL_2__15438_ gnd vdd FILL
XFILL_3__9085_ gnd vdd FILL
XFILL_0__13829_ gnd vdd FILL
XFILL_3__14989_ gnd vdd FILL
XFILL_1__14079_ gnd vdd FILL
XFILL_0__8327_ gnd vdd FILL
XFILL_1__7120_ gnd vdd FILL
XFILL_5__15549_ gnd vdd FILL
X_8955_ _8955_/A _9044_/A _8955_/C gnd _9047_/D vdd OAI21X1
XSFILL115160x21050 gnd vdd FILL
XFILL_2__15369_ gnd vdd FILL
XFILL_1__7051_ gnd vdd FILL
X_7906_ _7906_/Q _7778_/CLK _8418_/R vdd _7836_/Y gnd vdd DFFSR
XFILL_0__8258_ gnd vdd FILL
X_8886_ _8845_/B _7094_/B gnd _8887_/C vdd NAND2X1
XFILL_0__7209_ gnd vdd FILL
X_7837_ _7907_/Q gnd _7837_/Y vdd INVX1
XFILL_0__8189_ gnd vdd FILL
XFILL_4__7800_ gnd vdd FILL
XFILL111960x12050 gnd vdd FILL
XFILL_3__9987_ gnd vdd FILL
XFILL_4__8780_ gnd vdd FILL
XFILL112440x19050 gnd vdd FILL
X_7768_ _7768_/Q _7640_/CLK _7896_/R vdd _7768_/D gnd vdd DFFSR
XFILL_4__7731_ gnd vdd FILL
X_9507_ _9507_/A gnd _9509_/A vdd INVX1
XFILL112040x21050 gnd vdd FILL
XFILL_1__7953_ gnd vdd FILL
X_7699_ _7699_/A _7729_/B _7698_/Y gnd _7775_/D vdd OAI21X1
XFILL_3__8869_ gnd vdd FILL
X_9438_ _9438_/Q _7902_/CLK _7150_/R vdd _9360_/Y gnd vdd DFFSR
XFILL_6__8578_ gnd vdd FILL
XFILL_1__6904_ gnd vdd FILL
XFILL_1__7884_ gnd vdd FILL
XFILL_4__9401_ gnd vdd FILL
X_10320_ _14885_/A gnd _10320_/Y vdd INVX1
XFILL_4_BUFX2_insert500 gnd vdd FILL
XFILL_4__7593_ gnd vdd FILL
XFILL_4_BUFX2_insert511 gnd vdd FILL
XFILL_1__9623_ gnd vdd FILL
XSFILL114600x35050 gnd vdd FILL
X_9369_ _9367_/Y _9356_/A _9369_/C gnd _9441_/D vdd OAI21X1
XFILL_4_BUFX2_insert522 gnd vdd FILL
XFILL_4_BUFX2_insert533 gnd vdd FILL
X_10251_ _10333_/Q gnd _10253_/A vdd INVX1
XFILL_4_BUFX2_insert544 gnd vdd FILL
XFILL_4_BUFX2_insert555 gnd vdd FILL
XFILL_4_BUFX2_insert566 gnd vdd FILL
XSFILL69080x16050 gnd vdd FILL
XFILL_1__9554_ gnd vdd FILL
XFILL_4_BUFX2_insert577 gnd vdd FILL
XFILL_4_BUFX2_insert588 gnd vdd FILL
XFILL_4__9263_ gnd vdd FILL
XFILL_1__8505_ gnd vdd FILL
X_10182_ _10182_/A _10169_/A _10182_/C gnd _10182_/Y vdd OAI21X1
XFILL_4_BUFX2_insert599 gnd vdd FILL
XFILL_1__9485_ gnd vdd FILL
XFILL_4__8214_ gnd vdd FILL
XSFILL104280x25050 gnd vdd FILL
X_14990_ _12764_/A gnd _16216_/B vdd INVX2
XFILL_4__8145_ gnd vdd FILL
X_13941_ _13940_/Y _13941_/B gnd _13941_/Y vdd NOR2X1
XFILL_2__7160_ gnd vdd FILL
XFILL_1__8367_ gnd vdd FILL
XFILL_3_CLKBUF1_insert202 gnd vdd FILL
XFILL_4__8076_ gnd vdd FILL
XFILL_3_CLKBUF1_insert213 gnd vdd FILL
XFILL_3_CLKBUF1_insert224 gnd vdd FILL
XFILL_1__7318_ gnd vdd FILL
X_13872_ _13872_/A _13868_/Y gnd _13872_/Y vdd NOR2X1
XSFILL49240x45050 gnd vdd FILL
XFILL_2__7091_ gnd vdd FILL
X_15611_ _15369_/D _15611_/B _15351_/D _14141_/C gnd _15615_/A vdd OAI22X1
X_12823_ _12823_/A gnd _12823_/Y vdd INVX1
XFILL_1_BUFX2_insert401 gnd vdd FILL
XFILL_1__7249_ gnd vdd FILL
XFILL_1_BUFX2_insert412 gnd vdd FILL
XFILL_1_BUFX2_insert423 gnd vdd FILL
XFILL_1_BUFX2_insert434 gnd vdd FILL
XFILL_5__7840_ gnd vdd FILL
X_15542_ _15537_/Y _15542_/B _15542_/C gnd _15549_/B vdd NAND3X1
X_12754_ _12754_/A _12718_/B _12753_/Y gnd _12810_/D vdd OAI21X1
XFILL_1_BUFX2_insert445 gnd vdd FILL
XFILL_1_BUFX2_insert456 gnd vdd FILL
XFILL_3__10670_ gnd vdd FILL
XFILL_1_BUFX2_insert467 gnd vdd FILL
XFILL_1_BUFX2_insert478 gnd vdd FILL
XFILL_0__10490_ gnd vdd FILL
X_11705_ _11704_/Y _11074_/C _11743_/A gnd _11706_/C vdd OAI21X1
XFILL_4__8978_ gnd vdd FILL
XFILL_5__11230_ gnd vdd FILL
X_12685_ _12633_/A _12685_/CLK _12685_/R vdd _12685_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert489 gnd vdd FILL
XFILL_6__10781_ gnd vdd FILL
X_15473_ _15472_/Y _15473_/B gnd _15473_/Y vdd NOR2X1
XFILL_2__9801_ gnd vdd FILL
XFILL_4__11960_ gnd vdd FILL
XFILL_1__10800_ gnd vdd FILL
XFILL_2__11050_ gnd vdd FILL
XSFILL4200x62050 gnd vdd FILL
XFILL_5__9510_ gnd vdd FILL
XFILL_2__7993_ gnd vdd FILL
XFILL_6__12520_ gnd vdd FILL
XFILL_4__7929_ gnd vdd FILL
XFILL_1__11780_ gnd vdd FILL
X_11636_ _11615_/Y _11637_/B _11835_/C gnd _11636_/Y vdd AOI21X1
X_14424_ _9650_/A gnd _14426_/A vdd INVX1
XFILL_4__10911_ gnd vdd FILL
XFILL_3__12340_ gnd vdd FILL
XFILL_5__11161_ gnd vdd FILL
XFILL_2__10001_ gnd vdd FILL
XFILL_1_CLKBUF1_insert1080 gnd vdd FILL
XFILL_2__9732_ gnd vdd FILL
XFILL_2__6944_ gnd vdd FILL
XFILL_4__11891_ gnd vdd FILL
XFILL_0__12160_ gnd vdd FILL
XFILL_5__10112_ gnd vdd FILL
XSFILL69000x60050 gnd vdd FILL
XFILL_4__13630_ gnd vdd FILL
X_14355_ _14353_/Y _14354_/Y _14355_/C gnd _14356_/A vdd NAND3X1
X_11567_ _11856_/A _11856_/B _11857_/B gnd _12503_/B vdd OAI21X1
XFILL_3__12271_ gnd vdd FILL
XFILL_5__11092_ gnd vdd FILL
XFILL_2__9663_ gnd vdd FILL
XFILL_1__13450_ gnd vdd FILL
XFILL_0__11111_ gnd vdd FILL
XFILL_1__10662_ gnd vdd FILL
XFILL_0__12091_ gnd vdd FILL
XFILL_2__6875_ gnd vdd FILL
X_13306_ _13297_/C _13300_/B _13305_/Y gnd _13306_/Y vdd NOR3X1
XFILL_5__9372_ gnd vdd FILL
X_10518_ _10516_/Y _10581_/B _10517_/Y gnd _10518_/Y vdd OAI21X1
XFILL_5__10043_ gnd vdd FILL
XFILL_3__14010_ gnd vdd FILL
XFILL_6__12382_ gnd vdd FILL
XFILL_3__11222_ gnd vdd FILL
XFILL_5__14920_ gnd vdd FILL
X_14286_ _9385_/A _13883_/B _14285_/Y gnd _14286_/Y vdd AOI21X1
XFILL_2__8614_ gnd vdd FILL
XFILL_1__12401_ gnd vdd FILL
XSFILL59080x48050 gnd vdd FILL
XFILL_4__13561_ gnd vdd FILL
X_11498_ _11498_/A gnd _11513_/B vdd INVX2
XBUFX2_insert90 _12357_/Y gnd _9475_/B vdd BUFX2
XFILL_2__11952_ gnd vdd FILL
XFILL_2__14740_ gnd vdd FILL
XFILL_0__11042_ gnd vdd FILL
XFILL_4__10773_ gnd vdd FILL
XFILL_5__8323_ gnd vdd FILL
XFILL_1__13381_ gnd vdd FILL
XFILL_2__9594_ gnd vdd FILL
X_13237_ _13260_/B _13236_/Y _13289_/B gnd _13237_/Y vdd OAI21X1
X_16025_ _6974_/A gnd _16026_/C vdd INVX1
XFILL_4__15300_ gnd vdd FILL
XSFILL99480x53050 gnd vdd FILL
XFILL_6__11333_ gnd vdd FILL
XFILL_5__14851_ gnd vdd FILL
XFILL_4__12512_ gnd vdd FILL
X_10449_ _10450_/B _7889_/B gnd _10449_/Y vdd NAND2X1
XFILL_2__10903_ gnd vdd FILL
XSFILL74120x51050 gnd vdd FILL
XFILL_3__11153_ gnd vdd FILL
XFILL_4__16280_ gnd vdd FILL
XFILL_1__15120_ gnd vdd FILL
XFILL_1__12332_ gnd vdd FILL
XFILL_4__13492_ gnd vdd FILL
XFILL_2__11883_ gnd vdd FILL
XFILL_0__15850_ gnd vdd FILL
XFILL_2__14671_ gnd vdd FILL
XFILL_5__8254_ gnd vdd FILL
XFILL_5__13802_ gnd vdd FILL
X_13168_ _13166_/Y _13168_/B _13167_/Y gnd _13204_/D vdd OAI21X1
XFILL_4__15231_ gnd vdd FILL
XFILL_0__7560_ gnd vdd FILL
XFILL_3__10104_ gnd vdd FILL
XFILL_2__16410_ gnd vdd FILL
XFILL_4__12443_ gnd vdd FILL
XFILL_5__14782_ gnd vdd FILL
XFILL_2__13622_ gnd vdd FILL
XFILL_0__14801_ gnd vdd FILL
XFILL_1__15051_ gnd vdd FILL
XFILL_3__15961_ gnd vdd FILL
XFILL_5__11994_ gnd vdd FILL
XFILL_3__11084_ gnd vdd FILL
XFILL_2__10834_ gnd vdd FILL
XFILL_5__7205_ gnd vdd FILL
XFILL_2__8476_ gnd vdd FILL
XFILL_1__12263_ gnd vdd FILL
XFILL_0__15781_ gnd vdd FILL
X_12119_ _12123_/B _12119_/B gnd _12119_/Y vdd NAND2X1
XFILL_0__12993_ gnd vdd FILL
XFILL_5__13733_ gnd vdd FILL
XFILL_5__8185_ gnd vdd FILL
XFILL_5__10945_ gnd vdd FILL
XSFILL13800x66050 gnd vdd FILL
XFILL_1__14002_ gnd vdd FILL
X_13099_ _13099_/A _13099_/B _13098_/Y gnd _13181_/D vdd OAI21X1
XFILL_3__10035_ gnd vdd FILL
XFILL_0__7491_ gnd vdd FILL
XFILL_4__15162_ gnd vdd FILL
XFILL_6__11195_ gnd vdd FILL
XFILL_3__14912_ gnd vdd FILL
XFILL_2__7427_ gnd vdd FILL
XFILL_2__16341_ gnd vdd FILL
XFILL_4__12374_ gnd vdd FILL
XFILL_2__13553_ gnd vdd FILL
XFILL_1__11214_ gnd vdd FILL
XFILL_2__10765_ gnd vdd FILL
XFILL_3__15892_ gnd vdd FILL
XFILL_0__14732_ gnd vdd FILL
XFILL_0__9230_ gnd vdd FILL
XFILL_0__11944_ gnd vdd FILL
XFILL_1__12194_ gnd vdd FILL
XFILL_4__14113_ gnd vdd FILL
XFILL_2__12504_ gnd vdd FILL
XFILL_5__13664_ gnd vdd FILL
XFILL_4__11325_ gnd vdd FILL
XFILL_3__14843_ gnd vdd FILL
XFILL_2__7358_ gnd vdd FILL
XFILL_5__10876_ gnd vdd FILL
XFILL_4__15093_ gnd vdd FILL
XFILL_2__13484_ gnd vdd FILL
XFILL_1__11145_ gnd vdd FILL
XFILL_2__16272_ gnd vdd FILL
XFILL_5__15403_ gnd vdd FILL
XFILL_5__7067_ gnd vdd FILL
XFILL_0__14663_ gnd vdd FILL
XFILL_2__10696_ gnd vdd FILL
XFILL_5__12615_ gnd vdd FILL
XFILL_0__11875_ gnd vdd FILL
XFILL_0__9161_ gnd vdd FILL
XFILL_5__16383_ gnd vdd FILL
XFILL_4__14044_ gnd vdd FILL
XFILL_5__13595_ gnd vdd FILL
XFILL_2__15223_ gnd vdd FILL
XFILL_2__12435_ gnd vdd FILL
XFILL_0__16402_ gnd vdd FILL
XFILL_4__11256_ gnd vdd FILL
XFILL_0__13614_ gnd vdd FILL
XFILL_2__7289_ gnd vdd FILL
XFILL_3__14774_ gnd vdd FILL
XFILL_0__10826_ gnd vdd FILL
XFILL_3__11986_ gnd vdd FILL
XFILL_1__15953_ gnd vdd FILL
XFILL_0__8112_ gnd vdd FILL
XFILL_1__11076_ gnd vdd FILL
XFILL_0__14594_ gnd vdd FILL
XFILL_5__15334_ gnd vdd FILL
X_15809_ _15809_/A _15809_/B gnd _15810_/A vdd NOR2X1
XFILL_0__9092_ gnd vdd FILL
X_8740_ _8740_/A _8228_/B gnd _8741_/C vdd NAND2X1
XFILL_6__7880_ gnd vdd FILL
XFILL_3__9910_ gnd vdd FILL
XSFILL43880x61050 gnd vdd FILL
XFILL_2__9028_ gnd vdd FILL
XFILL_2_BUFX2_insert290 gnd vdd FILL
XFILL_2__15154_ gnd vdd FILL
XFILL_4__11187_ gnd vdd FILL
XFILL_3__13725_ gnd vdd FILL
XFILL_3__10937_ gnd vdd FILL
XFILL_2__12366_ gnd vdd FILL
XFILL_0__16333_ gnd vdd FILL
XFILL_1__14904_ gnd vdd FILL
XFILL_1__10027_ gnd vdd FILL
XFILL_0__13545_ gnd vdd FILL
XSFILL59160x28050 gnd vdd FILL
XFILL_0__10757_ gnd vdd FILL
XFILL_1__15884_ gnd vdd FILL
XFILL_5__15265_ gnd vdd FILL
XFILL_4__10138_ gnd vdd FILL
XFILL_6_BUFX2_insert628 gnd vdd FILL
XFILL_5__12477_ gnd vdd FILL
XFILL_2__11317_ gnd vdd FILL
XFILL_2__14105_ gnd vdd FILL
X_8671_ _8671_/Q _9716_/CLK _8682_/R vdd _8595_/Y gnd vdd DFFSR
XFILL_4__15995_ gnd vdd FILL
XFILL_3__13656_ gnd vdd FILL
XFILL_2__15085_ gnd vdd FILL
XFILL_1__14835_ gnd vdd FILL
XFILL_0__16264_ gnd vdd FILL
XFILL_2__12297_ gnd vdd FILL
XFILL_5__14216_ gnd vdd FILL
XFILL_0__13476_ gnd vdd FILL
XFILL_0__10688_ gnd vdd FILL
XFILL_5__7969_ gnd vdd FILL
X_7622_ _7622_/A _7577_/B _7622_/C gnd _7622_/Y vdd OAI21X1
XFILL111880x27050 gnd vdd FILL
XSFILL89800x10050 gnd vdd FILL
XFILL_5__11428_ gnd vdd FILL
XSFILL99000x76050 gnd vdd FILL
XFILL_5__15196_ gnd vdd FILL
XFILL_3__12607_ gnd vdd FILL
XFILL_2__14036_ gnd vdd FILL
XFILL_4__10069_ gnd vdd FILL
XFILL_4__14946_ gnd vdd FILL
XFILL_0__15215_ gnd vdd FILL
XFILL_1_BUFX2_insert990 gnd vdd FILL
XFILL_3__16375_ gnd vdd FILL
XFILL_2__11248_ gnd vdd FILL
XFILL_3__9772_ gnd vdd FILL
XFILL_3__13587_ gnd vdd FILL
XFILL_0__12427_ gnd vdd FILL
XFILL_3__10799_ gnd vdd FILL
XFILL_1__14766_ gnd vdd FILL
XFILL_0__16195_ gnd vdd FILL
XFILL_6__15506_ gnd vdd FILL
XFILL_1__11978_ gnd vdd FILL
XFILL_3__6984_ gnd vdd FILL
XSFILL23640x69050 gnd vdd FILL
XFILL_5__14147_ gnd vdd FILL
X_7553_ _7551_/Y _7568_/B _7553_/C gnd _7553_/Y vdd OAI21X1
XFILL_3__15326_ gnd vdd FILL
XSFILL108920x52050 gnd vdd FILL
XFILL_5__11359_ gnd vdd FILL
XFILL_4__14877_ gnd vdd FILL
XFILL_0__9994_ gnd vdd FILL
XFILL_3__8723_ gnd vdd FILL
XFILL_1__13717_ gnd vdd FILL
XFILL_1__10929_ gnd vdd FILL
XFILL112440x1050 gnd vdd FILL
XFILL_2__11179_ gnd vdd FILL
XFILL_0__15146_ gnd vdd FILL
XFILL_5__9639_ gnd vdd FILL
XFILL_0__12358_ gnd vdd FILL
XFILL_1__14697_ gnd vdd FILL
XFILL_6__12649_ gnd vdd FILL
XFILL_4__13828_ gnd vdd FILL
XFILL_5__14078_ gnd vdd FILL
X_7484_ _7425_/B _8636_/B gnd _7485_/C vdd NAND2X1
XFILL_3__15257_ gnd vdd FILL
XFILL_3__8654_ gnd vdd FILL
XFILL_1__13648_ gnd vdd FILL
XFILL_3__12469_ gnd vdd FILL
XFILL_0__11309_ gnd vdd FILL
XFILL_2__15987_ gnd vdd FILL
XSFILL38840x50050 gnd vdd FILL
XFILL_0__15077_ gnd vdd FILL
XFILL_5__13029_ gnd vdd FILL
XFILL_0__12289_ gnd vdd FILL
X_9223_ _9223_/A _9238_/B _9223_/C gnd _9223_/Y vdd OAI21X1
XFILL_3__14208_ gnd vdd FILL
XFILL_3__7605_ gnd vdd FILL
XFILL_4__13759_ gnd vdd FILL
XFILL_0__8876_ gnd vdd FILL
XFILL_1__16367_ gnd vdd FILL
XFILL_3__15188_ gnd vdd FILL
XFILL_0__14028_ gnd vdd FILL
XFILL_2__14938_ gnd vdd FILL
XFILL_3__8585_ gnd vdd FILL
XSFILL74120x3050 gnd vdd FILL
XFILL_1__13579_ gnd vdd FILL
XFILL_5_CLKBUF1_insert190 gnd vdd FILL
XFILL_6__14319_ gnd vdd FILL
X_9154_ _9170_/B _9282_/B gnd _9154_/Y vdd NAND2X1
XFILL_0__7827_ gnd vdd FILL
XFILL_3__14139_ gnd vdd FILL
XFILL_1__15318_ gnd vdd FILL
XFILL_2__14869_ gnd vdd FILL
XFILL_1__16298_ gnd vdd FILL
XSFILL43960x41050 gnd vdd FILL
X_8105_ _8167_/Q gnd _8107_/A vdd INVX1
XFILL_3_BUFX2_insert507 gnd vdd FILL
XFILL_4__15429_ gnd vdd FILL
XFILL_0__7758_ gnd vdd FILL
XFILL_3_BUFX2_insert518 gnd vdd FILL
X_9085_ _9116_/B _7293_/B gnd _9086_/C vdd NAND2X1
XFILL_3_BUFX2_insert529 gnd vdd FILL
XFILL_1__15249_ gnd vdd FILL
XSFILL84040x34050 gnd vdd FILL
XFILL_3__7467_ gnd vdd FILL
XFILL_0__15979_ gnd vdd FILL
XSFILL58200x44050 gnd vdd FILL
XFILL_1__9270_ gnd vdd FILL
X_8036_ _8036_/Q _8161_/CLK _7140_/R vdd _8036_/D gnd vdd DFFSR
XFILL_0__7689_ gnd vdd FILL
XFILL_3__9206_ gnd vdd FILL
XSFILL44040x50050 gnd vdd FILL
XFILL_1__8221_ gnd vdd FILL
XFILL_0__9428_ gnd vdd FILL
XFILL_3__9137_ gnd vdd FILL
XSFILL23720x49050 gnd vdd FILL
XSFILL8600x50 gnd vdd FILL
XFILL_0__9359_ gnd vdd FILL
X_9987_ _9996_/A _9347_/B gnd _9988_/C vdd NAND2X1
XFILL_1__7103_ gnd vdd FILL
XSFILL38920x30050 gnd vdd FILL
X_8938_ _8938_/Q _7007_/CLK _9332_/R vdd _8884_/Y gnd vdd DFFSR
XFILL_1__8083_ gnd vdd FILL
XFILL_3__8019_ gnd vdd FILL
XFILL_4__8901_ gnd vdd FILL
XSFILL64200x63050 gnd vdd FILL
XFILL_4__9881_ gnd vdd FILL
XFILL_1__7034_ gnd vdd FILL
X_8869_ _8867_/Y _8823_/B _8869_/C gnd _8933_/D vdd OAI21X1
XFILL_4__8832_ gnd vdd FILL
XFILL_0_BUFX2_insert408 gnd vdd FILL
XFILL_0_BUFX2_insert419 gnd vdd FILL
XSFILL3640x70050 gnd vdd FILL
XFILL_4__8763_ gnd vdd FILL
X_12470_ vdd _12029_/A gnd _12470_/Y vdd NAND2X1
XFILL_1__8985_ gnd vdd FILL
XFILL_4__7714_ gnd vdd FILL
XSFILL28840x82050 gnd vdd FILL
X_11421_ _11358_/A _11366_/B _11334_/A _11226_/B gnd _11421_/Y vdd OAI22X1
XFILL_4__8694_ gnd vdd FILL
XFILL_1__7936_ gnd vdd FILL
X_14140_ _8096_/A gnd _14141_/C vdd INVX1
XSFILL85000x42050 gnd vdd FILL
X_11352_ _11835_/C gnd _11352_/Y vdd INVX8
XFILL_1__7867_ gnd vdd FILL
X_10303_ _10304_/B _8255_/B gnd _10303_/Y vdd NAND2X1
XSFILL33960x73050 gnd vdd FILL
X_14071_ _14069_/Y _14071_/B _13461_/C _14071_/D gnd _14072_/B vdd OAI22X1
XFILL_4__7576_ gnd vdd FILL
XFILL_4_BUFX2_insert330 gnd vdd FILL
XFILL_4_BUFX2_insert341 gnd vdd FILL
XFILL_1__9606_ gnd vdd FILL
X_11283_ _11282_/Y _11094_/B gnd _11658_/A vdd NOR2X1
XFILL_4_BUFX2_insert352 gnd vdd FILL
XFILL_4_BUFX2_insert363 gnd vdd FILL
X_13022_ _13020_/Y vdd _13022_/C gnd _13070_/D vdd OAI21X1
XSFILL74040x66050 gnd vdd FILL
XFILL_1__7798_ gnd vdd FILL
X_10234_ _10325_/B _8314_/B gnd _10235_/C vdd NAND2X1
XFILL_4_BUFX2_insert374 gnd vdd FILL
XFILL_4_BUFX2_insert385 gnd vdd FILL
XFILL_4_BUFX2_insert396 gnd vdd FILL
XFILL_2__8330_ gnd vdd FILL
XFILL_1__9537_ gnd vdd FILL
XFILL_4__9246_ gnd vdd FILL
XSFILL13480x19050 gnd vdd FILL
X_10165_ _10219_/Q gnd _10165_/Y vdd INVX1
XFILL_2__8261_ gnd vdd FILL
XSFILL74280x9050 gnd vdd FILL
XFILL_1__9468_ gnd vdd FILL
XSFILL53880x24050 gnd vdd FILL
XFILL_6__10000_ gnd vdd FILL
XFILL_2__7212_ gnd vdd FILL
X_10096_ _14734_/A _8289_/CLK _7152_/R vdd _10054_/Y gnd vdd DFFSR
X_14973_ _7251_/A gnd _14973_/Y vdd INVX1
XFILL_2__8192_ gnd vdd FILL
XFILL_2__10550_ gnd vdd FILL
XSFILL3720x50050 gnd vdd FILL
XFILL_4__8128_ gnd vdd FILL
XFILL_1__9399_ gnd vdd FILL
XFILL_5__9990_ gnd vdd FILL
X_13924_ _13924_/A _13630_/B _14949_/C _13924_/D gnd _13925_/B vdd OAI22X1
XFILL_4__11110_ gnd vdd FILL
XFILL_5__10661_ gnd vdd FILL
XFILL_4__12090_ gnd vdd FILL
XFILL_3__11840_ gnd vdd FILL
XFILL_5__12400_ gnd vdd FILL
XFILL_4__8059_ gnd vdd FILL
XFILL_0__11660_ gnd vdd FILL
XFILL_4__11041_ gnd vdd FILL
X_13855_ _9998_/A gnd _13855_/Y vdd INVX1
XFILL_5__13380_ gnd vdd FILL
XFILL_2__12220_ gnd vdd FILL
XFILL_2__7074_ gnd vdd FILL
XFILL_3__11771_ gnd vdd FILL
XFILL_5__8872_ gnd vdd FILL
X_12806_ _12806_/Q _12538_/CLK _12689_/R vdd _12742_/Y gnd vdd DFFSR
XFILL_5__12331_ gnd vdd FILL
XFILL_0__11591_ gnd vdd FILL
XFILL_1_BUFX2_insert231 gnd vdd FILL
XFILL_3__13510_ gnd vdd FILL
X_13786_ _13786_/A _13782_/Y gnd _13787_/A vdd NOR2X1
XFILL_1_BUFX2_insert242 gnd vdd FILL
XFILL_1__11901_ gnd vdd FILL
XFILL_2__12151_ gnd vdd FILL
X_10998_ _10997_/Y gnd _11348_/A vdd INVX2
XFILL_0__13330_ gnd vdd FILL
XFILL_3__14490_ gnd vdd FILL
XFILL_1_BUFX2_insert253 gnd vdd FILL
XFILL_5__7823_ gnd vdd FILL
XFILL_0__10542_ gnd vdd FILL
XFILL_1__12881_ gnd vdd FILL
XFILL_4__14800_ gnd vdd FILL
XSFILL99480x48050 gnd vdd FILL
XFILL_5__15050_ gnd vdd FILL
X_15525_ _8343_/A gnd _15527_/D vdd INVX1
XFILL_1_BUFX2_insert264 gnd vdd FILL
X_12737_ _11882_/B gnd _12737_/Y vdd INVX1
XFILL_1_BUFX2_insert275 gnd vdd FILL
XFILL_5__12262_ gnd vdd FILL
XFILL_2__11102_ gnd vdd FILL
XFILL_1__14620_ gnd vdd FILL
XFILL_1_BUFX2_insert286 gnd vdd FILL
XFILL_3__13441_ gnd vdd FILL
XSFILL74120x46050 gnd vdd FILL
XFILL_4__15780_ gnd vdd FILL
XFILL_3__10653_ gnd vdd FILL
XFILL_2__12082_ gnd vdd FILL
XFILL_4__12992_ gnd vdd FILL
XFILL_1_BUFX2_insert297 gnd vdd FILL
XFILL_1__11832_ gnd vdd FILL
XFILL_0__13261_ gnd vdd FILL
XFILL_5__14001_ gnd vdd FILL
XFILL_5__7754_ gnd vdd FILL
XFILL_0_BUFX2_insert920 gnd vdd FILL
XFILL_5__11213_ gnd vdd FILL
XFILL_4__14731_ gnd vdd FILL
X_15456_ _15455_/Y _15456_/B _14402_/C gnd _12851_/B vdd AOI21X1
XFILL_0_BUFX2_insert931 gnd vdd FILL
XFILL_2__15910_ gnd vdd FILL
X_12668_ _12668_/Q _12669_/CLK _9050_/R vdd _12584_/Y gnd vdd DFFSR
XFILL_4__11943_ gnd vdd FILL
XFILL_0__15000_ gnd vdd FILL
XFILL_5__12193_ gnd vdd FILL
XFILL_3__16160_ gnd vdd FILL
XFILL_2__11033_ gnd vdd FILL
XFILL_1__14551_ gnd vdd FILL
XFILL_3__13372_ gnd vdd FILL
XFILL_0_BUFX2_insert942 gnd vdd FILL
XFILL_0__12212_ gnd vdd FILL
XFILL_2__7976_ gnd vdd FILL
XFILL_0_BUFX2_insert953 gnd vdd FILL
XFILL_1__11763_ gnd vdd FILL
XFILL_0_BUFX2_insert964 gnd vdd FILL
X_14407_ _14407_/A _14697_/B _14697_/C _14407_/D gnd _14411_/A vdd OAI22X1
XFILL_0_BUFX2_insert975 gnd vdd FILL
XFILL_5__11144_ gnd vdd FILL
XFILL_5__7685_ gnd vdd FILL
X_11619_ _11618_/B _11618_/A _11835_/C gnd _11619_/Y vdd AOI21X1
XFILL_3__15111_ gnd vdd FILL
XFILL_0__6991_ gnd vdd FILL
X_15387_ _15386_/Y _15387_/B gnd _15388_/C vdd NOR2X1
XFILL_3__12323_ gnd vdd FILL
XFILL_4__14662_ gnd vdd FILL
XFILL_1__13502_ gnd vdd FILL
XFILL_4__11874_ gnd vdd FILL
XFILL_2__6927_ gnd vdd FILL
XFILL_0_BUFX2_insert986 gnd vdd FILL
X_12599_ _12597_/Y vdd _12599_/C gnd _12673_/D vdd OAI21X1
XFILL_3__16091_ gnd vdd FILL
XFILL_2__15841_ gnd vdd FILL
XFILL_1__14482_ gnd vdd FILL
XFILL_0_BUFX2_insert997 gnd vdd FILL
XFILL_0__12143_ gnd vdd FILL
XFILL_5__9424_ gnd vdd FILL
XFILL_4__16401_ gnd vdd FILL
XFILL_1__11694_ gnd vdd FILL
XFILL_4__13613_ gnd vdd FILL
X_14338_ _7980_/A gnd _14338_/Y vdd INVX1
XFILL_0__8730_ gnd vdd FILL
XFILL_1__16221_ gnd vdd FILL
XFILL_3__15042_ gnd vdd FILL
XFILL_5__15952_ gnd vdd FILL
XFILL_5__11075_ gnd vdd FILL
XFILL_4__10825_ gnd vdd FILL
XFILL_4__14593_ gnd vdd FILL
XFILL_1__13433_ gnd vdd FILL
XFILL_2__9646_ gnd vdd FILL
XFILL_3__12254_ gnd vdd FILL
XFILL_2__6858_ gnd vdd FILL
XFILL_2__15772_ gnd vdd FILL
XSFILL54040x13050 gnd vdd FILL
XFILL_1__10645_ gnd vdd FILL
XFILL_5__9355_ gnd vdd FILL
XFILL_0__12074_ gnd vdd FILL
XFILL_2__12984_ gnd vdd FILL
XFILL_4__16332_ gnd vdd FILL
XFILL_6__15153_ gnd vdd FILL
XFILL_5__14903_ gnd vdd FILL
XFILL_5__10026_ gnd vdd FILL
XFILL_3__11205_ gnd vdd FILL
XFILL_4__13544_ gnd vdd FILL
XFILL_0__8661_ gnd vdd FILL
X_14269_ _10087_/Q gnd _14271_/D vdd INVX1
XFILL_3__12185_ gnd vdd FILL
XFILL_4__10756_ gnd vdd FILL
XFILL_2__14723_ gnd vdd FILL
XFILL_1__16152_ gnd vdd FILL
XFILL_5__15883_ gnd vdd FILL
XFILL_1__13364_ gnd vdd FILL
XFILL_0__15902_ gnd vdd FILL
XFILL_2__11935_ gnd vdd FILL
XFILL_0__11025_ gnd vdd FILL
XFILL_3__8370_ gnd vdd FILL
X_16008_ _14611_/Y _15394_/B _15726_/A _14619_/Y gnd _16009_/B vdd OAI22X1
XFILL_6__14104_ gnd vdd FILL
XFILL_1__10576_ gnd vdd FILL
XFILL_0__7612_ gnd vdd FILL
XFILL_5__9286_ gnd vdd FILL
XFILL_0__8592_ gnd vdd FILL
XFILL_5__14834_ gnd vdd FILL
XFILL_4__16263_ gnd vdd FILL
XFILL_3__11136_ gnd vdd FILL
XFILL_1__15103_ gnd vdd FILL
XFILL_3__7321_ gnd vdd FILL
XFILL_4__13475_ gnd vdd FILL
XFILL_1__12315_ gnd vdd FILL
XFILL_2__8528_ gnd vdd FILL
XFILL_4__10687_ gnd vdd FILL
XFILL_0__15833_ gnd vdd FILL
XFILL_2__11866_ gnd vdd FILL
XSFILL53960x50 gnd vdd FILL
XFILL_2__14654_ gnd vdd FILL
XFILL_1__16083_ gnd vdd FILL
XFILL_1__13295_ gnd vdd FILL
XFILL_5__8237_ gnd vdd FILL
XFILL_4__15214_ gnd vdd FILL
XFILL_0__7543_ gnd vdd FILL
XFILL_4__12426_ gnd vdd FILL
XFILL_2__13605_ gnd vdd FILL
XFILL_4__16194_ gnd vdd FILL
XFILL_3__15944_ gnd vdd FILL
XFILL_1__15034_ gnd vdd FILL
XFILL_5__11977_ gnd vdd FILL
XFILL_3__11067_ gnd vdd FILL
XFILL_5__14765_ gnd vdd FILL
XFILL_3__7252_ gnd vdd FILL
XFILL_2__8459_ gnd vdd FILL
XSFILL18680x32050 gnd vdd FILL
XFILL_1__12246_ gnd vdd FILL
XFILL_2__10817_ gnd vdd FILL
XFILL_2__14585_ gnd vdd FILL
XFILL_0__15764_ gnd vdd FILL
XFILL_2__11797_ gnd vdd FILL
XFILL_0__12976_ gnd vdd FILL
XSFILL74200x26050 gnd vdd FILL
X_9910_ _9917_/B _9782_/B gnd _9911_/C vdd NAND2X1
XFILL_5__10928_ gnd vdd FILL
XFILL_3__10018_ gnd vdd FILL
XFILL_5__13716_ gnd vdd FILL
XFILL_0__7474_ gnd vdd FILL
XFILL_4__15145_ gnd vdd FILL
XFILL_4__12357_ gnd vdd FILL
XFILL_2__16324_ gnd vdd FILL
XFILL_5__14696_ gnd vdd FILL
XFILL_3__7183_ gnd vdd FILL
XSFILL84360x70050 gnd vdd FILL
XFILL_0__14715_ gnd vdd FILL
XFILL_2__10748_ gnd vdd FILL
XFILL_2__13536_ gnd vdd FILL
XFILL_3__15875_ gnd vdd FILL
XFILL_5__7119_ gnd vdd FILL
XFILL_0__11927_ gnd vdd FILL
XFILL_1__12177_ gnd vdd FILL
XSFILL58520x80050 gnd vdd FILL
XFILL_0__15695_ gnd vdd FILL
XFILL_0__9213_ gnd vdd FILL
XFILL_5__8099_ gnd vdd FILL
XFILL_5__13647_ gnd vdd FILL
XFILL_4__11308_ gnd vdd FILL
XFILL_6__8981_ gnd vdd FILL
X_9841_ _9841_/Q _9834_/CLK _7793_/R vdd _9841_/D gnd vdd DFFSR
XFILL_3__14826_ gnd vdd FILL
XFILL_6__15986_ gnd vdd FILL
XFILL_4__15076_ gnd vdd FILL
XFILL_4__12288_ gnd vdd FILL
XFILL_1__11128_ gnd vdd FILL
XFILL_2__16255_ gnd vdd FILL
XFILL_2__10679_ gnd vdd FILL
XFILL_0__14646_ gnd vdd FILL
XFILL_2__13467_ gnd vdd FILL
XFILL_0__9144_ gnd vdd FILL
XFILL_6__7932_ gnd vdd FILL
XFILL_0__11858_ gnd vdd FILL
XFILL_4__14027_ gnd vdd FILL
XSFILL109560x13050 gnd vdd FILL
X_9772_ _9772_/A gnd _9774_/A vdd INVX1
XFILL_2__15206_ gnd vdd FILL
XFILL_5__13578_ gnd vdd FILL
XFILL_4__11239_ gnd vdd FILL
XFILL_5__16366_ gnd vdd FILL
XFILL_2__12418_ gnd vdd FILL
X_6984_ _6985_/B _7752_/B gnd _6984_/Y vdd NAND2X1
XFILL_3__14757_ gnd vdd FILL
XFILL_2__13398_ gnd vdd FILL
XFILL_2__16186_ gnd vdd FILL
XFILL_1__15936_ gnd vdd FILL
XFILL_3__11969_ gnd vdd FILL
XFILL_0__10809_ gnd vdd FILL
XFILL_1__11059_ gnd vdd FILL
XFILL_0__14577_ gnd vdd FILL
XFILL_5__15317_ gnd vdd FILL
XFILL112360x52050 gnd vdd FILL
XFILL_6_BUFX2_insert403 gnd vdd FILL
XFILL_5__12529_ gnd vdd FILL
X_8723_ _8723_/A _8753_/B _8722_/Y gnd _8799_/D vdd OAI21X1
XFILL_0__11789_ gnd vdd FILL
XSFILL64120x78050 gnd vdd FILL
XFILL_5__16297_ gnd vdd FILL
XFILL_3__13708_ gnd vdd FILL
XFILL_2__12349_ gnd vdd FILL
XFILL_0__16316_ gnd vdd FILL
XFILL_2__15137_ gnd vdd FILL
XFILL_6__9602_ gnd vdd FILL
XFILL_3__14688_ gnd vdd FILL
XFILL_0__13528_ gnd vdd FILL
XFILL_1__15867_ gnd vdd FILL
XFILL_5__15248_ gnd vdd FILL
X_8654_ _8655_/B _8654_/B gnd _8655_/C vdd NAND2X1
XFILL_3__13639_ gnd vdd FILL
XFILL_6_BUFX2_insert469 gnd vdd FILL
XFILL_4__15978_ gnd vdd FILL
XFILL_1__14818_ gnd vdd FILL
XFILL_2__15068_ gnd vdd FILL
XFILL_0__16247_ gnd vdd FILL
XFILL_0__13459_ gnd vdd FILL
X_7605_ _7605_/A gnd _7607_/A vdd INVX1
XFILL_1__15798_ gnd vdd FILL
XSFILL43960x36050 gnd vdd FILL
XFILL_5__15179_ gnd vdd FILL
X_8585_ _8577_/B _7177_/B gnd _8586_/C vdd NAND2X1
XFILL_2__14019_ gnd vdd FILL
XFILL_3__16358_ gnd vdd FILL
XFILL_4__14929_ gnd vdd FILL
XFILL_3__9755_ gnd vdd FILL
XFILL_3__6967_ gnd vdd FILL
XFILL_0__16178_ gnd vdd FILL
XFILL_4_BUFX2_insert1004 gnd vdd FILL
XFILL_1__14749_ gnd vdd FILL
XFILL_4_BUFX2_insert1015 gnd vdd FILL
XFILL_3__15309_ gnd vdd FILL
XFILL_4_BUFX2_insert1026 gnd vdd FILL
X_7536_ _7536_/Q _8560_/CLK _9313_/R vdd _7494_/Y gnd vdd DFFSR
XSFILL18760x12050 gnd vdd FILL
XFILL_4_BUFX2_insert1037 gnd vdd FILL
XFILL_3__8706_ gnd vdd FILL
XFILL_1__8770_ gnd vdd FILL
XFILL_0__9977_ gnd vdd FILL
XSFILL8600x22050 gnd vdd FILL
XFILL_4_BUFX2_insert1048 gnd vdd FILL
XSFILL44040x45050 gnd vdd FILL
XFILL_3__16289_ gnd vdd FILL
XFILL_0__15129_ gnd vdd FILL
XFILL_4_BUFX2_insert1059 gnd vdd FILL
XFILL_3__6898_ gnd vdd FILL
XFILL_4_BUFX2_insert80 gnd vdd FILL
XSFILL84440x50050 gnd vdd FILL
XFILL_1__7721_ gnd vdd FILL
XFILL_4_BUFX2_insert91 gnd vdd FILL
X_7467_ _7465_/Y _7470_/B _7467_/C gnd _7527_/D vdd OAI21X1
XFILL_3__8637_ gnd vdd FILL
XFILL_4__7430_ gnd vdd FILL
X_9206_ _9302_/Q gnd _9208_/A vdd INVX1
XSFILL84280x4050 gnd vdd FILL
XFILL_0__8859_ gnd vdd FILL
X_7398_ _7398_/Q _7282_/CLK _9054_/R vdd _7336_/Y gnd vdd DFFSR
XFILL_3__8568_ gnd vdd FILL
XFILL_4__7361_ gnd vdd FILL
XSFILL73480x74050 gnd vdd FILL
XFILL111800x66050 gnd vdd FILL
X_9137_ _9135_/Y _9112_/A _9137_/C gnd _9193_/D vdd OAI21X1
XFILL_4__9100_ gnd vdd FILL
XFILL_3_BUFX2_insert304 gnd vdd FILL
XFILL_1__7583_ gnd vdd FILL
XSFILL38920x25050 gnd vdd FILL
XFILL_3_BUFX2_insert315 gnd vdd FILL
XFILL112440x32050 gnd vdd FILL
XFILL_4__7292_ gnd vdd FILL
XFILL_3_BUFX2_insert326 gnd vdd FILL
XSFILL64200x58050 gnd vdd FILL
XFILL_2_BUFX2_insert1030 gnd vdd FILL
XFILL_3__8499_ gnd vdd FILL
XFILL_2_BUFX2_insert1041 gnd vdd FILL
XFILL_3_BUFX2_insert337 gnd vdd FILL
X_9068_ _9016_/A _8289_/CLK _7152_/R vdd _9068_/D gnd vdd DFFSR
XFILL_2_BUFX2_insert1052 gnd vdd FILL
XFILL_3_BUFX2_insert348 gnd vdd FILL
XSFILL79960x3050 gnd vdd FILL
XFILL_4__9031_ gnd vdd FILL
XFILL_3_BUFX2_insert359 gnd vdd FILL
XFILL_2_BUFX2_insert1063 gnd vdd FILL
XFILL_2_BUFX2_insert1085 gnd vdd FILL
X_8019_ _8019_/A gnd _8021_/A vdd INVX1
XSFILL39000x34050 gnd vdd FILL
XFILL_1__9253_ gnd vdd FILL
XSFILL3640x65050 gnd vdd FILL
XFILL_1__8204_ gnd vdd FILL
X_11970_ _11970_/A _11969_/A _11970_/C gnd _6865_/A vdd OAI21X1
XSFILL28840x77050 gnd vdd FILL
XSFILL28040x58050 gnd vdd FILL
X_10921_ _10920_/B _10906_/Y _10924_/A gnd _10922_/A vdd OAI21X1
XFILL_1__8135_ gnd vdd FILL
XFILL_4__9933_ gnd vdd FILL
X_13640_ _13640_/A _13824_/B _14575_/C _13640_/D gnd _13644_/B vdd OAI22X1
X_10852_ _14156_/A _9818_/CLK _8688_/R vdd _10852_/D gnd vdd DFFSR
XFILL_1__8066_ gnd vdd FILL
XSFILL44040x7050 gnd vdd FILL
XFILL_4_CLKBUF1_insert116 gnd vdd FILL
XFILL_4__9864_ gnd vdd FILL
XFILL_4_CLKBUF1_insert127 gnd vdd FILL
XSFILL33960x68050 gnd vdd FILL
X_10783_ _10783_/A _10773_/A _10782_/Y gnd _10851_/D vdd OAI21X1
X_13571_ _13571_/A _13570_/Y _13571_/C gnd _13571_/Y vdd NAND3X1
XFILL_4_CLKBUF1_insert138 gnd vdd FILL
XFILL_4_CLKBUF1_insert149 gnd vdd FILL
XSFILL7880x70050 gnd vdd FILL
X_15310_ _15310_/A _15303_/Y gnd _15338_/A vdd NOR2X1
XSFILL23400x26050 gnd vdd FILL
X_12522_ _12522_/A vdd _12521_/Y gnd _12522_/Y vdd OAI21X1
XFILL_4__9795_ gnd vdd FILL
XFILL_0_BUFX2_insert227 gnd vdd FILL
X_16290_ _16287_/Y _16290_/B _16289_/Y gnd _16296_/A vdd NAND3X1
XFILL_6_BUFX2_insert981 gnd vdd FILL
XFILL_2__7830_ gnd vdd FILL
XFILL_0_BUFX2_insert238 gnd vdd FILL
XFILL_0_BUFX2_insert249 gnd vdd FILL
XFILL_4__8746_ gnd vdd FILL
X_15241_ _15241_/A _15240_/Y _15234_/Y gnd _15241_/Y vdd NAND3X1
X_12453_ _12451_/Y vdd _12453_/C gnd _12539_/D vdd OAI21X1
XFILL_1__8968_ gnd vdd FILL
XSFILL89240x42050 gnd vdd FILL
XSFILL53880x19050 gnd vdd FILL
XFILL_2__7761_ gnd vdd FILL
XFILL_5__7470_ gnd vdd FILL
X_11404_ _11404_/A _11569_/B gnd _11404_/Y vdd NOR2X1
X_12384_ _12382_/Y _12395_/A _12384_/C gnd _12384_/Y vdd OAI21X1
XFILL_2__9500_ gnd vdd FILL
X_15172_ _15172_/A gnd _15390_/B vdd INVX8
XFILL_2__7692_ gnd vdd FILL
XFILL_4__7628_ gnd vdd FILL
XFILL_1__8899_ gnd vdd FILL
X_14123_ _14123_/A gnd _14125_/A vdd INVX1
X_11335_ _12204_/Y _12334_/Y _11202_/Y gnd _11336_/C vdd OAI21X1
XFILL_1__10430_ gnd vdd FILL
XSFILL28920x57050 gnd vdd FILL
XFILL_4__11590_ gnd vdd FILL
XSFILL94360x33050 gnd vdd FILL
XFILL_5__9140_ gnd vdd FILL
XFILL_5__11900_ gnd vdd FILL
XFILL_4__7559_ gnd vdd FILL
X_14054_ _13879_/B _14052_/Y _13857_/B _14053_/Y gnd _14055_/A vdd OAI22X1
X_11266_ _11266_/A _11076_/Y gnd _11732_/A vdd NOR2X1
XFILL_4__10541_ gnd vdd FILL
XFILL_5__12880_ gnd vdd FILL
XFILL_2__11720_ gnd vdd FILL
XFILL_2__9362_ gnd vdd FILL
XFILL_1__10361_ gnd vdd FILL
X_10217_ _10159_/A _7020_/CLK _9964_/R vdd _10217_/D gnd vdd DFFSR
X_13005_ _6888_/A gnd _13005_/Y vdd INVX1
XFILL_5__11831_ gnd vdd FILL
XFILL_4__13260_ gnd vdd FILL
XFILL_1__12100_ gnd vdd FILL
XFILL_2__8313_ gnd vdd FILL
X_11197_ _11197_/A _11191_/Y gnd _11419_/A vdd NOR2X1
XFILL_2__11651_ gnd vdd FILL
XFILL_2__9293_ gnd vdd FILL
XFILL_4__9229_ gnd vdd FILL
XFILL_1__13080_ gnd vdd FILL
XFILL_3__13990_ gnd vdd FILL
XFILL_0__12830_ gnd vdd FILL
XFILL_3_BUFX2_insert860 gnd vdd FILL
XFILL_1__10292_ gnd vdd FILL
XFILL_5__14550_ gnd vdd FILL
X_10148_ _10127_/A _8356_/B gnd _10148_/Y vdd NAND2X1
XFILL_4__12211_ gnd vdd FILL
XFILL_3_BUFX2_insert871 gnd vdd FILL
XFILL_5__11762_ gnd vdd FILL
XFILL_1__12031_ gnd vdd FILL
XFILL_2__14370_ gnd vdd FILL
XFILL_3_BUFX2_insert882 gnd vdd FILL
XFILL_2__8244_ gnd vdd FILL
XFILL_3_BUFX2_insert893 gnd vdd FILL
XFILL_2__11582_ gnd vdd FILL
XFILL_0__12761_ gnd vdd FILL
XFILL_5__13501_ gnd vdd FILL
XFILL_5__14481_ gnd vdd FILL
XSFILL34120x57050 gnd vdd FILL
XFILL_4__12142_ gnd vdd FILL
X_10079_ _13900_/A _9823_/CLK _9056_/R vdd _10079_/D gnd vdd DFFSR
X_14956_ _13621_/B _14956_/B _10869_/Q _14956_/D gnd _14956_/Y vdd AOI22X1
XFILL_2__13321_ gnd vdd FILL
XFILL_2__10533_ gnd vdd FILL
XFILL_0__14500_ gnd vdd FILL
XFILL_3__15660_ gnd vdd FILL
XFILL_5__11693_ gnd vdd FILL
XFILL_3__12872_ gnd vdd FILL
XFILL_0__11712_ gnd vdd FILL
XFILL_0__15480_ gnd vdd FILL
XFILL_5__16220_ gnd vdd FILL
XFILL_5__13432_ gnd vdd FILL
X_13907_ _13907_/A _13907_/B _13907_/C gnd _13908_/A vdd NAND3X1
XFILL_3__14611_ gnd vdd FILL
XFILL_0__7190_ gnd vdd FILL
XFILL_5__10644_ gnd vdd FILL
XSFILL89320x22050 gnd vdd FILL
XFILL_2__13252_ gnd vdd FILL
XFILL_2__16040_ gnd vdd FILL
XFILL_4__12073_ gnd vdd FILL
XFILL_3__11823_ gnd vdd FILL
X_14887_ _14885_/Y _14887_/B _13876_/C _14886_/Y gnd _14887_/Y vdd OAI22X1
XFILL_3__15591_ gnd vdd FILL
XFILL_0__14431_ gnd vdd FILL
XFILL_1__13982_ gnd vdd FILL
XFILL_0__11643_ gnd vdd FILL
XFILL_5__16151_ gnd vdd FILL
XFILL_5__13363_ gnd vdd FILL
XFILL_4__15901_ gnd vdd FILL
X_13838_ _13838_/A _13838_/B _13837_/Y gnd _13839_/B vdd NAND3X1
XFILL_2__12203_ gnd vdd FILL
XFILL_4__11024_ gnd vdd FILL
XFILL_5__10575_ gnd vdd FILL
XFILL_3__14542_ gnd vdd FILL
XFILL_2__7057_ gnd vdd FILL
XFILL112280x67050 gnd vdd FILL
XFILL_1__15721_ gnd vdd FILL
XFILL_3__11754_ gnd vdd FILL
XFILL_2__10395_ gnd vdd FILL
XFILL_0__14362_ gnd vdd FILL
XFILL_5__15102_ gnd vdd FILL
XFILL_5__8855_ gnd vdd FILL
XFILL_5__12314_ gnd vdd FILL
XFILL_0__11574_ gnd vdd FILL
XFILL_5__16082_ gnd vdd FILL
XFILL_5__13294_ gnd vdd FILL
X_13769_ _13769_/A _13769_/B _13769_/C gnd _13772_/C vdd NOR3X1
XFILL_2__12134_ gnd vdd FILL
XFILL_0__16101_ gnd vdd FILL
XFILL_4__15832_ gnd vdd FILL
XFILL_6__11865_ gnd vdd FILL
XSFILL94440x13050 gnd vdd FILL
XFILL_3__10705_ gnd vdd FILL
XFILL_0__13313_ gnd vdd FILL
XFILL_3__14473_ gnd vdd FILL
XFILL_3__7870_ gnd vdd FILL
XFILL_1__15652_ gnd vdd FILL
XFILL_5__7806_ gnd vdd FILL
XFILL_3__11685_ gnd vdd FILL
XFILL_0__10525_ gnd vdd FILL
XFILL_1__12864_ gnd vdd FILL
X_15508_ _16293_/A _7137_/Q _15380_/C _9879_/A gnd _15508_/Y vdd AOI22X1
XFILL_5__15033_ gnd vdd FILL
XFILL_0__14293_ gnd vdd FILL
XFILL_0__9900_ gnd vdd FILL
XFILL_6__10816_ gnd vdd FILL
XFILL_3__16212_ gnd vdd FILL
XFILL_5__12245_ gnd vdd FILL
XFILL_5__8786_ gnd vdd FILL
XFILL_3__13424_ gnd vdd FILL
XFILL_4__15763_ gnd vdd FILL
XFILL_3__10636_ gnd vdd FILL
XSFILL79240x74050 gnd vdd FILL
XFILL_1__14603_ gnd vdd FILL
XFILL_0__16032_ gnd vdd FILL
XFILL_4__12975_ gnd vdd FILL
XFILL_2__12065_ gnd vdd FILL
XFILL_1__11815_ gnd vdd FILL
XFILL_0__13244_ gnd vdd FILL
XFILL_0_BUFX2_insert750 gnd vdd FILL
XFILL_5__7737_ gnd vdd FILL
XFILL_1__15583_ gnd vdd FILL
XFILL_4__14714_ gnd vdd FILL
X_15439_ _15439_/A _15916_/B _15439_/C gnd _15440_/B vdd AOI21X1
XFILL_0_BUFX2_insert761 gnd vdd FILL
XFILL_4__11926_ gnd vdd FILL
XFILL_3__16143_ gnd vdd FILL
X_8370_ _8426_/Q gnd _8370_/Y vdd INVX1
XFILL_5__12176_ gnd vdd FILL
XFILL_2__11016_ gnd vdd FILL
XFILL_3__13355_ gnd vdd FILL
XFILL_4__15694_ gnd vdd FILL
XFILL_3__9540_ gnd vdd FILL
XFILL_0_BUFX2_insert772 gnd vdd FILL
XSFILL28840x7050 gnd vdd FILL
XFILL_2__7959_ gnd vdd FILL
XFILL_1__14534_ gnd vdd FILL
XFILL_0_BUFX2_insert783 gnd vdd FILL
XSFILL18680x27050 gnd vdd FILL
XFILL_1__11746_ gnd vdd FILL
XFILL_3__10567_ gnd vdd FILL
XSFILL114440x83050 gnd vdd FILL
XFILL_0_BUFX2_insert794 gnd vdd FILL
X_7321_ _7319_/Y _7336_/B _7320_/Y gnd _7393_/D vdd OAI21X1
XFILL_0__10387_ gnd vdd FILL
XFILL_5__11127_ gnd vdd FILL
XFILL_4__14645_ gnd vdd FILL
XFILL_0__9762_ gnd vdd FILL
XFILL_3__12306_ gnd vdd FILL
XFILL_0__6974_ gnd vdd FILL
XFILL_2__15824_ gnd vdd FILL
XFILL_3__16074_ gnd vdd FILL
XFILL_4__11857_ gnd vdd FILL
XFILL_3__9471_ gnd vdd FILL
XFILL_3__13286_ gnd vdd FILL
XFILL_1__14465_ gnd vdd FILL
XSFILL84360x65050 gnd vdd FILL
XFILL_5__9407_ gnd vdd FILL
XFILL_0__12126_ gnd vdd FILL
XFILL_3__10498_ gnd vdd FILL
XSFILL33720x30050 gnd vdd FILL
XFILL_1__11677_ gnd vdd FILL
XFILL_0__8713_ gnd vdd FILL
XFILL_3__15025_ gnd vdd FILL
XFILL_5__15935_ gnd vdd FILL
XFILL_4__10808_ gnd vdd FILL
XFILL_5__11058_ gnd vdd FILL
X_7252_ _7210_/A _7380_/B gnd _7253_/C vdd NAND2X1
XFILL_5__7599_ gnd vdd FILL
XFILL_1__16204_ gnd vdd FILL
XFILL_4__14576_ gnd vdd FILL
XFILL_1__13416_ gnd vdd FILL
XFILL_3__12237_ gnd vdd FILL
XFILL_2__9629_ gnd vdd FILL
XFILL_1__10628_ gnd vdd FILL
XFILL_4__11788_ gnd vdd FILL
XFILL_2__15755_ gnd vdd FILL
XSFILL59160x41050 gnd vdd FILL
XFILL_0__12057_ gnd vdd FILL
XFILL_1__14396_ gnd vdd FILL
XFILL_2__12967_ gnd vdd FILL
XFILL_5__9338_ gnd vdd FILL
XFILL_5__10009_ gnd vdd FILL
XFILL_4__16315_ gnd vdd FILL
XFILL_4__13527_ gnd vdd FILL
XFILL_0__8644_ gnd vdd FILL
X_7183_ _7184_/B _8207_/B gnd _7183_/Y vdd NAND2X1
XFILL_2__14706_ gnd vdd FILL
XFILL_5__15866_ gnd vdd FILL
XFILL_1__13347_ gnd vdd FILL
XFILL_3__8353_ gnd vdd FILL
XFILL_2__11918_ gnd vdd FILL
XFILL_3__12168_ gnd vdd FILL
XFILL_1__16135_ gnd vdd FILL
XFILL_0__11008_ gnd vdd FILL
XFILL_1__10559_ gnd vdd FILL
XFILL_2__15686_ gnd vdd FILL
XFILL_5__9269_ gnd vdd FILL
XFILL_2__12898_ gnd vdd FILL
XFILL_5__14817_ gnd vdd FILL
XFILL112360x47050 gnd vdd FILL
XFILL_4__16246_ gnd vdd FILL
XFILL_0__8575_ gnd vdd FILL
XFILL_3__7304_ gnd vdd FILL
XFILL_4__13458_ gnd vdd FILL
XFILL_3__11119_ gnd vdd FILL
XFILL_2__14637_ gnd vdd FILL
XFILL_3__12099_ gnd vdd FILL
XFILL_5__15797_ gnd vdd FILL
XFILL_1__16066_ gnd vdd FILL
XFILL_1__13278_ gnd vdd FILL
XFILL_0__15816_ gnd vdd FILL
XFILL_2__11849_ gnd vdd FILL
XFILL_4__12409_ gnd vdd FILL
XSFILL109400x72050 gnd vdd FILL
XFILL_3__15927_ gnd vdd FILL
XFILL_4__16177_ gnd vdd FILL
XFILL_1__15017_ gnd vdd FILL
XFILL_5__14748_ gnd vdd FILL
XFILL_4__13389_ gnd vdd FILL
XFILL_1__12229_ gnd vdd FILL
XFILL_3__7235_ gnd vdd FILL
XFILL_2__14568_ gnd vdd FILL
XFILL_1_BUFX2_insert6 gnd vdd FILL
XFILL_0__15747_ gnd vdd FILL
XFILL_0__12959_ gnd vdd FILL
XSFILL79320x54050 gnd vdd FILL
XFILL_4__15128_ gnd vdd FILL
XFILL_0__7457_ gnd vdd FILL
XFILL_2__16307_ gnd vdd FILL
XFILL_5__14679_ gnd vdd FILL
XFILL_2__13519_ gnd vdd FILL
XFILL_3__15858_ gnd vdd FILL
XFILL_3__7166_ gnd vdd FILL
XFILL_0__15678_ gnd vdd FILL
XFILL_2__14499_ gnd vdd FILL
XFILL_3__14809_ gnd vdd FILL
XFILL_4__15059_ gnd vdd FILL
X_9824_ _9748_/A _7530_/CLK _7523_/R vdd _9750_/Y gnd vdd DFFSR
XFILL_2__16238_ gnd vdd FILL
XSFILL114520x63050 gnd vdd FILL
XSFILL8600x17050 gnd vdd FILL
XFILL_0__14629_ gnd vdd FILL
XFILL_3__7097_ gnd vdd FILL
XFILL_3__15789_ gnd vdd FILL
XFILL_0__9127_ gnd vdd FILL
XSFILL33800x10050 gnd vdd FILL
XFILL_5__16349_ gnd vdd FILL
X_6967_ _6967_/A _6967_/B _6966_/Y gnd _6967_/Y vdd OAI21X1
X_9755_ _9737_/A _8987_/B gnd _9755_/Y vdd NAND2X1
XFILL_1__15919_ gnd vdd FILL
XFILL_2__16169_ gnd vdd FILL
XFILL_4__6930_ gnd vdd FILL
X_8706_ _8706_/A gnd _8706_/Y vdd INVX1
XFILL_6_BUFX2_insert244 gnd vdd FILL
XFILL_1__9940_ gnd vdd FILL
X_9686_ _9686_/Q _8818_/CLK _8278_/R vdd _9686_/D gnd vdd DFFSR
X_6898_ _6898_/A gnd memoryWriteData[28] vdd BUFX2
XFILL_4__6861_ gnd vdd FILL
XFILL_0__8009_ gnd vdd FILL
X_8637_ _8637_/A _8655_/B _8636_/Y gnd _8637_/Y vdd OAI21X1
XFILL_3__9807_ gnd vdd FILL
XFILL_1__9871_ gnd vdd FILL
XFILL_4__8600_ gnd vdd FILL
XFILL_5_BUFX2_insert900 gnd vdd FILL
XFILL_5_BUFX2_insert911 gnd vdd FILL
XFILL111960x20050 gnd vdd FILL
XFILL112440x27050 gnd vdd FILL
XFILL_3__7999_ gnd vdd FILL
XFILL_5_BUFX2_insert922 gnd vdd FILL
XFILL_1__8822_ gnd vdd FILL
XFILL_5_BUFX2_insert933 gnd vdd FILL
X_8568_ _8568_/A _8567_/B _8568_/C gnd _8662_/D vdd OAI21X1
XFILL_5_BUFX2_insert944 gnd vdd FILL
XFILL_5_BUFX2_insert955 gnd vdd FILL
XFILL_3__9738_ gnd vdd FILL
XFILL_4__8531_ gnd vdd FILL
XFILL_5_BUFX2_insert966 gnd vdd FILL
XFILL_5_BUFX2_insert977 gnd vdd FILL
XSFILL39000x29050 gnd vdd FILL
X_7519_ _7441_/A _7156_/CLK _7775_/R vdd _7519_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert988 gnd vdd FILL
XFILL_1__8753_ gnd vdd FILL
XFILL_5_BUFX2_insert999 gnd vdd FILL
XSFILL113720x15050 gnd vdd FILL
X_8499_ _8496_/A _9779_/B gnd _8500_/C vdd NAND2X1
XFILL_4__8462_ gnd vdd FILL
XFILL_3__9669_ gnd vdd FILL
XSFILL8600x8050 gnd vdd FILL
XFILL_1__7704_ gnd vdd FILL
X_11120_ _12171_/Y _12290_/Y gnd _11120_/Y vdd NOR2X1
XFILL_4__8393_ gnd vdd FILL
XSFILL94280x48050 gnd vdd FILL
XSFILL114600x43050 gnd vdd FILL
XFILL_1__7635_ gnd vdd FILL
XFILL_3_BUFX2_insert101 gnd vdd FILL
XFILL_4__7344_ gnd vdd FILL
X_11051_ _11731_/B _11050_/Y gnd _11055_/A vdd NOR2X1
XSFILL69080x24050 gnd vdd FILL
XFILL_1__7566_ gnd vdd FILL
X_10002_ _10054_/B _7954_/B gnd _10002_/Y vdd NAND2X1
XFILL_4__9014_ gnd vdd FILL
XFILL_1__7497_ gnd vdd FILL
XFILL_2_BUFX2_insert801 gnd vdd FILL
X_14810_ _14810_/A _14810_/B gnd _14811_/C vdd NOR2X1
XFILL_2_BUFX2_insert812 gnd vdd FILL
XFILL_2_BUFX2_insert823 gnd vdd FILL
X_15790_ _15045_/D _15790_/B _15789_/Y gnd _15790_/Y vdd OAI21X1
XFILL_1__9236_ gnd vdd FILL
XFILL_2_BUFX2_insert834 gnd vdd FILL
XFILL_2_BUFX2_insert845 gnd vdd FILL
XFILL_2_BUFX2_insert856 gnd vdd FILL
X_14741_ _14741_/A _14740_/Y gnd _14741_/Y vdd NOR2X1
X_11953_ _13145_/A gnd _11955_/A vdd INVX1
XSFILL23800x42050 gnd vdd FILL
XFILL_2_BUFX2_insert867 gnd vdd FILL
XFILL_1__9167_ gnd vdd FILL
XFILL_2_BUFX2_insert878 gnd vdd FILL
XFILL_2_BUFX2_insert889 gnd vdd FILL
XSFILL89240x37050 gnd vdd FILL
X_10904_ _10898_/Y _10920_/B gnd _16450_/A vdd NOR2X1
XFILL_5__6970_ gnd vdd FILL
XFILL_1__8118_ gnd vdd FILL
X_14672_ _9839_/Q _14712_/B _14672_/C gnd _14680_/B vdd AOI21X1
X_11884_ _11884_/A gnd _11884_/Y vdd INVX1
XFILL_4__9916_ gnd vdd FILL
XFILL_1__9098_ gnd vdd FILL
XFILL_2__9980_ gnd vdd FILL
X_16411_ _16268_/A gnd _16413_/A vdd INVX1
X_13623_ _8959_/A gnd _13623_/Y vdd INVX1
XFILL_5__10360_ gnd vdd FILL
XSFILL38840x2050 gnd vdd FILL
X_10835_ _10869_/Q gnd _10837_/A vdd INVX1
XFILL_2__10180_ gnd vdd FILL
XFILL_5__8640_ gnd vdd FILL
XBUFX2_insert800 _13334_/Y gnd _9398_/A vdd BUFX2
XFILL_4__9847_ gnd vdd FILL
XSFILL94360x28050 gnd vdd FILL
X_16342_ _16342_/A gnd _16344_/A vdd INVX1
XBUFX2_insert811 _13329_/Y gnd _8996_/A vdd BUFX2
XBUFX2_insert822 _13287_/Y gnd _7472_/A vdd BUFX2
X_13554_ _14456_/C _15163_/B _14030_/C _13554_/D gnd _13558_/A vdd OAI22X1
X_10766_ _10846_/Q gnd _10766_/Y vdd INVX1
XBUFX2_insert833 _15046_/Y gnd _15841_/C vdd BUFX2
XFILL_5__10291_ gnd vdd FILL
XFILL_0__10310_ gnd vdd FILL
XFILL_2__8862_ gnd vdd FILL
XBUFX2_insert844 _12375_/Y gnd _7061_/B vdd BUFX2
XFILL_3__11470_ gnd vdd FILL
X_12505_ _12409_/A gnd _12505_/Y vdd INVX1
XFILL_5__12030_ gnd vdd FILL
XBUFX2_insert855 _13269_/Y gnd _7124_/A vdd BUFX2
XFILL_0__11290_ gnd vdd FILL
XFILL_5__8571_ gnd vdd FILL
XFILL_4__9778_ gnd vdd FILL
XBUFX2_insert866 _13438_/Y gnd _14557_/C vdd BUFX2
X_16273_ _16272_/Y _16271_/Y gnd _16273_/Y vdd NOR2X1
XFILL_3__10421_ gnd vdd FILL
XFILL_4__12760_ gnd vdd FILL
XBUFX2_insert877 _15019_/Y gnd _16026_/D vdd BUFX2
XFILL_1__11600_ gnd vdd FILL
XFILL_2__7813_ gnd vdd FILL
X_13485_ _13485_/A _14956_/D _14065_/C _15122_/A gnd _13489_/A vdd AOI22X1
X_10697_ _10697_/A _10681_/A _10696_/Y gnd _10697_/Y vdd OAI21X1
XBUFX2_insert888 _13432_/Y gnd _14377_/B vdd BUFX2
XFILL_0__10241_ gnd vdd FILL
XFILL_1__12580_ gnd vdd FILL
XFILL_4__8729_ gnd vdd FILL
XBUFX2_insert899 _15072_/Y gnd _15563_/C vdd BUFX2
XFILL_6__10532_ gnd vdd FILL
X_15224_ _15045_/D gnd _15383_/D vdd INVX8
X_12436_ _12436_/A gnd _12436_/Y vdd INVX1
XFILL_4__11711_ gnd vdd FILL
XFILL_3__13140_ gnd vdd FILL
XFILL_2__7744_ gnd vdd FILL
XFILL_1__11531_ gnd vdd FILL
XFILL_2__13870_ gnd vdd FILL
XFILL_0__10172_ gnd vdd FILL
XFILL_5__7453_ gnd vdd FILL
X_15155_ _15155_/A _15154_/Y gnd _15156_/B vdd NOR2X1
XFILL_4__14430_ gnd vdd FILL
X_12367_ _11912_/B gnd _12367_/Y vdd INVX1
XFILL_4__11642_ gnd vdd FILL
XFILL_1__14250_ gnd vdd FILL
XFILL_5__13981_ gnd vdd FILL
XFILL_3__10283_ gnd vdd FILL
XFILL_1__11462_ gnd vdd FILL
XFILL_2__7675_ gnd vdd FILL
XFILL_0__14980_ gnd vdd FILL
X_14106_ _14106_/A _14106_/B _14106_/C gnd _14121_/A vdd NAND3X1
XFILL_5__15720_ gnd vdd FILL
X_11318_ _11637_/B _11433_/C _11318_/C gnd _11513_/A vdd AOI21X1
XSFILL59080x56050 gnd vdd FILL
XFILL_3__12022_ gnd vdd FILL
XFILL_2__9414_ gnd vdd FILL
X_15086_ _15726_/A gnd _15086_/Y vdd INVX8
XFILL_4__14361_ gnd vdd FILL
XSFILL89320x17050 gnd vdd FILL
X_12298_ _12298_/A _12298_/B _12297_/Y gnd _12298_/Y vdd NAND3X1
XFILL_2__15540_ gnd vdd FILL
XFILL_1__10413_ gnd vdd FILL
XFILL_4__11573_ gnd vdd FILL
XFILL_5__9123_ gnd vdd FILL
XFILL_2__12752_ gnd vdd FILL
XFILL_1__14181_ gnd vdd FILL
XFILL_0__13931_ gnd vdd FILL
XFILL_4__16100_ gnd vdd FILL
XFILL_1__11393_ gnd vdd FILL
XFILL_4__13312_ gnd vdd FILL
X_14037_ _8418_/Q _14037_/B _14037_/C _6938_/A gnd _14037_/Y vdd AOI22X1
X_11249_ _11025_/A _12129_/Y gnd _11249_/Y vdd XOR2X1
XFILL_5__15651_ gnd vdd FILL
XFILL_4__10524_ gnd vdd FILL
XFILL_5__12863_ gnd vdd FILL
XFILL_2__9345_ gnd vdd FILL
XFILL_1__13132_ gnd vdd FILL
XFILL_2__11703_ gnd vdd FILL
XFILL_4__14292_ gnd vdd FILL
XFILL_2__15471_ gnd vdd FILL
XFILL_0__13862_ gnd vdd FILL
XFILL_0__8360_ gnd vdd FILL
XFILL_5__14602_ gnd vdd FILL
XFILL_4__16031_ gnd vdd FILL
XSFILL109880x44050 gnd vdd FILL
XFILL_5__11814_ gnd vdd FILL
XFILL_4__13243_ gnd vdd FILL
XFILL_5__15582_ gnd vdd FILL
XFILL_2__14422_ gnd vdd FILL
XFILL_2__9276_ gnd vdd FILL
XFILL_5__8005_ gnd vdd FILL
XFILL_2__11634_ gnd vdd FILL
XFILL_0__15601_ gnd vdd FILL
XFILL_3__13973_ gnd vdd FILL
XFILL_1__10275_ gnd vdd FILL
XFILL_0__7311_ gnd vdd FILL
XFILL_0__13793_ gnd vdd FILL
XFILL_3_BUFX2_insert690 gnd vdd FILL
XFILL_3__15712_ gnd vdd FILL
XFILL_5__14533_ gnd vdd FILL
XFILL_5__11745_ gnd vdd FILL
XFILL_2__8227_ gnd vdd FILL
X_15988_ _15988_/A _15987_/Y gnd _15994_/A vdd NOR2X1
XFILL_1__12014_ gnd vdd FILL
XFILL_4__13174_ gnd vdd FILL
XSFILL79240x69050 gnd vdd FILL
XFILL_0__15532_ gnd vdd FILL
XFILL_2__14353_ gnd vdd FILL
XFILL_4__10386_ gnd vdd FILL
XFILL_2__11565_ gnd vdd FILL
XFILL_0__12744_ gnd vdd FILL
XFILL_0__7242_ gnd vdd FILL
XFILL_6__15823_ gnd vdd FILL
XFILL_5__14464_ gnd vdd FILL
XFILL_4__12125_ gnd vdd FILL
X_14939_ _14939_/A _14931_/Y _14938_/Y gnd _14952_/B vdd NAND3X1
XFILL_2__13304_ gnd vdd FILL
X_7870_ _7918_/Q gnd _7872_/A vdd INVX1
XFILL_3__15643_ gnd vdd FILL
XFILL_5__11676_ gnd vdd FILL
XFILL_2__10516_ gnd vdd FILL
XFILL_3__12855_ gnd vdd FILL
XFILL_0__15463_ gnd vdd FILL
XFILL_2__11496_ gnd vdd FILL
XFILL_2__14284_ gnd vdd FILL
XFILL_5__16203_ gnd vdd FILL
XFILL_5__13415_ gnd vdd FILL
XSFILL114440x78050 gnd vdd FILL
XFILL_5__10627_ gnd vdd FILL
XFILL_0__7173_ gnd vdd FILL
XFILL_2__16023_ gnd vdd FILL
XFILL_2__7109_ gnd vdd FILL
XFILL_4__12056_ gnd vdd FILL
XFILL_5__14395_ gnd vdd FILL
XFILL_3__11806_ gnd vdd FILL
XFILL_2__13235_ gnd vdd FILL
XFILL_2__10447_ gnd vdd FILL
XFILL_3__15574_ gnd vdd FILL
XFILL_0__14414_ gnd vdd FILL
XFILL_3__12786_ gnd vdd FILL
XFILL_3__8971_ gnd vdd FILL
XFILL_2__8089_ gnd vdd FILL
XFILL_5__8907_ gnd vdd FILL
XFILL_0__11626_ gnd vdd FILL
XSFILL33720x25050 gnd vdd FILL
XFILL_0__15394_ gnd vdd FILL
XFILL_1__13965_ gnd vdd FILL
XFILL_5__13346_ gnd vdd FILL
XFILL_6__11917_ gnd vdd FILL
X_9540_ _9584_/Q gnd _9540_/Y vdd INVX1
XFILL_5__9887_ gnd vdd FILL
XFILL_4__11007_ gnd vdd FILL
XFILL_5__16134_ gnd vdd FILL
XFILL_5__10558_ gnd vdd FILL
XFILL_6__15685_ gnd vdd FILL
XFILL_3__14525_ gnd vdd FILL
XFILL_2__13166_ gnd vdd FILL
XFILL_1__15704_ gnd vdd FILL
XFILL_3__11737_ gnd vdd FILL
XFILL_2__10378_ gnd vdd FILL
XFILL_0__14345_ gnd vdd FILL
XFILL_1__12916_ gnd vdd FILL
XSFILL59160x36050 gnd vdd FILL
XFILL_5__8838_ gnd vdd FILL
XFILL_0__11557_ gnd vdd FILL
XFILL_6__14636_ gnd vdd FILL
XFILL_5__16065_ gnd vdd FILL
XFILL_1__13896_ gnd vdd FILL
X_9471_ _9561_/Q gnd _9471_/Y vdd INVX1
XFILL_5__13277_ gnd vdd FILL
XFILL_2__12117_ gnd vdd FILL
XFILL_4__15815_ gnd vdd FILL
XFILL_3__14456_ gnd vdd FILL
XFILL_5__10489_ gnd vdd FILL
XFILL_0__10508_ gnd vdd FILL
XFILL_1__15635_ gnd vdd FILL
XFILL_2__13097_ gnd vdd FILL
XFILL_3__7853_ gnd vdd FILL
XFILL_3__11668_ gnd vdd FILL
XFILL_1__12847_ gnd vdd FILL
XFILL_0__14276_ gnd vdd FILL
X_8422_ _8422_/Q _8947_/CLK _8038_/R vdd _8422_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert229 gnd vdd FILL
XFILL_5__12228_ gnd vdd FILL
XFILL_5__15016_ gnd vdd FILL
XFILL_5__8769_ gnd vdd FILL
XFILL_0__11488_ gnd vdd FILL
XFILL_3__13407_ gnd vdd FILL
XFILL_0__16015_ gnd vdd FILL
XFILL_2__12048_ gnd vdd FILL
XFILL_4__15746_ gnd vdd FILL
XFILL_3__10619_ gnd vdd FILL
XFILL_4__12958_ gnd vdd FILL
XFILL_0__13227_ gnd vdd FILL
XFILL_6__9301_ gnd vdd FILL
XFILL_3__14387_ gnd vdd FILL
XSFILL109960x24050 gnd vdd FILL
XFILL_1__12778_ gnd vdd FILL
XFILL_1__15566_ gnd vdd FILL
XFILL_0__10439_ gnd vdd FILL
XFILL_3__11599_ gnd vdd FILL
XFILL_0_BUFX2_insert580 gnd vdd FILL
XFILL_4__11909_ gnd vdd FILL
X_8353_ _8333_/B _9633_/B gnd _8354_/C vdd NAND2X1
XFILL_0_BUFX2_insert591 gnd vdd FILL
XFILL_5__12159_ gnd vdd FILL
XFILL_3__16126_ gnd vdd FILL
XFILL_3__13338_ gnd vdd FILL
XFILL_4__15677_ gnd vdd FILL
XFILL_6__14498_ gnd vdd FILL
XFILL_3__9523_ gnd vdd FILL
XFILL_4_BUFX2_insert907 gnd vdd FILL
XFILL_1__14517_ gnd vdd FILL
XFILL_4__12889_ gnd vdd FILL
XFILL_1__11729_ gnd vdd FILL
XFILL_4_BUFX2_insert918 gnd vdd FILL
XFILL_0__13158_ gnd vdd FILL
XFILL_6__16237_ gnd vdd FILL
X_7304_ _7388_/Q gnd _7304_/Y vdd INVX1
XFILL_1__15497_ gnd vdd FILL
XFILL_6__13449_ gnd vdd FILL
XFILL_4_BUFX2_insert929 gnd vdd FILL
XFILL_0__9745_ gnd vdd FILL
XFILL_4__14628_ gnd vdd FILL
X_8284_ _8200_/A _9436_/CLK _9454_/R vdd _8202_/Y gnd vdd DFFSR
XFILL_0__6957_ gnd vdd FILL
XFILL_2__15807_ gnd vdd FILL
XFILL_3__16057_ gnd vdd FILL
XFILL_3__13269_ gnd vdd FILL
XFILL_0__12109_ gnd vdd FILL
XFILL_1__14448_ gnd vdd FILL
XFILL_0__13089_ gnd vdd FILL
XFILL_2__13999_ gnd vdd FILL
XFILL_5__15918_ gnd vdd FILL
XFILL_3__15008_ gnd vdd FILL
X_7235_ _7233_/Y _7166_/B _7235_/C gnd _7279_/D vdd OAI21X1
XFILL_4__14559_ gnd vdd FILL
XFILL_0__9676_ gnd vdd FILL
XFILL_3__8405_ gnd vdd FILL
XFILL_0__6888_ gnd vdd FILL
XFILL_2__15738_ gnd vdd FILL
XFILL_1__14379_ gnd vdd FILL
XFILL_3__9385_ gnd vdd FILL
XFILL_1__7420_ gnd vdd FILL
XFILL_0__8627_ gnd vdd FILL
XFILL_6__16099_ gnd vdd FILL
XFILL_5__15849_ gnd vdd FILL
X_7166_ _7164_/Y _7166_/B _7165_/Y gnd _7256_/D vdd OAI21X1
XFILL_3__8336_ gnd vdd FILL
XFILL_1__16118_ gnd vdd FILL
XFILL_2__15669_ gnd vdd FILL
XFILL_4__16229_ gnd vdd FILL
XFILL_1__7351_ gnd vdd FILL
X_7097_ _7068_/B _8889_/B gnd _7098_/C vdd NAND2X1
XFILL_3__8267_ gnd vdd FILL
XFILL_1__16049_ gnd vdd FILL
XFILL_4__7060_ gnd vdd FILL
XFILL_2_BUFX2_insert108 gnd vdd FILL
XFILL_0__7509_ gnd vdd FILL
XFILL_0__8489_ gnd vdd FILL
XFILL_3__7218_ gnd vdd FILL
XFILL_3__8198_ gnd vdd FILL
XFILL_1__9021_ gnd vdd FILL
XSFILL23720x57050 gnd vdd FILL
XFILL_1_BUFX2_insert808 gnd vdd FILL
X_9807_ _9805_/Y _9789_/B _9807_/C gnd _9843_/D vdd OAI21X1
XFILL_1_BUFX2_insert819 gnd vdd FILL
X_7999_ _7937_/B _7231_/B gnd _8000_/C vdd NAND2X1
XFILL_4__7962_ gnd vdd FILL
XFILL_6__8878_ gnd vdd FILL
X_9738_ _9738_/A _9737_/A _9738_/C gnd _9738_/Y vdd OAI21X1
XFILL_4__6913_ gnd vdd FILL
XBUFX2_insert107 _10925_/Y gnd _11900_/A vdd BUFX2
XFILL_4__7893_ gnd vdd FILL
XFILL_6__7829_ gnd vdd FILL
X_10620_ _15130_/B gnd _10622_/A vdd INVX1
XFILL_1__9923_ gnd vdd FILL
XFILL_4__9632_ gnd vdd FILL
X_9669_ _9625_/B _7877_/B gnd _9670_/C vdd NAND2X1
XFILL_4__6844_ gnd vdd FILL
X_10551_ _10551_/A _10535_/A _10551_/C gnd _10551_/Y vdd OAI21X1
XFILL_5_BUFX2_insert730 gnd vdd FILL
XFILL_1__9854_ gnd vdd FILL
XSFILL69080x19050 gnd vdd FILL
XFILL_5_BUFX2_insert741 gnd vdd FILL
XFILL_5_BUFX2_insert752 gnd vdd FILL
X_13270_ _13270_/A gnd _13284_/B vdd INVX1
X_10482_ _10442_/A _7129_/CLK _8542_/R vdd _10482_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert763 gnd vdd FILL
XSFILL109480x3050 gnd vdd FILL
XFILL_5_BUFX2_insert774 gnd vdd FILL
XFILL_5_BUFX2_insert785 gnd vdd FILL
XFILL_1__9785_ gnd vdd FILL
XFILL_4__8514_ gnd vdd FILL
XFILL_1__6997_ gnd vdd FILL
XFILL_4__9494_ gnd vdd FILL
XFILL_5_BUFX2_insert796 gnd vdd FILL
X_12221_ _6871_/A _12237_/B _12269_/C gnd gnd _12222_/C vdd AOI22X1
XFILL_1__8736_ gnd vdd FILL
XFILL_4__8445_ gnd vdd FILL
X_12152_ _12150_/B _12859_/A gnd _12153_/C vdd NAND2X1
XSFILL23800x37050 gnd vdd FILL
XFILL_2__7460_ gnd vdd FILL
XSFILL104360x50 gnd vdd FILL
X_11103_ _12310_/Y gnd _11103_/Y vdd INVX1
XSFILL33960x81050 gnd vdd FILL
XFILL_4__8376_ gnd vdd FILL
X_12083_ _11999_/A _12083_/B _11999_/C gnd _12086_/A vdd NAND3X1
XFILL_1__7618_ gnd vdd FILL
XFILL_1__8598_ gnd vdd FILL
XFILL_4__7327_ gnd vdd FILL
X_15911_ _10293_/A _15178_/C gnd _15917_/A vdd NAND2X1
X_11034_ _11785_/A _11034_/B _11034_/C gnd _11041_/A vdd AOI21X1
XSFILL89640x53050 gnd vdd FILL
XFILL_2__9130_ gnd vdd FILL
XFILL_1__7549_ gnd vdd FILL
XSFILL13480x27050 gnd vdd FILL
X_15842_ _15842_/A _14370_/D _15842_/C _15644_/D gnd _15843_/A vdd OAI22X1
XFILL_4__10240_ gnd vdd FILL
XFILL_2_BUFX2_insert620 gnd vdd FILL
XFILL_3__10970_ gnd vdd FILL
XFILL_1__10060_ gnd vdd FILL
XFILL_2_BUFX2_insert631 gnd vdd FILL
XFILL_0__10790_ gnd vdd FILL
XFILL_2_BUFX2_insert642 gnd vdd FILL
XFILL_5__11530_ gnd vdd FILL
XFILL_4__7189_ gnd vdd FILL
XFILL_1__9219_ gnd vdd FILL
XFILL_2__8012_ gnd vdd FILL
XFILL_2_BUFX2_insert653 gnd vdd FILL
X_15773_ _7084_/A gnd _15773_/Y vdd INVX1
XFILL_4__10171_ gnd vdd FILL
X_12985_ vdd _12985_/B gnd _12986_/C vdd NAND2X1
XFILL_2_BUFX2_insert664 gnd vdd FILL
XFILL_2__11350_ gnd vdd FILL
XFILL_2_BUFX2_insert675 gnd vdd FILL
XFILL_5__9810_ gnd vdd FILL
X_14724_ _8772_/A gnd _14725_/B vdd INVX1
XFILL_2_BUFX2_insert686 gnd vdd FILL
XFILL_2__10301_ gnd vdd FILL
X_11936_ _11934_/B _11936_/B gnd _11937_/C vdd NAND2X1
XFILL_2_BUFX2_insert697 gnd vdd FILL
XFILL_5__11461_ gnd vdd FILL
XFILL_3__12640_ gnd vdd FILL
XSFILL28920x70050 gnd vdd FILL
XFILL_2__11281_ gnd vdd FILL
XFILL_5__9741_ gnd vdd FILL
XFILL_0__12460_ gnd vdd FILL
XFILL_5__10412_ gnd vdd FILL
XFILL_5__6953_ gnd vdd FILL
XFILL_2__13020_ gnd vdd FILL
XFILL_5__14180_ gnd vdd FILL
X_14655_ _8943_/Q _14482_/B _13854_/B _9281_/A gnd _14655_/Y vdd AOI22X1
XFILL_4__13930_ gnd vdd FILL
XFILL_2__10232_ gnd vdd FILL
XFILL_5_BUFX2_insert13 gnd vdd FILL
X_11867_ _12077_/A _12065_/A gnd _11868_/B vdd NOR2X1
XFILL_5__11392_ gnd vdd FILL
XFILL_3__12571_ gnd vdd FILL
XFILL_0__11411_ gnd vdd FILL
XFILL_5_BUFX2_insert24 gnd vdd FILL
XFILL_5_BUFX2_insert35 gnd vdd FILL
XFILL_1__10962_ gnd vdd FILL
XFILL_1__13750_ gnd vdd FILL
XFILL_0__12391_ gnd vdd FILL
X_13606_ _14615_/B gnd _13853_/B vdd INVX4
XFILL_5__13131_ gnd vdd FILL
XFILL_5__9672_ gnd vdd FILL
XFILL_6__11702_ gnd vdd FILL
XFILL_5_BUFX2_insert46 gnd vdd FILL
XFILL_5__6884_ gnd vdd FILL
XFILL_3__14310_ gnd vdd FILL
X_10818_ _10773_/A _6978_/B gnd _10818_/Y vdd NAND2X1
XFILL_6__15470_ gnd vdd FILL
XFILL_5_BUFX2_insert57 gnd vdd FILL
XFILL_4__13861_ gnd vdd FILL
X_14586_ _14456_/C _15997_/C _14849_/B _15996_/B gnd _14586_/Y vdd OAI22X1
XFILL_3__11522_ gnd vdd FILL
XFILL_2__8914_ gnd vdd FILL
XFILL_1__12701_ gnd vdd FILL
XFILL_0__14130_ gnd vdd FILL
XFILL_5_BUFX2_insert68 gnd vdd FILL
XFILL_2__10163_ gnd vdd FILL
XFILL_3__15290_ gnd vdd FILL
X_11798_ _11796_/Y _11797_/Y _11798_/C gnd _11798_/Y vdd OAI21X1
XFILL_5_BUFX2_insert79 gnd vdd FILL
XBUFX2_insert630 _13465_/Y gnd _13850_/B vdd BUFX2
XFILL_1__13681_ gnd vdd FILL
XFILL_2__9894_ gnd vdd FILL
XFILL_5__8623_ gnd vdd FILL
XFILL_0__11342_ gnd vdd FILL
XSFILL99480x56050 gnd vdd FILL
XFILL_1__10893_ gnd vdd FILL
XFILL_6__14421_ gnd vdd FILL
XBUFX2_insert641 _12438_/Y gnd _9172_/B vdd BUFX2
X_16325_ gnd gnd gnd _16325_/Y vdd NAND2X1
XBUFX2_insert652 _12429_/Y gnd _7499_/B vdd BUFX2
XSFILL49320x28050 gnd vdd FILL
XFILL_4__15600_ gnd vdd FILL
X_13537_ _13537_/A gnd _13537_/Y vdd INVX1
XFILL_3__14241_ gnd vdd FILL
XFILL_5__10274_ gnd vdd FILL
X_10749_ _10809_/A _7037_/B gnd _10749_/Y vdd NAND2X1
XBUFX2_insert663 _11364_/Y gnd _11509_/B vdd BUFX2
XFILL_1__12632_ gnd vdd FILL
XFILL_4__13792_ gnd vdd FILL
XFILL_2__8845_ gnd vdd FILL
XFILL_3__11453_ gnd vdd FILL
XFILL_1__15420_ gnd vdd FILL
XSFILL59480x72050 gnd vdd FILL
XFILL_0__14061_ gnd vdd FILL
XBUFX2_insert674 _15064_/Y gnd _15792_/B vdd BUFX2
XFILL_2__14971_ gnd vdd FILL
XFILL_5__12013_ gnd vdd FILL
XBUFX2_insert685 _13459_/Y gnd _13461_/C vdd BUFX2
XFILL_0__11273_ gnd vdd FILL
XBUFX2_insert696 _13362_/Y gnd _10505_/A vdd BUFX2
XFILL_4__15531_ gnd vdd FILL
XFILL_6__11564_ gnd vdd FILL
X_16256_ _14904_/A _16099_/B _16099_/C _16255_/Y gnd _16257_/A vdd OAI22X1
XFILL_4__12743_ gnd vdd FILL
XFILL_3__10404_ gnd vdd FILL
X_13468_ _8950_/A gnd _13468_/Y vdd INVX1
XFILL_0__7860_ gnd vdd FILL
XFILL_3__14172_ gnd vdd FILL
XFILL_2__13922_ gnd vdd FILL
XFILL_0__13012_ gnd vdd FILL
XFILL_1__15351_ gnd vdd FILL
XFILL_5__7505_ gnd vdd FILL
XFILL_2__8776_ gnd vdd FILL
XFILL_3__11384_ gnd vdd FILL
X_15207_ _15207_/A _15187_/Y _15206_/Y gnd _15208_/B vdd NOR3X1
XFILL_5__8485_ gnd vdd FILL
X_12419_ _12419_/A _12642_/A gnd _12420_/C vdd NAND2X1
XSFILL53960x12050 gnd vdd FILL
XSFILL13800x69050 gnd vdd FILL
X_16187_ _16187_/A gnd _16187_/Y vdd INVX1
XFILL_3__13123_ gnd vdd FILL
XFILL_4__15462_ gnd vdd FILL
XFILL_6__14283_ gnd vdd FILL
X_13399_ _13395_/Y _14865_/B _13587_/C _13399_/D gnd _13399_/Y vdd OAI22X1
XFILL_2__7727_ gnd vdd FILL
XFILL_1__11514_ gnd vdd FILL
XFILL_1__14302_ gnd vdd FILL
XFILL_2__13853_ gnd vdd FILL
XSFILL28600x29050 gnd vdd FILL
XFILL_1__15282_ gnd vdd FILL
XFILL_5__7436_ gnd vdd FILL
XFILL_6__16022_ gnd vdd FILL
XFILL_1__12494_ gnd vdd FILL
XFILL_0__10155_ gnd vdd FILL
XFILL_6__13234_ gnd vdd FILL
XFILL_0__9530_ gnd vdd FILL
X_15138_ _8408_/Q _15978_/B _15978_/C _8536_/Q gnd _15143_/B vdd AOI22X1
XFILL_4__14413_ gnd vdd FILL
XFILL_4__11625_ gnd vdd FILL
XFILL112280x80050 gnd vdd FILL
XFILL_4__15393_ gnd vdd FILL
XFILL_1__14233_ gnd vdd FILL
XFILL_3__10266_ gnd vdd FILL
XFILL_5__13964_ gnd vdd FILL
XFILL_1__11445_ gnd vdd FILL
XSFILL54040x21050 gnd vdd FILL
XFILL_2__13784_ gnd vdd FILL
XFILL_5__15703_ gnd vdd FILL
X_7020_ _7020_/Q _7020_/CLK _9580_/R vdd _6970_/Y gnd vdd DFFSR
XFILL_0__14963_ gnd vdd FILL
XFILL_5__7367_ gnd vdd FILL
XFILL_2__10996_ gnd vdd FILL
XFILL_3__12005_ gnd vdd FILL
X_15069_ _14986_/A _16037_/B _15024_/C gnd _15069_/Y vdd NAND3X1
XFILL_4__14344_ gnd vdd FILL
XFILL_5__12915_ gnd vdd FILL
XFILL_2__15523_ gnd vdd FILL
XFILL_4__11556_ gnd vdd FILL
XFILL_2__12735_ gnd vdd FILL
XFILL_1__14164_ gnd vdd FILL
XFILL_3__10197_ gnd vdd FILL
XFILL_5__9106_ gnd vdd FILL
XFILL_5__13895_ gnd vdd FILL
XFILL_3__9170_ gnd vdd FILL
XFILL_2__7589_ gnd vdd FILL
XFILL_0__13914_ gnd vdd FILL
XFILL_1__11376_ gnd vdd FILL
XFILL_6__12116_ gnd vdd FILL
XFILL_0__14894_ gnd vdd FILL
XFILL_4__10507_ gnd vdd FILL
XFILL_5__7298_ gnd vdd FILL
XFILL_5__15634_ gnd vdd FILL
XSFILL43880x64050 gnd vdd FILL
XFILL_3__8121_ gnd vdd FILL
XFILL_5__12846_ gnd vdd FILL
XFILL_1__13115_ gnd vdd FILL
XFILL_0__9392_ gnd vdd FILL
XFILL_4__14275_ gnd vdd FILL
XFILL_4__11487_ gnd vdd FILL
XFILL_2__15454_ gnd vdd FILL
XFILL_5__9037_ gnd vdd FILL
XFILL_0__13845_ gnd vdd FILL
XFILL_1__14095_ gnd vdd FILL
XFILL_4__16014_ gnd vdd FILL
XFILL_4__13226_ gnd vdd FILL
XFILL_0__8343_ gnd vdd FILL
XFILL_5__12777_ gnd vdd FILL
XFILL_4__10438_ gnd vdd FILL
XFILL_5__15565_ gnd vdd FILL
XFILL_2__14405_ gnd vdd FILL
X_8971_ _8971_/A gnd _8971_/Y vdd INVX1
XSFILL18680x40050 gnd vdd FILL
XSFILL99560x36050 gnd vdd FILL
XFILL_1__13046_ gnd vdd FILL
XFILL_2__9259_ gnd vdd FILL
XFILL_3__13956_ gnd vdd FILL
XFILL_2__11617_ gnd vdd FILL
XFILL_2__15385_ gnd vdd FILL
XFILL_1__10258_ gnd vdd FILL
XFILL_0__13776_ gnd vdd FILL
XFILL_2__12597_ gnd vdd FILL
XSFILL74200x34050 gnd vdd FILL
XFILL_6__9850_ gnd vdd FILL
XFILL_5__14516_ gnd vdd FILL
XFILL_0__10988_ gnd vdd FILL
X_7922_ _7922_/Q _7662_/CLK _8166_/R vdd _7922_/D gnd vdd DFFSR
XFILL_4__13157_ gnd vdd FILL
XFILL_3__12907_ gnd vdd FILL
XFILL_5__11728_ gnd vdd FILL
XFILL_0__8274_ gnd vdd FILL
XFILL_4__10369_ gnd vdd FILL
XFILL_2__14336_ gnd vdd FILL
XFILL_5__15496_ gnd vdd FILL
XFILL_0__12727_ gnd vdd FILL
XFILL_3__13887_ gnd vdd FILL
XFILL_0__15515_ gnd vdd FILL
XFILL_2__11548_ gnd vdd FILL
XFILL_1__10189_ gnd vdd FILL
XFILL_0__7225_ gnd vdd FILL
XFILL_4__12108_ gnd vdd FILL
XSFILL49000x10050 gnd vdd FILL
XFILL_3__15626_ gnd vdd FILL
X_7853_ _7800_/B _7853_/B gnd _7854_/C vdd NAND2X1
XFILL_5__11659_ gnd vdd FILL
XFILL_5__14447_ gnd vdd FILL
XFILL_4__13088_ gnd vdd FILL
XFILL_3__12838_ gnd vdd FILL
XFILL112440x4050 gnd vdd FILL
XFILL_0__15446_ gnd vdd FILL
XFILL_2__14267_ gnd vdd FILL
XFILL_0__12658_ gnd vdd FILL
XFILL_2__11479_ gnd vdd FILL
XFILL_1__14997_ gnd vdd FILL
XFILL_5__9939_ gnd vdd FILL
XFILL_2__16006_ gnd vdd FILL
XFILL_4__12039_ gnd vdd FILL
XFILL_0_CLKBUF1_insert208 gnd vdd FILL
XFILL_2__13218_ gnd vdd FILL
XFILL_3__15557_ gnd vdd FILL
X_7784_ _7724_/A _7016_/CLK _8424_/R vdd _7784_/D gnd vdd DFFSR
XFILL_5__14378_ gnd vdd FILL
XFILL_3__12769_ gnd vdd FILL
XFILL_0_CLKBUF1_insert219 gnd vdd FILL
XFILL_0__11609_ gnd vdd FILL
XFILL_3__8954_ gnd vdd FILL
XFILL_2__14198_ gnd vdd FILL
XFILL_0__15377_ gnd vdd FILL
XFILL_1__13948_ gnd vdd FILL
XFILL_0__12589_ gnd vdd FILL
XFILL112360x60050 gnd vdd FILL
XFILL_5__16117_ gnd vdd FILL
XFILL_5__13329_ gnd vdd FILL
XFILL_3__14508_ gnd vdd FILL
XFILL_0__7087_ gnd vdd FILL
X_9523_ _9529_/A _9907_/B gnd _9524_/C vdd NAND2X1
XFILL_2__13149_ gnd vdd FILL
XFILL_0__14328_ gnd vdd FILL
XFILL_3__15488_ gnd vdd FILL
XFILL_3__8885_ gnd vdd FILL
XSFILL74120x6050 gnd vdd FILL
XFILL_1__13879_ gnd vdd FILL
XFILL_1__6920_ gnd vdd FILL
X_9454_ _9454_/Q _7662_/CLK _9454_/R vdd _9454_/D gnd vdd DFFSR
XFILL_5__16048_ gnd vdd FILL
XFILL_6__8594_ gnd vdd FILL
XFILL_3__14439_ gnd vdd FILL
XFILL_1__15618_ gnd vdd FILL
XFILL_3__7836_ gnd vdd FILL
XFILL_0__14259_ gnd vdd FILL
XSFILL114120x55050 gnd vdd FILL
XSFILL43960x44050 gnd vdd FILL
XFILL_6__7545_ gnd vdd FILL
X_8405_ _8403_/Y _8365_/A _8404_/Y gnd _8437_/D vdd OAI21X1
XFILL_4__15729_ gnd vdd FILL
XFILL_1__6851_ gnd vdd FILL
X_9385_ _9385_/A gnd _9387_/A vdd INVX1
XFILL_1__15549_ gnd vdd FILL
XFILL_4_BUFX2_insert704 gnd vdd FILL
X_8336_ _8334_/Y _8321_/B _8336_/C gnd _8414_/D vdd OAI21X1
XFILL_4_BUFX2_insert715 gnd vdd FILL
XFILL_3__16109_ gnd vdd FILL
XSFILL18760x20050 gnd vdd FILL
XFILL_4_BUFX2_insert726 gnd vdd FILL
XFILL_3__9506_ gnd vdd FILL
XSFILL8600x30050 gnd vdd FILL
XFILL_0__7989_ gnd vdd FILL
XSFILL44040x53050 gnd vdd FILL
XFILL_4_BUFX2_insert737 gnd vdd FILL
XFILL_4_BUFX2_insert748 gnd vdd FILL
XFILL_3__7698_ gnd vdd FILL
XFILL_0__9728_ gnd vdd FILL
XFILL_1__8521_ gnd vdd FILL
XFILL_4_BUFX2_insert759 gnd vdd FILL
X_8267_ _8249_/A _7243_/B gnd _8267_/Y vdd NAND2X1
XFILL_4__8230_ gnd vdd FILL
XFILL_6__9146_ gnd vdd FILL
X_7218_ _7274_/Q gnd _7220_/A vdd INVX1
XFILL_0__9659_ gnd vdd FILL
XFILL_1__8452_ gnd vdd FILL
XSFILL23880x11050 gnd vdd FILL
XFILL112040x19050 gnd vdd FILL
X_8198_ _8237_/A _7558_/B gnd _8199_/C vdd NAND2X1
XFILL_3__9368_ gnd vdd FILL
XSFILL78920x17050 gnd vdd FILL
X_7149_ _7149_/Q _8947_/CLK _9069_/R vdd _7101_/Y gnd vdd DFFSR
XFILL_3__8319_ gnd vdd FILL
XFILL_1__8383_ gnd vdd FILL
XSFILL38920x33050 gnd vdd FILL
XFILL_4__7112_ gnd vdd FILL
XFILL112440x40050 gnd vdd FILL
XFILL_4__8092_ gnd vdd FILL
XSFILL64200x66050 gnd vdd FILL
XFILL_3__9299_ gnd vdd FILL
XFILL_1__7334_ gnd vdd FILL
XFILL_4__7043_ gnd vdd FILL
XSFILL94680x59050 gnd vdd FILL
XSFILL3640x73050 gnd vdd FILL
XSFILL68840x69050 gnd vdd FILL
XFILL_1__9004_ gnd vdd FILL
XFILL_1_BUFX2_insert605 gnd vdd FILL
X_12770_ _12770_/A gnd _12770_/Y vdd INVX1
XFILL_1_BUFX2_insert616 gnd vdd FILL
XFILL_1__7196_ gnd vdd FILL
XSFILL3720x1050 gnd vdd FILL
XFILL_6__9979_ gnd vdd FILL
XFILL_1_BUFX2_insert627 gnd vdd FILL
XSFILL94280x61050 gnd vdd FILL
XFILL_4__8994_ gnd vdd FILL
XFILL_1_BUFX2_insert638 gnd vdd FILL
X_11721_ _11743_/A _11704_/C _11721_/C gnd _11727_/C vdd NAND3X1
XFILL_1_BUFX2_insert649 gnd vdd FILL
XFILL_4__7945_ gnd vdd FILL
X_14440_ _6962_/A gnd _15870_/D vdd INVX1
X_11652_ _11448_/B gnd _11654_/B vdd INVX1
XSFILL89880x50 gnd vdd FILL
XFILL_2__6960_ gnd vdd FILL
XSFILL103640x80050 gnd vdd FILL
X_10603_ _14454_/A _9195_/CLK _9963_/R vdd _10551_/Y gnd vdd DFFSR
XFILL_4__7876_ gnd vdd FILL
XFILL_1__9906_ gnd vdd FILL
X_14371_ _8297_/Q gnd _15842_/C vdd INVX1
X_11583_ _11583_/A _11153_/Y _11129_/Y gnd _11589_/C vdd OAI21X1
XFILL_4__9615_ gnd vdd FILL
XFILL_2__6891_ gnd vdd FILL
X_16110_ _16109_/Y _16110_/B gnd _16110_/Y vdd NOR2X1
X_13322_ _13321_/Y gnd _13322_/Y vdd INVX1
X_10534_ _10534_/A gnd _10536_/A vdd INVX1
XFILL_2__8630_ gnd vdd FILL
XFILL_5_BUFX2_insert560 gnd vdd FILL
XFILL_4__9546_ gnd vdd FILL
XFILL_5_BUFX2_insert571 gnd vdd FILL
XFILL_5_BUFX2_insert582 gnd vdd FILL
XSFILL49640x64050 gnd vdd FILL
X_16041_ _16041_/A _15683_/B _15376_/B _14641_/Y gnd _16041_/Y vdd OAI22X1
X_13253_ _13253_/A _13252_/Y gnd _13297_/A vdd NAND2X1
X_10465_ _10465_/Q _8560_/CLK _9313_/R vdd _10465_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert593 gnd vdd FILL
XFILL_1__9768_ gnd vdd FILL
XSFILL89240x50050 gnd vdd FILL
XSFILL18760x1050 gnd vdd FILL
XSFILL74120x50 gnd vdd FILL
XFILL_6__10300_ gnd vdd FILL
XFILL_5__8270_ gnd vdd FILL
X_12204_ _12204_/A _12179_/A _12204_/C gnd _12204_/Y vdd OAI21X1
XFILL_4__9477_ gnd vdd FILL
XFILL_3__10120_ gnd vdd FILL
XFILL_1__8719_ gnd vdd FILL
X_13184_ _11914_/A _13184_/CLK _8033_/R vdd _13184_/D gnd vdd DFFSR
X_10396_ _10396_/A _10395_/A _10396_/C gnd _10466_/D vdd OAI21X1
XFILL_5__7221_ gnd vdd FILL
XFILL_2__8492_ gnd vdd FILL
X_12135_ _12135_/A _12134_/A _12135_/C gnd _12135_/Y vdd OAI21X1
XFILL_4__11410_ gnd vdd FILL
XFILL_5__10961_ gnd vdd FILL
XFILL_3__10051_ gnd vdd FILL
XFILL_4__12390_ gnd vdd FILL
XFILL_2__7443_ gnd vdd FILL
XFILL_1__11230_ gnd vdd FILL
XSFILL94360x41050 gnd vdd FILL
XFILL_2__10781_ gnd vdd FILL
XFILL_2_CLKBUF1_insert130 gnd vdd FILL
XFILL_4__8359_ gnd vdd FILL
XFILL_0__11960_ gnd vdd FILL
XFILL_2_CLKBUF1_insert141 gnd vdd FILL
XFILL_5__12700_ gnd vdd FILL
XFILL_2_CLKBUF1_insert152 gnd vdd FILL
XFILL_5__13680_ gnd vdd FILL
X_12066_ _12066_/A _12066_/B _12066_/C gnd _13137_/B vdd NAND3X1
XFILL_4__11341_ gnd vdd FILL
XFILL_2__12520_ gnd vdd FILL
XFILL_5__10892_ gnd vdd FILL
XFILL_2_CLKBUF1_insert163 gnd vdd FILL
XFILL_0__10911_ gnd vdd FILL
XFILL_2__7374_ gnd vdd FILL
XFILL_1__11161_ gnd vdd FILL
XFILL_2_CLKBUF1_insert174 gnd vdd FILL
XFILL_2_CLKBUF1_insert185 gnd vdd FILL
XFILL_5__12631_ gnd vdd FILL
XFILL_2_CLKBUF1_insert196 gnd vdd FILL
XFILL_0__11891_ gnd vdd FILL
XFILL_5__7083_ gnd vdd FILL
X_11017_ _11384_/A _12138_/Y gnd _11383_/A vdd AND2X2
XFILL_3__13810_ gnd vdd FILL
XFILL_4__14060_ gnd vdd FILL
XFILL_2__9113_ gnd vdd FILL
XFILL_1__10112_ gnd vdd FILL
XFILL_4__11272_ gnd vdd FILL
XFILL_0__13630_ gnd vdd FILL
XFILL_2__12451_ gnd vdd FILL
XFILL_3__14790_ gnd vdd FILL
XFILL_1__11092_ gnd vdd FILL
X_15825_ _15824_/Y _15819_/Y gnd _15825_/Y vdd NOR2X1
XFILL_4__13011_ gnd vdd FILL
XFILL_5__15350_ gnd vdd FILL
XFILL_3__13741_ gnd vdd FILL
XSFILL74120x49050 gnd vdd FILL
XFILL_2_BUFX2_insert450 gnd vdd FILL
XFILL_2__11402_ gnd vdd FILL
XFILL_2__9044_ gnd vdd FILL
XFILL_3__10953_ gnd vdd FILL
XFILL_1__10043_ gnd vdd FILL
XFILL_2__15170_ gnd vdd FILL
XFILL_2__12382_ gnd vdd FILL
XFILL_1__14920_ gnd vdd FILL
XFILL_2_BUFX2_insert461 gnd vdd FILL
XBUFX2_insert7 _13280_/Y gnd _7366_/B vdd BUFX2
XFILL_0__13561_ gnd vdd FILL
XFILL_2_BUFX2_insert472 gnd vdd FILL
XFILL_5__14301_ gnd vdd FILL
XFILL_5__11513_ gnd vdd FILL
XFILL_0__10773_ gnd vdd FILL
XFILL_2_BUFX2_insert483 gnd vdd FILL
XFILL_5__15281_ gnd vdd FILL
X_15756_ _15544_/A _15755_/Y _14278_/B _15756_/D gnd _15756_/Y vdd OAI22X1
XFILL_0__15300_ gnd vdd FILL
XFILL_5__12493_ gnd vdd FILL
XFILL_4__10154_ gnd vdd FILL
XFILL_2_BUFX2_insert494 gnd vdd FILL
XFILL_2__14121_ gnd vdd FILL
X_12968_ _12968_/A vdd _12967_/Y gnd _13052_/D vdd OAI21X1
XFILL_0__12512_ gnd vdd FILL
XFILL_3__13672_ gnd vdd FILL
XSFILL84120x1050 gnd vdd FILL
XFILL_2__11333_ gnd vdd FILL
XFILL_1__14851_ gnd vdd FILL
XFILL_3__10884_ gnd vdd FILL
XFILL_0__16280_ gnd vdd FILL
X_14707_ _8432_/Q gnd _14708_/A vdd INVX1
XFILL_0__13492_ gnd vdd FILL
XFILL_5__14232_ gnd vdd FILL
XFILL_3__15411_ gnd vdd FILL
X_11919_ _11919_/A _11900_/A _11919_/C gnd _6848_/A vdd OAI21X1
XFILL_5__7985_ gnd vdd FILL
XFILL_5__11444_ gnd vdd FILL
XFILL_3__12623_ gnd vdd FILL
X_15687_ _15687_/A _14207_/Y _14208_/A _16018_/C gnd _15687_/Y vdd OAI22X1
XFILL_1__13802_ gnd vdd FILL
XFILL_0__15231_ gnd vdd FILL
XFILL_2__14052_ gnd vdd FILL
XFILL_3__16391_ gnd vdd FILL
XFILL_4__14962_ gnd vdd FILL
XFILL_2__11264_ gnd vdd FILL
X_12899_ vdd _12899_/B gnd _12900_/C vdd NAND2X1
XFILL_0__12443_ gnd vdd FILL
XFILL_5__6936_ gnd vdd FILL
XFILL_1__11994_ gnd vdd FILL
XFILL_5__9724_ gnd vdd FILL
XFILL_1__14782_ gnd vdd FILL
X_14638_ _8558_/Q gnd _14638_/Y vdd INVX1
XFILL_5__14163_ gnd vdd FILL
XFILL_3__15342_ gnd vdd FILL
XFILL_2__13003_ gnd vdd FILL
XFILL_4__13913_ gnd vdd FILL
XFILL_5__11375_ gnd vdd FILL
XFILL_4__14893_ gnd vdd FILL
XFILL112280x75050 gnd vdd FILL
XFILL_0__15162_ gnd vdd FILL
XFILL_1__13733_ gnd vdd FILL
XSFILL54040x16050 gnd vdd FILL
XFILL_2__11195_ gnd vdd FILL
XFILL_1__10945_ gnd vdd FILL
XFILL_5__9655_ gnd vdd FILL
XFILL_0__12374_ gnd vdd FILL
XFILL_5__13114_ gnd vdd FILL
XFILL_5__6867_ gnd vdd FILL
XFILL_0__8961_ gnd vdd FILL
X_14569_ _14560_/Y _14561_/Y _14568_/Y gnd _14570_/A vdd NAND3X1
XFILL_3__11505_ gnd vdd FILL
XFILL_5__14094_ gnd vdd FILL
XFILL_4__13844_ gnd vdd FILL
XFILL_2__10146_ gnd vdd FILL
XFILL_0__14113_ gnd vdd FILL
XFILL_3__15273_ gnd vdd FILL
XFILL_3__12485_ gnd vdd FILL
XBUFX2_insert460 _15044_/Y gnd _15197_/C vdd BUFX2
XFILL_2__9877_ gnd vdd FILL
XFILL_5__8606_ gnd vdd FILL
XFILL_0__11325_ gnd vdd FILL
XBUFX2_insert471 _13318_/Y gnd _8333_/B vdd BUFX2
XFILL_1__13664_ gnd vdd FILL
X_16308_ _16308_/A _16307_/Y gnd _16308_/Y vdd NAND2X1
XFILL_1__10876_ gnd vdd FILL
XFILL_0__15093_ gnd vdd FILL
XBUFX2_insert482 _14979_/Y gnd _14989_/A vdd BUFX2
XFILL_5__13045_ gnd vdd FILL
XFILL_3__14224_ gnd vdd FILL
XFILL_5__10257_ gnd vdd FILL
XSFILL79240x82050 gnd vdd FILL
XFILL_1__15403_ gnd vdd FILL
XBUFX2_insert493 _13471_/Y gnd _14593_/C vdd BUFX2
XFILL_4__13775_ gnd vdd FILL
XSFILL43880x59050 gnd vdd FILL
XFILL_0__8892_ gnd vdd FILL
XFILL_3__7621_ gnd vdd FILL
XFILL_3__11436_ gnd vdd FILL
XFILL_2__8828_ gnd vdd FILL
XFILL_1__12615_ gnd vdd FILL
XFILL_0__14044_ gnd vdd FILL
XFILL_2__14954_ gnd vdd FILL
XFILL_1__16383_ gnd vdd FILL
XFILL_1__13595_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1075 gnd vdd FILL
XFILL_0__11256_ gnd vdd FILL
X_16239_ _10573_/A gnd _16239_/Y vdd INVX1
XFILL_0__7843_ gnd vdd FILL
XFILL_4__12726_ gnd vdd FILL
XFILL_4__15514_ gnd vdd FILL
X_9170_ _9170_/A _9170_/B _9170_/C gnd _9204_/D vdd OAI21X1
XFILL_5__10188_ gnd vdd FILL
XFILL_3__14155_ gnd vdd FILL
XFILL_2__13905_ gnd vdd FILL
XFILL_3__7552_ gnd vdd FILL
XFILL_2__8759_ gnd vdd FILL
XFILL_1__15334_ gnd vdd FILL
XSFILL18680x35050 gnd vdd FILL
XFILL_3__11367_ gnd vdd FILL
XSFILL8520x45050 gnd vdd FILL
XFILL_2__14885_ gnd vdd FILL
X_8121_ _8142_/A _8377_/B gnd _8122_/C vdd NAND2X1
XSFILL74200x29050 gnd vdd FILL
XFILL_5__8468_ gnd vdd FILL
XFILL_0__11187_ gnd vdd FILL
XFILL_3__13106_ gnd vdd FILL
XFILL_4__12657_ gnd vdd FILL
XFILL_3__10318_ gnd vdd FILL
XFILL_4__15445_ gnd vdd FILL
XSFILL84360x73050 gnd vdd FILL
XFILL_2__13836_ gnd vdd FILL
XFILL_5__14996_ gnd vdd FILL
XFILL_3__14086_ gnd vdd FILL
XFILL_0__10138_ gnd vdd FILL
XFILL_3__7483_ gnd vdd FILL
XFILL_1__12477_ gnd vdd FILL
XFILL_3__11298_ gnd vdd FILL
XFILL_1__15265_ gnd vdd FILL
XFILL_5__7419_ gnd vdd FILL
XFILL_0__9513_ gnd vdd FILL
XFILL_6__10429_ gnd vdd FILL
XFILL_5__8399_ gnd vdd FILL
XFILL_0__15995_ gnd vdd FILL
XFILL_4__11608_ gnd vdd FILL
X_8052_ _8052_/Q _8297_/CLK _7796_/R vdd _8052_/D gnd vdd DFFSR
XFILL_4__15376_ gnd vdd FILL
XFILL_3__13037_ gnd vdd FILL
XFILL_5__13947_ gnd vdd FILL
XFILL_3__9222_ gnd vdd FILL
XFILL_4__12588_ gnd vdd FILL
XFILL_3__10249_ gnd vdd FILL
XFILL_1__14216_ gnd vdd FILL
XFILL_1__11428_ gnd vdd FILL
XFILL_2__13767_ gnd vdd FILL
XFILL_1_BUFX2_insert11 gnd vdd FILL
XFILL_2__10979_ gnd vdd FILL
XFILL_1__15196_ gnd vdd FILL
XFILL_0__10069_ gnd vdd FILL
XFILL_0__14946_ gnd vdd FILL
X_7003_ _6917_/A _8792_/CLK _9048_/R vdd _6919_/Y gnd vdd DFFSR
XFILL_4__14327_ gnd vdd FILL
XFILL_1_BUFX2_insert22 gnd vdd FILL
XFILL_2__15506_ gnd vdd FILL
XFILL_4__11539_ gnd vdd FILL
XSFILL109560x16050 gnd vdd FILL
XFILL_1_BUFX2_insert33 gnd vdd FILL
XFILL_5__13878_ gnd vdd FILL
XFILL_2__12718_ gnd vdd FILL
XFILL_3__9153_ gnd vdd FILL
XFILL_1__14147_ gnd vdd FILL
XFILL_1_BUFX2_insert44 gnd vdd FILL
XFILL_1__11359_ gnd vdd FILL
XFILL_1_BUFX2_insert55 gnd vdd FILL
XSFILL38840x48050 gnd vdd FILL
XFILL_2__13698_ gnd vdd FILL
XFILL_0__14877_ gnd vdd FILL
XFILL112360x55050 gnd vdd FILL
XFILL_5__15617_ gnd vdd FILL
XFILL_1_BUFX2_insert66 gnd vdd FILL
XFILL_4__14258_ gnd vdd FILL
XFILL_3__8104_ gnd vdd FILL
XFILL_6__13079_ gnd vdd FILL
XFILL_1_BUFX2_insert77 gnd vdd FILL
XFILL_0__9375_ gnd vdd FILL
XFILL_5__12829_ gnd vdd FILL
XFILL_1_BUFX2_insert88 gnd vdd FILL
XFILL_2__15437_ gnd vdd FILL
XFILL_2__12649_ gnd vdd FILL
XFILL_3__14988_ gnd vdd FILL
XFILL_1__14078_ gnd vdd FILL
XFILL_3__9084_ gnd vdd FILL
XFILL_0__13828_ gnd vdd FILL
XFILL_1_BUFX2_insert99 gnd vdd FILL
XFILL_4__13209_ gnd vdd FILL
XFILL_0__8326_ gnd vdd FILL
XSFILL109400x80050 gnd vdd FILL
XFILL_5__15548_ gnd vdd FILL
XFILL_4__14189_ gnd vdd FILL
XFILL_1__13029_ gnd vdd FILL
X_8954_ _9044_/A _6906_/B gnd _8955_/C vdd NAND2X1
XFILL_3__13939_ gnd vdd FILL
XFILL_2__15368_ gnd vdd FILL
XSFILL79320x62050 gnd vdd FILL
XFILL_0__13759_ gnd vdd FILL
XFILL_1__7050_ gnd vdd FILL
XSFILL43960x39050 gnd vdd FILL
XSFILL114920x69050 gnd vdd FILL
X_7905_ _7831_/A _9188_/CLK _9441_/R vdd _7833_/Y gnd vdd DFFSR
XFILL_0__8257_ gnd vdd FILL
XFILL_2__14319_ gnd vdd FILL
XFILL_5__15479_ gnd vdd FILL
X_8885_ _8939_/Q gnd _8887_/A vdd INVX1
XFILL_2__15299_ gnd vdd FILL
XFILL_0__7208_ gnd vdd FILL
XSFILL18760x15050 gnd vdd FILL
XSFILL114520x71050 gnd vdd FILL
X_7836_ _7836_/A _7800_/B _7836_/C gnd _7836_/Y vdd OAI21X1
XFILL_0__8188_ gnd vdd FILL
XFILL_3__15609_ gnd vdd FILL
XSFILL8600x25050 gnd vdd FILL
XSFILL44040x48050 gnd vdd FILL
XFILL_3__9986_ gnd vdd FILL
XFILL_0__15429_ gnd vdd FILL
XFILL_4__7730_ gnd vdd FILL
X_7767_ _7673_/A _8663_/CLK _7131_/R vdd _7675_/Y gnd vdd DFFSR
X_9506_ _9506_/A _9533_/B _9506_/C gnd _9572_/D vdd OAI21X1
XFILL_1__7952_ gnd vdd FILL
X_7698_ _7729_/B _7314_/B gnd _7698_/Y vdd NAND2X1
XFILL_3__8868_ gnd vdd FILL
XFILL111800x69050 gnd vdd FILL
XFILL_1__6903_ gnd vdd FILL
X_9437_ _9437_/Q _9707_/CLK _8819_/R vdd _9357_/Y gnd vdd DFFSR
XFILL_4__9400_ gnd vdd FILL
XFILL_3__7819_ gnd vdd FILL
XFILL_1__7883_ gnd vdd FILL
XSFILL38920x28050 gnd vdd FILL
XFILL112440x35050 gnd vdd FILL
XFILL_4__7592_ gnd vdd FILL
XFILL_4_BUFX2_insert501 gnd vdd FILL
XFILL_1__9622_ gnd vdd FILL
XFILL_4_BUFX2_insert512 gnd vdd FILL
X_9368_ _9356_/A _8472_/B gnd _9369_/C vdd NAND2X1
XFILL_4_BUFX2_insert523 gnd vdd FILL
X_10250_ _10248_/Y _10304_/B _10250_/C gnd _10332_/D vdd OAI21X1
XSFILL89160x65050 gnd vdd FILL
XFILL_4_BUFX2_insert534 gnd vdd FILL
XFILL_4_BUFX2_insert545 gnd vdd FILL
XSFILL39000x37050 gnd vdd FILL
X_8319_ _8409_/Q gnd _8319_/Y vdd INVX1
XFILL_4_BUFX2_insert556 gnd vdd FILL
XFILL_1__9553_ gnd vdd FILL
X_9299_ _9333_/Q gnd _9299_/Y vdd INVX1
XFILL_4_BUFX2_insert567 gnd vdd FILL
XSFILL79400x42050 gnd vdd FILL
XFILL_4__9262_ gnd vdd FILL
XFILL_4_BUFX2_insert578 gnd vdd FILL
XSFILL3640x68050 gnd vdd FILL
XFILL_1__8504_ gnd vdd FILL
X_10181_ _10169_/A _9413_/B gnd _10182_/C vdd NAND2X1
XFILL_4_BUFX2_insert589 gnd vdd FILL
XFILL_1__9484_ gnd vdd FILL
XFILL_4__8213_ gnd vdd FILL
XSFILL94280x56050 gnd vdd FILL
XSFILL114600x51050 gnd vdd FILL
XFILL_4__8144_ gnd vdd FILL
X_13940_ _13940_/A _14901_/B _14711_/B _13940_/D gnd _13940_/Y vdd OAI22X1
XSFILL69080x32050 gnd vdd FILL
XFILL_1__8366_ gnd vdd FILL
XFILL_3_CLKBUF1_insert203 gnd vdd FILL
XFILL_4__8075_ gnd vdd FILL
XFILL_3_CLKBUF1_insert214 gnd vdd FILL
X_13871_ _13871_/A _13869_/Y _13871_/C _13871_/D gnd _13872_/A vdd OAI22X1
XFILL_1__7317_ gnd vdd FILL
XFILL_2__7090_ gnd vdd FILL
X_15610_ _15610_/A _15610_/B _14791_/C gnd _15610_/Y vdd AOI21X1
X_12822_ _12788_/A _12692_/CLK _12692_/R vdd _12822_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert402 gnd vdd FILL
XFILL_1__7248_ gnd vdd FILL
XFILL_1_BUFX2_insert413 gnd vdd FILL
XFILL_1_BUFX2_insert424 gnd vdd FILL
X_15541_ _15541_/A _15541_/B gnd _15542_/C vdd NOR2X1
X_12753_ _12718_/B memoryOutData[19] gnd _12753_/Y vdd NAND2X1
XFILL_1_BUFX2_insert435 gnd vdd FILL
XFILL_1_BUFX2_insert446 gnd vdd FILL
XFILL_1__7179_ gnd vdd FILL
XSFILL89240x45050 gnd vdd FILL
XFILL_1_BUFX2_insert457 gnd vdd FILL
XFILL_1_BUFX2_insert468 gnd vdd FILL
X_11704_ _12258_/Y _11071_/Y _11704_/C gnd _11704_/Y vdd OAI21X1
XFILL_4__8977_ gnd vdd FILL
XFILL_1_BUFX2_insert479 gnd vdd FILL
X_15472_ _15472_/A _15468_/Y _15471_/Y gnd _15472_/Y vdd NAND3X1
XFILL_2__9800_ gnd vdd FILL
X_12684_ _12407_/B _12809_/CLK _12809_/R vdd _12684_/D gnd vdd DFFSR
XFILL_2__7992_ gnd vdd FILL
XFILL_4__7928_ gnd vdd FILL
X_14423_ _14412_/Y _14423_/B gnd _14450_/B vdd NOR2X1
XFILL_4__10910_ gnd vdd FILL
XFILL_2__10000_ gnd vdd FILL
XFILL_5__11160_ gnd vdd FILL
X_11635_ _11632_/Y _11635_/B gnd _11638_/A vdd NOR2X1
XFILL_1_CLKBUF1_insert1081 gnd vdd FILL
XFILL_2__9731_ gnd vdd FILL
XFILL_4__11890_ gnd vdd FILL
XFILL_2__6943_ gnd vdd FILL
XSFILL94360x36050 gnd vdd FILL
XFILL_5__10111_ gnd vdd FILL
XFILL_4__7859_ gnd vdd FILL
X_14354_ _10412_/A _14389_/B _14868_/D _9192_/Q gnd _14354_/Y vdd AOI22X1
XFILL_5__11091_ gnd vdd FILL
X_11566_ _11565_/Y _11563_/Y _11558_/Y gnd _11857_/B vdd AOI21X1
XFILL_2__9662_ gnd vdd FILL
XFILL_3__12270_ gnd vdd FILL
XFILL_0__11110_ gnd vdd FILL
XFILL_1__10661_ gnd vdd FILL
XFILL_2__6874_ gnd vdd FILL
X_13305_ _13305_/A _13305_/B _13308_/B gnd _13305_/Y vdd OAI21X1
XFILL_0__12090_ gnd vdd FILL
XFILL_5__9371_ gnd vdd FILL
XSFILL69160x12050 gnd vdd FILL
XFILL_5__10042_ gnd vdd FILL
X_10517_ _10581_/B _7317_/B gnd _10517_/Y vdd NAND2X1
XFILL_2__8613_ gnd vdd FILL
XFILL_4__13560_ gnd vdd FILL
XFILL_3__11221_ gnd vdd FILL
X_14285_ _14284_/Y _14768_/D gnd _14285_/Y vdd NOR2X1
XFILL_5_BUFX2_insert390 gnd vdd FILL
XFILL_1__12400_ gnd vdd FILL
X_11497_ _11176_/Y _11423_/B _11497_/C gnd _11503_/C vdd OAI21X1
XFILL_4__10772_ gnd vdd FILL
XFILL_5__8322_ gnd vdd FILL
XFILL_2__11951_ gnd vdd FILL
XFILL_1__13380_ gnd vdd FILL
XFILL_4__9529_ gnd vdd FILL
XFILL_2__9593_ gnd vdd FILL
XFILL_0__11041_ gnd vdd FILL
XBUFX2_insert80 _15015_/Y gnd _15449_/C vdd BUFX2
X_16024_ _16024_/A _15197_/B _15197_/C _16024_/D gnd _16024_/Y vdd OAI22X1
XBUFX2_insert91 _12357_/Y gnd _9859_/B vdd BUFX2
X_13236_ _13230_/Y _13236_/B _13235_/Y gnd _13236_/Y vdd OAI21X1
XFILL_4__12511_ gnd vdd FILL
XFILL_5__14850_ gnd vdd FILL
X_10448_ _14918_/A gnd _10450_/A vdd INVX1
XSFILL104360x21050 gnd vdd FILL
XFILL_2__10902_ gnd vdd FILL
XFILL_1__12331_ gnd vdd FILL
XFILL_3__11152_ gnd vdd FILL
XFILL_4__13491_ gnd vdd FILL
XFILL_2__14670_ gnd vdd FILL
XFILL_5__8253_ gnd vdd FILL
XFILL_2__11882_ gnd vdd FILL
XFILL_5__13801_ gnd vdd FILL
XFILL_4__15230_ gnd vdd FILL
XSFILL104600x83050 gnd vdd FILL
X_13167_ _13168_/B _13167_/B gnd _13167_/Y vdd NAND2X1
XFILL_4__12442_ gnd vdd FILL
XFILL_3__10103_ gnd vdd FILL
X_10379_ _10379_/A gnd _10379_/Y vdd INVX1
XFILL_2__13621_ gnd vdd FILL
XFILL_5__14781_ gnd vdd FILL
XFILL_5__7204_ gnd vdd FILL
XFILL_0__14800_ gnd vdd FILL
XFILL_2__8475_ gnd vdd FILL
XFILL_1__15050_ gnd vdd FILL
XFILL_3__15960_ gnd vdd FILL
XFILL_5__11993_ gnd vdd FILL
XFILL_1__12262_ gnd vdd FILL
XFILL_3__11083_ gnd vdd FILL
XFILL_2__10833_ gnd vdd FILL
XFILL_5__8184_ gnd vdd FILL
XFILL_0__15780_ gnd vdd FILL
X_12118_ _11890_/A gnd _12120_/A vdd INVX1
XFILL_0__12992_ gnd vdd FILL
XSFILL59080x64050 gnd vdd FILL
XFILL_5__13732_ gnd vdd FILL
XFILL_4__15161_ gnd vdd FILL
XSFILL89320x25050 gnd vdd FILL
XFILL_2__16340_ gnd vdd FILL
XFILL_5__10944_ gnd vdd FILL
XFILL_2__7426_ gnd vdd FILL
X_13098_ _13099_/B _13098_/B gnd _13098_/Y vdd NAND2X1
XFILL_1__14001_ gnd vdd FILL
XFILL_4__12373_ gnd vdd FILL
XFILL_3__10034_ gnd vdd FILL
XFILL_0__7490_ gnd vdd FILL
XFILL_3__14911_ gnd vdd FILL
XFILL_1__11213_ gnd vdd FILL
XFILL_2__13552_ gnd vdd FILL
XFILL_3__15891_ gnd vdd FILL
XFILL_2__10764_ gnd vdd FILL
XFILL_0__11943_ gnd vdd FILL
XFILL_0__14731_ gnd vdd FILL
XFILL_1__12193_ gnd vdd FILL
XFILL_6__10145_ gnd vdd FILL
XFILL_4__14112_ gnd vdd FILL
XFILL_5__16451_ gnd vdd FILL
X_12049_ _12485_/B _12105_/B _12001_/C gnd gnd _12049_/Y vdd AOI22X1
XFILL_4__11324_ gnd vdd FILL
XFILL_3__14842_ gnd vdd FILL
XFILL_2__12503_ gnd vdd FILL
XFILL_5__13663_ gnd vdd FILL
XFILL_5__10875_ gnd vdd FILL
XFILL_4__15092_ gnd vdd FILL
XFILL_2__7357_ gnd vdd FILL
XFILL_1__11144_ gnd vdd FILL
XFILL_2__16271_ gnd vdd FILL
XFILL_2__13483_ gnd vdd FILL
XFILL_0__11874_ gnd vdd FILL
XFILL_5__15402_ gnd vdd FILL
XFILL_5__7066_ gnd vdd FILL
XFILL_0__14662_ gnd vdd FILL
XFILL_2__10695_ gnd vdd FILL
XFILL_5__12614_ gnd vdd FILL
XFILL_4__14043_ gnd vdd FILL
XSFILL109080x33050 gnd vdd FILL
XFILL_0__9160_ gnd vdd FILL
XFILL_6__14953_ gnd vdd FILL
XFILL_5__16382_ gnd vdd FILL
XFILL_2__15222_ gnd vdd FILL
XSFILL94440x16050 gnd vdd FILL
XFILL_4__11255_ gnd vdd FILL
XFILL_2__12434_ gnd vdd FILL
XFILL_5__13594_ gnd vdd FILL
XFILL_0__16401_ gnd vdd FILL
XFILL_3__14773_ gnd vdd FILL
XFILL_0__13613_ gnd vdd FILL
XFILL_3__11985_ gnd vdd FILL
XFILL_2__7288_ gnd vdd FILL
XFILL_1__15952_ gnd vdd FILL
XFILL_1__11075_ gnd vdd FILL
XFILL_0__10825_ gnd vdd FILL
XFILL_0__14593_ gnd vdd FILL
XFILL_0__8111_ gnd vdd FILL
XFILL_6__13904_ gnd vdd FILL
XSFILL13800x82050 gnd vdd FILL
XFILL_5__15333_ gnd vdd FILL
X_15808_ _15392_/C _15806_/Y _15808_/C _15070_/C gnd _15809_/B vdd OAI22X1
XFILL_0__9091_ gnd vdd FILL
XFILL_2__9027_ gnd vdd FILL
XFILL_3__13724_ gnd vdd FILL
XFILL_3__10936_ gnd vdd FILL
XFILL_2_BUFX2_insert280 gnd vdd FILL
XFILL_2__15153_ gnd vdd FILL
XFILL_4__11186_ gnd vdd FILL
XFILL_1__14903_ gnd vdd FILL
XFILL_1__10026_ gnd vdd FILL
XFILL_2__12365_ gnd vdd FILL
XFILL_0__16332_ gnd vdd FILL
XSFILL94280x2050 gnd vdd FILL
XFILL_2_BUFX2_insert291 gnd vdd FILL
XFILL_0__13544_ gnd vdd FILL
XFILL_0__10756_ gnd vdd FILL
XFILL_1__15883_ gnd vdd FILL
XFILL_6_BUFX2_insert607 gnd vdd FILL
X_15739_ _15175_/B _10409_/A _14289_/D _15357_/B gnd _15739_/Y vdd AOI22X1
X_8670_ _8670_/Q _7781_/CLK _8670_/R vdd _8670_/D gnd vdd DFFSR
XFILL_4__10137_ gnd vdd FILL
XFILL_5__12476_ gnd vdd FILL
XFILL_5__15264_ gnd vdd FILL
XFILL_2__14104_ gnd vdd FILL
XFILL_6_BUFX2_insert618 gnd vdd FILL
XFILL_3__13655_ gnd vdd FILL
XFILL_2__11316_ gnd vdd FILL
XFILL_4__15994_ gnd vdd FILL
XFILL_1__14834_ gnd vdd FILL
XFILL_2__15084_ gnd vdd FILL
XFILL_0__13475_ gnd vdd FILL
XFILL_0__16263_ gnd vdd FILL
XFILL_2__12296_ gnd vdd FILL
XFILL_0__10687_ gnd vdd FILL
XFILL_5__14215_ gnd vdd FILL
XFILL_5__7968_ gnd vdd FILL
XFILL_5__11427_ gnd vdd FILL
XFILL_3__12606_ gnd vdd FILL
XFILL_6__13766_ gnd vdd FILL
X_7621_ _7577_/B _6981_/B gnd _7622_/C vdd NAND2X1
XFILL_5__15195_ gnd vdd FILL
XFILL_1_BUFX2_insert980 gnd vdd FILL
XFILL_2__14035_ gnd vdd FILL
XFILL_4__10068_ gnd vdd FILL
XFILL_4__14945_ gnd vdd FILL
XFILL_3__16374_ gnd vdd FILL
XFILL_3__13586_ gnd vdd FILL
XFILL_1_BUFX2_insert991 gnd vdd FILL
XFILL_0__15214_ gnd vdd FILL
XFILL_0__12426_ gnd vdd FILL
XFILL_3__9771_ gnd vdd FILL
XFILL_6__8500_ gnd vdd FILL
XFILL_2__11247_ gnd vdd FILL
XFILL_0__16194_ gnd vdd FILL
XFILL_3__10798_ gnd vdd FILL
XFILL_5__6919_ gnd vdd FILL
XFILL_3__6983_ gnd vdd FILL
XFILL_1__14765_ gnd vdd FILL
XFILL_6__12717_ gnd vdd FILL
XFILL_1__11977_ gnd vdd FILL
X_7552_ _7568_/B _9344_/B gnd _7553_/C vdd NAND2X1
XFILL_3__15325_ gnd vdd FILL
XFILL_5__14146_ gnd vdd FILL
XFILL_5__11358_ gnd vdd FILL
XFILL_0__9993_ gnd vdd FILL
XFILL_3__8722_ gnd vdd FILL
XFILL_4__14876_ gnd vdd FILL
XFILL_1__13716_ gnd vdd FILL
XFILL_2__11178_ gnd vdd FILL
XFILL_0__15145_ gnd vdd FILL
XFILL_2__9929_ gnd vdd FILL
XFILL_1__10928_ gnd vdd FILL
XFILL_0__12357_ gnd vdd FILL
XFILL_5__9638_ gnd vdd FILL
XFILL_5__10309_ gnd vdd FILL
XFILL_1__14696_ gnd vdd FILL
XFILL_5__14077_ gnd vdd FILL
X_7483_ _7533_/Q gnd _7483_/Y vdd INVX1
XFILL_4__13827_ gnd vdd FILL
XFILL_3__15256_ gnd vdd FILL
XFILL_5__11289_ gnd vdd FILL
XFILL_2__10129_ gnd vdd FILL
XFILL_3__8653_ gnd vdd FILL
XSFILL19160x60050 gnd vdd FILL
XFILL_3__12468_ gnd vdd FILL
XBUFX2_insert290 _15059_/Y gnd _15940_/B vdd BUFX2
XFILL_0__11308_ gnd vdd FILL
XFILL_2__15986_ gnd vdd FILL
XFILL_1__13647_ gnd vdd FILL
XFILL_0__15076_ gnd vdd FILL
XFILL_0__12288_ gnd vdd FILL
XFILL_5__13028_ gnd vdd FILL
XFILL_6__15367_ gnd vdd FILL
XFILL_3__14207_ gnd vdd FILL
X_9222_ _9238_/B _7558_/B gnd _9223_/C vdd NAND2X1
XFILL_0__8875_ gnd vdd FILL
XFILL_3__7604_ gnd vdd FILL
XFILL_3__11419_ gnd vdd FILL
XFILL_3__15187_ gnd vdd FILL
XFILL_4__13758_ gnd vdd FILL
XFILL_0__14027_ gnd vdd FILL
XFILL_2__14937_ gnd vdd FILL
XFILL_3__8584_ gnd vdd FILL
XFILL_3__12399_ gnd vdd FILL
XFILL_0__11239_ gnd vdd FILL
XFILL_1__16366_ gnd vdd FILL
XFILL_5_CLKBUF1_insert180 gnd vdd FILL
XFILL_1__13578_ gnd vdd FILL
XFILL_5_CLKBUF1_insert191 gnd vdd FILL
X_9153_ _9199_/Q gnd _9155_/A vdd INVX1
XFILL_0__7826_ gnd vdd FILL
XFILL_4__12709_ gnd vdd FILL
XFILL_3__14138_ gnd vdd FILL
XSFILL109400x75050 gnd vdd FILL
XFILL_1__15317_ gnd vdd FILL
XFILL_4__13689_ gnd vdd FILL
XFILL_2__14868_ gnd vdd FILL
XFILL_1__12529_ gnd vdd FILL
XSFILL8680x3050 gnd vdd FILL
XFILL_6__7244_ gnd vdd FILL
X_8104_ _8102_/Y _8142_/A _8104_/C gnd _8104_/Y vdd OAI21X1
XFILL_1__16297_ gnd vdd FILL
XSFILL79320x57050 gnd vdd FILL
XFILL_0__7757_ gnd vdd FILL
XFILL_3_BUFX2_insert508 gnd vdd FILL
XSFILL89400x3050 gnd vdd FILL
X_9084_ _9176_/Q gnd _9084_/Y vdd INVX1
XFILL_4__15428_ gnd vdd FILL
XFILL_2__13819_ gnd vdd FILL
XFILL_5__14979_ gnd vdd FILL
XFILL_3__14069_ gnd vdd FILL
XFILL_1__15248_ gnd vdd FILL
XFILL_3_BUFX2_insert519 gnd vdd FILL
XFILL_3__7466_ gnd vdd FILL
XFILL_2__14799_ gnd vdd FILL
XFILL_0__15978_ gnd vdd FILL
X_8035_ _8035_/Q _7791_/CLK _9711_/R vdd _7967_/Y gnd vdd DFFSR
XFILL_0__7688_ gnd vdd FILL
XFILL_4__15359_ gnd vdd FILL
XSFILL114520x66050 gnd vdd FILL
XFILL_1__15179_ gnd vdd FILL
XFILL_0__14929_ gnd vdd FILL
XFILL_1__8220_ gnd vdd FILL
XFILL_0__9427_ gnd vdd FILL
XFILL_3__9136_ gnd vdd FILL
XFILL_0__9358_ gnd vdd FILL
X_9986_ _9986_/A gnd _9988_/A vdd INVX1
XFILL_1__7102_ gnd vdd FILL
XFILL_0__9289_ gnd vdd FILL
X_8937_ _8879_/A _8169_/CLK _8937_/R vdd _8881_/Y gnd vdd DFFSR
XFILL_1__8082_ gnd vdd FILL
XFILL_3__8018_ gnd vdd FILL
XFILL_4__8900_ gnd vdd FILL
XFILL_4__9880_ gnd vdd FILL
XFILL_1__7033_ gnd vdd FILL
XFILL_4__8831_ gnd vdd FILL
X_8868_ _8823_/B _8868_/B gnd _8869_/C vdd NAND2X1
X_7819_ _7901_/Q gnd _7819_/Y vdd INVX1
XSFILL49160x76050 gnd vdd FILL
XFILL_0_BUFX2_insert409 gnd vdd FILL
XFILL_4__8762_ gnd vdd FILL
X_8799_ _8799_/Q _7007_/CLK _9332_/R vdd _8799_/D gnd vdd DFFSR
XFILL_6__9678_ gnd vdd FILL
XFILL_1__8984_ gnd vdd FILL
XSFILL39400x53050 gnd vdd FILL
XFILL_4__7713_ gnd vdd FILL
X_11420_ _11415_/C _11419_/Y _11414_/C gnd _11420_/Y vdd NAND3X1
XFILL_6__8629_ gnd vdd FILL
XFILL_1__7935_ gnd vdd FILL
X_11351_ _11338_/A _11348_/A gnd _11351_/Y vdd AND2X2
XSFILL69080x27050 gnd vdd FILL
XFILL_1__7866_ gnd vdd FILL
X_10302_ _10302_/A gnd _10302_/Y vdd INVX1
XFILL_4_BUFX2_insert320 gnd vdd FILL
XFILL_4__7575_ gnd vdd FILL
X_14070_ _8034_/Q gnd _14071_/D vdd INVX1
XFILL_1__9605_ gnd vdd FILL
XFILL_4_BUFX2_insert331 gnd vdd FILL
X_11282_ _12278_/Y gnd _11282_/Y vdd INVX1
XFILL_4_BUFX2_insert342 gnd vdd FILL
XFILL_4_BUFX2_insert353 gnd vdd FILL
X_13021_ vdd _13021_/B gnd _13022_/C vdd NAND2X1
XFILL_4_BUFX2_insert364 gnd vdd FILL
XFILL_4_BUFX2_insert375 gnd vdd FILL
X_10233_ _13497_/A gnd _10235_/A vdd INVX1
XFILL_1__9536_ gnd vdd FILL
XFILL_4_BUFX2_insert386 gnd vdd FILL
XFILL_4_BUFX2_insert397 gnd vdd FILL
XFILL_4__9245_ gnd vdd FILL
X_10164_ _10162_/Y _10160_/A _10164_/C gnd _10218_/D vdd OAI21X1
XSFILL23800x45050 gnd vdd FILL
XFILL_2__8260_ gnd vdd FILL
XFILL_1__9467_ gnd vdd FILL
XFILL112120x12050 gnd vdd FILL
X_10095_ _14660_/A _8815_/CLK _9056_/R vdd _10095_/D gnd vdd DFFSR
XFILL_2__7211_ gnd vdd FILL
X_14972_ _8821_/Q gnd _14974_/D vdd INVX1
XSFILL74040x82050 gnd vdd FILL
XFILL_4__8127_ gnd vdd FILL
XFILL_2__8191_ gnd vdd FILL
XFILL_1__9398_ gnd vdd FILL
X_13923_ _7953_/A gnd _13924_/D vdd INVX1
XFILL_5__10660_ gnd vdd FILL
XFILL_1__8349_ gnd vdd FILL
XFILL_4__8058_ gnd vdd FILL
X_13854_ _9310_/Q _13854_/B _13592_/D _7054_/A gnd _13854_/Y vdd AOI22X1
XFILL_4__11040_ gnd vdd FILL
XFILL_2__7073_ gnd vdd FILL
XFILL_3__11770_ gnd vdd FILL
XFILL_5__8871_ gnd vdd FILL
X_12805_ _11882_/B _7005_/CLK _12799_/R vdd _12739_/Y gnd vdd DFFSR
XFILL_5__12330_ gnd vdd FILL
XFILL_0__11590_ gnd vdd FILL
XFILL_6__11881_ gnd vdd FILL
X_13785_ _13785_/A _13843_/C _13871_/D _13783_/Y gnd _13786_/A vdd OAI22X1
XFILL_1__11900_ gnd vdd FILL
XFILL_2__12150_ gnd vdd FILL
XFILL_1_BUFX2_insert232 gnd vdd FILL
X_10997_ _10996_/Y _10997_/B gnd _10997_/Y vdd NOR2X1
XFILL_5__7822_ gnd vdd FILL
XFILL_1_BUFX2_insert243 gnd vdd FILL
XFILL_0__10541_ gnd vdd FILL
XFILL_1_BUFX2_insert254 gnd vdd FILL
X_15524_ _15524_/A _14018_/D _13999_/Y _15351_/A gnd _15528_/B vdd OAI22X1
XFILL_1__12880_ gnd vdd FILL
X_12736_ _12736_/A _12723_/A _12736_/C gnd _12736_/Y vdd OAI21X1
XFILL_1_BUFX2_insert265 gnd vdd FILL
XFILL_5__12261_ gnd vdd FILL
XFILL_6__10832_ gnd vdd FILL
XFILL_3__13440_ gnd vdd FILL
XFILL_2__11101_ gnd vdd FILL
XFILL_1_BUFX2_insert276 gnd vdd FILL
XFILL_2__12081_ gnd vdd FILL
XFILL_3__10652_ gnd vdd FILL
XFILL_4__12991_ gnd vdd FILL
XSFILL104360x16050 gnd vdd FILL
XFILL_0__13260_ gnd vdd FILL
XFILL_1_BUFX2_insert287 gnd vdd FILL
XFILL_1__11831_ gnd vdd FILL
XFILL_5__14000_ gnd vdd FILL
XFILL_1_BUFX2_insert298 gnd vdd FILL
XFILL_5__7753_ gnd vdd FILL
XFILL_5__11212_ gnd vdd FILL
XFILL_0_BUFX2_insert910 gnd vdd FILL
XFILL_6__13551_ gnd vdd FILL
X_15455_ _15440_/Y _15455_/B gnd _15455_/Y vdd NOR2X1
X_12667_ _12667_/Q _12667_/CLK _12809_/R vdd _12667_/D gnd vdd DFFSR
XFILL_4__11942_ gnd vdd FILL
XFILL_0_BUFX2_insert921 gnd vdd FILL
XFILL_4__14730_ gnd vdd FILL
XFILL_5__12192_ gnd vdd FILL
XFILL_2__11032_ gnd vdd FILL
XFILL_3__13371_ gnd vdd FILL
XFILL_0__12211_ gnd vdd FILL
XFILL_0_BUFX2_insert932 gnd vdd FILL
XFILL_2__7975_ gnd vdd FILL
XFILL_1__14550_ gnd vdd FILL
XFILL_0_BUFX2_insert943 gnd vdd FILL
X_14406_ _8938_/Q gnd _14407_/A vdd INVX1
XFILL_1__11762_ gnd vdd FILL
XFILL_0_BUFX2_insert954 gnd vdd FILL
XFILL_5__7684_ gnd vdd FILL
XFILL_5__11143_ gnd vdd FILL
X_11618_ _11618_/A _11618_/B gnd _11628_/A vdd OR2X2
XFILL_3__15110_ gnd vdd FILL
XFILL_0_BUFX2_insert965 gnd vdd FILL
X_15386_ _13859_/Y _15386_/B _15386_/C _15386_/D gnd _15386_/Y vdd OAI22X1
XFILL_3__12322_ gnd vdd FILL
XFILL_0__6990_ gnd vdd FILL
XFILL_4__11873_ gnd vdd FILL
XFILL_2__6926_ gnd vdd FILL
X_12598_ vdd memoryOutData[10] gnd _12599_/C vdd NAND2X1
XSFILL59080x59050 gnd vdd FILL
XFILL_0_BUFX2_insert976 gnd vdd FILL
XFILL_3__16090_ gnd vdd FILL
XFILL_2__15840_ gnd vdd FILL
XFILL_4__14661_ gnd vdd FILL
XFILL_1__13501_ gnd vdd FILL
XFILL_5__9423_ gnd vdd FILL
XSFILL9480x42050 gnd vdd FILL
XFILL_0__12142_ gnd vdd FILL
XFILL_0_BUFX2_insert987 gnd vdd FILL
XFILL_1__14481_ gnd vdd FILL
XSFILL99480x64050 gnd vdd FILL
XFILL_0_BUFX2_insert998 gnd vdd FILL
XFILL_1__11693_ gnd vdd FILL
XFILL_4__16400_ gnd vdd FILL
XFILL_6__12433_ gnd vdd FILL
X_14337_ _9004_/A gnd _15805_/D vdd INVX1
XFILL_4__13612_ gnd vdd FILL
XFILL_3__15041_ gnd vdd FILL
XFILL_5__15951_ gnd vdd FILL
X_11549_ _11549_/A _11546_/Y _11548_/Y gnd _12077_/A vdd NAND3X1
XFILL_5__11074_ gnd vdd FILL
XFILL_4__10824_ gnd vdd FILL
XFILL_4__14592_ gnd vdd FILL
XFILL_1__16220_ gnd vdd FILL
XFILL_2__9645_ gnd vdd FILL
XFILL_3__12253_ gnd vdd FILL
XFILL_1__13432_ gnd vdd FILL
XFILL_2__6857_ gnd vdd FILL
XFILL_2__15771_ gnd vdd FILL
XFILL_1__10644_ gnd vdd FILL
XFILL_5__9354_ gnd vdd FILL
XFILL_0__12073_ gnd vdd FILL
XFILL_2__12983_ gnd vdd FILL
XFILL_5__14902_ gnd vdd FILL
XFILL_5__10025_ gnd vdd FILL
XFILL_4__16331_ gnd vdd FILL
XFILL_3__11204_ gnd vdd FILL
XFILL_4__13543_ gnd vdd FILL
XFILL_0__8660_ gnd vdd FILL
X_14268_ _14268_/A _14865_/B _14320_/C _14268_/D gnd _14268_/Y vdd OAI22X1
XFILL_4__10755_ gnd vdd FILL
XFILL_2__14722_ gnd vdd FILL
XFILL_5__15882_ gnd vdd FILL
XFILL_0__15901_ gnd vdd FILL
XFILL_2__11934_ gnd vdd FILL
XFILL_3__12184_ gnd vdd FILL
XFILL_0__11024_ gnd vdd FILL
XFILL_1__16151_ gnd vdd FILL
XFILL_1__10575_ gnd vdd FILL
XFILL_1__13363_ gnd vdd FILL
X_16007_ _14614_/Y _15386_/C _15180_/C _14638_/Y gnd _16007_/Y vdd OAI22X1
X_13219_ _13251_/B _13219_/B _13295_/C gnd _13226_/B vdd AOI21X1
XFILL_0__7611_ gnd vdd FILL
XFILL_5__9285_ gnd vdd FILL
XSFILL13800x77050 gnd vdd FILL
XFILL_5__14833_ gnd vdd FILL
XFILL_0__8591_ gnd vdd FILL
X_14199_ _7269_/Q gnd _14199_/Y vdd INVX1
XFILL_2__8527_ gnd vdd FILL
XFILL_3__7320_ gnd vdd FILL
XFILL_4__13474_ gnd vdd FILL
XFILL_6__12295_ gnd vdd FILL
XFILL_3__11135_ gnd vdd FILL
XFILL_1__15102_ gnd vdd FILL
XFILL_4__16262_ gnd vdd FILL
XFILL_4__10686_ gnd vdd FILL
XFILL_1__12314_ gnd vdd FILL
XFILL_2__14653_ gnd vdd FILL
XFILL_1__13294_ gnd vdd FILL
XFILL_0__15832_ gnd vdd FILL
XFILL_5__8236_ gnd vdd FILL
XFILL_2__11865_ gnd vdd FILL
XFILL_1__16082_ gnd vdd FILL
XSFILL38760x81050 gnd vdd FILL
XFILL_4__15213_ gnd vdd FILL
XFILL_4__12425_ gnd vdd FILL
XFILL_0__7542_ gnd vdd FILL
XFILL_6__11246_ gnd vdd FILL
XFILL_2__13604_ gnd vdd FILL
XFILL_4__16193_ gnd vdd FILL
XFILL_5__14764_ gnd vdd FILL
XFILL_2__10816_ gnd vdd FILL
XFILL_5__11976_ gnd vdd FILL
XFILL_2__8458_ gnd vdd FILL
XFILL_1__15033_ gnd vdd FILL
XFILL_3__15943_ gnd vdd FILL
XFILL_1__12245_ gnd vdd FILL
XFILL_3__11066_ gnd vdd FILL
XFILL_3__7251_ gnd vdd FILL
XFILL_2__14584_ gnd vdd FILL
XSFILL113960x74050 gnd vdd FILL
XFILL_0__15763_ gnd vdd FILL
XFILL_2__11796_ gnd vdd FILL
XFILL_0__12975_ gnd vdd FILL
XFILL_5__13715_ gnd vdd FILL
XFILL_4__15144_ gnd vdd FILL
XFILL_5__10927_ gnd vdd FILL
XFILL_4__12356_ gnd vdd FILL
XFILL_3__10017_ gnd vdd FILL
XFILL_2__16323_ gnd vdd FILL
XFILL_0__7473_ gnd vdd FILL
XFILL_5__14695_ gnd vdd FILL
XFILL_2__13535_ gnd vdd FILL
XFILL_3__7182_ gnd vdd FILL
XFILL_5__7118_ gnd vdd FILL
XFILL_0__14714_ gnd vdd FILL
XFILL_2__8389_ gnd vdd FILL
XFILL_2__10747_ gnd vdd FILL
XFILL_1__12176_ gnd vdd FILL
XFILL_3__15874_ gnd vdd FILL
XFILL_0__11926_ gnd vdd FILL
XFILL_0__9212_ gnd vdd FILL
XFILL_0__15694_ gnd vdd FILL
XFILL_5__8098_ gnd vdd FILL
XFILL_4__11307_ gnd vdd FILL
XSFILL43880x72050 gnd vdd FILL
XFILL_5__13646_ gnd vdd FILL
XFILL_4__15075_ gnd vdd FILL
X_9840_ _9796_/A _9328_/CLK _7152_/R vdd _9798_/Y gnd vdd DFFSR
XFILL_3__14825_ gnd vdd FILL
XFILL_4__12287_ gnd vdd FILL
XFILL_1__11127_ gnd vdd FILL
XFILL_2__16254_ gnd vdd FILL
XFILL_2__13466_ gnd vdd FILL
XFILL_2__10678_ gnd vdd FILL
XFILL_0__14645_ gnd vdd FILL
XFILL_5__7049_ gnd vdd FILL
XFILL_0__11857_ gnd vdd FILL
XFILL_0__9143_ gnd vdd FILL
XFILL_4__14026_ gnd vdd FILL
XSFILL59160x39050 gnd vdd FILL
XFILL_2__15205_ gnd vdd FILL
XFILL_5__16365_ gnd vdd FILL
XFILL_4__11238_ gnd vdd FILL
XFILL_5__10789_ gnd vdd FILL
XFILL_2__12417_ gnd vdd FILL
X_9771_ _9771_/A _9770_/A _9771_/C gnd _9831_/D vdd OAI21X1
XFILL_5__13577_ gnd vdd FILL
XFILL_3__14756_ gnd vdd FILL
XFILL_2__16185_ gnd vdd FILL
XFILL_1__15935_ gnd vdd FILL
XFILL_3__11968_ gnd vdd FILL
XFILL_0__10808_ gnd vdd FILL
XFILL_1__11058_ gnd vdd FILL
X_6983_ _7025_/Q gnd _6985_/A vdd INVX1
XFILL_2__13397_ gnd vdd FILL
XSFILL74200x42050 gnd vdd FILL
XFILL_0__14576_ gnd vdd FILL
XFILL_5__15316_ gnd vdd FILL
XFILL_0__11788_ gnd vdd FILL
XFILL_5__12528_ gnd vdd FILL
XFILL111880x38050 gnd vdd FILL
X_8722_ _8753_/B _7186_/B gnd _8722_/Y vdd NAND2X1
XFILL_3__10919_ gnd vdd FILL
XFILL_1__10009_ gnd vdd FILL
XFILL_5__16296_ gnd vdd FILL
XFILL_2__15136_ gnd vdd FILL
XFILL_3__13707_ gnd vdd FILL
XFILL_4__11169_ gnd vdd FILL
XFILL_2__12348_ gnd vdd FILL
XFILL_0__16315_ gnd vdd FILL
XFILL_3__14687_ gnd vdd FILL
XFILL_0__13527_ gnd vdd FILL
XFILL_3__11899_ gnd vdd FILL
XFILL_1__15866_ gnd vdd FILL
XFILL_5__15247_ gnd vdd FILL
X_8653_ _8653_/A gnd _8655_/A vdd INVX1
XFILL_3__13638_ gnd vdd FILL
XFILL_5__12459_ gnd vdd FILL
XFILL_4__15977_ gnd vdd FILL
XFILL_1__14817_ gnd vdd FILL
XFILL_2__15067_ gnd vdd FILL
XFILL_6_BUFX2_insert459 gnd vdd FILL
XFILL_0__13458_ gnd vdd FILL
XFILL_2__12279_ gnd vdd FILL
XFILL_0__16246_ gnd vdd FILL
XFILL_1__15797_ gnd vdd FILL
X_7604_ _7604_/A _7570_/A _7604_/C gnd _7604_/Y vdd OAI21X1
XFILL_5__15178_ gnd vdd FILL
XFILL_2__14018_ gnd vdd FILL
XFILL_3__16357_ gnd vdd FILL
XFILL_4__14928_ gnd vdd FILL
X_8584_ _8668_/Q gnd _8584_/Y vdd INVX1
XFILL_3__9754_ gnd vdd FILL
XFILL_3__13569_ gnd vdd FILL
XFILL_3__6966_ gnd vdd FILL
XSFILL38840x61050 gnd vdd FILL
XFILL_0__12409_ gnd vdd FILL
XFILL_1__14748_ gnd vdd FILL
XFILL_0__16177_ gnd vdd FILL
XFILL_0__13389_ gnd vdd FILL
XFILL_4_BUFX2_insert1005 gnd vdd FILL
XFILL_4_BUFX2_insert1016 gnd vdd FILL
XFILL_5__14129_ gnd vdd FILL
XFILL_3__8705_ gnd vdd FILL
XFILL_3__15308_ gnd vdd FILL
XFILL_0__9976_ gnd vdd FILL
X_7535_ _7535_/Q _7535_/CLK _7523_/R vdd _7535_/D gnd vdd DFFSR
XFILL_4__14859_ gnd vdd FILL
XFILL_3__16288_ gnd vdd FILL
XFILL_4_BUFX2_insert1027 gnd vdd FILL
XFILL_4_BUFX2_insert1038 gnd vdd FILL
XFILL_3__9685_ gnd vdd FILL
XFILL_0__15128_ gnd vdd FILL
XFILL_4_BUFX2_insert1049 gnd vdd FILL
XFILL_3__6897_ gnd vdd FILL
XFILL_1__14679_ gnd vdd FILL
XFILL_6__15419_ gnd vdd FILL
XSFILL95000x21050 gnd vdd FILL
XFILL_1__7720_ gnd vdd FILL
XFILL_4_BUFX2_insert70 gnd vdd FILL
XFILL_6__9394_ gnd vdd FILL
XFILL_3__15239_ gnd vdd FILL
XFILL_4_BUFX2_insert81 gnd vdd FILL
X_7466_ _7470_/B _9770_/B gnd _7467_/C vdd NAND2X1
XFILL_3__8636_ gnd vdd FILL
XFILL_4_BUFX2_insert92 gnd vdd FILL
XFILL_2__15969_ gnd vdd FILL
XSFILL43960x52050 gnd vdd FILL
XFILL_0__15059_ gnd vdd FILL
XFILL_6__8345_ gnd vdd FILL
X_9205_ _9205_/Q _9205_/CLK _7285_/R vdd _9205_/D gnd vdd DFFSR
XFILL_0__8858_ gnd vdd FILL
X_7397_ _7397_/Q _7406_/CLK _9692_/R vdd _7397_/D gnd vdd DFFSR
XFILL_3__8567_ gnd vdd FILL
XFILL_4__7360_ gnd vdd FILL
XFILL_1__16349_ gnd vdd FILL
XFILL_0__7809_ gnd vdd FILL
X_9136_ _9112_/A _7856_/B gnd _9137_/C vdd NAND2X1
XSFILL44040x61050 gnd vdd FILL
XFILL_1__7582_ gnd vdd FILL
XFILL_0__8789_ gnd vdd FILL
XFILL_3_BUFX2_insert305 gnd vdd FILL
XFILL_2_BUFX2_insert1020 gnd vdd FILL
XFILL_3_BUFX2_insert316 gnd vdd FILL
XFILL111960x18050 gnd vdd FILL
XFILL_3__8498_ gnd vdd FILL
XFILL_4__7291_ gnd vdd FILL
XFILL_2_BUFX2_insert1031 gnd vdd FILL
XFILL_3_BUFX2_insert327 gnd vdd FILL
X_9067_ _9067_/Q _7147_/CLK _7133_/R vdd _9015_/Y gnd vdd DFFSR
XSFILL53640x7050 gnd vdd FILL
XFILL_2_BUFX2_insert1042 gnd vdd FILL
XFILL_3_BUFX2_insert338 gnd vdd FILL
XFILL_4__9030_ gnd vdd FILL
XFILL_2_BUFX2_insert1053 gnd vdd FILL
XFILL_3__7449_ gnd vdd FILL
XFILL_3_BUFX2_insert349 gnd vdd FILL
XFILL_2_BUFX2_insert1064 gnd vdd FILL
XFILL_1__9252_ gnd vdd FILL
XFILL112040x27050 gnd vdd FILL
X_8018_ _8018_/A _8006_/B _8017_/Y gnd _8052_/D vdd OAI21X1
XFILL_2_BUFX2_insert1086 gnd vdd FILL
XFILL_1__8203_ gnd vdd FILL
XSFILL23320x62050 gnd vdd FILL
XFILL_6__7089_ gnd vdd FILL
XSFILL38920x41050 gnd vdd FILL
XFILL_3__9119_ gnd vdd FILL
XSFILL64200x74050 gnd vdd FILL
X_10920_ _10906_/Y _10920_/B gnd _10920_/Y vdd NOR2X1
XFILL_1__8134_ gnd vdd FILL
X_9969_ _9969_/Q _8433_/CLK _7921_/R vdd _9969_/D gnd vdd DFFSR
XFILL_4__9932_ gnd vdd FILL
XSFILL39000x50050 gnd vdd FILL
X_10851_ _15583_/A _7530_/CLK _7523_/R vdd _10851_/D gnd vdd DFFSR
XFILL_1__8065_ gnd vdd FILL
XSFILL3640x81050 gnd vdd FILL
XSFILL14280x78050 gnd vdd FILL
XSFILL68840x77050 gnd vdd FILL
XFILL_0_BUFX2_insert1090 gnd vdd FILL
XFILL_4_CLKBUF1_insert117 gnd vdd FILL
XFILL_4__9863_ gnd vdd FILL
XFILL_4_CLKBUF1_insert128 gnd vdd FILL
X_13570_ _9816_/Q _13751_/B _14283_/C _9852_/A gnd _13570_/Y vdd AOI22X1
XSFILL29080x38050 gnd vdd FILL
XSFILL109480x6050 gnd vdd FILL
X_10782_ _10773_/A _9246_/B gnd _10782_/Y vdd NAND2X1
XFILL_4_CLKBUF1_insert139 gnd vdd FILL
X_12521_ vdd _12521_/B gnd _12521_/Y vdd NAND2X1
XFILL_6_BUFX2_insert960 gnd vdd FILL
XFILL_4__9794_ gnd vdd FILL
XFILL_6_BUFX2_insert971 gnd vdd FILL
XFILL_0_BUFX2_insert228 gnd vdd FILL
XFILL_0_BUFX2_insert239 gnd vdd FILL
XFILL_4__8745_ gnd vdd FILL
X_15240_ _15239_/Y _15236_/Y gnd _15240_/Y vdd NOR2X1
X_12452_ vdd _12005_/A gnd _12453_/C vdd NAND2X1
XFILL_1__8967_ gnd vdd FILL
XFILL_2__7760_ gnd vdd FILL
XSFILL18840x50 gnd vdd FILL
X_11403_ _11403_/A _11402_/Y gnd _11569_/B vdd NAND2X1
X_15171_ _15169_/Y _15170_/Y gnd _15171_/Y vdd NOR2X1
X_12383_ _12371_/A _12676_/Q gnd _12384_/C vdd NAND2X1
XFILL_2__7691_ gnd vdd FILL
XFILL_4__7627_ gnd vdd FILL
XFILL_1__8898_ gnd vdd FILL
X_14122_ _14122_/A _14122_/B _14791_/C gnd _12991_/B vdd AOI21X1
X_11334_ _11334_/A _11359_/B gnd _11337_/A vdd NOR2X1
XFILL_1__7849_ gnd vdd FILL
XFILL_4__7558_ gnd vdd FILL
X_14053_ _8090_/A gnd _14053_/Y vdd INVX1
XFILL_4__10540_ gnd vdd FILL
X_11265_ _12254_/Y gnd _11266_/A vdd INVX1
XFILL_2__9361_ gnd vdd FILL
XFILL_1__10360_ gnd vdd FILL
X_13004_ _13002_/Y vdd _13004_/C gnd _13064_/D vdd OAI21X1
X_10216_ _10216_/Q _8680_/CLK _8034_/R vdd _10158_/Y gnd vdd DFFSR
XFILL_6__12080_ gnd vdd FILL
XFILL_4__7489_ gnd vdd FILL
XFILL_5__11830_ gnd vdd FILL
XFILL_2__8312_ gnd vdd FILL
XFILL_1__9519_ gnd vdd FILL
X_11196_ _11196_/A _12326_/Y _11196_/C gnd _11197_/A vdd OAI21X1
XFILL_4__9228_ gnd vdd FILL
XFILL_2__9292_ gnd vdd FILL
XFILL_5__8021_ gnd vdd FILL
XFILL_2__11650_ gnd vdd FILL
XFILL_6__11031_ gnd vdd FILL
XFILL_1__10291_ gnd vdd FILL
XFILL_3_BUFX2_insert850 gnd vdd FILL
XFILL_4__12210_ gnd vdd FILL
X_10147_ _10213_/Q gnd _10147_/Y vdd INVX1
XFILL_3_BUFX2_insert861 gnd vdd FILL
XSFILL28920x73050 gnd vdd FILL
XFILL_3_BUFX2_insert872 gnd vdd FILL
XFILL_1__12030_ gnd vdd FILL
XFILL_2__8243_ gnd vdd FILL
XFILL_5__11761_ gnd vdd FILL
XFILL_0__12760_ gnd vdd FILL
XFILL_3_BUFX2_insert883 gnd vdd FILL
XFILL_2__11581_ gnd vdd FILL
XFILL_4__9159_ gnd vdd FILL
XFILL_3_BUFX2_insert894 gnd vdd FILL
XFILL_5__13500_ gnd vdd FILL
XFILL_4__12141_ gnd vdd FILL
X_14955_ _8659_/A _13864_/B _14954_/Y gnd _14964_/A vdd AOI21X1
XFILL_2__13320_ gnd vdd FILL
X_10078_ _9998_/A _7269_/CLK _9061_/R vdd _10000_/Y gnd vdd DFFSR
XFILL_5__14480_ gnd vdd FILL
XFILL_5__11692_ gnd vdd FILL
XFILL_2__10532_ gnd vdd FILL
XFILL_3__12871_ gnd vdd FILL
XFILL_0__11711_ gnd vdd FILL
XFILL_3__14610_ gnd vdd FILL
XFILL_5__13431_ gnd vdd FILL
X_13906_ _13906_/A _13906_/B gnd _13907_/C vdd NOR2X1
XFILL_5__10643_ gnd vdd FILL
XFILL_4__12072_ gnd vdd FILL
XFILL_2__7125_ gnd vdd FILL
XFILL_3__11822_ gnd vdd FILL
X_14886_ _9936_/A gnd _14886_/Y vdd INVX1
XFILL_2__13251_ gnd vdd FILL
XFILL_3__15590_ gnd vdd FILL
XFILL_0__11642_ gnd vdd FILL
XFILL_0__14430_ gnd vdd FILL
XFILL_1__13981_ gnd vdd FILL
XSFILL48840x24050 gnd vdd FILL
XFILL_4__15900_ gnd vdd FILL
X_13837_ _13837_/A _13833_/Y gnd _13837_/Y vdd NOR2X1
XSFILL99480x59050 gnd vdd FILL
XFILL_4__11023_ gnd vdd FILL
XFILL_5__16150_ gnd vdd FILL
XFILL_5__10574_ gnd vdd FILL
XFILL_5__13362_ gnd vdd FILL
XSFILL74120x57050 gnd vdd FILL
XFILL_3__14541_ gnd vdd FILL
XFILL_2__12202_ gnd vdd FILL
XFILL_2__7056_ gnd vdd FILL
XFILL_1__15720_ gnd vdd FILL
XFILL_3__11753_ gnd vdd FILL
XFILL_2__10394_ gnd vdd FILL
XFILL_0__14361_ gnd vdd FILL
XFILL_0__11573_ gnd vdd FILL
XFILL_5__15101_ gnd vdd FILL
XFILL_5__12313_ gnd vdd FILL
XFILL_5__8854_ gnd vdd FILL
XFILL_5__13293_ gnd vdd FILL
X_13768_ _14045_/A _13767_/Y _14174_/C _13768_/D gnd _13769_/B vdd OAI22X1
XFILL_4__15831_ gnd vdd FILL
XFILL_5__16081_ gnd vdd FILL
XFILL_3__10704_ gnd vdd FILL
XFILL_0__13312_ gnd vdd FILL
XFILL_3__14472_ gnd vdd FILL
XFILL_2__12133_ gnd vdd FILL
XFILL_0__16100_ gnd vdd FILL
XFILL_1__15651_ gnd vdd FILL
XFILL_0__10524_ gnd vdd FILL
XFILL_3__11684_ gnd vdd FILL
XFILL_5__7805_ gnd vdd FILL
XFILL_1__12863_ gnd vdd FILL
XFILL_0__14292_ gnd vdd FILL
X_12719_ _12719_/A gnd _12721_/A vdd INVX1
XFILL_3__16211_ gnd vdd FILL
X_15507_ _9751_/A _15390_/B _15507_/C gnd _15510_/C vdd AOI21X1
XFILL_5__15032_ gnd vdd FILL
XFILL_5__8785_ gnd vdd FILL
XSFILL53960x15050 gnd vdd FILL
XFILL_3__13423_ gnd vdd FILL
XFILL_5__12244_ gnd vdd FILL
XFILL_3__10635_ gnd vdd FILL
XFILL_1__14602_ gnd vdd FILL
XFILL_4__15762_ gnd vdd FILL
X_13699_ _13699_/A gnd _15283_/D vdd INVX1
XFILL_0__13243_ gnd vdd FILL
XFILL_0__16031_ gnd vdd FILL
XFILL_4__12974_ gnd vdd FILL
XFILL_2__12064_ gnd vdd FILL
XFILL_1__11814_ gnd vdd FILL
XFILL_5__7736_ gnd vdd FILL
XFILL_1__15582_ gnd vdd FILL
XFILL_0_BUFX2_insert740 gnd vdd FILL
X_15438_ _13924_/A _16151_/B _16247_/C _13919_/Y gnd _15439_/C vdd OAI22X1
XFILL_0_BUFX2_insert751 gnd vdd FILL
XFILL_5__12175_ gnd vdd FILL
XFILL_4__14713_ gnd vdd FILL
XFILL_3__16142_ gnd vdd FILL
XFILL_3__13354_ gnd vdd FILL
XFILL_4__11925_ gnd vdd FILL
XFILL_0_BUFX2_insert762 gnd vdd FILL
XFILL_2__11015_ gnd vdd FILL
XFILL112280x83050 gnd vdd FILL
XFILL_0_BUFX2_insert773 gnd vdd FILL
XFILL_1__14533_ gnd vdd FILL
XFILL_4__15693_ gnd vdd FILL
XFILL_3__10566_ gnd vdd FILL
XFILL_2__7958_ gnd vdd FILL
XSFILL54040x24050 gnd vdd FILL
XFILL_0__13174_ gnd vdd FILL
XFILL_1__11745_ gnd vdd FILL
X_7320_ _7336_/B _9624_/B gnd _7320_/Y vdd NAND2X1
XFILL_0__10386_ gnd vdd FILL
XFILL_5__11126_ gnd vdd FILL
XFILL_0_BUFX2_insert784 gnd vdd FILL
X_15369_ _15369_/A _13833_/B _13835_/Y _15369_/D gnd _15369_/Y vdd OAI22X1
XFILL_0__9761_ gnd vdd FILL
XFILL_0_BUFX2_insert795 gnd vdd FILL
XFILL_3__12305_ gnd vdd FILL
XFILL_0__6973_ gnd vdd FILL
XFILL_6__10677_ gnd vdd FILL
XFILL_4__14644_ gnd vdd FILL
XFILL_2__15823_ gnd vdd FILL
XFILL_2__6909_ gnd vdd FILL
XFILL_3__16073_ gnd vdd FILL
XFILL_3__13285_ gnd vdd FILL
XFILL_0__12125_ gnd vdd FILL
XFILL_3__9470_ gnd vdd FILL
XFILL_4__11856_ gnd vdd FILL
XFILL_3__10497_ gnd vdd FILL
XFILL_1__14464_ gnd vdd FILL
XFILL_6__15204_ gnd vdd FILL
XFILL_5__9406_ gnd vdd FILL
XFILL_2__7889_ gnd vdd FILL
XFILL_0__8712_ gnd vdd FILL
XFILL_1__11676_ gnd vdd FILL
XFILL_5__15934_ gnd vdd FILL
XFILL_3__15024_ gnd vdd FILL
XFILL_5__7598_ gnd vdd FILL
XFILL_5__11057_ gnd vdd FILL
X_7251_ _7251_/A gnd _7253_/A vdd INVX1
XFILL_4__10807_ gnd vdd FILL
XFILL_1__16203_ gnd vdd FILL
XFILL_2__9628_ gnd vdd FILL
XFILL_3__12236_ gnd vdd FILL
XFILL_4__14575_ gnd vdd FILL
XFILL_1__13415_ gnd vdd FILL
XFILL_4__11787_ gnd vdd FILL
XFILL_2__15754_ gnd vdd FILL
XFILL_1__10627_ gnd vdd FILL
XFILL_0__12056_ gnd vdd FILL
XFILL_2__12966_ gnd vdd FILL
XFILL_5__10008_ gnd vdd FILL
XFILL_1__14395_ gnd vdd FILL
XFILL_5__9337_ gnd vdd FILL
XFILL_4__16314_ gnd vdd FILL
XFILL_0__8643_ gnd vdd FILL
X_7182_ _7262_/Q gnd _7182_/Y vdd INVX1
XFILL_2__14705_ gnd vdd FILL
XFILL_4__13526_ gnd vdd FILL
XFILL_5__15865_ gnd vdd FILL
XFILL_3__8352_ gnd vdd FILL
XSFILL18680x43050 gnd vdd FILL
XFILL_2__11917_ gnd vdd FILL
XFILL_3__12167_ gnd vdd FILL
XFILL_0__11007_ gnd vdd FILL
XFILL_1__16134_ gnd vdd FILL
XFILL_1__13346_ gnd vdd FILL
XFILL_2__15685_ gnd vdd FILL
XFILL_1__10558_ gnd vdd FILL
XFILL_2__12897_ gnd vdd FILL
XSFILL74200x37050 gnd vdd FILL
XFILL_5__9268_ gnd vdd FILL
XFILL_6__8061_ gnd vdd FILL
XFILL_6__15066_ gnd vdd FILL
XFILL_5__14816_ gnd vdd FILL
XFILL_3__11118_ gnd vdd FILL
XFILL_0__8574_ gnd vdd FILL
XFILL_4__16245_ gnd vdd FILL
XFILL_3__7303_ gnd vdd FILL
XSFILL84360x81050 gnd vdd FILL
XFILL_2__14636_ gnd vdd FILL
XFILL_4__13457_ gnd vdd FILL
XFILL_5__15796_ gnd vdd FILL
XFILL_4__10669_ gnd vdd FILL
XFILL_5__8219_ gnd vdd FILL
XFILL_3__12098_ gnd vdd FILL
XFILL_0__15815_ gnd vdd FILL
XFILL_1__16065_ gnd vdd FILL
XFILL_2__11848_ gnd vdd FILL
XFILL_1__13277_ gnd vdd FILL
XFILL_6__14017_ gnd vdd FILL
XFILL_1__10489_ gnd vdd FILL
XSFILL49000x13050 gnd vdd FILL
XFILL_4__12408_ gnd vdd FILL
XFILL_5__14747_ gnd vdd FILL
XFILL_3__15926_ gnd vdd FILL
XFILL_5__11959_ gnd vdd FILL
XFILL_4__16176_ gnd vdd FILL
XFILL_4__13388_ gnd vdd FILL
XFILL_1__15016_ gnd vdd FILL
XFILL_3__7234_ gnd vdd FILL
XFILL_3__11049_ gnd vdd FILL
XFILL_2__14567_ gnd vdd FILL
XFILL_1__12228_ gnd vdd FILL
XFILL_1_BUFX2_insert7 gnd vdd FILL
XFILL_0__15746_ gnd vdd FILL
XFILL112440x7050 gnd vdd FILL
XFILL_2__11779_ gnd vdd FILL
XFILL_0__12958_ gnd vdd FILL
XFILL_0__7456_ gnd vdd FILL
XFILL_4__12339_ gnd vdd FILL
XFILL_2__16306_ gnd vdd FILL
XFILL_4__15127_ gnd vdd FILL
XFILL_5__14678_ gnd vdd FILL
XFILL_2__13518_ gnd vdd FILL
XFILL_3__7165_ gnd vdd FILL
XFILL_3__15857_ gnd vdd FILL
XFILL_2__14498_ gnd vdd FILL
XFILL_0__11909_ gnd vdd FILL
XSFILL38840x56050 gnd vdd FILL
XFILL_1__12159_ gnd vdd FILL
XFILL_0__15677_ gnd vdd FILL
XFILL_5__13629_ gnd vdd FILL
XFILL112360x63050 gnd vdd FILL
XFILL_0__12889_ gnd vdd FILL
X_9823_ _9745_/A _9823_/CLK _9823_/R vdd _9823_/D gnd vdd DFFSR
XFILL_2__16237_ gnd vdd FILL
XFILL_3__14808_ gnd vdd FILL
XFILL_4__15058_ gnd vdd FILL
XFILL_2__13449_ gnd vdd FILL
XFILL_0__14628_ gnd vdd FILL
XFILL_3__7096_ gnd vdd FILL
XFILL_3__15788_ gnd vdd FILL
XFILL_0__9126_ gnd vdd FILL
XSFILL74120x9050 gnd vdd FILL
XFILL_4__14009_ gnd vdd FILL
XFILL_5__16348_ gnd vdd FILL
XFILL_6__15899_ gnd vdd FILL
X_9754_ _9826_/Q gnd _9756_/A vdd INVX1
X_6966_ _6967_/B _7094_/B gnd _6966_/Y vdd NAND2X1
XFILL_1__15918_ gnd vdd FILL
XFILL_2__16168_ gnd vdd FILL
XFILL_3__14739_ gnd vdd FILL
XFILL_0__14559_ gnd vdd FILL
X_8705_ _8703_/Y _8740_/A _8705_/C gnd _8705_/Y vdd OAI21X1
XSFILL114120x58050 gnd vdd FILL
XFILL_6_BUFX2_insert234 gnd vdd FILL
XFILL_2__15119_ gnd vdd FILL
XFILL_5__16279_ gnd vdd FILL
X_9685_ _9685_/A _9675_/A _9685_/C gnd _9717_/D vdd OAI21X1
XFILL_4__6860_ gnd vdd FILL
XFILL_2__16099_ gnd vdd FILL
XFILL_1__15849_ gnd vdd FILL
X_6897_ _6897_/A gnd memoryWriteData[27] vdd BUFX2
XFILL_0__8008_ gnd vdd FILL
XSFILL18760x23050 gnd vdd FILL
X_8636_ _8655_/B _8636_/B gnd _8636_/Y vdd NAND2X1
XFILL_1__9870_ gnd vdd FILL
XFILL_3__16409_ gnd vdd FILL
XSFILL8600x33050 gnd vdd FILL
XFILL_3__9806_ gnd vdd FILL
XFILL_0__16229_ gnd vdd FILL
XSFILL44040x56050 gnd vdd FILL
XFILL_5_BUFX2_insert901 gnd vdd FILL
XFILL_3__7998_ gnd vdd FILL
XSFILL59640x35050 gnd vdd FILL
XFILL_5_BUFX2_insert912 gnd vdd FILL
XSFILL84440x61050 gnd vdd FILL
XFILL_5_BUFX2_insert923 gnd vdd FILL
XFILL_5_BUFX2_insert934 gnd vdd FILL
X_8567_ _8567_/A _8567_/B gnd _8568_/C vdd NAND2X1
XFILL_4__8530_ gnd vdd FILL
XFILL_3__6949_ gnd vdd FILL
XFILL_3__9737_ gnd vdd FILL
XFILL_5_BUFX2_insert945 gnd vdd FILL
XFILL_5_BUFX2_insert956 gnd vdd FILL
XFILL_5_BUFX2_insert967 gnd vdd FILL
X_7518_ _7518_/Q _9817_/CLK _8542_/R vdd _7440_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert978 gnd vdd FILL
XFILL_1__8752_ gnd vdd FILL
XFILL_5_BUFX2_insert989 gnd vdd FILL
XFILL_4__8461_ gnd vdd FILL
XFILL_3__9668_ gnd vdd FILL
X_8498_ _8498_/A gnd _8500_/A vdd INVX1
XFILL_1__7703_ gnd vdd FILL
X_7449_ _7449_/A _7457_/A _7448_/Y gnd _7521_/D vdd OAI21X1
XSFILL38920x36050 gnd vdd FILL
XSFILL38120x17050 gnd vdd FILL
XFILL_3__8619_ gnd vdd FILL
XFILL_3__9599_ gnd vdd FILL
XFILL112440x43050 gnd vdd FILL
XFILL_4__8392_ gnd vdd FILL
XSFILL64200x69050 gnd vdd FILL
XFILL_1__7634_ gnd vdd FILL
XFILL_4__7343_ gnd vdd FILL
XSFILL89160x73050 gnd vdd FILL
XFILL_3_BUFX2_insert102 gnd vdd FILL
X_11050_ _12250_/Y _12141_/Y gnd _11050_/Y vdd XOR2X1
X_9119_ _9117_/Y _9170_/B _9119_/C gnd _9119_/Y vdd OAI21X1
XFILL_1__7565_ gnd vdd FILL
X_10001_ _13900_/A gnd _10001_/Y vdd INVX1
XSFILL3640x76050 gnd vdd FILL
XFILL_4__9013_ gnd vdd FILL
XSFILL3720x4050 gnd vdd FILL
XFILL_1__7496_ gnd vdd FILL
XCLKBUF1_insert1080 clk gnd CLKBUF1_insert150/A vdd CLKBUF1
XFILL_2_BUFX2_insert802 gnd vdd FILL
XSFILL94280x64050 gnd vdd FILL
XFILL_1__9235_ gnd vdd FILL
XFILL_2_BUFX2_insert813 gnd vdd FILL
XFILL_2_BUFX2_insert824 gnd vdd FILL
XFILL_2_BUFX2_insert835 gnd vdd FILL
X_14740_ _14738_/Y _14740_/B _14740_/C gnd _14740_/Y vdd NAND3X1
XFILL_2_BUFX2_insert846 gnd vdd FILL
X_11952_ _11952_/A _11909_/A _11952_/C gnd _6859_/A vdd OAI21X1
XSFILL69080x40050 gnd vdd FILL
XFILL_2_BUFX2_insert857 gnd vdd FILL
XFILL_1__9166_ gnd vdd FILL
XFILL_2_BUFX2_insert868 gnd vdd FILL
XFILL_2_BUFX2_insert879 gnd vdd FILL
X_10903_ _10903_/A _10903_/B gnd _10920_/B vdd NAND2X1
XSFILL33960x79050 gnd vdd FILL
XFILL_1__8117_ gnd vdd FILL
XFILL_0_BUFX2_insert90 gnd vdd FILL
X_14671_ _16048_/A _14721_/A gnd _14672_/C vdd NOR2X1
X_11883_ _11883_/A _11874_/B _11882_/Y gnd _13246_/A vdd OAI21X1
XFILL_1__9097_ gnd vdd FILL
XFILL_4__9915_ gnd vdd FILL
X_16410_ _16410_/A gnd _16410_/C gnd _16410_/Y vdd OAI21X1
X_13622_ _13622_/A _13621_/Y _13622_/C gnd _13636_/A vdd NAND3X1
X_10834_ _10834_/A _10822_/B _10833_/Y gnd _10868_/D vdd OAI21X1
X_16341_ _16341_/A gnd _16341_/C gnd _16423_/D vdd OAI21X1
XFILL_4__9846_ gnd vdd FILL
XBUFX2_insert801 _15091_/Y gnd _15178_/C vdd BUFX2
X_13553_ _9980_/A gnd _13554_/D vdd INVX1
XBUFX2_insert812 _13329_/Y gnd _9044_/A vdd BUFX2
X_10765_ _10763_/Y _10831_/B _10765_/C gnd _10845_/D vdd OAI21X1
XFILL_5__10290_ gnd vdd FILL
XBUFX2_insert823 _13287_/Y gnd _7416_/B vdd BUFX2
XSFILL18760x4050 gnd vdd FILL
XFILL_2__8861_ gnd vdd FILL
XBUFX2_insert834 _15046_/Y gnd _15351_/A vdd BUFX2
X_12504_ _12504_/A vdd _12503_/Y gnd _12504_/Y vdd OAI21X1
XBUFX2_insert845 _12375_/Y gnd _7317_/B vdd BUFX2
XFILL_5__8570_ gnd vdd FILL
XBUFX2_insert856 _13314_/Y gnd _8208_/B vdd BUFX2
XFILL_4__6989_ gnd vdd FILL
XFILL_4__9777_ gnd vdd FILL
X_16272_ _16272_/A _15958_/B _15010_/A _16272_/D gnd _16272_/Y vdd OAI22X1
XFILL_2__7812_ gnd vdd FILL
X_13484_ _13630_/B gnd _13484_/Y vdd INVX8
XFILL_3__10420_ gnd vdd FILL
XBUFX2_insert867 _13438_/Y gnd _14413_/A vdd BUFX2
X_10696_ _10681_/A _8008_/B gnd _10696_/Y vdd NAND2X1
XFILL_0__10240_ gnd vdd FILL
XSFILL3720x56050 gnd vdd FILL
XBUFX2_insert878 _15019_/Y gnd _15633_/D vdd BUFX2
XFILL_1__9999_ gnd vdd FILL
XFILL_4__8728_ gnd vdd FILL
X_15223_ _7002_/Q _15382_/B _16096_/C _7298_/A gnd _15223_/Y vdd AOI22X1
XBUFX2_insert889 _13432_/Y gnd _14636_/C vdd BUFX2
X_12435_ _12433_/Y _12395_/A _12435_/C gnd _12435_/Y vdd OAI21X1
XFILL_4__11710_ gnd vdd FILL
XFILL_2__7743_ gnd vdd FILL
XFILL_1__11530_ gnd vdd FILL
XFILL_0__10171_ gnd vdd FILL
XFILL_5__7452_ gnd vdd FILL
XSFILL94360x44050 gnd vdd FILL
X_15154_ _15153_/Y _16151_/B _16309_/A _13554_/D gnd _15154_/Y vdd OAI22X1
XFILL_4__8659_ gnd vdd FILL
X_12366_ _12364_/Y _12407_/A _12366_/C gnd _12366_/Y vdd OAI21X1
XFILL_4__11641_ gnd vdd FILL
XFILL_5__13980_ gnd vdd FILL
XFILL_3__10282_ gnd vdd FILL
XFILL_2__7674_ gnd vdd FILL
XFILL_1__11461_ gnd vdd FILL
X_14105_ _14105_/A _14105_/B gnd _14106_/A vdd NOR2X1
X_11317_ _11303_/B _11533_/A _11317_/C gnd _11318_/C vdd OAI21X1
XFILL_3__12021_ gnd vdd FILL
XFILL_2__9413_ gnd vdd FILL
XFILL_4__14360_ gnd vdd FILL
X_15085_ _15085_/A _15084_/Y _15085_/C gnd _15103_/C vdd NAND3X1
XFILL_6__10393_ gnd vdd FILL
XFILL_4__11572_ gnd vdd FILL
X_12297_ _6890_/A _12289_/B _12289_/C _12297_/D gnd _12297_/Y vdd AOI22X1
XFILL_2__12751_ gnd vdd FILL
XFILL_5__9122_ gnd vdd FILL
XFILL_1__10412_ gnd vdd FILL
XFILL_1__14180_ gnd vdd FILL
XFILL_1__11392_ gnd vdd FILL
XFILL_0__13930_ gnd vdd FILL
X_14036_ _14032_/Y _14035_/Y _14036_/C gnd _14048_/B vdd NAND3X1
XFILL_4__13311_ gnd vdd FILL
XFILL_5__15650_ gnd vdd FILL
XFILL_4__10523_ gnd vdd FILL
X_11248_ _12238_/Y _11030_/A gnd _11787_/C vdd XOR2X1
XFILL_2__9344_ gnd vdd FILL
XFILL_4__14291_ gnd vdd FILL
XFILL_2__11702_ gnd vdd FILL
XFILL_5__12862_ gnd vdd FILL
XFILL_1__13131_ gnd vdd FILL
XFILL_2__15470_ gnd vdd FILL
XFILL_0__13861_ gnd vdd FILL
XFILL_5__14601_ gnd vdd FILL
XSFILL74280x11050 gnd vdd FILL
XFILL_4__13242_ gnd vdd FILL
XFILL_4__16030_ gnd vdd FILL
XFILL_5__11813_ gnd vdd FILL
XFILL_2__14421_ gnd vdd FILL
XFILL_5__15581_ gnd vdd FILL
X_11179_ _12189_/Y gnd _11179_/Y vdd INVX1
XFILL_2__9275_ gnd vdd FILL
XFILL_5__8004_ gnd vdd FILL
XFILL_2__11633_ gnd vdd FILL
XFILL_0__15600_ gnd vdd FILL
XFILL_3__13972_ gnd vdd FILL
XFILL_1__10274_ gnd vdd FILL
XFILL_0__7310_ gnd vdd FILL
XFILL_3_BUFX2_insert680 gnd vdd FILL
XFILL_0__13792_ gnd vdd FILL
XFILL_5__14532_ gnd vdd FILL
XFILL_3_BUFX2_insert691 gnd vdd FILL
XFILL_3__15711_ gnd vdd FILL
XFILL_2__8226_ gnd vdd FILL
XFILL_4__13173_ gnd vdd FILL
XFILL_5__11744_ gnd vdd FILL
X_15987_ _16026_/D _14554_/Y _15899_/C _14550_/Y gnd _15987_/Y vdd OAI22X1
XFILL_1__12013_ gnd vdd FILL
XFILL_2__14352_ gnd vdd FILL
XFILL_4__10385_ gnd vdd FILL
XFILL_0__15531_ gnd vdd FILL
XSFILL109480x39050 gnd vdd FILL
XFILL_2__11564_ gnd vdd FILL
XFILL_0__12743_ gnd vdd FILL
XFILL_4__12124_ gnd vdd FILL
XFILL_0__7241_ gnd vdd FILL
XFILL_2__13303_ gnd vdd FILL
XFILL_5__14463_ gnd vdd FILL
X_14938_ _14934_/Y _14938_/B gnd _14938_/Y vdd NOR2X1
XFILL_3__15642_ gnd vdd FILL
XFILL_3__12854_ gnd vdd FILL
XFILL_5__11675_ gnd vdd FILL
XFILL_2__10515_ gnd vdd FILL
XFILL112280x78050 gnd vdd FILL
XFILL_2__14283_ gnd vdd FILL
XFILL_5__16202_ gnd vdd FILL
XFILL_2__11495_ gnd vdd FILL
XFILL_0__15462_ gnd vdd FILL
XSFILL54040x19050 gnd vdd FILL
XFILL_5__13414_ gnd vdd FILL
XFILL_2__16022_ gnd vdd FILL
XFILL_0__7172_ gnd vdd FILL
XFILL_5__10626_ gnd vdd FILL
XFILL_6__12965_ gnd vdd FILL
XFILL_2__7108_ gnd vdd FILL
XFILL_4__12055_ gnd vdd FILL
XFILL_3__11805_ gnd vdd FILL
XFILL_2__13234_ gnd vdd FILL
X_14869_ _14867_/Y _14869_/B _14869_/C gnd _14880_/B vdd NAND3X1
XFILL_5__14394_ gnd vdd FILL
XFILL_3__12785_ gnd vdd FILL
XFILL_2__10446_ gnd vdd FILL
XFILL_3__8970_ gnd vdd FILL
XFILL_2__8088_ gnd vdd FILL
XFILL_3__15573_ gnd vdd FILL
XFILL_0__14413_ gnd vdd FILL
XFILL_5__8906_ gnd vdd FILL
XFILL_0__11625_ gnd vdd FILL
XFILL_1__13964_ gnd vdd FILL
XFILL_0__15393_ gnd vdd FILL
XFILL_4__11006_ gnd vdd FILL
XFILL_5__16133_ gnd vdd FILL
XFILL_5__13345_ gnd vdd FILL
XFILL_5__9886_ gnd vdd FILL
XFILL_2__7039_ gnd vdd FILL
XFILL_1__15703_ gnd vdd FILL
XFILL_5__10557_ gnd vdd FILL
XSFILL28600x50050 gnd vdd FILL
XFILL_3__14524_ gnd vdd FILL
XFILL_3__11736_ gnd vdd FILL
XFILL_2__13165_ gnd vdd FILL
XFILL_1__12915_ gnd vdd FILL
XFILL_2__10377_ gnd vdd FILL
XFILL_0__14344_ gnd vdd FILL
XFILL_0__11556_ gnd vdd FILL
XFILL_5__8837_ gnd vdd FILL
XFILL_1__13895_ gnd vdd FILL
XFILL_4__15814_ gnd vdd FILL
XFILL_5__16064_ gnd vdd FILL
XFILL_5__13276_ gnd vdd FILL
XFILL_3__14455_ gnd vdd FILL
XFILL_5__10488_ gnd vdd FILL
XFILL_2__12116_ gnd vdd FILL
X_9470_ _9470_/A _9514_/A _9469_/Y gnd _9560_/D vdd OAI21X1
XFILL_0__10507_ gnd vdd FILL
XFILL_1__15634_ gnd vdd FILL
XFILL_3__7852_ gnd vdd FILL
XFILL_3__11667_ gnd vdd FILL
XFILL_1__12846_ gnd vdd FILL
XFILL_2__13096_ gnd vdd FILL
XSFILL18680x38050 gnd vdd FILL
XSFILL73720x25050 gnd vdd FILL
XFILL_5__15015_ gnd vdd FILL
XFILL_0__11487_ gnd vdd FILL
XFILL_0__14275_ gnd vdd FILL
XFILL_5__8768_ gnd vdd FILL
X_8421_ _8421_/Q _8046_/CLK _9692_/R vdd _8421_/D gnd vdd DFFSR
XFILL_3__13406_ gnd vdd FILL
XFILL_5__12227_ gnd vdd FILL
XFILL_3__10618_ gnd vdd FILL
XFILL_6__11778_ gnd vdd FILL
XFILL_4__15745_ gnd vdd FILL
XFILL_0__16014_ gnd vdd FILL
XFILL_2__12047_ gnd vdd FILL
XFILL_3__14386_ gnd vdd FILL
XFILL_4__12957_ gnd vdd FILL
XSFILL84360x76050 gnd vdd FILL
XFILL_0__13226_ gnd vdd FILL
XFILL_0__10438_ gnd vdd FILL
XFILL_1__15565_ gnd vdd FILL
XFILL_3__11598_ gnd vdd FILL
XFILL_1__12777_ gnd vdd FILL
XFILL_5__7719_ gnd vdd FILL
XFILL_0_BUFX2_insert570 gnd vdd FILL
XFILL_0__9813_ gnd vdd FILL
XFILL_0_BUFX2_insert581 gnd vdd FILL
XFILL_6__7492_ gnd vdd FILL
XFILL_3__13337_ gnd vdd FILL
XFILL_0_BUFX2_insert592 gnd vdd FILL
XFILL_4__11908_ gnd vdd FILL
X_8352_ _8420_/Q gnd _8354_/A vdd INVX1
XFILL_5__12158_ gnd vdd FILL
XFILL_3__16125_ gnd vdd FILL
XFILL_3__9522_ gnd vdd FILL
XFILL_5__8699_ gnd vdd FILL
XFILL_3__10549_ gnd vdd FILL
XFILL_4__15676_ gnd vdd FILL
XFILL_1__14516_ gnd vdd FILL
XFILL_4__12888_ gnd vdd FILL
XSFILL59160x52050 gnd vdd FILL
XFILL_0__13157_ gnd vdd FILL
XFILL_1__11728_ gnd vdd FILL
XSFILL89400x13050 gnd vdd FILL
XFILL_0__10369_ gnd vdd FILL
XFILL_4_BUFX2_insert908 gnd vdd FILL
XFILL_1__15496_ gnd vdd FILL
XFILL_0__9744_ gnd vdd FILL
XFILL_4_BUFX2_insert919 gnd vdd FILL
XFILL_5__11109_ gnd vdd FILL
X_7303_ _7303_/A _7369_/B _7302_/Y gnd _7387_/D vdd OAI21X1
XFILL_4__14627_ gnd vdd FILL
XFILL_5__12089_ gnd vdd FILL
XFILL_0__6956_ gnd vdd FILL
XFILL_3__16056_ gnd vdd FILL
XSFILL109560x19050 gnd vdd FILL
X_8283_ _8283_/Q _8551_/CLK _7015_/R vdd _8199_/Y gnd vdd DFFSR
XFILL_3__13268_ gnd vdd FILL
XFILL_0__12108_ gnd vdd FILL
XFILL_2__15806_ gnd vdd FILL
XFILL_4__11839_ gnd vdd FILL
XFILL_1__14447_ gnd vdd FILL
XFILL_0__13088_ gnd vdd FILL
XFILL_6__9162_ gnd vdd FILL
XFILL_2__13998_ gnd vdd FILL
XFILL_1__11659_ gnd vdd FILL
XFILL_5__15917_ gnd vdd FILL
XFILL111880x51050 gnd vdd FILL
XFILL_3__15007_ gnd vdd FILL
XFILL112360x58050 gnd vdd FILL
XFILL_0__9675_ gnd vdd FILL
XFILL_3__8404_ gnd vdd FILL
X_7234_ _7166_/B _7490_/B gnd _7235_/C vdd NAND2X1
XFILL_3__12219_ gnd vdd FILL
XFILL_4__14558_ gnd vdd FILL
XFILL_0__6887_ gnd vdd FILL
XFILL_3__9384_ gnd vdd FILL
XFILL_0__12039_ gnd vdd FILL
XFILL_6__8113_ gnd vdd FILL
XFILL_2__15737_ gnd vdd FILL
XFILL_1__14378_ gnd vdd FILL
XFILL_0__8626_ gnd vdd FILL
XFILL_5__15848_ gnd vdd FILL
X_7165_ _7166_/B _7293_/B gnd _7165_/Y vdd NAND2X1
XFILL_4__13509_ gnd vdd FILL
XSFILL109400x83050 gnd vdd FILL
XFILL_3__8335_ gnd vdd FILL
XFILL_1__16117_ gnd vdd FILL
XFILL_1__13329_ gnd vdd FILL
XFILL_2__15668_ gnd vdd FILL
XFILL_4__14489_ gnd vdd FILL
XSFILL79320x65050 gnd vdd FILL
XFILL_1__7350_ gnd vdd FILL
XFILL_4__16228_ gnd vdd FILL
XFILL_2__14619_ gnd vdd FILL
X_7096_ _7148_/Q gnd _7096_/Y vdd INVX1
XFILL_5__15779_ gnd vdd FILL
XFILL_3__8266_ gnd vdd FILL
XFILL_1__16048_ gnd vdd FILL
XFILL_2__15599_ gnd vdd FILL
XFILL_0__7508_ gnd vdd FILL
XFILL_2_BUFX2_insert109 gnd vdd FILL
XFILL_3__15909_ gnd vdd FILL
XFILL_0__8488_ gnd vdd FILL
XFILL_3__7217_ gnd vdd FILL
XFILL_4__16159_ gnd vdd FILL
XSFILL18760x18050 gnd vdd FILL
XSFILL8600x28050 gnd vdd FILL
XFILL_0__15729_ gnd vdd FILL
XFILL_3__8197_ gnd vdd FILL
XFILL_1__9020_ gnd vdd FILL
XFILL_0__7439_ gnd vdd FILL
XSFILL33800x21050 gnd vdd FILL
XSFILL84440x56050 gnd vdd FILL
X_9806_ _9789_/B _8014_/B gnd _9807_/C vdd NAND2X1
XFILL_1_BUFX2_insert809 gnd vdd FILL
XSFILL85080x22050 gnd vdd FILL
X_7998_ _8046_/Q gnd _7998_/Y vdd INVX1
XFILL_3__7079_ gnd vdd FILL
XFILL_4__7961_ gnd vdd FILL
XFILL_0__9109_ gnd vdd FILL
X_9737_ _9737_/A _9737_/B gnd _9738_/C vdd NAND2X1
X_6949_ _6947_/Y _6948_/A _6949_/C gnd _7013_/D vdd OAI21X1
XFILL111960x31050 gnd vdd FILL
XFILL_4__6912_ gnd vdd FILL
XFILL112440x38050 gnd vdd FILL
XFILL_4__7892_ gnd vdd FILL
XBUFX2_insert108 _10925_/Y gnd _11975_/A vdd BUFX2
XFILL_1__9922_ gnd vdd FILL
XSFILL23720x73050 gnd vdd FILL
X_9668_ _9712_/Q gnd _9668_/Y vdd INVX1
XFILL_4__6843_ gnd vdd FILL
XFILL_4__9631_ gnd vdd FILL
X_10550_ _10535_/A _9782_/B gnd _10551_/C vdd NAND2X1
XFILL_1__9853_ gnd vdd FILL
X_8619_ _8619_/A _8619_/B _8618_/Y gnd _8679_/D vdd OAI21X1
XFILL_5_BUFX2_insert720 gnd vdd FILL
X_9599_ _9689_/Q gnd _9599_/Y vdd INVX1
XFILL_5_BUFX2_insert731 gnd vdd FILL
XFILL_5_BUFX2_insert742 gnd vdd FILL
XFILL_5_BUFX2_insert753 gnd vdd FILL
X_10481_ _10481_/Q _7786_/CLK _7153_/R vdd _10481_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert764 gnd vdd FILL
XFILL_1__9784_ gnd vdd FILL
XFILL_1__6996_ gnd vdd FILL
XFILL_4__8513_ gnd vdd FILL
XFILL_5_BUFX2_insert775 gnd vdd FILL
XFILL_5_BUFX2_insert786 gnd vdd FILL
X_12220_ _12224_/A _12792_/Q _12224_/C gnd _12222_/B vdd NAND3X1
XFILL_4__9493_ gnd vdd FILL
XFILL_5_BUFX2_insert797 gnd vdd FILL
XSFILL114600x54050 gnd vdd FILL
XFILL_1__8735_ gnd vdd FILL
XFILL_4__8444_ gnd vdd FILL
XSFILL84520x36050 gnd vdd FILL
X_12151_ _12151_/A gnd _12153_/A vdd INVX1
XSFILL69080x35050 gnd vdd FILL
XFILL_4__8375_ gnd vdd FILL
X_11102_ _12186_/Y gnd _11102_/Y vdd INVX1
X_12082_ _12082_/A _12082_/B _12081_/Y gnd _13149_/B vdd NAND3X1
XFILL_1__7617_ gnd vdd FILL
XFILL_1__8597_ gnd vdd FILL
XFILL_4__7326_ gnd vdd FILL
X_15910_ _15910_/A _15910_/B gnd _15929_/B vdd NOR2X1
X_11033_ _11025_/A _11032_/Y gnd _11785_/A vdd NOR2X1
XFILL_1__7548_ gnd vdd FILL
XSFILL23800x53050 gnd vdd FILL
X_15841_ _14365_/A _15958_/B _15841_/C _15841_/D gnd _15841_/Y vdd OAI22X1
XFILL_1__7479_ gnd vdd FILL
XFILL_2_BUFX2_insert610 gnd vdd FILL
XFILL_2_BUFX2_insert621 gnd vdd FILL
XFILL112120x20050 gnd vdd FILL
XFILL_2_BUFX2_insert632 gnd vdd FILL
XFILL_4__7188_ gnd vdd FILL
XFILL_1__9218_ gnd vdd FILL
XFILL_2__8011_ gnd vdd FILL
XFILL_2_BUFX2_insert643 gnd vdd FILL
XFILL_4__10170_ gnd vdd FILL
X_12984_ _6881_/A gnd _12984_/Y vdd INVX1
X_15772_ _15916_/B _10668_/A _7656_/Q _15662_/A gnd _15772_/Y vdd AOI22X1
XFILL_2_BUFX2_insert654 gnd vdd FILL
XFILL_2_BUFX2_insert665 gnd vdd FILL
XFILL_2_BUFX2_insert676 gnd vdd FILL
X_11935_ _11935_/A gnd _11937_/A vdd INVX1
XFILL_2_BUFX2_insert687 gnd vdd FILL
X_14723_ _9712_/Q gnd _14725_/C vdd INVX1
XFILL_1__9149_ gnd vdd FILL
XFILL_2__10300_ gnd vdd FILL
XFILL_2_BUFX2_insert698 gnd vdd FILL
XFILL_5__11460_ gnd vdd FILL
XFILL_2__11280_ gnd vdd FILL
XFILL_5__9740_ gnd vdd FILL
XSFILL13480x43050 gnd vdd FILL
XSFILL94360x39050 gnd vdd FILL
XFILL_5__6952_ gnd vdd FILL
XFILL_5__10411_ gnd vdd FILL
X_14654_ _14654_/A _14653_/Y gnd _14654_/Y vdd NOR2X1
X_11866_ _12101_/A _12093_/A gnd _11866_/Y vdd NOR2X1
XFILL_5__11391_ gnd vdd FILL
XFILL_3__12570_ gnd vdd FILL
XFILL_2__10231_ gnd vdd FILL
XFILL_0__11410_ gnd vdd FILL
XFILL_5_BUFX2_insert14 gnd vdd FILL
XFILL_1__10961_ gnd vdd FILL
X_13605_ _10457_/Q _14389_/B _13605_/C gnd _13610_/A vdd AOI21X1
XFILL_0__12390_ gnd vdd FILL
XFILL_5_BUFX2_insert25 gnd vdd FILL
XSFILL69160x15050 gnd vdd FILL
XFILL_5_BUFX2_insert36 gnd vdd FILL
XFILL_5__13130_ gnd vdd FILL
XFILL_5__9671_ gnd vdd FILL
X_10817_ _16071_/A gnd _10819_/A vdd INVX1
XFILL_5__6883_ gnd vdd FILL
X_14585_ _8045_/Q gnd _15996_/B vdd INVX1
XFILL_5_BUFX2_insert47 gnd vdd FILL
XFILL_3__11521_ gnd vdd FILL
XFILL_1__12700_ gnd vdd FILL
XFILL_4__13860_ gnd vdd FILL
X_11797_ _11795_/Y _11034_/B _11751_/C gnd _11797_/Y vdd OAI21X1
XFILL_2__8913_ gnd vdd FILL
XFILL_2__9893_ gnd vdd FILL
XBUFX2_insert620 _13430_/Y gnd _13619_/B vdd BUFX2
XFILL_2__10162_ gnd vdd FILL
XFILL_5_BUFX2_insert58 gnd vdd FILL
XFILL_0__11341_ gnd vdd FILL
XFILL_1__13680_ gnd vdd FILL
XFILL_5_BUFX2_insert69 gnd vdd FILL
XFILL_5__8622_ gnd vdd FILL
XBUFX2_insert631 _13465_/Y gnd _14711_/B vdd BUFX2
X_16324_ _16324_/A gnd _16326_/A vdd INVX1
XFILL_1__10892_ gnd vdd FILL
X_13536_ _13534_/Y _14865_/B _14320_/C _13536_/D gnd _13540_/B vdd OAI22X1
XFILL_3__14240_ gnd vdd FILL
XFILL_5__10273_ gnd vdd FILL
XBUFX2_insert642 _13424_/Y gnd _14934_/B vdd BUFX2
X_10748_ _13568_/C gnd _10750_/A vdd INVX1
XBUFX2_insert653 _12429_/Y gnd _9803_/B vdd BUFX2
XFILL_3__11452_ gnd vdd FILL
XSFILL104360x24050 gnd vdd FILL
XFILL_1__12631_ gnd vdd FILL
XFILL_4__13791_ gnd vdd FILL
XFILL_2__8844_ gnd vdd FILL
XFILL_0__14060_ gnd vdd FILL
XFILL_2__14970_ gnd vdd FILL
XBUFX2_insert664 _11364_/Y gnd _11848_/A vdd BUFX2
XBUFX2_insert675 _13541_/Y gnd _13771_/D vdd BUFX2
XFILL_0__11272_ gnd vdd FILL
XSFILL104520x7050 gnd vdd FILL
XFILL_5__12012_ gnd vdd FILL
XBUFX2_insert686 _13459_/Y gnd _14949_/C vdd BUFX2
X_16255_ _8820_/Q gnd _16255_/Y vdd INVX1
XFILL_3__10403_ gnd vdd FILL
X_13467_ _13467_/A _14987_/B _14640_/C _13464_/Y gnd _13467_/Y vdd OAI22X1
XFILL_4__15530_ gnd vdd FILL
X_10679_ _10677_/Y _10678_/A _10679_/C gnd _10731_/D vdd OAI21X1
XFILL_4__12742_ gnd vdd FILL
XFILL_3__14171_ gnd vdd FILL
XBUFX2_insert697 _12420_/Y gnd _8642_/B vdd BUFX2
XFILL_2__13921_ gnd vdd FILL
XFILL_0__13011_ gnd vdd FILL
XFILL_1__15350_ gnd vdd FILL
XFILL_2__8775_ gnd vdd FILL
XFILL_3__11383_ gnd vdd FILL
X_15206_ _15201_/Y _15206_/B gnd _15206_/Y vdd NAND2X1
XSFILL8040x65050 gnd vdd FILL
XFILL_5__7504_ gnd vdd FILL
XFILL_5__8484_ gnd vdd FILL
X_12418_ _12418_/A gnd _12418_/Y vdd INVX1
X_16186_ _14796_/D _15203_/B _16186_/C gnd _16186_/Y vdd OAI21X1
XFILL_3__13122_ gnd vdd FILL
XSFILL59080x67050 gnd vdd FILL
X_13398_ _13398_/A _13377_/Y gnd _14865_/B vdd NAND2X1
XFILL_2__7726_ gnd vdd FILL
XFILL_1__14301_ gnd vdd FILL
XFILL_4__15461_ gnd vdd FILL
XFILL_2__13852_ gnd vdd FILL
XFILL_1__11513_ gnd vdd FILL
XFILL_5__7435_ gnd vdd FILL
XFILL_0__10154_ gnd vdd FILL
XFILL_1__15281_ gnd vdd FILL
XFILL_1__12493_ gnd vdd FILL
X_15137_ _7256_/Q _15177_/B gnd _15143_/A vdd NAND2X1
X_12349_ _12349_/A gnd _12349_/Y vdd INVX1
XFILL_4__14412_ gnd vdd FILL
XFILL_4__11624_ gnd vdd FILL
XFILL_5__13963_ gnd vdd FILL
XFILL_1__14232_ gnd vdd FILL
XFILL_4__15392_ gnd vdd FILL
XFILL_3__10265_ gnd vdd FILL
XFILL_2__13783_ gnd vdd FILL
XFILL_1__11444_ gnd vdd FILL
XFILL_5__15702_ gnd vdd FILL
XFILL_0__14962_ gnd vdd FILL
XFILL_5__7366_ gnd vdd FILL
XFILL_2__10995_ gnd vdd FILL
X_15068_ _16232_/B _16035_/B gnd _15068_/Y vdd NAND2X1
XFILL_3__12004_ gnd vdd FILL
XFILL_5__12914_ gnd vdd FILL
XFILL_2__15522_ gnd vdd FILL
XFILL_4__14343_ gnd vdd FILL
XFILL_4__11555_ gnd vdd FILL
XFILL_2__12734_ gnd vdd FILL
XFILL_5__13894_ gnd vdd FILL
XSFILL94440x19050 gnd vdd FILL
XFILL_2__7588_ gnd vdd FILL
XFILL_1__14163_ gnd vdd FILL
XFILL_3__10196_ gnd vdd FILL
XFILL_5__9105_ gnd vdd FILL
XFILL_0__13913_ gnd vdd FILL
X_14019_ _14019_/A _14018_/Y gnd _14022_/C vdd NOR2X1
XFILL_1__11375_ gnd vdd FILL
XFILL_5__7297_ gnd vdd FILL
XFILL_4__10506_ gnd vdd FILL
XFILL_5__15633_ gnd vdd FILL
XFILL_0__14893_ gnd vdd FILL
XFILL_5__12845_ gnd vdd FILL
XFILL_3__8120_ gnd vdd FILL
XFILL_6__13095_ gnd vdd FILL
XFILL_0__9391_ gnd vdd FILL
XFILL_1__13114_ gnd vdd FILL
XFILL_4__11486_ gnd vdd FILL
XFILL_2__15453_ gnd vdd FILL
XFILL_4__14274_ gnd vdd FILL
XFILL_5__9036_ gnd vdd FILL
XFILL_0__13844_ gnd vdd FILL
XSFILL94280x5050 gnd vdd FILL
XFILL_1__14094_ gnd vdd FILL
XFILL_4__16013_ gnd vdd FILL
XFILL_0__8342_ gnd vdd FILL
XFILL_4__13225_ gnd vdd FILL
XFILL_4__10437_ gnd vdd FILL
XFILL_5__15564_ gnd vdd FILL
XFILL_2__14404_ gnd vdd FILL
XFILL_5__12776_ gnd vdd FILL
X_8970_ _8968_/Y _8969_/A _8969_/Y gnd _9052_/D vdd OAI21X1
XFILL_2__9258_ gnd vdd FILL
XFILL_2__11616_ gnd vdd FILL
XFILL_2__15384_ gnd vdd FILL
XFILL_1__13045_ gnd vdd FILL
XFILL_1__10257_ gnd vdd FILL
XFILL_3__13955_ gnd vdd FILL
XFILL_2__12596_ gnd vdd FILL
XFILL_0__13775_ gnd vdd FILL
XFILL_5__14515_ gnd vdd FILL
XFILL_4__13156_ gnd vdd FILL
XFILL_5__11727_ gnd vdd FILL
XFILL_2__8209_ gnd vdd FILL
X_7921_ _7921_/Q _8433_/CLK _7921_/R vdd _7881_/Y gnd vdd DFFSR
XFILL_0__8273_ gnd vdd FILL
XFILL_4__10368_ gnd vdd FILL
XFILL_2__14335_ gnd vdd FILL
XFILL_3__12906_ gnd vdd FILL
XFILL_5__15495_ gnd vdd FILL
XFILL_0__15514_ gnd vdd FILL
XFILL_2__11547_ gnd vdd FILL
XFILL_0__12726_ gnd vdd FILL
XFILL_3__13886_ gnd vdd FILL
XFILL_1__10188_ gnd vdd FILL
XFILL_0__7224_ gnd vdd FILL
XFILL_4__12107_ gnd vdd FILL
XFILL_5__14446_ gnd vdd FILL
XFILL_3__15625_ gnd vdd FILL
XFILL_4__13087_ gnd vdd FILL
X_7852_ _7852_/A gnd _7852_/Y vdd INVX1
XFILL_5__11658_ gnd vdd FILL
XFILL_4__10299_ gnd vdd FILL
XFILL_3__12837_ gnd vdd FILL
XFILL_2__14266_ gnd vdd FILL
XFILL_2__11478_ gnd vdd FILL
XFILL_0__15445_ gnd vdd FILL
XFILL_0__12657_ gnd vdd FILL
XSFILL59160x47050 gnd vdd FILL
XFILL_1__14996_ gnd vdd FILL
XFILL_5__9938_ gnd vdd FILL
XFILL_2__16005_ gnd vdd FILL
XFILL_4__12038_ gnd vdd FILL
XFILL_6__15736_ gnd vdd FILL
XFILL_2__13217_ gnd vdd FILL
XFILL_5__14377_ gnd vdd FILL
XFILL_2__10429_ gnd vdd FILL
XFILL_3__12768_ gnd vdd FILL
XFILL_3__15556_ gnd vdd FILL
XFILL_5__11589_ gnd vdd FILL
X_7783_ _7721_/A _8679_/CLK _9959_/R vdd _7783_/D gnd vdd DFFSR
XFILL_2__14197_ gnd vdd FILL
XSFILL74200x50050 gnd vdd FILL
XFILL_0__11608_ gnd vdd FILL
XFILL_1__13947_ gnd vdd FILL
XFILL_3__8953_ gnd vdd FILL
XFILL_0_CLKBUF1_insert209 gnd vdd FILL
XFILL_0__15376_ gnd vdd FILL
XFILL_5__16116_ gnd vdd FILL
XFILL_0__12588_ gnd vdd FILL
XFILL_5__13328_ gnd vdd FILL
XFILL_5__9869_ gnd vdd FILL
XFILL111880x46050 gnd vdd FILL
X_9522_ _9578_/Q gnd _9522_/Y vdd INVX1
XFILL_3__14507_ gnd vdd FILL
XFILL_0__7086_ gnd vdd FILL
XFILL_3__11719_ gnd vdd FILL
XFILL_2__13148_ gnd vdd FILL
XFILL_3__12699_ gnd vdd FILL
XFILL_0__14327_ gnd vdd FILL
XFILL_3__15487_ gnd vdd FILL
XFILL_1__13878_ gnd vdd FILL
XFILL_3__8884_ gnd vdd FILL
XFILL_0__11539_ gnd vdd FILL
XFILL_5__16047_ gnd vdd FILL
XFILL_5__13259_ gnd vdd FILL
X_9453_ _9453_/Q _9453_/CLK _9453_/R vdd _9405_/Y gnd vdd DFFSR
XFILL_6__15598_ gnd vdd FILL
XSFILL109400x78050 gnd vdd FILL
XFILL_1__15617_ gnd vdd FILL
XFILL_3__14438_ gnd vdd FILL
XFILL_2__13079_ gnd vdd FILL
XFILL_4__13989_ gnd vdd FILL
XFILL_3__7835_ gnd vdd FILL
XFILL_1__12829_ gnd vdd FILL
XFILL_0__14258_ gnd vdd FILL
XSFILL8680x6050 gnd vdd FILL
XFILL_6__14549_ gnd vdd FILL
X_8404_ _8365_/A _7380_/B gnd _8404_/Y vdd NAND2X1
XFILL_4__15728_ gnd vdd FILL
XFILL_1__6850_ gnd vdd FILL
XSFILL54040x8050 gnd vdd FILL
X_9384_ _9382_/Y _9359_/A _9384_/C gnd _9446_/D vdd OAI21X1
XFILL_3__14369_ gnd vdd FILL
XSFILL89400x6050 gnd vdd FILL
XFILL_0__13209_ gnd vdd FILL
XFILL_1__15548_ gnd vdd FILL
XFILL_0__14189_ gnd vdd FILL
XFILL_4_BUFX2_insert705 gnd vdd FILL
X_8335_ _8321_/B _8719_/B gnd _8336_/C vdd NAND2X1
XFILL_3__16108_ gnd vdd FILL
XFILL_4__15659_ gnd vdd FILL
XFILL_3__9505_ gnd vdd FILL
XFILL_4_BUFX2_insert716 gnd vdd FILL
XFILL_0__7988_ gnd vdd FILL
XFILL_4_BUFX2_insert727 gnd vdd FILL
XFILL_4_BUFX2_insert738 gnd vdd FILL
XFILL_1__15479_ gnd vdd FILL
XFILL_6__9214_ gnd vdd FILL
XFILL_3__7697_ gnd vdd FILL
XFILL_4_BUFX2_insert749 gnd vdd FILL
XFILL_1__8520_ gnd vdd FILL
XFILL_0__9727_ gnd vdd FILL
XFILL_0__6939_ gnd vdd FILL
XSFILL33800x16050 gnd vdd FILL
X_8266_ _8266_/A gnd _8268_/A vdd INVX1
XFILL_3__16039_ gnd vdd FILL
XSFILL43960x60050 gnd vdd FILL
XFILL_1__8451_ gnd vdd FILL
XFILL_0__9658_ gnd vdd FILL
X_7217_ _7217_/A _7202_/B _7216_/Y gnd _7217_/Y vdd OAI21X1
XFILL_3__9367_ gnd vdd FILL
X_8197_ _8283_/Q gnd _8197_/Y vdd INVX1
XFILL_0__8609_ gnd vdd FILL
XFILL_1__8382_ gnd vdd FILL
X_7148_ _7148_/Q _9958_/CLK _8929_/R vdd _7098_/Y gnd vdd DFFSR
XFILL_4__7111_ gnd vdd FILL
XFILL_3__8318_ gnd vdd FILL
XFILL_4__8091_ gnd vdd FILL
XFILL_3__9298_ gnd vdd FILL
XFILL_1__7333_ gnd vdd FILL
X_7079_ _7100_/A _7079_/B gnd _7080_/C vdd NAND2X1
XFILL_3__8249_ gnd vdd FILL
XFILL_4__7042_ gnd vdd FILL
XSFILL23720x68050 gnd vdd FILL
XFILL_5_BUFX2_insert1090 gnd vdd FILL
XFILL_1__9003_ gnd vdd FILL
XFILL_1_BUFX2_insert606 gnd vdd FILL
XFILL_1__7195_ gnd vdd FILL
XSFILL64200x82050 gnd vdd FILL
XFILL_1_BUFX2_insert617 gnd vdd FILL
XFILL_1_BUFX2_insert628 gnd vdd FILL
X_11720_ _11720_/A _11720_/B gnd _11721_/C vdd NAND2X1
XFILL_4__8993_ gnd vdd FILL
XFILL_1_BUFX2_insert639 gnd vdd FILL
XFILL_4__7944_ gnd vdd FILL
X_11651_ _11281_/Y gnd _11651_/Y vdd INVX1
X_10602_ _15878_/A _9194_/CLK _7796_/R vdd _10602_/D gnd vdd DFFSR
X_14370_ _14370_/A _14045_/A _13467_/A _14370_/D gnd _14374_/A vdd OAI22X1
XFILL_4__7875_ gnd vdd FILL
XFILL_1__9905_ gnd vdd FILL
XSFILL84120x33050 gnd vdd FILL
X_11582_ _11406_/Y _11626_/C _11582_/C gnd _11583_/A vdd AOI21X1
XFILL_4__9614_ gnd vdd FILL
XFILL_2__6890_ gnd vdd FILL
X_13321_ _13220_/A _13239_/B gnd _13321_/Y vdd NOR2X1
X_10533_ _10531_/Y _10511_/A _10533_/C gnd _10597_/D vdd OAI21X1
XFILL_5_BUFX2_insert550 gnd vdd FILL
XFILL_5_BUFX2_insert561 gnd vdd FILL
XFILL_5_BUFX2_insert572 gnd vdd FILL
X_16040_ _7918_/Q gnd _16041_/A vdd INVX1
XFILL_4__9545_ gnd vdd FILL
X_13252_ _13252_/A _13249_/Y gnd _13252_/Y vdd NOR2X1
XFILL_5_BUFX2_insert583 gnd vdd FILL
X_10464_ _13972_/A _8815_/CLK _8047_/R vdd _10464_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert594 gnd vdd FILL
XFILL_1__9767_ gnd vdd FILL
XSFILL88760x36050 gnd vdd FILL
XFILL_1__6979_ gnd vdd FILL
X_12203_ _12179_/A _12910_/A gnd _12204_/C vdd NAND2X1
XFILL_4__9476_ gnd vdd FILL
X_13183_ _13103_/A _9060_/CLK _9060_/R vdd _13183_/D gnd vdd DFFSR
XFILL_1__8718_ gnd vdd FILL
X_10395_ _10395_/A _7579_/B gnd _10396_/C vdd NAND2X1
XSFILL49240x59050 gnd vdd FILL
XSFILL23400x50050 gnd vdd FILL
XFILL_2__8491_ gnd vdd FILL
XFILL_5__7220_ gnd vdd FILL
X_12134_ _12134_/A _12841_/A gnd _12135_/C vdd NAND2X1
XFILL_5__10960_ gnd vdd FILL
XFILL_3__10050_ gnd vdd FILL
XSFILL38840x8050 gnd vdd FILL
XFILL_2__7442_ gnd vdd FILL
XFILL_1__8649_ gnd vdd FILL
XFILL_2_CLKBUF1_insert120 gnd vdd FILL
XFILL_4__8358_ gnd vdd FILL
XFILL_2__10780_ gnd vdd FILL
XFILL_2_CLKBUF1_insert131 gnd vdd FILL
XFILL_2_CLKBUF1_insert142 gnd vdd FILL
X_12065_ _12065_/A _12093_/B _12061_/C gnd gnd _12066_/C vdd AOI22X1
XFILL_4__11340_ gnd vdd FILL
XFILL_2_CLKBUF1_insert153 gnd vdd FILL
XFILL_2__7373_ gnd vdd FILL
XFILL_2_CLKBUF1_insert164 gnd vdd FILL
XFILL_5__10891_ gnd vdd FILL
XFILL_1__11160_ gnd vdd FILL
XFILL_0__10910_ gnd vdd FILL
XFILL_4__7309_ gnd vdd FILL
XFILL_2_CLKBUF1_insert175 gnd vdd FILL
XFILL_5__7082_ gnd vdd FILL
X_11016_ _11012_/Y _11008_/Y _11015_/Y gnd _11016_/Y vdd OAI21X1
XFILL_5__12630_ gnd vdd FILL
XFILL_2_CLKBUF1_insert186 gnd vdd FILL
XFILL_2__9112_ gnd vdd FILL
XFILL_0__11890_ gnd vdd FILL
XFILL_1__10111_ gnd vdd FILL
XFILL_4__11271_ gnd vdd FILL
XFILL_2_CLKBUF1_insert197 gnd vdd FILL
XFILL_2__12450_ gnd vdd FILL
XFILL_1__11091_ gnd vdd FILL
XFILL_4__13010_ gnd vdd FILL
XFILL_6__13920_ gnd vdd FILL
XSFILL84200x13050 gnd vdd FILL
X_15824_ _15822_/Y _15824_/B _15824_/C gnd _15824_/Y vdd NAND3X1
XSFILL28920x81050 gnd vdd FILL
XFILL_2__11401_ gnd vdd FILL
XFILL_2__9043_ gnd vdd FILL
XFILL_3__10952_ gnd vdd FILL
XFILL_1__10042_ gnd vdd FILL
XFILL_3__13740_ gnd vdd FILL
XFILL_2_BUFX2_insert440 gnd vdd FILL
XSFILL104360x19050 gnd vdd FILL
XFILL_2_BUFX2_insert451 gnd vdd FILL
XFILL_2__12381_ gnd vdd FILL
XFILL_2_BUFX2_insert462 gnd vdd FILL
XFILL_5__14300_ gnd vdd FILL
XFILL_0__13560_ gnd vdd FILL
XFILL_0__10772_ gnd vdd FILL
XSFILL69000x74050 gnd vdd FILL
XBUFX2_insert8 _13280_/Y gnd _7336_/B vdd BUFX2
XFILL_2_BUFX2_insert473 gnd vdd FILL
XFILL_5__11512_ gnd vdd FILL
XFILL_4__10153_ gnd vdd FILL
XFILL_2__14120_ gnd vdd FILL
XFILL_5__15280_ gnd vdd FILL
X_12967_ vdd _12967_/B gnd _12967_/Y vdd NAND2X1
X_15755_ _7721_/A gnd _15755_/Y vdd INVX1
XFILL_3__13671_ gnd vdd FILL
XFILL_5__12492_ gnd vdd FILL
XFILL_2_BUFX2_insert484 gnd vdd FILL
XFILL_2__11332_ gnd vdd FILL
XFILL_1__14850_ gnd vdd FILL
XFILL_0__12511_ gnd vdd FILL
XFILL_3__10883_ gnd vdd FILL
XFILL_2_BUFX2_insert495 gnd vdd FILL
XFILL_5__14231_ gnd vdd FILL
X_14706_ _10736_/Q gnd _16106_/B vdd INVX1
X_11918_ _11900_/A _12027_/B gnd _11919_/C vdd NAND2X1
XFILL_0__13491_ gnd vdd FILL
XFILL_3__12622_ gnd vdd FILL
XFILL_3__15410_ gnd vdd FILL
XFILL_5__7984_ gnd vdd FILL
XFILL_5__11443_ gnd vdd FILL
XFILL_1__13801_ gnd vdd FILL
X_15686_ _15686_/A _15407_/B _15407_/C _14175_/Y gnd _15688_/A vdd OAI22X1
XFILL_2__14051_ gnd vdd FILL
XFILL_4__14961_ gnd vdd FILL
X_12898_ _12898_/A gnd _12900_/A vdd INVX1
XFILL_3__16390_ gnd vdd FILL
XFILL_0__15230_ gnd vdd FILL
XFILL_2__11263_ gnd vdd FILL
XFILL_6__15521_ gnd vdd FILL
XFILL_0__12442_ gnd vdd FILL
XSFILL48840x32050 gnd vdd FILL
XFILL_5__9723_ gnd vdd FILL
XFILL_1__14781_ gnd vdd FILL
XFILL_6__12733_ gnd vdd FILL
XSFILL99480x67050 gnd vdd FILL
XFILL_5__6935_ gnd vdd FILL
XFILL_1__11993_ gnd vdd FILL
XSFILL64040x3050 gnd vdd FILL
X_14637_ _14636_/Y _14637_/B gnd _14645_/A vdd NOR2X1
XFILL_5__14162_ gnd vdd FILL
XFILL_4__13912_ gnd vdd FILL
X_11849_ _11849_/A _11849_/B _11848_/Y gnd _12440_/A vdd NAND3X1
XFILL_2__13002_ gnd vdd FILL
XSFILL74120x65050 gnd vdd FILL
XFILL_3__15341_ gnd vdd FILL
XFILL_5__11374_ gnd vdd FILL
XFILL_1__13732_ gnd vdd FILL
XFILL_4__14892_ gnd vdd FILL
XFILL_1__10944_ gnd vdd FILL
XFILL_0__12373_ gnd vdd FILL
XFILL_0__15161_ gnd vdd FILL
XFILL_2__11194_ gnd vdd FILL
XFILL_5__9654_ gnd vdd FILL
XFILL_5__13113_ gnd vdd FILL
XFILL_0__8960_ gnd vdd FILL
X_14568_ _14568_/A _14567_/Y gnd _14568_/Y vdd NOR2X1
XFILL_5__6866_ gnd vdd FILL
XFILL_3__11504_ gnd vdd FILL
XFILL_5__10325_ gnd vdd FILL
XFILL_4__13843_ gnd vdd FILL
XFILL_5__14093_ gnd vdd FILL
XFILL_3__15272_ gnd vdd FILL
XFILL_1__16451_ gnd vdd FILL
XFILL_3__12484_ gnd vdd FILL
XFILL_2__10145_ gnd vdd FILL
XBUFX2_insert450 _13276_/Y gnd _7202_/B vdd BUFX2
XFILL_0__11324_ gnd vdd FILL
XFILL_0__14112_ gnd vdd FILL
XFILL_1__13663_ gnd vdd FILL
XSFILL3400x28050 gnd vdd FILL
XFILL_2__9876_ gnd vdd FILL
XFILL_5__8605_ gnd vdd FILL
XBUFX2_insert461 _15044_/Y gnd _15760_/A vdd BUFX2
XFILL_1__10875_ gnd vdd FILL
X_16307_ _16307_/A _16306_/Y gnd _16307_/Y vdd NOR2X1
XFILL_0__15092_ gnd vdd FILL
XFILL_6__11615_ gnd vdd FILL
XFILL_5__10256_ gnd vdd FILL
XFILL_6__15383_ gnd vdd FILL
XFILL_3__14223_ gnd vdd FILL
XBUFX2_insert472 _15041_/Y gnd _15708_/C vdd BUFX2
XFILL_5__13044_ gnd vdd FILL
X_13519_ _13518_/Y _13519_/B gnd _13532_/A vdd NAND2X1
XFILL_1__15402_ gnd vdd FILL
X_14499_ _14499_/A _14483_/Y gnd _14500_/A vdd NOR2X1
XFILL_0__8891_ gnd vdd FILL
XBUFX2_insert483 _14979_/Y gnd _15313_/B vdd BUFX2
XFILL_3__7620_ gnd vdd FILL
XFILL_3__11435_ gnd vdd FILL
XFILL_4__13774_ gnd vdd FILL
XFILL_1__12614_ gnd vdd FILL
XBUFX2_insert494 BUFX2_insert494/A gnd _9964_/R vdd BUFX2
XFILL_2__8827_ gnd vdd FILL
XFILL_1__16382_ gnd vdd FILL
XFILL_0__14043_ gnd vdd FILL
XFILL_2__14953_ gnd vdd FILL
XFILL_0__11255_ gnd vdd FILL
XFILL_1__13594_ gnd vdd FILL
XFILL_6__14334_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1076 gnd vdd FILL
X_16238_ _14855_/Y _15203_/B _16237_/Y gnd _16238_/Y vdd OAI21X1
XFILL_0__7842_ gnd vdd FILL
XFILL_4__15513_ gnd vdd FILL
XFILL_4__12725_ gnd vdd FILL
XFILL_5__10187_ gnd vdd FILL
XFILL_3__14154_ gnd vdd FILL
XFILL_3__7551_ gnd vdd FILL
XFILL_1__15333_ gnd vdd FILL
XFILL_2__13904_ gnd vdd FILL
XFILL_3__11366_ gnd vdd FILL
XFILL_2__8758_ gnd vdd FILL
XSFILL54040x32050 gnd vdd FILL
XFILL_2__14884_ gnd vdd FILL
XFILL_0__11186_ gnd vdd FILL
X_8120_ _8120_/A gnd _8122_/A vdd INVX1
XFILL_3__13105_ gnd vdd FILL
XFILL_5__8467_ gnd vdd FILL
XFILL_3__10317_ gnd vdd FILL
X_16169_ _9802_/A gnd _16170_/B vdd INVX1
XFILL_6__11477_ gnd vdd FILL
XFILL_4__15444_ gnd vdd FILL
XFILL_4__12656_ gnd vdd FILL
XFILL_2__13835_ gnd vdd FILL
XFILL_5__14995_ gnd vdd FILL
XFILL_2__7709_ gnd vdd FILL
XFILL_3__14085_ gnd vdd FILL
XFILL_0__10137_ gnd vdd FILL
XFILL_3__7482_ gnd vdd FILL
XFILL_3__11297_ gnd vdd FILL
XFILL_1__15264_ gnd vdd FILL
XFILL_0__9512_ gnd vdd FILL
XFILL_1__12476_ gnd vdd FILL
XFILL_5__7418_ gnd vdd FILL
XFILL_5__8398_ gnd vdd FILL
XFILL_0__15994_ gnd vdd FILL
X_8051_ _8013_/A _8051_/CLK _8051_/R vdd _8051_/D gnd vdd DFFSR
XFILL_6__14196_ gnd vdd FILL
XFILL_3__13036_ gnd vdd FILL
XFILL_4__11607_ gnd vdd FILL
XFILL_5__13946_ gnd vdd FILL
XFILL_3__9221_ gnd vdd FILL
XSFILL43880x75050 gnd vdd FILL
XFILL_3__10248_ gnd vdd FILL
XFILL_4__15375_ gnd vdd FILL
XFILL_1__14215_ gnd vdd FILL
XFILL_4__12587_ gnd vdd FILL
XFILL_2__13766_ gnd vdd FILL
XFILL_1__11427_ gnd vdd FILL
XFILL_2__10978_ gnd vdd FILL
XFILL_1__15195_ gnd vdd FILL
XFILL_0__10068_ gnd vdd FILL
XFILL_0__14945_ gnd vdd FILL
XSFILL109320x3050 gnd vdd FILL
XFILL_5__7349_ gnd vdd FILL
X_7002_ _7002_/Q _8541_/CLK _7258_/R vdd _7002_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert12 gnd vdd FILL
XFILL_4__14326_ gnd vdd FILL
XFILL_2__12717_ gnd vdd FILL
XFILL_5__13877_ gnd vdd FILL
XFILL_3__9152_ gnd vdd FILL
XFILL_2__15505_ gnd vdd FILL
XFILL_4__11538_ gnd vdd FILL
XSFILL48920x12050 gnd vdd FILL
XFILL_1_BUFX2_insert23 gnd vdd FILL
XFILL_1_BUFX2_insert34 gnd vdd FILL
XSFILL18680x51050 gnd vdd FILL
XFILL_1__14146_ gnd vdd FILL
XFILL_3__10179_ gnd vdd FILL
XFILL_1_BUFX2_insert45 gnd vdd FILL
XFILL_2__13697_ gnd vdd FILL
XSFILL49400x19050 gnd vdd FILL
XFILL_1__11358_ gnd vdd FILL
XFILL_0__14876_ gnd vdd FILL
XFILL_5__15616_ gnd vdd FILL
XSFILL74200x45050 gnd vdd FILL
XFILL_1_BUFX2_insert56 gnd vdd FILL
XFILL_3__8103_ gnd vdd FILL
XFILL_0__9374_ gnd vdd FILL
XFILL_5__12828_ gnd vdd FILL
XSFILL89800x24050 gnd vdd FILL
XFILL_4__14257_ gnd vdd FILL
XFILL_1_BUFX2_insert67 gnd vdd FILL
XFILL_2__12648_ gnd vdd FILL
XFILL_1_BUFX2_insert78 gnd vdd FILL
XFILL_1__10309_ gnd vdd FILL
XFILL_2__15436_ gnd vdd FILL
XFILL_4__11469_ gnd vdd FILL
XFILL_3__9083_ gnd vdd FILL
XFILL_5__9019_ gnd vdd FILL
XFILL_0__13827_ gnd vdd FILL
XFILL_1_BUFX2_insert89 gnd vdd FILL
XFILL_3__14987_ gnd vdd FILL
XFILL_1__14077_ gnd vdd FILL
XFILL_6__9901_ gnd vdd FILL
XFILL_6__12029_ gnd vdd FILL
XFILL_1__11289_ gnd vdd FILL
XFILL_0__8325_ gnd vdd FILL
XSFILL49000x21050 gnd vdd FILL
XFILL_4__13208_ gnd vdd FILL
XFILL_5__15547_ gnd vdd FILL
XFILL_5__12759_ gnd vdd FILL
X_8953_ _9047_/Q gnd _8955_/A vdd INVX1
XFILL_2__15367_ gnd vdd FILL
XFILL_4__14188_ gnd vdd FILL
XFILL_3__13938_ gnd vdd FILL
XFILL_1__13028_ gnd vdd FILL
XFILL_2__12579_ gnd vdd FILL
XFILL_0__13758_ gnd vdd FILL
XFILL_0__8256_ gnd vdd FILL
XSFILL109560x32050 gnd vdd FILL
X_7904_ _7828_/A _9568_/CLK _7648_/R vdd _7830_/Y gnd vdd DFFSR
XFILL_4__13139_ gnd vdd FILL
XFILL_2__14318_ gnd vdd FILL
XFILL_5__15478_ gnd vdd FILL
X_8884_ _8884_/A _8854_/B _8883_/Y gnd _8884_/Y vdd OAI21X1
XFILL_3__13869_ gnd vdd FILL
XFILL_0__12709_ gnd vdd FILL
XFILL_2__15298_ gnd vdd FILL
XSFILL38040x45050 gnd vdd FILL
XSFILL38840x64050 gnd vdd FILL
XFILL_0__7207_ gnd vdd FILL
XFILL112360x71050 gnd vdd FILL
XSFILL54120x12050 gnd vdd FILL
XFILL_0__13689_ gnd vdd FILL
XFILL_5__14429_ gnd vdd FILL
XFILL_6__6975_ gnd vdd FILL
X_7835_ _7800_/B _7579_/B gnd _7836_/C vdd NAND2X1
XFILL_3__15608_ gnd vdd FILL
XFILL_0__8187_ gnd vdd FILL
XFILL_2__14249_ gnd vdd FILL
XFILL_0__15428_ gnd vdd FILL
XFILL_3__9985_ gnd vdd FILL
XFILL_1__14979_ gnd vdd FILL
XFILL_3__15539_ gnd vdd FILL
X_7766_ _7766_/Q _8818_/CLK _8278_/R vdd _7766_/D gnd vdd DFFSR
XSFILL39000x50 gnd vdd FILL
XFILL_0__15359_ gnd vdd FILL
X_9505_ _9533_/B _9633_/B gnd _9506_/C vdd NAND2X1
XSFILL43960x55050 gnd vdd FILL
XFILL_6__8645_ gnd vdd FILL
XFILL_1__7951_ gnd vdd FILL
XFILL_0__7069_ gnd vdd FILL
X_7697_ _7697_/A gnd _7699_/A vdd INVX1
XFILL_3__8867_ gnd vdd FILL
XFILL_1__6902_ gnd vdd FILL
X_9436_ _9352_/A _9436_/CLK _9454_/R vdd _9436_/D gnd vdd DFFSR
XSFILL18760x31050 gnd vdd FILL
XFILL_1__7882_ gnd vdd FILL
XSFILL8600x41050 gnd vdd FILL
XSFILL44040x64050 gnd vdd FILL
XFILL_3__7818_ gnd vdd FILL
XFILL_4__7591_ gnd vdd FILL
XFILL_1__9621_ gnd vdd FILL
X_9367_ _9367_/A gnd _9367_/Y vdd INVX1
XFILL_4_BUFX2_insert502 gnd vdd FILL
XFILL_4_BUFX2_insert513 gnd vdd FILL
XFILL_4_BUFX2_insert524 gnd vdd FILL
XFILL_3__7749_ gnd vdd FILL
XFILL_4_BUFX2_insert535 gnd vdd FILL
X_8318_ _8318_/A _8315_/B _8318_/C gnd _8408_/D vdd OAI21X1
XFILL_1__9552_ gnd vdd FILL
XFILL_4_BUFX2_insert546 gnd vdd FILL
XSFILL23880x22050 gnd vdd FILL
XFILL_4__9261_ gnd vdd FILL
XFILL_4_BUFX2_insert557 gnd vdd FILL
X_9298_ _9296_/Y _9282_/A _9298_/C gnd _9332_/D vdd OAI21X1
XFILL_4_BUFX2_insert568 gnd vdd FILL
XFILL_1__8503_ gnd vdd FILL
XFILL_4_BUFX2_insert579 gnd vdd FILL
X_10180_ _14732_/A gnd _10182_/A vdd INVX1
XFILL_1__9483_ gnd vdd FILL
X_8249_ _8249_/A _8377_/B gnd _8250_/C vdd NAND2X1
XFILL_4__8212_ gnd vdd FILL
XSFILL89560x79050 gnd vdd FILL
XFILL_3__9419_ gnd vdd FILL
XSFILL38920x44050 gnd vdd FILL
XFILL112440x51050 gnd vdd FILL
XSFILL64200x77050 gnd vdd FILL
XSFILL39560x10050 gnd vdd FILL
XFILL_4__8143_ gnd vdd FILL
XFILL_1__8365_ gnd vdd FILL
XFILL_4__8074_ gnd vdd FILL
XFILL_3_CLKBUF1_insert204 gnd vdd FILL
XFILL_3_CLKBUF1_insert215 gnd vdd FILL
X_13870_ _10334_/Q gnd _13871_/C vdd INVX1
XFILL_1__7316_ gnd vdd FILL
XSFILL109480x9050 gnd vdd FILL
XSFILL18840x11050 gnd vdd FILL
X_12821_ _12785_/A _12692_/CLK _12692_/R vdd _12821_/D gnd vdd DFFSR
XSFILL94280x72050 gnd vdd FILL
XFILL_1__7247_ gnd vdd FILL
XSFILL29480x62050 gnd vdd FILL
XFILL_1_BUFX2_insert403 gnd vdd FILL
XFILL_1_BUFX2_insert414 gnd vdd FILL
X_12752_ _11881_/A gnd _12754_/A vdd INVX1
XFILL_1_BUFX2_insert425 gnd vdd FILL
X_15540_ _15070_/C _14056_/Y _16199_/C _14030_/D gnd _15541_/B vdd OAI22X1
XFILL_1__7178_ gnd vdd FILL
XFILL_1_BUFX2_insert436 gnd vdd FILL
XFILL_1_BUFX2_insert447 gnd vdd FILL
XFILL_1_BUFX2_insert458 gnd vdd FILL
X_11703_ _11739_/B _11392_/Y _11703_/C gnd _11704_/C vdd OAI21X1
XFILL_4__8976_ gnd vdd FILL
X_15471_ _15471_/A _15469_/Y gnd _15471_/Y vdd NOR2X1
XFILL_1_BUFX2_insert469 gnd vdd FILL
X_12683_ _12683_/Q _12669_/CLK _12795_/R vdd _12683_/D gnd vdd DFFSR
XSFILL58920x50 gnd vdd FILL
XFILL_2__7991_ gnd vdd FILL
XFILL_4__7927_ gnd vdd FILL
X_14422_ _14413_/Y _14414_/Y _14422_/C gnd _14423_/B vdd NAND3X1
X_11634_ _11634_/A _11484_/B _11634_/C gnd _11635_/B vdd OAI21X1
XFILL_2__9730_ gnd vdd FILL
XFILL_2__6942_ gnd vdd FILL
XFILL_1_CLKBUF1_insert1082 gnd vdd FILL
XFILL_5__10110_ gnd vdd FILL
X_14353_ _14353_/A _7400_/Q _7852_/A _13865_/B gnd _14353_/Y vdd AOI22X1
XFILL_4__7858_ gnd vdd FILL
XFILL_5__11090_ gnd vdd FILL
X_11565_ _11565_/A _11521_/A gnd _11565_/Y vdd NOR2X1
XFILL_2__6873_ gnd vdd FILL
XFILL_2__9661_ gnd vdd FILL
XSFILL89240x61050 gnd vdd FILL
XSFILL53880x38050 gnd vdd FILL
XFILL_1__10660_ gnd vdd FILL
X_13304_ _13252_/A _13303_/Y gnd _13308_/B vdd NOR2X1
XFILL_6__11400_ gnd vdd FILL
XFILL_5__9370_ gnd vdd FILL
XFILL_5__10041_ gnd vdd FILL
X_10516_ _10592_/Q gnd _10516_/Y vdd INVX1
XFILL_3__11220_ gnd vdd FILL
X_14284_ _9641_/A gnd _14284_/Y vdd INVX1
XFILL_2__8612_ gnd vdd FILL
XFILL_5_BUFX2_insert380 gnd vdd FILL
XFILL_4__10771_ gnd vdd FILL
X_11496_ _11495_/Y _11494_/Y gnd _11497_/C vdd AND2X2
XSFILL3720x64050 gnd vdd FILL
XFILL_2__11950_ gnd vdd FILL
XFILL_5_BUFX2_insert391 gnd vdd FILL
XBUFX2_insert70 _13393_/Y gnd _13601_/B vdd BUFX2
XFILL_2__9592_ gnd vdd FILL
XFILL_0__11040_ gnd vdd FILL
XFILL_5__8321_ gnd vdd FILL
XFILL_4__9528_ gnd vdd FILL
XBUFX2_insert81 _13372_/Y gnd _14946_/A vdd BUFX2
XSFILL28680x14050 gnd vdd FILL
X_13235_ _13220_/A _13305_/A _13235_/C gnd _13235_/Y vdd OAI21X1
X_16023_ _7406_/Q gnd _16024_/A vdd INVX1
XBUFX2_insert92 _12357_/Y gnd _9347_/B vdd BUFX2
X_10447_ _10445_/Y _10443_/A _10447_/C gnd _10483_/D vdd OAI21X1
XFILL_4__12510_ gnd vdd FILL
XFILL_2__10901_ gnd vdd FILL
XFILL_3__11151_ gnd vdd FILL
XSFILL28920x76050 gnd vdd FILL
XFILL_4__13490_ gnd vdd FILL
XFILL_1__12330_ gnd vdd FILL
XFILL_5__8252_ gnd vdd FILL
XFILL_2__11881_ gnd vdd FILL
XSFILL94360x52050 gnd vdd FILL
XFILL_5__13800_ gnd vdd FILL
X_13166_ _11974_/A gnd _13166_/Y vdd INVX1
XFILL_3__10102_ gnd vdd FILL
XFILL_6__11262_ gnd vdd FILL
XFILL_4__12441_ gnd vdd FILL
X_10378_ _10378_/A _10405_/B _10377_/Y gnd _10378_/Y vdd OAI21X1
XFILL_2__13620_ gnd vdd FILL
XFILL_5__14780_ gnd vdd FILL
XFILL_2__8474_ gnd vdd FILL
XFILL_5__11992_ gnd vdd FILL
XFILL_3__11082_ gnd vdd FILL
XFILL_2__10832_ gnd vdd FILL
XFILL_5__7203_ gnd vdd FILL
XFILL_6__13001_ gnd vdd FILL
XFILL_1__12261_ gnd vdd FILL
XFILL_5__8183_ gnd vdd FILL
X_12117_ _12117_/A _12117_/B _12117_/C gnd _12117_/Y vdd OAI21X1
XFILL_5__13731_ gnd vdd FILL
XFILL_0__12991_ gnd vdd FILL
XFILL_5__10943_ gnd vdd FILL
XFILL_2__7425_ gnd vdd FILL
XFILL_4__12372_ gnd vdd FILL
X_13097_ _13097_/A gnd _13099_/A vdd INVX1
XFILL_1__14000_ gnd vdd FILL
XFILL_3__10033_ gnd vdd FILL
XFILL_4__15160_ gnd vdd FILL
XFILL_3__14910_ gnd vdd FILL
XFILL_2__13551_ gnd vdd FILL
XFILL_1__11212_ gnd vdd FILL
XFILL_2__10763_ gnd vdd FILL
XFILL_0__14730_ gnd vdd FILL
XFILL_3__15890_ gnd vdd FILL
XFILL_0__11942_ gnd vdd FILL
XFILL_1__12192_ gnd vdd FILL
XFILL_5__16450_ gnd vdd FILL
X_12048_ _12084_/A _11879_/B _12084_/C gnd _12050_/B vdd NAND3X1
XFILL_4__14111_ gnd vdd FILL
XFILL_2__12502_ gnd vdd FILL
XFILL_5__13662_ gnd vdd FILL
XFILL_4__11323_ gnd vdd FILL
XFILL_3__14841_ gnd vdd FILL
XFILL_2__7356_ gnd vdd FILL
XFILL_5__10874_ gnd vdd FILL
XFILL_2__16270_ gnd vdd FILL
XFILL_4__15091_ gnd vdd FILL
XFILL_1__11143_ gnd vdd FILL
XFILL_2__13482_ gnd vdd FILL
XFILL_5__15401_ gnd vdd FILL
XFILL_5__7065_ gnd vdd FILL
XFILL_2__10694_ gnd vdd FILL
XFILL_0__14661_ gnd vdd FILL
XFILL_0__11873_ gnd vdd FILL
XFILL_5__12613_ gnd vdd FILL
XFILL_2__15221_ gnd vdd FILL
XFILL_4__14042_ gnd vdd FILL
XFILL_5__16381_ gnd vdd FILL
XFILL_4__11254_ gnd vdd FILL
XFILL_5__13593_ gnd vdd FILL
XFILL_0__16400_ gnd vdd FILL
XFILL_2__12433_ gnd vdd FILL
XFILL_0__13612_ gnd vdd FILL
XFILL_3__11984_ gnd vdd FILL
XFILL_2__7287_ gnd vdd FILL
XFILL_1__15951_ gnd vdd FILL
XFILL_1__11074_ gnd vdd FILL
XFILL_3__14772_ gnd vdd FILL
XFILL_0__8110_ gnd vdd FILL
XFILL_0__10824_ gnd vdd FILL
XFILL_0__14592_ gnd vdd FILL
XFILL_5__15332_ gnd vdd FILL
X_15807_ _9192_/Q gnd _15808_/C vdd INVX1
XFILL_0__9090_ gnd vdd FILL
XFILL_2__9026_ gnd vdd FILL
XFILL_2_BUFX2_insert270 gnd vdd FILL
XFILL_3__13723_ gnd vdd FILL
XFILL_4__11185_ gnd vdd FILL
XFILL_2__15152_ gnd vdd FILL
XFILL_3__10935_ gnd vdd FILL
XFILL_2__12364_ gnd vdd FILL
XFILL_0__16331_ gnd vdd FILL
XFILL_2_BUFX2_insert281 gnd vdd FILL
XSFILL109480x47050 gnd vdd FILL
X_13999_ _7959_/A gnd _13999_/Y vdd INVX1
XFILL_1__14902_ gnd vdd FILL
XFILL_1__10025_ gnd vdd FILL
XFILL_2_BUFX2_insert292 gnd vdd FILL
XFILL_0__13543_ gnd vdd FILL
XFILL_1__15882_ gnd vdd FILL
XFILL_0__10755_ gnd vdd FILL
XFILL_4__10136_ gnd vdd FILL
X_15738_ _10343_/Q _16166_/A gnd _15740_/B vdd NAND2X1
XFILL_2__14103_ gnd vdd FILL
XFILL_5__15263_ gnd vdd FILL
XSFILL38760x79050 gnd vdd FILL
XFILL_5__12475_ gnd vdd FILL
XFILL_2__11315_ gnd vdd FILL
XFILL_4__15993_ gnd vdd FILL
XFILL_3__13654_ gnd vdd FILL
XFILL_1__14833_ gnd vdd FILL
XFILL_2__15083_ gnd vdd FILL
XFILL_2__12295_ gnd vdd FILL
XSFILL54040x27050 gnd vdd FILL
XFILL_0__16262_ gnd vdd FILL
XFILL_0__10686_ gnd vdd FILL
XFILL_5__14214_ gnd vdd FILL
XFILL_0__13474_ gnd vdd FILL
X_7620_ _7620_/A gnd _7622_/A vdd INVX1
XFILL_5__7967_ gnd vdd FILL
XFILL_5__11426_ gnd vdd FILL
XFILL_3__12605_ gnd vdd FILL
XFILL_5__15194_ gnd vdd FILL
X_15669_ _9829_/Q _15390_/B gnd _15679_/A vdd NAND2X1
XFILL_1_BUFX2_insert970 gnd vdd FILL
XFILL_2__14034_ gnd vdd FILL
XFILL_4__10067_ gnd vdd FILL
XFILL_4__14944_ gnd vdd FILL
XSFILL94440x32050 gnd vdd FILL
XFILL_0__15213_ gnd vdd FILL
XFILL_2__11246_ gnd vdd FILL
XFILL_3__16373_ gnd vdd FILL
XFILL_3__9770_ gnd vdd FILL
XFILL_3__13585_ gnd vdd FILL
XFILL_0__12425_ gnd vdd FILL
XFILL_3__6982_ gnd vdd FILL
XFILL_3__10797_ gnd vdd FILL
XFILL_1_BUFX2_insert981 gnd vdd FILL
XFILL_1__14764_ gnd vdd FILL
XFILL_1_BUFX2_insert992 gnd vdd FILL
XFILL_1__11976_ gnd vdd FILL
XFILL_0__16193_ gnd vdd FILL
XFILL_5__6918_ gnd vdd FILL
XFILL_5__14145_ gnd vdd FILL
X_7551_ _7641_/Q gnd _7551_/Y vdd INVX1
XFILL_3__15324_ gnd vdd FILL
XFILL_5__11357_ gnd vdd FILL
XFILL_4__14875_ gnd vdd FILL
XFILL_0__9992_ gnd vdd FILL
XFILL_1__13715_ gnd vdd FILL
XFILL_3__8721_ gnd vdd FILL
XFILL_2__9928_ gnd vdd FILL
XFILL_1__10927_ gnd vdd FILL
XFILL_0__15144_ gnd vdd FILL
XFILL_2__11177_ gnd vdd FILL
XFILL_5__9637_ gnd vdd FILL
XFILL_0__12356_ gnd vdd FILL
XFILL_1__14695_ gnd vdd FILL
XFILL_5__6849_ gnd vdd FILL
XFILL_5__10308_ gnd vdd FILL
XFILL_4__13826_ gnd vdd FILL
XFILL_5__14076_ gnd vdd FILL
XFILL_2__10128_ gnd vdd FILL
XFILL_3__15255_ gnd vdd FILL
XBUFX2_insert280 _13419_/Y gnd _13617_/D vdd BUFX2
X_7482_ _7482_/A _7457_/A _7482_/C gnd _7532_/D vdd OAI21X1
XFILL_3__12467_ gnd vdd FILL
XFILL_5__11288_ gnd vdd FILL
XFILL_3__8652_ gnd vdd FILL
XFILL_2__9859_ gnd vdd FILL
XFILL_1__13646_ gnd vdd FILL
XSFILL18680x46050 gnd vdd FILL
XFILL_0__11307_ gnd vdd FILL
XFILL_2__15985_ gnd vdd FILL
XFILL_0__15075_ gnd vdd FILL
XBUFX2_insert291 _13356_/Y gnd _10325_/B vdd BUFX2
XFILL_0__12287_ gnd vdd FILL
XFILL_6__8361_ gnd vdd FILL
XFILL_5__13027_ gnd vdd FILL
X_9221_ _9221_/A gnd _9223_/A vdd INVX1
XFILL_6__12578_ gnd vdd FILL
XFILL_5__10239_ gnd vdd FILL
XFILL_3__14206_ gnd vdd FILL
XFILL_0__8874_ gnd vdd FILL
XFILL_3__11418_ gnd vdd FILL
XFILL_4__13757_ gnd vdd FILL
XFILL_3__7603_ gnd vdd FILL
XFILL_4__10969_ gnd vdd FILL
XFILL_3__12398_ gnd vdd FILL
XFILL_3__15186_ gnd vdd FILL
XFILL_2__10059_ gnd vdd FILL
XFILL_1__16365_ gnd vdd FILL
XFILL_0__14026_ gnd vdd FILL
XFILL_2__14936_ gnd vdd FILL
XFILL_3__8583_ gnd vdd FILL
XFILL_6__7312_ gnd vdd FILL
XFILL_5__8519_ gnd vdd FILL
XFILL_1__13577_ gnd vdd FILL
XFILL_0__11238_ gnd vdd FILL
XFILL_1__10789_ gnd vdd FILL
XFILL_5_CLKBUF1_insert170 gnd vdd FILL
XFILL_0__7825_ gnd vdd FILL
XFILL_5_CLKBUF1_insert181 gnd vdd FILL
XFILL_4__12708_ gnd vdd FILL
X_9152_ _9150_/Y _9151_/A _9152_/C gnd _9198_/D vdd OAI21X1
XFILL_5__9499_ gnd vdd FILL
XSFILL49000x16050 gnd vdd FILL
XFILL_5_CLKBUF1_insert192 gnd vdd FILL
XFILL_1__15316_ gnd vdd FILL
XFILL_3__14137_ gnd vdd FILL
XFILL_3__11349_ gnd vdd FILL
XFILL_1__12528_ gnd vdd FILL
XFILL_4__13688_ gnd vdd FILL
XSFILL89400x21050 gnd vdd FILL
XFILL_2__14867_ gnd vdd FILL
XSFILL59160x60050 gnd vdd FILL
XFILL_1__16296_ gnd vdd FILL
XFILL_0__11169_ gnd vdd FILL
X_8103_ _8142_/A _9383_/B gnd _8104_/C vdd NAND2X1
XFILL_0__7756_ gnd vdd FILL
XSFILL109560x27050 gnd vdd FILL
XFILL_4__15427_ gnd vdd FILL
XFILL_4__12639_ gnd vdd FILL
XFILL_3__14068_ gnd vdd FILL
XFILL_5__14978_ gnd vdd FILL
X_9083_ _9081_/Y _9116_/B _9082_/Y gnd _9083_/Y vdd OAI21X1
XFILL_2__13818_ gnd vdd FILL
XFILL_1__15247_ gnd vdd FILL
XFILL_3__7465_ gnd vdd FILL
XFILL_3_BUFX2_insert509 gnd vdd FILL
XFILL_1__12459_ gnd vdd FILL
XFILL_0__15977_ gnd vdd FILL
XSFILL38840x59050 gnd vdd FILL
XFILL_2__14798_ gnd vdd FILL
XFILL112360x66050 gnd vdd FILL
XFILL_3__13019_ gnd vdd FILL
X_8034_ _8034_/Q _7382_/CLK _8034_/R vdd _7964_/Y gnd vdd DFFSR
XFILL_5__13929_ gnd vdd FILL
XFILL_4__15358_ gnd vdd FILL
XFILL_0__7687_ gnd vdd FILL
XFILL_1__15178_ gnd vdd FILL
XFILL_2__13749_ gnd vdd FILL
XSFILL94520x12050 gnd vdd FILL
XFILL_0__14928_ gnd vdd FILL
XFILL_0__9426_ gnd vdd FILL
XFILL_4__14309_ gnd vdd FILL
XFILL_1__14129_ gnd vdd FILL
XFILL_3__9135_ gnd vdd FILL
XFILL_4__15289_ gnd vdd FILL
XFILL_0__14859_ gnd vdd FILL
XSFILL79320x73050 gnd vdd FILL
XFILL_0__9357_ gnd vdd FILL
X_9985_ _9983_/Y _9985_/B _9984_/Y gnd _9985_/Y vdd OAI21X1
XFILL_2__15419_ gnd vdd FILL
XFILL_1__7101_ gnd vdd FILL
XFILL_2__16399_ gnd vdd FILL
X_8936_ _8936_/Q _7400_/CLK _9704_/R vdd _8936_/D gnd vdd DFFSR
XFILL_0__9288_ gnd vdd FILL
XFILL_1__8081_ gnd vdd FILL
XFILL_3__8017_ gnd vdd FILL
XSFILL18760x26050 gnd vdd FILL
XSFILL114520x82050 gnd vdd FILL
XSFILL8600x36050 gnd vdd FILL
XSFILL44040x59050 gnd vdd FILL
XSFILL18200x69050 gnd vdd FILL
XFILL_1__7032_ gnd vdd FILL
XFILL_0__8239_ gnd vdd FILL
X_8867_ _8933_/Q gnd _8867_/Y vdd INVX1
XFILL_4__8830_ gnd vdd FILL
XFILL_6__9746_ gnd vdd FILL
X_7818_ _7816_/Y _7824_/B _7818_/C gnd _7900_/D vdd OAI21X1
XSFILL23880x17050 gnd vdd FILL
X_8798_ _8718_/A _7902_/CLK _7150_/R vdd _8798_/D gnd vdd DFFSR
XFILL_4__8761_ gnd vdd FILL
X_7749_ _7729_/B _9797_/B gnd _7749_/Y vdd NAND2X1
XFILL_1__8983_ gnd vdd FILL
XFILL_4__7712_ gnd vdd FILL
XSFILL38920x39050 gnd vdd FILL
XFILL112440x46050 gnd vdd FILL
XFILL_3__9899_ gnd vdd FILL
XFILL_1__7934_ gnd vdd FILL
XSFILL23720x81050 gnd vdd FILL
X_11350_ _11350_/A _11348_/Y gnd _11354_/C vdd NOR2X1
X_9419_ _9420_/B _9803_/B gnd _9420_/C vdd NAND2X1
XFILL_1__7865_ gnd vdd FILL
X_10301_ _10299_/Y _10318_/A _10301_/C gnd _10349_/D vdd OAI21X1
XFILL_4__7574_ gnd vdd FILL
XSFILL3640x79050 gnd vdd FILL
XFILL_4_BUFX2_insert310 gnd vdd FILL
XFILL_1__9604_ gnd vdd FILL
XFILL_4_BUFX2_insert321 gnd vdd FILL
X_11281_ _11280_/Y _11065_/Y _11278_/Y gnd _11281_/Y vdd AOI21X1
XFILL_4_BUFX2_insert332 gnd vdd FILL
XSFILL3720x7050 gnd vdd FILL
XFILL_4_BUFX2_insert343 gnd vdd FILL
XFILL_4_BUFX2_insert354 gnd vdd FILL
X_13020_ _6893_/A gnd _13020_/Y vdd INVX1
X_10232_ _10232_/A _10280_/B _10232_/C gnd _10232_/Y vdd OAI21X1
XSFILL114600x62050 gnd vdd FILL
XFILL_4_BUFX2_insert365 gnd vdd FILL
XFILL_1__9535_ gnd vdd FILL
XFILL_4_BUFX2_insert376 gnd vdd FILL
XFILL_4_BUFX2_insert387 gnd vdd FILL
XFILL_4__9244_ gnd vdd FILL
XFILL_4_BUFX2_insert398 gnd vdd FILL
X_10163_ _10160_/A _9907_/B gnd _10164_/C vdd NAND2X1
XSFILL69080x43050 gnd vdd FILL
XFILL_1__9466_ gnd vdd FILL
XFILL_2__7210_ gnd vdd FILL
X_10094_ _10094_/Q _7269_/CLK _9061_/R vdd _10094_/D gnd vdd DFFSR
X_14971_ _14971_/A _13420_/C _14030_/C _14969_/Y gnd _14975_/B vdd OAI22X1
XFILL_1__9397_ gnd vdd FILL
XFILL_2__8190_ gnd vdd FILL
XFILL_4__8126_ gnd vdd FILL
X_13922_ _13922_/A gnd _13924_/A vdd INVX1
XFILL_1__8348_ gnd vdd FILL
XFILL_4__8057_ gnd vdd FILL
X_13853_ _8718_/A _13853_/B _13853_/C _6926_/A gnd _13853_/Y vdd AOI22X1
XSFILL23800x61050 gnd vdd FILL
XFILL_2__7072_ gnd vdd FILL
XSFILL89240x56050 gnd vdd FILL
XSFILL18760x7050 gnd vdd FILL
XFILL_6__10900_ gnd vdd FILL
XFILL_5__8870_ gnd vdd FILL
X_12804_ _11879_/B _12669_/CLK _12795_/R vdd _12736_/Y gnd vdd DFFSR
X_13784_ _7388_/Q gnd _13785_/A vdd INVX1
X_10996_ _12207_/Y _12338_/Y gnd _10996_/Y vdd NOR2X1
XFILL_0__10540_ gnd vdd FILL
XFILL_1_BUFX2_insert233 gnd vdd FILL
XFILL_5__7821_ gnd vdd FILL
XFILL_1_BUFX2_insert244 gnd vdd FILL
X_15523_ _15523_/A _15522_/Y gnd _15535_/A vdd NAND2X1
X_12735_ _12723_/A memoryOutData[13] gnd _12736_/C vdd NAND2X1
XFILL_1_BUFX2_insert255 gnd vdd FILL
XFILL_5__12260_ gnd vdd FILL
XFILL_2__11100_ gnd vdd FILL
XFILL_3__10651_ gnd vdd FILL
XFILL_1_BUFX2_insert266 gnd vdd FILL
XFILL_2__12080_ gnd vdd FILL
XFILL_1__11830_ gnd vdd FILL
XFILL_1_BUFX2_insert277 gnd vdd FILL
XFILL_4__12990_ gnd vdd FILL
XSFILL94360x47050 gnd vdd FILL
XFILL_1_BUFX2_insert288 gnd vdd FILL
XFILL_4__8959_ gnd vdd FILL
XFILL_0_BUFX2_insert900 gnd vdd FILL
XSFILL33960x1050 gnd vdd FILL
XFILL_5__7752_ gnd vdd FILL
XFILL_5__11211_ gnd vdd FILL
X_12666_ _12576_/A _12809_/CLK _12799_/R vdd _12666_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert299 gnd vdd FILL
XFILL_0_BUFX2_insert911 gnd vdd FILL
X_15454_ _15454_/A _15454_/B _15441_/Y gnd _15455_/B vdd NAND3X1
XFILL_4__11941_ gnd vdd FILL
XFILL_3__13370_ gnd vdd FILL
XFILL_5__12191_ gnd vdd FILL
XFILL_2__11031_ gnd vdd FILL
XFILL_0_BUFX2_insert922 gnd vdd FILL
XFILL_0__12210_ gnd vdd FILL
XFILL_2__7974_ gnd vdd FILL
XFILL_1__11761_ gnd vdd FILL
XFILL_0_BUFX2_insert933 gnd vdd FILL
X_14405_ _9266_/A gnd _14407_/D vdd INVX1
X_11617_ _11617_/A _11617_/B _11616_/Y gnd _11618_/A vdd OAI21X1
XFILL_0_BUFX2_insert944 gnd vdd FILL
XFILL_0_BUFX2_insert955 gnd vdd FILL
XFILL_5__7683_ gnd vdd FILL
XFILL_3__12321_ gnd vdd FILL
XFILL_5__11142_ gnd vdd FILL
XFILL_0_BUFX2_insert966 gnd vdd FILL
X_15385_ _8718_/A gnd _15386_/D vdd INVX1
X_12597_ _12673_/Q gnd _12597_/Y vdd INVX1
XFILL_4__14660_ gnd vdd FILL
XFILL_1__13500_ gnd vdd FILL
XFILL_4__11872_ gnd vdd FILL
XFILL_2__6925_ gnd vdd FILL
XFILL_1__14480_ gnd vdd FILL
XFILL_5__9422_ gnd vdd FILL
XFILL_0__12141_ gnd vdd FILL
XFILL_0_BUFX2_insert977 gnd vdd FILL
XFILL_0_BUFX2_insert988 gnd vdd FILL
XFILL_1__11692_ gnd vdd FILL
XFILL_4__13611_ gnd vdd FILL
XFILL_0_BUFX2_insert999 gnd vdd FILL
X_14336_ _14336_/A _14830_/B _14051_/C _14335_/Y gnd _14340_/B vdd OAI22X1
X_11548_ _11660_/A _11534_/Y _11547_/Y gnd _11548_/Y vdd NAND3X1
XFILL_3__15040_ gnd vdd FILL
XFILL_5__15950_ gnd vdd FILL
XSFILL104360x32050 gnd vdd FILL
XFILL_3__12252_ gnd vdd FILL
XFILL_5__11073_ gnd vdd FILL
XFILL_4__10823_ gnd vdd FILL
XFILL_4__14591_ gnd vdd FILL
XFILL_2__6856_ gnd vdd FILL
XFILL_1__13431_ gnd vdd FILL
XFILL_2__9644_ gnd vdd FILL
XSFILL34680x28050 gnd vdd FILL
XFILL_0__12072_ gnd vdd FILL
XFILL_2__15770_ gnd vdd FILL
XFILL_2__12982_ gnd vdd FILL
XFILL_1__10643_ gnd vdd FILL
XFILL_5__9353_ gnd vdd FILL
XFILL_4__16330_ gnd vdd FILL
XFILL_5__10024_ gnd vdd FILL
XSFILL74280x14050 gnd vdd FILL
XFILL_5__14901_ gnd vdd FILL
X_14267_ _8167_/Q gnd _14268_/D vdd INVX1
XFILL_3__11203_ gnd vdd FILL
XFILL_4__13542_ gnd vdd FILL
X_11479_ _11466_/Y _11479_/B _11478_/Y gnd _12521_/B vdd NAND3X1
XFILL_5__15881_ gnd vdd FILL
XFILL_0__15900_ gnd vdd FILL
XFILL_2__11933_ gnd vdd FILL
XFILL_4__10754_ gnd vdd FILL
XFILL_2__14721_ gnd vdd FILL
XFILL_3__12183_ gnd vdd FILL
XFILL_0__11023_ gnd vdd FILL
XFILL_1__16150_ gnd vdd FILL
XFILL_1__13362_ gnd vdd FILL
XFILL_1__10574_ gnd vdd FILL
X_13218_ _13218_/A _13231_/B gnd _13251_/B vdd NAND2X1
XFILL_0__7610_ gnd vdd FILL
X_16006_ _16006_/A _16006_/B _14597_/C gnd _12893_/B vdd AOI21X1
XFILL_5__14832_ gnd vdd FILL
XFILL_5__9284_ gnd vdd FILL
XSFILL33400x3050 gnd vdd FILL
XFILL_0__8590_ gnd vdd FILL
XSFILL59080x75050 gnd vdd FILL
X_14198_ _7141_/Q gnd _14198_/Y vdd INVX1
XFILL_3__11134_ gnd vdd FILL
XFILL_1__15101_ gnd vdd FILL
XFILL_4__16261_ gnd vdd FILL
XFILL_2__8526_ gnd vdd FILL
XFILL_4__13473_ gnd vdd FILL
XFILL_1__12313_ gnd vdd FILL
XFILL_4__10685_ gnd vdd FILL
XFILL_0__15831_ gnd vdd FILL
XFILL_2__11864_ gnd vdd FILL
XFILL_2__14652_ gnd vdd FILL
XFILL_1__16081_ gnd vdd FILL
XFILL_1__13293_ gnd vdd FILL
XSFILL99480x80050 gnd vdd FILL
XFILL_5__8235_ gnd vdd FILL
X_13149_ _13149_/A _13149_/B gnd _13150_/C vdd NAND2X1
XFILL_4__15212_ gnd vdd FILL
XFILL_4__12424_ gnd vdd FILL
XSFILL3800x39050 gnd vdd FILL
XFILL_5__14763_ gnd vdd FILL
XFILL_2__10815_ gnd vdd FILL
XFILL_2__13603_ gnd vdd FILL
XFILL_5__11975_ gnd vdd FILL
XFILL_4__16192_ gnd vdd FILL
XFILL_1__15032_ gnd vdd FILL
XFILL_3__15942_ gnd vdd FILL
XFILL_3__11065_ gnd vdd FILL
XFILL_3__7250_ gnd vdd FILL
XFILL_2__14583_ gnd vdd FILL
XFILL_2__8457_ gnd vdd FILL
XFILL_1__12244_ gnd vdd FILL
XFILL_0__15762_ gnd vdd FILL
XFILL_2__11795_ gnd vdd FILL
XFILL_0__12974_ gnd vdd FILL
XFILL_5__13714_ gnd vdd FILL
XFILL_5__10926_ gnd vdd FILL
XFILL_3__10016_ gnd vdd FILL
XFILL_0__7472_ gnd vdd FILL
XFILL_4__15143_ gnd vdd FILL
XFILL_2__16322_ gnd vdd FILL
XFILL_4__12355_ gnd vdd FILL
XFILL_5__14694_ gnd vdd FILL
XSFILL13560x31050 gnd vdd FILL
XSFILL94440x27050 gnd vdd FILL
XFILL_2__13534_ gnd vdd FILL
XFILL_3__7181_ gnd vdd FILL
XFILL_0__14713_ gnd vdd FILL
XFILL_2__8388_ gnd vdd FILL
XFILL_3__15873_ gnd vdd FILL
XFILL_2__10746_ gnd vdd FILL
XFILL_5__7117_ gnd vdd FILL
XFILL_0__11925_ gnd vdd FILL
XFILL_1__12175_ gnd vdd FILL
XFILL_0__9211_ gnd vdd FILL
XFILL_0__15693_ gnd vdd FILL
XFILL_5__8097_ gnd vdd FILL
XFILL_5__13645_ gnd vdd FILL
XFILL_4__11306_ gnd vdd FILL
XSFILL78760x81050 gnd vdd FILL
XFILL_3__14824_ gnd vdd FILL
XFILL_4__15074_ gnd vdd FILL
XFILL_2__7339_ gnd vdd FILL
XFILL_2__13465_ gnd vdd FILL
XFILL_1__11126_ gnd vdd FILL
XFILL_2__16253_ gnd vdd FILL
XFILL_4__12286_ gnd vdd FILL
XFILL_2__10677_ gnd vdd FILL
XFILL_0__14644_ gnd vdd FILL
XFILL_5__7048_ gnd vdd FILL
XFILL_0__9142_ gnd vdd FILL
XFILL_0__11856_ gnd vdd FILL
XFILL_5__16364_ gnd vdd FILL
XFILL_4__14025_ gnd vdd FILL
X_9770_ _9770_/A _9770_/B gnd _9771_/C vdd NAND2X1
XFILL_2__15204_ gnd vdd FILL
XFILL_2__12416_ gnd vdd FILL
XFILL_5__13576_ gnd vdd FILL
XFILL_4__11237_ gnd vdd FILL
XFILL_5__10788_ gnd vdd FILL
XFILL_2__16184_ gnd vdd FILL
X_6982_ _6982_/A _6982_/B _6981_/Y gnd _7024_/D vdd OAI21X1
XFILL_3__14755_ gnd vdd FILL
XFILL_0__10807_ gnd vdd FILL
XFILL_3__11967_ gnd vdd FILL
XFILL_2__13396_ gnd vdd FILL
XFILL_1__15934_ gnd vdd FILL
XFILL_1__11057_ gnd vdd FILL
XFILL_0__14575_ gnd vdd FILL
XFILL_5__15315_ gnd vdd FILL
XSFILL104440x12050 gnd vdd FILL
XFILL_5__12527_ gnd vdd FILL
X_8721_ _8799_/Q gnd _8723_/A vdd INVX1
XFILL_0__11787_ gnd vdd FILL
XFILL_6__14866_ gnd vdd FILL
XFILL_2__9009_ gnd vdd FILL
XFILL_5__16295_ gnd vdd FILL
XFILL_3__13706_ gnd vdd FILL
XFILL_2__15135_ gnd vdd FILL
XFILL_4__11168_ gnd vdd FILL
XFILL_3__10918_ gnd vdd FILL
XFILL_2__12347_ gnd vdd FILL
XFILL_1__10008_ gnd vdd FILL
XFILL_0__16314_ gnd vdd FILL
XSFILL8680x10050 gnd vdd FILL
XFILL_3__14686_ gnd vdd FILL
XFILL_0__13526_ gnd vdd FILL
XFILL_3__11898_ gnd vdd FILL
XFILL_1__15865_ gnd vdd FILL
XFILL_6__13817_ gnd vdd FILL
XFILL_5__15246_ gnd vdd FILL
XFILL_4__10119_ gnd vdd FILL
XFILL_5__8999_ gnd vdd FILL
X_8652_ _8650_/Y _8655_/B _8652_/C gnd _8652_/Y vdd OAI21X1
XFILL_5__12458_ gnd vdd FILL
XFILL_4__15976_ gnd vdd FILL
XFILL_3__13637_ gnd vdd FILL
XSFILL74600x56050 gnd vdd FILL
XFILL_2__15066_ gnd vdd FILL
XFILL_6_BUFX2_insert449 gnd vdd FILL
XFILL_4__11099_ gnd vdd FILL
XFILL_1__14816_ gnd vdd FILL
XFILL_2__12278_ gnd vdd FILL
XFILL_0__16245_ gnd vdd FILL
XSFILL59160x55050 gnd vdd FILL
XFILL_0__13457_ gnd vdd FILL
XFILL_1__15796_ gnd vdd FILL
XSFILL89400x16050 gnd vdd FILL
XFILL_0__10669_ gnd vdd FILL
XFILL_5__11409_ gnd vdd FILL
X_7603_ _7570_/A _9011_/B gnd _7604_/C vdd NAND2X1
XFILL_5__15177_ gnd vdd FILL
XFILL_2__14017_ gnd vdd FILL
XFILL_4__14927_ gnd vdd FILL
XFILL_5__12389_ gnd vdd FILL
XFILL_3__16356_ gnd vdd FILL
X_8583_ _8583_/A _8619_/B _8582_/Y gnd _8583_/Y vdd OAI21X1
XFILL_2__11229_ gnd vdd FILL
XFILL_0__12408_ gnd vdd FILL
XFILL_3__9753_ gnd vdd FILL
XFILL_1__14747_ gnd vdd FILL
XFILL_3__13568_ gnd vdd FILL
XFILL_3__6965_ gnd vdd FILL
XFILL_1__11959_ gnd vdd FILL
XFILL_0__16176_ gnd vdd FILL
XFILL_5__14128_ gnd vdd FILL
XFILL_0__13388_ gnd vdd FILL
XFILL_6__9462_ gnd vdd FILL
X_7534_ _7534_/Q _7534_/CLK _8430_/R vdd _7534_/D gnd vdd DFFSR
XFILL_3__15307_ gnd vdd FILL
XFILL_6__13679_ gnd vdd FILL
XFILL_4_BUFX2_insert1006 gnd vdd FILL
XFILL_3__8704_ gnd vdd FILL
XFILL_4__14858_ gnd vdd FILL
XFILL_0__9975_ gnd vdd FILL
XFILL_3__12519_ gnd vdd FILL
XFILL_4_BUFX2_insert1017 gnd vdd FILL
XFILL_4_BUFX2_insert1028 gnd vdd FILL
XFILL_3__16287_ gnd vdd FILL
XFILL_0__15127_ gnd vdd FILL
XFILL_4_BUFX2_insert1039 gnd vdd FILL
XFILL_3__9684_ gnd vdd FILL
XFILL_3__6896_ gnd vdd FILL
XFILL_0__12339_ gnd vdd FILL
XFILL_1__14678_ gnd vdd FILL
XFILL_3__13499_ gnd vdd FILL
XFILL_4_BUFX2_insert60 gnd vdd FILL
XSFILL13640x11050 gnd vdd FILL
XFILL_4__13809_ gnd vdd FILL
XFILL_5__14059_ gnd vdd FILL
XFILL_4_BUFX2_insert71 gnd vdd FILL
XFILL_3__15238_ gnd vdd FILL
X_7465_ _7527_/Q gnd _7465_/Y vdd INVX1
XFILL_3__8635_ gnd vdd FILL
XFILL_1__13629_ gnd vdd FILL
XFILL_4_BUFX2_insert82 gnd vdd FILL
XFILL_4__14789_ gnd vdd FILL
XFILL_4_BUFX2_insert93 gnd vdd FILL
XFILL_0__15058_ gnd vdd FILL
XFILL_2__15968_ gnd vdd FILL
X_9204_ _9204_/Q _9194_/CLK _9460_/R vdd _9204_/D gnd vdd DFFSR
XSFILL79320x68050 gnd vdd FILL
XFILL_0__8857_ gnd vdd FILL
XFILL_3__15169_ gnd vdd FILL
X_7396_ _7328_/A _7642_/CLK _8676_/R vdd _7396_/D gnd vdd DFFSR
XFILL_0__14009_ gnd vdd FILL
XFILL_1__16348_ gnd vdd FILL
XFILL_2__14919_ gnd vdd FILL
XFILL_3__8566_ gnd vdd FILL
XFILL_2__15899_ gnd vdd FILL
XFILL_0__7808_ gnd vdd FILL
X_9135_ _9193_/Q gnd _9135_/Y vdd INVX1
XFILL_1__7581_ gnd vdd FILL
XFILL_0__8788_ gnd vdd FILL
XFILL_1__16279_ gnd vdd FILL
XFILL_4__7290_ gnd vdd FILL
XFILL_3_BUFX2_insert306 gnd vdd FILL
XFILL_2_BUFX2_insert1010 gnd vdd FILL
XFILL_3__8497_ gnd vdd FILL
XFILL_3_BUFX2_insert317 gnd vdd FILL
XFILL_2_BUFX2_insert1021 gnd vdd FILL
XFILL_0__7739_ gnd vdd FILL
XFILL_3_BUFX2_insert328 gnd vdd FILL
XFILL_2_BUFX2_insert1032 gnd vdd FILL
X_9066_ _9066_/Q _7156_/CLK _7391_/R vdd _9066_/D gnd vdd DFFSR
XSFILL33800x24050 gnd vdd FILL
XFILL_2_BUFX2_insert1043 gnd vdd FILL
XFILL_3_BUFX2_insert339 gnd vdd FILL
XFILL_3__7448_ gnd vdd FILL
XFILL_2_BUFX2_insert1054 gnd vdd FILL
XFILL_1__9251_ gnd vdd FILL
XFILL_2_BUFX2_insert1065 gnd vdd FILL
X_8017_ _8006_/B _9041_/B gnd _8017_/Y vdd NAND2X1
XSFILL28760x2050 gnd vdd FILL
XFILL_2_BUFX2_insert1087 gnd vdd FILL
XFILL_3__7379_ gnd vdd FILL
XFILL_1__8202_ gnd vdd FILL
XFILL_0__9409_ gnd vdd FILL
XFILL_3__9118_ gnd vdd FILL
XFILL111960x34050 gnd vdd FILL
XFILL_1__8133_ gnd vdd FILL
X_9968_ _9924_/A _7268_/CLK _9313_/R vdd _9968_/D gnd vdd DFFSR
XSFILL23720x76050 gnd vdd FILL
XFILL_4__9931_ gnd vdd FILL
X_10850_ _10778_/A _7778_/CLK _8418_/R vdd _10850_/D gnd vdd DFFSR
XFILL_1__8064_ gnd vdd FILL
X_8919_ _8919_/Q _6999_/CLK _7011_/R vdd _8919_/D gnd vdd DFFSR
XSFILL48680x80050 gnd vdd FILL
X_9899_ _9897_/Y _9902_/B _9898_/Y gnd _9959_/D vdd OAI21X1
XSFILL79400x48050 gnd vdd FILL
XFILL_4__9862_ gnd vdd FILL
XFILL_4_CLKBUF1_insert118 gnd vdd FILL
XFILL_0_BUFX2_insert1091 gnd vdd FILL
X_10781_ _15583_/A gnd _10783_/A vdd INVX1
XFILL_4_CLKBUF1_insert129 gnd vdd FILL
X_12520_ _11969_/B gnd _12522_/A vdd INVX1
XFILL_6_BUFX2_insert950 gnd vdd FILL
XFILL_4__9793_ gnd vdd FILL
XSFILL114600x57050 gnd vdd FILL
XFILL_0_BUFX2_insert229 gnd vdd FILL
XFILL_4__8744_ gnd vdd FILL
X_12451_ _12355_/A gnd _12451_/Y vdd INVX1
XSFILL69080x38050 gnd vdd FILL
XFILL_1__8966_ gnd vdd FILL
X_11402_ _11139_/Y gnd _11402_/Y vdd INVX1
X_15170_ _15677_/A _13596_/Y _13632_/Y _15170_/D gnd _15170_/Y vdd OAI22X1
X_12382_ _12382_/A gnd _12382_/Y vdd INVX1
XFILL_2__7690_ gnd vdd FILL
XFILL_4__7626_ gnd vdd FILL
XFILL_1__8897_ gnd vdd FILL
X_14121_ _14121_/A _14120_/Y gnd _14122_/A vdd NOR2X1
X_11333_ _11414_/A gnd _11359_/B vdd INVX2
XFILL_1__7848_ gnd vdd FILL
X_14052_ _9826_/Q gnd _14052_/Y vdd INVX1
XFILL_4__7557_ gnd vdd FILL
X_11264_ _11448_/A _11448_/B gnd _11431_/C vdd NAND2X1
XFILL_2__9360_ gnd vdd FILL
X_13003_ vdd _13003_/B gnd _13004_/C vdd NAND2X1
X_10215_ _10215_/Q _8680_/CLK _8034_/R vdd _10215_/D gnd vdd DFFSR
XFILL_4__7488_ gnd vdd FILL
XFILL_2__8311_ gnd vdd FILL
XFILL_1__9518_ gnd vdd FILL
X_11195_ _11195_/A _11173_/Y _11194_/Y gnd _11196_/C vdd OAI21X1
XFILL_2__9291_ gnd vdd FILL
XFILL_4__9227_ gnd vdd FILL
XFILL_5__8020_ gnd vdd FILL
XFILL_3_BUFX2_insert840 gnd vdd FILL
XFILL_1__10290_ gnd vdd FILL
X_10146_ _10146_/A _10169_/A _10145_/Y gnd _10146_/Y vdd OAI21X1
XFILL_3_BUFX2_insert851 gnd vdd FILL
XFILL_2__8242_ gnd vdd FILL
XFILL_5__11760_ gnd vdd FILL
XFILL_3_BUFX2_insert862 gnd vdd FILL
XFILL_2__11580_ gnd vdd FILL
XFILL_3_BUFX2_insert873 gnd vdd FILL
XFILL_4__9158_ gnd vdd FILL
XFILL_3_BUFX2_insert884 gnd vdd FILL
XFILL_3_BUFX2_insert895 gnd vdd FILL
X_10077_ _9995_/A _7261_/CLK _8669_/R vdd _9997_/Y gnd vdd DFFSR
XFILL_4__12140_ gnd vdd FILL
X_14954_ _16314_/B _14643_/C gnd _14954_/Y vdd NOR2X1
XFILL_2__10531_ gnd vdd FILL
XFILL_5__11691_ gnd vdd FILL
XFILL_3__12870_ gnd vdd FILL
XFILL_4__8109_ gnd vdd FILL
XFILL_0__11710_ gnd vdd FILL
XFILL_4__9089_ gnd vdd FILL
XFILL_5__13430_ gnd vdd FILL
X_13905_ _13905_/A _14697_/B _14752_/C _15429_/C gnd _13906_/A vdd OAI22X1
XSFILL69160x18050 gnd vdd FILL
XFILL_4__12071_ gnd vdd FILL
XFILL_2__7124_ gnd vdd FILL
XFILL_6__12981_ gnd vdd FILL
XFILL_5__10642_ gnd vdd FILL
XFILL_2__13250_ gnd vdd FILL
X_14885_ _14885_/A gnd _14885_/Y vdd INVX1
XFILL_3__11821_ gnd vdd FILL
XFILL_1__13980_ gnd vdd FILL
XFILL_0__11641_ gnd vdd FILL
XSFILL84200x21050 gnd vdd FILL
XFILL_6__11932_ gnd vdd FILL
XFILL_4__11022_ gnd vdd FILL
XFILL_5__13361_ gnd vdd FILL
X_13836_ _13835_/Y _13836_/B _14862_/C _15341_/A gnd _13837_/A vdd OAI22X1
XFILL_2__12201_ gnd vdd FILL
XFILL_5__10573_ gnd vdd FILL
XFILL_2__7055_ gnd vdd FILL
XFILL_3__14540_ gnd vdd FILL
XSFILL104360x27050 gnd vdd FILL
XFILL_3__11752_ gnd vdd FILL
XFILL_5__15100_ gnd vdd FILL
XFILL_2__10393_ gnd vdd FILL
XFILL_0__14360_ gnd vdd FILL
XFILL_5__12312_ gnd vdd FILL
XFILL_5__8853_ gnd vdd FILL
XFILL_0__11572_ gnd vdd FILL
XSFILL69000x82050 gnd vdd FILL
XFILL_4__15830_ gnd vdd FILL
XFILL_6__14651_ gnd vdd FILL
XFILL_5__16080_ gnd vdd FILL
XFILL_5__13292_ gnd vdd FILL
XFILL_3__10703_ gnd vdd FILL
X_10979_ vdd _10979_/B gnd _10980_/C vdd NAND2X1
X_13767_ _7260_/Q gnd _13767_/Y vdd INVX1
XFILL_2__12132_ gnd vdd FILL
XFILL_0__13311_ gnd vdd FILL
XFILL_3__14471_ gnd vdd FILL
XFILL_1__15650_ gnd vdd FILL
XFILL_3__11683_ gnd vdd FILL
XFILL_0__10523_ gnd vdd FILL
XFILL_5__7804_ gnd vdd FILL
XFILL_1__12862_ gnd vdd FILL
XFILL_6__13602_ gnd vdd FILL
X_15506_ _15506_/A _16208_/B _15322_/A _14008_/Y gnd _15507_/C vdd OAI22X1
XFILL_5__15031_ gnd vdd FILL
XFILL_0__14291_ gnd vdd FILL
X_12718_ _12718_/A _12718_/B _12718_/C gnd _12798_/D vdd OAI21X1
XFILL_3__16210_ gnd vdd FILL
XFILL_5__12243_ gnd vdd FILL
XFILL_5__8784_ gnd vdd FILL
XFILL_1__14601_ gnd vdd FILL
XFILL_3__10634_ gnd vdd FILL
XFILL_3__13422_ gnd vdd FILL
XFILL_6__11794_ gnd vdd FILL
XFILL_4__15761_ gnd vdd FILL
XFILL_0__16030_ gnd vdd FILL
XFILL_4__12973_ gnd vdd FILL
XFILL_2__12063_ gnd vdd FILL
X_13698_ _13698_/A _13698_/B _13697_/Y gnd _13698_/Y vdd NAND3X1
XFILL_1__11813_ gnd vdd FILL
XFILL_0__13242_ gnd vdd FILL
XFILL_1__15581_ gnd vdd FILL
XFILL_5__7735_ gnd vdd FILL
XSFILL99480x75050 gnd vdd FILL
XFILL_0_BUFX2_insert730 gnd vdd FILL
XFILL_0_BUFX2_insert741 gnd vdd FILL
XFILL_4__14712_ gnd vdd FILL
X_15437_ _15437_/A _15175_/B _15437_/C gnd _15437_/Y vdd AOI21X1
XFILL_6__10745_ gnd vdd FILL
X_12649_ vdd memoryOutData[27] gnd _12649_/Y vdd NAND2X1
XSFILL74120x73050 gnd vdd FILL
XFILL_4__11924_ gnd vdd FILL
XFILL_5__12174_ gnd vdd FILL
XFILL_2__11014_ gnd vdd FILL
XFILL_3__16141_ gnd vdd FILL
XFILL_3__13353_ gnd vdd FILL
XFILL_0_BUFX2_insert752 gnd vdd FILL
XFILL_4__15692_ gnd vdd FILL
XFILL_1__14532_ gnd vdd FILL
XFILL_3__10565_ gnd vdd FILL
XFILL_0_BUFX2_insert763 gnd vdd FILL
XFILL_2__7957_ gnd vdd FILL
XFILL_1__11744_ gnd vdd FILL
XFILL_0_BUFX2_insert774 gnd vdd FILL
XFILL_0__13173_ gnd vdd FILL
XFILL_0__10385_ gnd vdd FILL
XFILL_6__13464_ gnd vdd FILL
XFILL_0_BUFX2_insert785 gnd vdd FILL
XFILL_5__11125_ gnd vdd FILL
XFILL_6__16252_ gnd vdd FILL
XFILL_0__6972_ gnd vdd FILL
X_15368_ _13799_/Y _15924_/B _16000_/A _13798_/A gnd _15370_/A vdd OAI22X1
XFILL_4__14643_ gnd vdd FILL
XFILL_0__9760_ gnd vdd FILL
XFILL_3__12304_ gnd vdd FILL
XFILL_3__13284_ gnd vdd FILL
XFILL_2__15822_ gnd vdd FILL
XFILL_2__6908_ gnd vdd FILL
XFILL_3__16072_ gnd vdd FILL
XFILL_0_BUFX2_insert796 gnd vdd FILL
XFILL_4__11855_ gnd vdd FILL
XFILL_3__10496_ gnd vdd FILL
XFILL_1__14463_ gnd vdd FILL
XFILL_5__9405_ gnd vdd FILL
XFILL_0__12124_ gnd vdd FILL
XFILL_1__11675_ gnd vdd FILL
XFILL_2__7888_ gnd vdd FILL
X_14319_ _7724_/A gnd _14320_/B vdd INVX1
XFILL_0__8711_ gnd vdd FILL
XFILL_4__10806_ gnd vdd FILL
XFILL_1__16202_ gnd vdd FILL
XFILL_5__15933_ gnd vdd FILL
XFILL_3__15023_ gnd vdd FILL
XFILL_5__7597_ gnd vdd FILL
XFILL_3__12235_ gnd vdd FILL
XFILL_5__11056_ gnd vdd FILL
X_7250_ _7250_/A _7250_/B _7249_/Y gnd _7284_/D vdd OAI21X1
XFILL_4__14574_ gnd vdd FILL
XSFILL109480x60050 gnd vdd FILL
X_15299_ _15677_/A _15299_/B _13743_/Y _15677_/D gnd _15302_/B vdd OAI22X1
XFILL_1__13414_ gnd vdd FILL
XFILL_2__9627_ gnd vdd FILL
XFILL_1__10626_ gnd vdd FILL
XFILL_2__6839_ gnd vdd FILL
XFILL_4__11786_ gnd vdd FILL
XFILL_2__15753_ gnd vdd FILL
XSFILL53400x74050 gnd vdd FILL
XFILL_5__9336_ gnd vdd FILL
XFILL_2__12965_ gnd vdd FILL
XFILL_0__12055_ gnd vdd FILL
XFILL_1__14394_ gnd vdd FILL
XSFILL94280x8050 gnd vdd FILL
XFILL_5__10007_ gnd vdd FILL
XFILL_6__12346_ gnd vdd FILL
XFILL_4__16313_ gnd vdd FILL
XFILL_0__8642_ gnd vdd FILL
XFILL_4__13525_ gnd vdd FILL
X_7181_ _7181_/A _7181_/B _7180_/Y gnd _7261_/D vdd OAI21X1
XFILL_2__14704_ gnd vdd FILL
XFILL_3__12166_ gnd vdd FILL
XFILL_5__15864_ gnd vdd FILL
XFILL_1__16133_ gnd vdd FILL
XFILL_1__13345_ gnd vdd FILL
XFILL_2__11916_ gnd vdd FILL
XSFILL54040x40050 gnd vdd FILL
XFILL_3__8351_ gnd vdd FILL
XFILL_0__11006_ gnd vdd FILL
XFILL_2__15684_ gnd vdd FILL
XFILL_2__12896_ gnd vdd FILL
XFILL_1__10557_ gnd vdd FILL
XFILL_5__9267_ gnd vdd FILL
XFILL_4__16244_ gnd vdd FILL
XFILL_5__14815_ gnd vdd FILL
XFILL_3__11117_ gnd vdd FILL
XFILL_0__8573_ gnd vdd FILL
XFILL_2__8509_ gnd vdd FILL
XFILL_4__13456_ gnd vdd FILL
XFILL_5__15795_ gnd vdd FILL
XFILL_3__7302_ gnd vdd FILL
XFILL_2__14635_ gnd vdd FILL
XFILL_3__12097_ gnd vdd FILL
XFILL_4__10668_ gnd vdd FILL
XFILL_0__15814_ gnd vdd FILL
XFILL_1__16064_ gnd vdd FILL
XFILL_2__11847_ gnd vdd FILL
XFILL_1__13276_ gnd vdd FILL
XFILL_5__8218_ gnd vdd FILL
XFILL_2__9489_ gnd vdd FILL
XFILL_1__10488_ gnd vdd FILL
XFILL_4__12407_ gnd vdd FILL
XFILL_5__14746_ gnd vdd FILL
XSFILL43880x83050 gnd vdd FILL
XFILL_3__15925_ gnd vdd FILL
XFILL_4__16175_ gnd vdd FILL
XFILL_5__11958_ gnd vdd FILL
XFILL_1__15015_ gnd vdd FILL
XFILL_3__11048_ gnd vdd FILL
XFILL_3__7233_ gnd vdd FILL
XFILL_4__13387_ gnd vdd FILL
XFILL_1__12227_ gnd vdd FILL
XFILL_2__14566_ gnd vdd FILL
XSFILL58680x43050 gnd vdd FILL
XFILL_2__11778_ gnd vdd FILL
XFILL_0__15745_ gnd vdd FILL
XFILL_5__8149_ gnd vdd FILL
XFILL_0__12957_ gnd vdd FILL
XFILL_5__10909_ gnd vdd FILL
XFILL_1_BUFX2_insert8 gnd vdd FILL
XFILL_0__7455_ gnd vdd FILL
XFILL_6__11159_ gnd vdd FILL
XFILL_4__15126_ gnd vdd FILL
XFILL_2__16305_ gnd vdd FILL
XFILL_4__12338_ gnd vdd FILL
XFILL_5__14677_ gnd vdd FILL
XFILL_5__11889_ gnd vdd FILL
XFILL_3__15856_ gnd vdd FILL
XFILL_3__7164_ gnd vdd FILL
XFILL_2__13517_ gnd vdd FILL
XFILL_2__14497_ gnd vdd FILL
XFILL_0__11908_ gnd vdd FILL
XFILL_1__12158_ gnd vdd FILL
XSFILL49400x27050 gnd vdd FILL
XFILL_0__15676_ gnd vdd FILL
XSFILL74200x53050 gnd vdd FILL
X_9822_ _9742_/A _7790_/CLK _9566_/R vdd _9822_/D gnd vdd DFFSR
XFILL_5__13628_ gnd vdd FILL
XFILL_0__12888_ gnd vdd FILL
XFILL111880x49050 gnd vdd FILL
XFILL_5__16416_ gnd vdd FILL
XFILL_3__14807_ gnd vdd FILL
XFILL_4__15057_ gnd vdd FILL
XFILL_2__16236_ gnd vdd FILL
XFILL_2__13448_ gnd vdd FILL
XFILL_4__12269_ gnd vdd FILL
XFILL_1__11109_ gnd vdd FILL
XFILL_3__7095_ gnd vdd FILL
XFILL_0__14627_ gnd vdd FILL
XFILL_3__15787_ gnd vdd FILL
XFILL_0__9125_ gnd vdd FILL
XFILL_1__12089_ gnd vdd FILL
XFILL_3__12999_ gnd vdd FILL
XFILL_0__11839_ gnd vdd FILL
XFILL_4__14008_ gnd vdd FILL
XFILL_5__16347_ gnd vdd FILL
XFILL_6__8893_ gnd vdd FILL
X_9753_ _9751_/Y _9741_/B _9753_/C gnd _9825_/D vdd OAI21X1
XFILL_5__13559_ gnd vdd FILL
X_6965_ _7019_/Q gnd _6967_/A vdd INVX1
XFILL_3__14738_ gnd vdd FILL
XFILL_1__15917_ gnd vdd FILL
XFILL_2__16167_ gnd vdd FILL
XFILL_2__13379_ gnd vdd FILL
XFILL_0__14558_ gnd vdd FILL
XSFILL8680x9050 gnd vdd FILL
X_8704_ _8740_/A _9344_/B gnd _8705_/C vdd NAND2X1
XFILL_6__7844_ gnd vdd FILL
XFILL_5__16278_ gnd vdd FILL
XSFILL64680x62050 gnd vdd FILL
X_9684_ _9675_/A _9556_/B gnd _9685_/C vdd NAND2X1
XFILL_2__15118_ gnd vdd FILL
XFILL_2__16098_ gnd vdd FILL
X_6896_ _6896_/A gnd memoryWriteData[26] vdd BUFX2
XFILL_3__14669_ gnd vdd FILL
XFILL_0__13509_ gnd vdd FILL
XSFILL38840x72050 gnd vdd FILL
XFILL_1__15848_ gnd vdd FILL
XFILL_0__8007_ gnd vdd FILL
XFILL_0__14489_ gnd vdd FILL
XFILL_5__15229_ gnd vdd FILL
X_8635_ _8685_/Q gnd _8637_/A vdd INVX1
XFILL_3__16408_ gnd vdd FILL
XSFILL54120x20050 gnd vdd FILL
XFILL_3__9805_ gnd vdd FILL
XFILL_0__16228_ gnd vdd FILL
XFILL_2__15049_ gnd vdd FILL
XFILL_4__15959_ gnd vdd FILL
XFILL_5_BUFX2_insert902 gnd vdd FILL
XFILL_3__7997_ gnd vdd FILL
XFILL_1__15779_ gnd vdd FILL
XFILL_5_BUFX2_insert913 gnd vdd FILL
XFILL_3__16339_ gnd vdd FILL
X_8566_ _8662_/Q gnd _8568_/A vdd INVX1
XFILL_5_BUFX2_insert924 gnd vdd FILL
XSFILL33800x19050 gnd vdd FILL
XFILL_5_BUFX2_insert935 gnd vdd FILL
XFILL_3__9736_ gnd vdd FILL
XFILL_3__6948_ gnd vdd FILL
XFILL_5_BUFX2_insert946 gnd vdd FILL
XFILL_0__16159_ gnd vdd FILL
XSFILL43960x63050 gnd vdd FILL
XFILL_5_BUFX2_insert957 gnd vdd FILL
X_7517_ _7435_/A _7261_/CLK _8669_/R vdd _7517_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert968 gnd vdd FILL
XFILL_1__8751_ gnd vdd FILL
XFILL_5_BUFX2_insert979 gnd vdd FILL
X_8497_ _8495_/Y _8496_/A _8497_/C gnd _8553_/D vdd OAI21X1
XFILL_4__8460_ gnd vdd FILL
XFILL_3__9667_ gnd vdd FILL
XFILL_3__6879_ gnd vdd FILL
XFILL_0__8909_ gnd vdd FILL
XFILL_1__7702_ gnd vdd FILL
X_7448_ _7457_/A _8088_/B gnd _7448_/Y vdd NAND2X1
XSFILL44040x72050 gnd vdd FILL
XFILL_0__9889_ gnd vdd FILL
XFILL_3__8618_ gnd vdd FILL
XFILL_3__9598_ gnd vdd FILL
XFILL_4__8391_ gnd vdd FILL
XSFILL64920x4050 gnd vdd FILL
XFILL_1__7633_ gnd vdd FILL
X_7379_ _7413_/Q gnd _7381_/A vdd INVX1
XFILL_4__7342_ gnd vdd FILL
XFILL_3_BUFX2_insert103 gnd vdd FILL
X_9118_ _9086_/B _9374_/B gnd _9119_/C vdd NAND2X1
XFILL_1__7564_ gnd vdd FILL
XFILL112040x38050 gnd vdd FILL
X_10000_ _9998_/Y _9975_/B _9999_/Y gnd _10000_/Y vdd OAI21X1
X_9049_ _8959_/A _8921_/CLK _9049_/R vdd _8961_/Y gnd vdd DFFSR
XFILL_1__7495_ gnd vdd FILL
XFILL_4__9012_ gnd vdd FILL
XCLKBUF1_insert1081 clk gnd CLKBUF1_insert218/A vdd CLKBUF1
XSFILL79800x64050 gnd vdd FILL
XFILL_1__9234_ gnd vdd FILL
XFILL_2_BUFX2_insert803 gnd vdd FILL
XFILL_2_BUFX2_insert814 gnd vdd FILL
XFILL_2_BUFX2_insert825 gnd vdd FILL
XFILL_2_BUFX2_insert836 gnd vdd FILL
XSFILL39000x61050 gnd vdd FILL
XFILL_2_BUFX2_insert847 gnd vdd FILL
XFILL_1__9165_ gnd vdd FILL
X_11951_ _11909_/A _12406_/A gnd _11952_/C vdd NAND2X1
XFILL_2_BUFX2_insert858 gnd vdd FILL
XFILL_2_BUFX2_insert869 gnd vdd FILL
X_10902_ _10984_/Q gnd _10903_/B vdd INVX1
XFILL_1__8116_ gnd vdd FILL
X_11882_ _11874_/B _11882_/B gnd _11882_/Y vdd NAND2X1
X_14670_ _9025_/A gnd _16048_/A vdd INVX1
XFILL_0_BUFX2_insert80 gnd vdd FILL
XFILL_0_BUFX2_insert91 gnd vdd FILL
XFILL_1__9096_ gnd vdd FILL
XFILL_4__9914_ gnd vdd FILL
XSFILL94280x80050 gnd vdd FILL
X_13621_ _10239_/A _13621_/B _14867_/C _9945_/Q gnd _13621_/Y vdd AOI22X1
X_10833_ _10822_/B _9041_/B gnd _10833_/Y vdd NAND2X1
X_16340_ gnd gnd gnd _16341_/C vdd NAND2X1
X_10764_ _10831_/B _9100_/B gnd _10765_/C vdd NAND2X1
XBUFX2_insert802 _15091_/Y gnd _16166_/A vdd BUFX2
X_13552_ _13552_/A gnd _15163_/B vdd INVX1
XBUFX2_insert813 _13329_/Y gnd _9005_/A vdd BUFX2
XFILL_2__8860_ gnd vdd FILL
XBUFX2_insert824 _13287_/Y gnd _7470_/B vdd BUFX2
XBUFX2_insert835 _13324_/Y gnd _8589_/B vdd BUFX2
X_12503_ vdd _12503_/B gnd _12503_/Y vdd NAND2X1
XFILL_4__9776_ gnd vdd FILL
XFILL112120x18050 gnd vdd FILL
XFILL_4__6988_ gnd vdd FILL
XBUFX2_insert846 _12375_/Y gnd _8853_/B vdd BUFX2
X_13483_ _13482_/Y _13483_/B gnd _13489_/C vdd NOR2X1
X_16271_ _16270_/Y _15527_/A _14999_/A _16269_/Y gnd _16271_/Y vdd OAI22X1
XFILL_2__7811_ gnd vdd FILL
XBUFX2_insert857 _13314_/Y gnd _8187_/B vdd BUFX2
X_10695_ _10737_/Q gnd _10697_/A vdd INVX1
XBUFX2_insert868 _13379_/Y gnd _14626_/A vdd BUFX2
XFILL_4__8727_ gnd vdd FILL
XBUFX2_insert879 _15019_/Y gnd _15761_/D vdd BUFX2
XFILL_1__9998_ gnd vdd FILL
X_12434_ _12407_/A _12693_/Q gnd _12435_/C vdd NAND2X1
X_15222_ _15197_/B gnd _16096_/C vdd INVX4
XFILL_2__7742_ gnd vdd FILL
XFILL_0__10170_ gnd vdd FILL
XFILL_5__7451_ gnd vdd FILL
XFILL_4__8658_ gnd vdd FILL
X_12365_ _12407_/A _12588_/A gnd _12366_/C vdd NAND2X1
X_15153_ _13568_/C gnd _15153_/Y vdd INVX1
XFILL_4__11640_ gnd vdd FILL
XFILL_3__10281_ gnd vdd FILL
XFILL_4__7609_ gnd vdd FILL
XFILL_2__7673_ gnd vdd FILL
XFILL_1__11460_ gnd vdd FILL
X_11316_ _11313_/Y _11437_/C gnd _11317_/C vdd AND2X2
X_14104_ _14104_/A _14934_/B _14317_/C _15595_/A gnd _14105_/A vdd OAI22X1
XFILL_4__8589_ gnd vdd FILL
XFILL_3__12020_ gnd vdd FILL
X_15084_ _9977_/A _15696_/A gnd _15084_/Y vdd NAND2X1
XFILL_2__9412_ gnd vdd FILL
X_12296_ _12216_/B _12297_/D _12300_/C gnd _12298_/B vdd NAND3X1
XFILL_2__12750_ gnd vdd FILL
XFILL_1__10411_ gnd vdd FILL
XFILL_4__11571_ gnd vdd FILL
XFILL_5__9121_ gnd vdd FILL
X_14035_ _9954_/Q _13751_/C _14035_/C gnd _14035_/Y vdd AOI21X1
XFILL_1__11391_ gnd vdd FILL
XFILL_6__12131_ gnd vdd FILL
XFILL_4__13310_ gnd vdd FILL
XSFILL84200x16050 gnd vdd FILL
X_11247_ _11245_/Y _11247_/B gnd _11247_/Y vdd NAND2X1
XFILL_4__10522_ gnd vdd FILL
XFILL_5__12861_ gnd vdd FILL
XFILL_2__11701_ gnd vdd FILL
XFILL_2__9343_ gnd vdd FILL
XFILL_1__13130_ gnd vdd FILL
XFILL_4__14290_ gnd vdd FILL
XSFILL94360x60050 gnd vdd FILL
XFILL_0__13860_ gnd vdd FILL
XFILL_5__14600_ gnd vdd FILL
XFILL_5__11812_ gnd vdd FILL
XFILL_4__13241_ gnd vdd FILL
X_11178_ _11494_/A gnd _11492_/B vdd INVX2
XFILL_5__15580_ gnd vdd FILL
XFILL_4__10453_ gnd vdd FILL
XFILL_2__14420_ gnd vdd FILL
XFILL_2__11632_ gnd vdd FILL
XFILL_2__9274_ gnd vdd FILL
XFILL_5__8003_ gnd vdd FILL
XFILL_3__13971_ gnd vdd FILL
XFILL_1__10273_ gnd vdd FILL
XFILL_3_BUFX2_insert670 gnd vdd FILL
XFILL_0__13791_ gnd vdd FILL
XFILL_5__14531_ gnd vdd FILL
X_10129_ _13892_/A gnd _10129_/Y vdd INVX1
XFILL_3__15710_ gnd vdd FILL
XFILL_3_BUFX2_insert681 gnd vdd FILL
XFILL_5__11743_ gnd vdd FILL
XFILL_4__10384_ gnd vdd FILL
X_15986_ _15986_/A _15197_/B _15197_/C _14589_/Y gnd _15988_/A vdd OAI22X1
XFILL_2__8225_ gnd vdd FILL
XFILL_1__12012_ gnd vdd FILL
XFILL_4__13172_ gnd vdd FILL
XFILL_2__14351_ gnd vdd FILL
XFILL_3_BUFX2_insert692 gnd vdd FILL
XFILL_0__15530_ gnd vdd FILL
XFILL_2__11563_ gnd vdd FILL
XFILL_0__12742_ gnd vdd FILL
XFILL_0__7240_ gnd vdd FILL
XFILL_2__13302_ gnd vdd FILL
XFILL_5__14462_ gnd vdd FILL
X_14937_ _14937_/A _13843_/C _14815_/C _14937_/D gnd _14938_/B vdd OAI22X1
XSFILL99400x4050 gnd vdd FILL
XFILL_4__12123_ gnd vdd FILL
XSFILL74120x68050 gnd vdd FILL
XFILL_3__15641_ gnd vdd FILL
XFILL_5__11674_ gnd vdd FILL
XFILL_2__10514_ gnd vdd FILL
XFILL_3__12853_ gnd vdd FILL
XFILL_2__14282_ gnd vdd FILL
XSFILL89720x47050 gnd vdd FILL
XFILL_2__11494_ gnd vdd FILL
XFILL_0__15461_ gnd vdd FILL
XFILL_5__16201_ gnd vdd FILL
XFILL_5__13413_ gnd vdd FILL
XFILL_5__10625_ gnd vdd FILL
XFILL_0__7171_ gnd vdd FILL
XFILL_2__7107_ gnd vdd FILL
XFILL_2__13233_ gnd vdd FILL
X_14868_ _14868_/A _10739_/Q _9203_/Q _14868_/D gnd _14869_/B vdd AOI22X1
XFILL_2__16021_ gnd vdd FILL
XFILL_4__12054_ gnd vdd FILL
XFILL_5__14393_ gnd vdd FILL
XFILL_3__11804_ gnd vdd FILL
XFILL_2__10445_ gnd vdd FILL
XFILL_2__8087_ gnd vdd FILL
XFILL_3__15572_ gnd vdd FILL
XFILL_0__14412_ gnd vdd FILL
XFILL_3__12784_ gnd vdd FILL
XFILL_5__8905_ gnd vdd FILL
XFILL_0__11624_ gnd vdd FILL
XFILL_1__13963_ gnd vdd FILL
XFILL_0__15392_ gnd vdd FILL
XFILL_5__16132_ gnd vdd FILL
XFILL_5__13344_ gnd vdd FILL
X_13819_ _7133_/Q gnd _13821_/D vdd INVX1
XFILL_5__9885_ gnd vdd FILL
XFILL_4__11005_ gnd vdd FILL
XFILL_5__10556_ gnd vdd FILL
XFILL_3__14523_ gnd vdd FILL
XFILL_2__7038_ gnd vdd FILL
XFILL_1__15702_ gnd vdd FILL
X_14799_ _14567_/D _16194_/B _14797_/Y _13846_/A gnd _14799_/Y vdd OAI22X1
XFILL_2__13164_ gnd vdd FILL
XFILL_1__12914_ gnd vdd FILL
XSFILL59720x5050 gnd vdd FILL
XFILL_3__11735_ gnd vdd FILL
XFILL_2__10376_ gnd vdd FILL
XSFILL109480x55050 gnd vdd FILL
XFILL_0__14343_ gnd vdd FILL
XFILL_5__8836_ gnd vdd FILL
XFILL_1__13894_ gnd vdd FILL
XFILL_0__11555_ gnd vdd FILL
XSFILL13800x8050 gnd vdd FILL
XFILL_5__16063_ gnd vdd FILL
XFILL_5__13275_ gnd vdd FILL
XFILL_2__12115_ gnd vdd FILL
XFILL_4__15813_ gnd vdd FILL
XFILL_3__14454_ gnd vdd FILL
XFILL_5__10487_ gnd vdd FILL
XFILL_1__12845_ gnd vdd FILL
XFILL_0__10506_ gnd vdd FILL
XFILL_1__15633_ gnd vdd FILL
XFILL_2__13095_ gnd vdd FILL
XSFILL54040x35050 gnd vdd FILL
XFILL_3__7851_ gnd vdd FILL
XFILL_3__11666_ gnd vdd FILL
XFILL_5__15014_ gnd vdd FILL
XFILL_0__14274_ gnd vdd FILL
XFILL_5__8767_ gnd vdd FILL
X_8420_ _8420_/Q _9306_/CLK _9306_/R vdd _8354_/Y gnd vdd DFFSR
XFILL_6__7560_ gnd vdd FILL
XFILL_5__12226_ gnd vdd FILL
XFILL_0__11486_ gnd vdd FILL
XFILL_3__13405_ gnd vdd FILL
XFILL_4__15744_ gnd vdd FILL
XFILL_0__16013_ gnd vdd FILL
XFILL_2__12046_ gnd vdd FILL
XFILL_3__10617_ gnd vdd FILL
XFILL_4__12956_ gnd vdd FILL
XFILL_0__13225_ gnd vdd FILL
XFILL_1__15564_ gnd vdd FILL
XFILL_3__14385_ gnd vdd FILL
XFILL_3__11597_ gnd vdd FILL
XFILL_1__12776_ gnd vdd FILL
XFILL_5__7718_ gnd vdd FILL
XFILL_0__10437_ gnd vdd FILL
XFILL_6__16304_ gnd vdd FILL
XFILL_2__8989_ gnd vdd FILL
XFILL_0_BUFX2_insert560 gnd vdd FILL
XFILL_0__9812_ gnd vdd FILL
XFILL_4__11907_ gnd vdd FILL
XFILL_5__12157_ gnd vdd FILL
XFILL_3__16124_ gnd vdd FILL
XFILL_0_BUFX2_insert571 gnd vdd FILL
X_8351_ _8349_/Y _8315_/B _8351_/C gnd _8351_/Y vdd OAI21X1
XFILL_5__8698_ gnd vdd FILL
XFILL_0_BUFX2_insert582 gnd vdd FILL
XFILL_3__13336_ gnd vdd FILL
XSFILL43880x78050 gnd vdd FILL
XFILL_4__15675_ gnd vdd FILL
XFILL_3__9521_ gnd vdd FILL
XFILL_4__12887_ gnd vdd FILL
XFILL_1__14515_ gnd vdd FILL
XFILL_0_BUFX2_insert593 gnd vdd FILL
XFILL_1__11727_ gnd vdd FILL
XFILL_3__10548_ gnd vdd FILL
XFILL_0__13156_ gnd vdd FILL
XFILL_1__15495_ gnd vdd FILL
XFILL_0__10368_ gnd vdd FILL
XFILL_4_BUFX2_insert909 gnd vdd FILL
XSFILL109320x6050 gnd vdd FILL
XFILL_5__11108_ gnd vdd FILL
X_7302_ _7369_/B _7558_/B gnd _7302_/Y vdd NAND2X1
XFILL_0__9743_ gnd vdd FILL
XFILL_4__14626_ gnd vdd FILL
X_8282_ _8282_/Q _7389_/CLK _8285_/R vdd _8282_/D gnd vdd DFFSR
XFILL_5__12088_ gnd vdd FILL
XFILL_2__15805_ gnd vdd FILL
XFILL_3__16055_ gnd vdd FILL
XFILL_0__6955_ gnd vdd FILL
XFILL_4__11838_ gnd vdd FILL
XFILL_3__13267_ gnd vdd FILL
XSFILL18680x54050 gnd vdd FILL
XFILL_0__12107_ gnd vdd FILL
XSFILL48920x15050 gnd vdd FILL
XFILL_1__14446_ gnd vdd FILL
XFILL_1__11658_ gnd vdd FILL
XFILL_0__10299_ gnd vdd FILL
XSFILL74200x48050 gnd vdd FILL
XFILL_0__13087_ gnd vdd FILL
XFILL_2__13997_ gnd vdd FILL
XFILL_5__15916_ gnd vdd FILL
XFILL_3__15006_ gnd vdd FILL
X_7233_ _7279_/Q gnd _7233_/Y vdd INVX1
XFILL_5__11039_ gnd vdd FILL
XFILL_4__14557_ gnd vdd FILL
XFILL_0__9674_ gnd vdd FILL
XFILL_0__6886_ gnd vdd FILL
XFILL_3__12218_ gnd vdd FILL
XFILL_3__8403_ gnd vdd FILL
XFILL_4__11769_ gnd vdd FILL
XFILL_2__15736_ gnd vdd FILL
XFILL_3__9383_ gnd vdd FILL
XFILL_0__12038_ gnd vdd FILL
XFILL_1__14377_ gnd vdd FILL
XFILL_1__11589_ gnd vdd FILL
XFILL_6__15117_ gnd vdd FILL
XFILL_0__8625_ gnd vdd FILL
XFILL_4__13508_ gnd vdd FILL
XFILL_5__15847_ gnd vdd FILL
X_7164_ _7256_/Q gnd _7164_/Y vdd INVX1
XFILL_1__13328_ gnd vdd FILL
XFILL_3__8334_ gnd vdd FILL
XFILL_4__14488_ gnd vdd FILL
XFILL_1__16116_ gnd vdd FILL
XFILL_3__12149_ gnd vdd FILL
XFILL_2__15667_ gnd vdd FILL
XFILL_2__12879_ gnd vdd FILL
XFILL_4__16227_ gnd vdd FILL
XFILL_4__13439_ gnd vdd FILL
X_7095_ _7095_/A _7095_/B _7094_/Y gnd _7147_/D vdd OAI21X1
XFILL_2__14618_ gnd vdd FILL
XFILL_5__15778_ gnd vdd FILL
XFILL_1__16047_ gnd vdd FILL
XFILL_1__13259_ gnd vdd FILL
XFILL_3__8265_ gnd vdd FILL
XFILL_2__15598_ gnd vdd FILL
XFILL112360x74050 gnd vdd FILL
XFILL_0__13989_ gnd vdd FILL
XFILL_0__7507_ gnd vdd FILL
XFILL_0__8487_ gnd vdd FILL
XFILL_3__15908_ gnd vdd FILL
XFILL_5__14729_ gnd vdd FILL
XSFILL54120x15050 gnd vdd FILL
XFILL_4__16158_ gnd vdd FILL
XFILL_3__7216_ gnd vdd FILL
XFILL_3__8196_ gnd vdd FILL
XFILL_2__14549_ gnd vdd FILL
XFILL_0__15728_ gnd vdd FILL
XFILL_0__7438_ gnd vdd FILL
XFILL_4__15109_ gnd vdd FILL
XFILL_6__9994_ gnd vdd FILL
XFILL_4__16089_ gnd vdd FILL
XFILL_3__15839_ gnd vdd FILL
XFILL_0__15659_ gnd vdd FILL
XSFILL43960x58050 gnd vdd FILL
X_9805_ _9843_/Q gnd _9805_/Y vdd INVX1
XFILL_0__7369_ gnd vdd FILL
XFILL_2__16219_ gnd vdd FILL
XFILL_3__7078_ gnd vdd FILL
X_7997_ _7995_/Y _7997_/B _7997_/C gnd _8045_/D vdd OAI21X1
XFILL_4__7960_ gnd vdd FILL
XFILL_0__9108_ gnd vdd FILL
XSFILL18760x34050 gnd vdd FILL
X_6948_ _6948_/A _7972_/B gnd _6949_/C vdd NAND2X1
X_9736_ _9820_/Q gnd _9738_/A vdd INVX1
XSFILL8600x44050 gnd vdd FILL
XFILL_4__6911_ gnd vdd FILL
XSFILL44040x67050 gnd vdd FILL
XFILL_0__9039_ gnd vdd FILL
XSFILL59640x46050 gnd vdd FILL
XFILL_4__7891_ gnd vdd FILL
XSFILL48840x6050 gnd vdd FILL
XBUFX2_insert109 _10925_/Y gnd _11969_/A vdd BUFX2
XFILL_1__9921_ gnd vdd FILL
X_9667_ _9665_/Y _9597_/A _9666_/Y gnd _9711_/D vdd OAI21X1
X_6879_ _6879_/A gnd memoryWriteData[9] vdd BUFX2
XFILL_4__9630_ gnd vdd FILL
XFILL_4__6842_ gnd vdd FILL
X_8618_ _8619_/B _9770_/B gnd _8618_/Y vdd NAND2X1
XFILL_5_BUFX2_insert710 gnd vdd FILL
XFILL_1__9852_ gnd vdd FILL
XSFILL23880x25050 gnd vdd FILL
XFILL_5_BUFX2_insert721 gnd vdd FILL
X_9598_ _9596_/Y _9597_/A _9598_/C gnd _9598_/Y vdd OAI21X1
XFILL_5_BUFX2_insert732 gnd vdd FILL
X_10480_ _16105_/A _7268_/CLK _8688_/R vdd _10438_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert743 gnd vdd FILL
XFILL_6__7689_ gnd vdd FILL
X_8549_ _8549_/Q _8165_/CLK _8165_/R vdd _8549_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert754 gnd vdd FILL
XFILL_1__9783_ gnd vdd FILL
XFILL_4__8512_ gnd vdd FILL
XFILL_5_BUFX2_insert765 gnd vdd FILL
XFILL_3__9719_ gnd vdd FILL
XSFILL38920x47050 gnd vdd FILL
XFILL_5_BUFX2_insert776 gnd vdd FILL
XFILL112440x54050 gnd vdd FILL
XFILL_1__6995_ gnd vdd FILL
XFILL_4__9492_ gnd vdd FILL
XFILL_5_BUFX2_insert787 gnd vdd FILL
XFILL_5_BUFX2_insert798 gnd vdd FILL
XFILL_1__8734_ gnd vdd FILL
XFILL_4__8443_ gnd vdd FILL
X_12150_ _12150_/A _12150_/B _12150_/C gnd _12150_/Y vdd OAI21X1
XFILL_6__9359_ gnd vdd FILL
X_11101_ _11290_/A _11544_/A gnd _11542_/A vdd NOR2X1
XFILL_4__8374_ gnd vdd FILL
X_12081_ _12081_/A _12073_/B _12073_/C gnd gnd _12081_/Y vdd AOI22X1
XFILL_1__7616_ gnd vdd FILL
XFILL_1__8596_ gnd vdd FILL
XFILL_4__7325_ gnd vdd FILL
X_11032_ _12129_/Y gnd _11032_/Y vdd INVX1
XSFILL94280x75050 gnd vdd FILL
XSFILL114600x70050 gnd vdd FILL
XFILL_1__7547_ gnd vdd FILL
XSFILL29480x65050 gnd vdd FILL
XSFILL84520x52050 gnd vdd FILL
X_15840_ _15833_/Y _15840_/B gnd _15851_/A vdd NAND2X1
XSFILL69880x70050 gnd vdd FILL
XSFILL69080x51050 gnd vdd FILL
XSFILL99320x12050 gnd vdd FILL
XFILL_1__7478_ gnd vdd FILL
XFILL_2_BUFX2_insert600 gnd vdd FILL
XFILL_2_BUFX2_insert611 gnd vdd FILL
XFILL_2_BUFX2_insert622 gnd vdd FILL
XFILL_4__7187_ gnd vdd FILL
XFILL_2__8010_ gnd vdd FILL
XFILL_1__9217_ gnd vdd FILL
XFILL_2_BUFX2_insert633 gnd vdd FILL
X_15771_ _8808_/Q _15821_/B _15978_/C _8492_/A gnd _15777_/A vdd AOI22X1
XFILL_2_BUFX2_insert644 gnd vdd FILL
X_12983_ _12983_/A vdd _12983_/C gnd _13057_/D vdd OAI21X1
XSFILL73560x76050 gnd vdd FILL
XFILL_2_BUFX2_insert655 gnd vdd FILL
XFILL_2_BUFX2_insert666 gnd vdd FILL
XSFILL23800x3050 gnd vdd FILL
X_14722_ _14721_/Y _14722_/B gnd _14730_/B vdd NOR2X1
X_11934_ _11934_/A _11934_/B _11933_/Y gnd _6853_/A vdd OAI21X1
XFILL_2_BUFX2_insert677 gnd vdd FILL
XFILL_1__9148_ gnd vdd FILL
XFILL_2_BUFX2_insert688 gnd vdd FILL
XFILL_2_BUFX2_insert699 gnd vdd FILL
XFILL_5__6951_ gnd vdd FILL
XFILL_5__10410_ gnd vdd FILL
X_14653_ _14651_/Y _14441_/B _14377_/B _16069_/C gnd _14653_/Y vdd OAI22X1
XFILL_1__9079_ gnd vdd FILL
XFILL_2__10230_ gnd vdd FILL
X_11865_ _11865_/A _11865_/B _11858_/Y gnd _11865_/Y vdd NAND3X1
XFILL_5__11390_ gnd vdd FILL
XSFILL89240x64050 gnd vdd FILL
XFILL_1__10960_ gnd vdd FILL
XFILL_5_BUFX2_insert15 gnd vdd FILL
XFILL_5_BUFX2_insert26 gnd vdd FILL
X_13604_ _13603_/Y _13857_/B gnd _13605_/C vdd NOR2X1
XFILL_5__9670_ gnd vdd FILL
X_10816_ _10814_/Y _10789_/B _10816_/C gnd _10862_/D vdd OAI21X1
XFILL_5__6882_ gnd vdd FILL
X_14584_ _14584_/A gnd _15997_/C vdd INVX1
XFILL_5_BUFX2_insert37 gnd vdd FILL
XFILL_3__11520_ gnd vdd FILL
X_11796_ _11795_/Y _11034_/B gnd _11796_/Y vdd AND2X2
XFILL_2__8912_ gnd vdd FILL
XFILL_5_BUFX2_insert48 gnd vdd FILL
XFILL_2__10161_ gnd vdd FILL
XFILL_2__9892_ gnd vdd FILL
XFILL_5_BUFX2_insert59 gnd vdd FILL
XBUFX2_insert610 _15035_/Y gnd _15187_/A vdd BUFX2
XFILL_5__8621_ gnd vdd FILL
XFILL_0__11340_ gnd vdd FILL
X_16323_ _16321_/Y gnd _16323_/C gnd _16323_/Y vdd OAI21X1
XFILL_1__10891_ gnd vdd FILL
XBUFX2_insert621 _13430_/Y gnd _13434_/B vdd BUFX2
XBUFX2_insert632 _12354_/Y gnd _8576_/B vdd BUFX2
X_13535_ _8152_/Q gnd _13536_/D vdd INVX1
XFILL_5__10272_ gnd vdd FILL
XBUFX2_insert643 _13424_/Y gnd _13775_/B vdd BUFX2
XFILL_3__11451_ gnd vdd FILL
X_10747_ _10745_/Y _10809_/A _10747_/C gnd _10839_/D vdd OAI21X1
XFILL_1__12630_ gnd vdd FILL
XFILL_4__13790_ gnd vdd FILL
XFILL_2__8843_ gnd vdd FILL
XBUFX2_insert654 _12429_/Y gnd _8011_/B vdd BUFX2
XSFILL94360x55050 gnd vdd FILL
XFILL_5__12011_ gnd vdd FILL
XFILL_4__9759_ gnd vdd FILL
XFILL_0__11271_ gnd vdd FILL
XBUFX2_insert665 _11364_/Y gnd _11732_/B vdd BUFX2
X_16254_ _15841_/C _14923_/D _16254_/C _15813_/C gnd _16257_/B vdd OAI22X1
XBUFX2_insert676 _13541_/Y gnd _14403_/C vdd BUFX2
X_10678_ _10678_/A _9782_/B gnd _10679_/C vdd NAND2X1
XFILL_4__12741_ gnd vdd FILL
X_13466_ _13423_/A _13398_/A _13465_/C gnd _13467_/A vdd NAND3X1
XBUFX2_insert687 _13459_/Y gnd _14849_/B vdd BUFX2
XFILL_3__10402_ gnd vdd FILL
XFILL_3__14170_ gnd vdd FILL
XSFILL84600x32050 gnd vdd FILL
XFILL_0__13010_ gnd vdd FILL
XBUFX2_insert698 _12420_/Y gnd _7490_/B vdd BUFX2
XFILL_2__13920_ gnd vdd FILL
XFILL_3__11382_ gnd vdd FILL
XFILL_5__7503_ gnd vdd FILL
XFILL_2__8774_ gnd vdd FILL
XFILL_6__13301_ gnd vdd FILL
X_15205_ _15203_/Y _15205_/B gnd _15206_/B vdd NOR2X1
XSFILL69160x31050 gnd vdd FILL
X_12417_ _12415_/Y _12380_/A _12417_/C gnd _12417_/Y vdd OAI21X1
XFILL_5__8483_ gnd vdd FILL
X_16185_ _9418_/A _15202_/B _15071_/C gnd _16186_/C vdd NAND3X1
XFILL_3__13121_ gnd vdd FILL
XFILL_1__14300_ gnd vdd FILL
XFILL_4__15460_ gnd vdd FILL
XSFILL103720x74050 gnd vdd FILL
X_13397_ _13423_/A _13423_/B _13718_/B gnd _13587_/C vdd NAND3X1
XFILL_2__7725_ gnd vdd FILL
XFILL_1__11512_ gnd vdd FILL
XFILL_2__13851_ gnd vdd FILL
XFILL_0__10153_ gnd vdd FILL
XFILL_1__15280_ gnd vdd FILL
XFILL_5__7434_ gnd vdd FILL
XFILL_1__12492_ gnd vdd FILL
XFILL_6__10444_ gnd vdd FILL
XSFILL7960x72050 gnd vdd FILL
XFILL_4__14411_ gnd vdd FILL
X_15136_ _15136_/A _15130_/Y _15136_/C gnd _15144_/B vdd NAND3X1
X_12348_ _12346_/Y _12395_/A _12348_/C gnd _12348_/Y vdd OAI21X1
XFILL_4__11623_ gnd vdd FILL
XFILL_5__13962_ gnd vdd FILL
XFILL_4__15391_ gnd vdd FILL
XFILL_1__14231_ gnd vdd FILL
XFILL_3__10264_ gnd vdd FILL
XFILL_1__11443_ gnd vdd FILL
XFILL_2__13782_ gnd vdd FILL
XFILL_0__14961_ gnd vdd FILL
XFILL_2__10994_ gnd vdd FILL
XFILL_5__15701_ gnd vdd FILL
XFILL_5__7365_ gnd vdd FILL
XSFILL74280x22050 gnd vdd FILL
X_15067_ _15067_/A _15067_/B _15062_/Y gnd _15075_/A vdd NOR3X1
XFILL_3__12003_ gnd vdd FILL
XFILL_4__14342_ gnd vdd FILL
XFILL_5__12913_ gnd vdd FILL
X_12279_ _12239_/A gnd _12239_/C gnd _12279_/Y vdd NAND3X1
XFILL_2__15521_ gnd vdd FILL
XFILL_5__13893_ gnd vdd FILL
XFILL_4__11554_ gnd vdd FILL
XFILL_2__12733_ gnd vdd FILL
XFILL_5__9104_ gnd vdd FILL
XFILL_1__14162_ gnd vdd FILL
XFILL_3__10195_ gnd vdd FILL
XFILL_0__13912_ gnd vdd FILL
XFILL_2__7587_ gnd vdd FILL
XFILL_1__11374_ gnd vdd FILL
X_14018_ _13836_/B _14018_/B _14872_/C _14018_/D gnd _14018_/Y vdd OAI22X1
XFILL_0__14892_ gnd vdd FILL
XSFILL59080x83050 gnd vdd FILL
XFILL_5__7296_ gnd vdd FILL
XFILL_5__12844_ gnd vdd FILL
XFILL_4__10505_ gnd vdd FILL
XFILL_5__15632_ gnd vdd FILL
XSFILL89320x44050 gnd vdd FILL
XFILL_0__9390_ gnd vdd FILL
XFILL_1__13113_ gnd vdd FILL
XFILL_4__14273_ gnd vdd FILL
XFILL_2__15452_ gnd vdd FILL
XFILL_4__11485_ gnd vdd FILL
XFILL_1__10325_ gnd vdd FILL
XFILL_0__13843_ gnd vdd FILL
XFILL_5__9035_ gnd vdd FILL
XFILL_1__14093_ gnd vdd FILL
XFILL_4__16012_ gnd vdd FILL
XFILL_0__8341_ gnd vdd FILL
XFILL_4__13224_ gnd vdd FILL
XSFILL3800x47050 gnd vdd FILL
XFILL_5__12775_ gnd vdd FILL
XFILL_4__10436_ gnd vdd FILL
XFILL_5__15563_ gnd vdd FILL
XFILL_2__14403_ gnd vdd FILL
XFILL_1__13044_ gnd vdd FILL
XFILL_2__9257_ gnd vdd FILL
XFILL_3__13954_ gnd vdd FILL
XFILL_2__11615_ gnd vdd FILL
XFILL_1__10256_ gnd vdd FILL
XFILL_2__15383_ gnd vdd FILL
XFILL_2__12595_ gnd vdd FILL
XFILL_0__13774_ gnd vdd FILL
XFILL_5__14514_ gnd vdd FILL
X_7920_ _7876_/A _7664_/CLK _7920_/R vdd _7878_/Y gnd vdd DFFSR
XFILL_5__11726_ gnd vdd FILL
XFILL_0__8272_ gnd vdd FILL
XFILL_2__8208_ gnd vdd FILL
X_15969_ _8813_/Q _15821_/B _15969_/C _7739_/A gnd _15969_/Y vdd AOI22X1
XFILL_4__13155_ gnd vdd FILL
XSFILL94440x35050 gnd vdd FILL
XFILL_5__15494_ gnd vdd FILL
XFILL_3__12905_ gnd vdd FILL
XFILL_4__10367_ gnd vdd FILL
XFILL_0__15513_ gnd vdd FILL
XFILL_2__14334_ gnd vdd FILL
XFILL_2__11546_ gnd vdd FILL
XFILL_0__12725_ gnd vdd FILL
XFILL_3__13885_ gnd vdd FILL
XSFILL58840x1050 gnd vdd FILL
XFILL_0__7223_ gnd vdd FILL
XFILL_1__10187_ gnd vdd FILL
XFILL_4__12106_ gnd vdd FILL
XFILL_5__14445_ gnd vdd FILL
XFILL_6__6991_ gnd vdd FILL
XFILL_3__15624_ gnd vdd FILL
X_7851_ _7851_/A _7800_/B _7850_/Y gnd _7851_/Y vdd OAI21X1
XFILL_5__11657_ gnd vdd FILL
XFILL_3__12836_ gnd vdd FILL
XFILL_4__13086_ gnd vdd FILL
XFILL_6__13996_ gnd vdd FILL
XFILL_2__8139_ gnd vdd FILL
XSFILL69240x11050 gnd vdd FILL
XFILL_2__14265_ gnd vdd FILL
XFILL_4__10298_ gnd vdd FILL
XFILL_2__11477_ gnd vdd FILL
XFILL_0__15444_ gnd vdd FILL
XFILL_0__12656_ gnd vdd FILL
XFILL_5__9937_ gnd vdd FILL
XFILL_1__14995_ gnd vdd FILL
XFILL_2__16004_ gnd vdd FILL
XFILL_4__12037_ gnd vdd FILL
XFILL_5__14376_ gnd vdd FILL
X_7782_ _7782_/Q _8921_/CLK _9049_/R vdd _7720_/Y gnd vdd DFFSR
XFILL_2__10428_ gnd vdd FILL
XFILL_2__13216_ gnd vdd FILL
XFILL_3__15555_ gnd vdd FILL
XFILL_5__11588_ gnd vdd FILL
XFILL_3__12767_ gnd vdd FILL
XFILL_2__14196_ gnd vdd FILL
XSFILL18680x49050 gnd vdd FILL
XFILL_0__11607_ gnd vdd FILL
XFILL_3__8952_ gnd vdd FILL
XFILL_0__15375_ gnd vdd FILL
XFILL_1__13946_ gnd vdd FILL
XSFILL104440x20050 gnd vdd FILL
XFILL_5__13327_ gnd vdd FILL
XFILL_0__12587_ gnd vdd FILL
XFILL_5__9868_ gnd vdd FILL
XFILL_5__16115_ gnd vdd FILL
X_9521_ _9519_/Y _9529_/A _9521_/C gnd _9577_/D vdd OAI21X1
XFILL_5__10539_ gnd vdd FILL
XFILL_3__14506_ gnd vdd FILL
XFILL_0__7085_ gnd vdd FILL
XFILL_2__13147_ gnd vdd FILL
XFILL_3__11718_ gnd vdd FILL
XFILL_2__10359_ gnd vdd FILL
XFILL_0__14326_ gnd vdd FILL
XFILL_3__15486_ gnd vdd FILL
XFILL_3__12698_ gnd vdd FILL
XFILL_3__8883_ gnd vdd FILL
XFILL_0__11538_ gnd vdd FILL
XFILL_1__13877_ gnd vdd FILL
XFILL_5__16046_ gnd vdd FILL
XSFILL99160x47050 gnd vdd FILL
XFILL_5__13258_ gnd vdd FILL
X_9452_ _9400_/A _7020_/CLK _9964_/R vdd _9452_/D gnd vdd DFFSR
XFILL_5__9799_ gnd vdd FILL
XFILL_3__14437_ gnd vdd FILL
XFILL_1__15616_ gnd vdd FILL
XFILL_3__7834_ gnd vdd FILL
XFILL_4__13988_ gnd vdd FILL
XFILL_3__11649_ gnd vdd FILL
XFILL_0__14257_ gnd vdd FILL
XSFILL59160x63050 gnd vdd FILL
XFILL_1__12828_ gnd vdd FILL
XFILL_5__12209_ gnd vdd FILL
X_8403_ _8437_/Q gnd _8403_/Y vdd INVX1
XFILL_0__11469_ gnd vdd FILL
X_9383_ _9359_/A _9383_/B gnd _9384_/C vdd NAND2X1
XFILL_4__15727_ gnd vdd FILL
XFILL_2__12029_ gnd vdd FILL
XFILL_0__13208_ gnd vdd FILL
XFILL_3__14368_ gnd vdd FILL
XFILL_1__12759_ gnd vdd FILL
XFILL_1__15547_ gnd vdd FILL
XFILL_3__7765_ gnd vdd FILL
XFILL111880x62050 gnd vdd FILL
XFILL_0__14188_ gnd vdd FILL
XFILL_0_BUFX2_insert390 gnd vdd FILL
X_8334_ _8414_/Q gnd _8334_/Y vdd INVX1
XFILL_3__16107_ gnd vdd FILL
XFILL_3__13319_ gnd vdd FILL
XFILL112360x69050 gnd vdd FILL
XFILL_4__15658_ gnd vdd FILL
XFILL_3__9504_ gnd vdd FILL
XFILL_4_BUFX2_insert706 gnd vdd FILL
XFILL_4_BUFX2_insert717 gnd vdd FILL
XFILL_0__7987_ gnd vdd FILL
XFILL_0__13139_ gnd vdd FILL
XFILL_4_BUFX2_insert728 gnd vdd FILL
XFILL_3__14299_ gnd vdd FILL
XFILL_3__7696_ gnd vdd FILL
XFILL_1__15478_ gnd vdd FILL
XFILL_4__14609_ gnd vdd FILL
XFILL_4_BUFX2_insert739 gnd vdd FILL
XFILL_0__9726_ gnd vdd FILL
XFILL_3__16038_ gnd vdd FILL
XFILL_0__6938_ gnd vdd FILL
X_8265_ _8263_/Y _8187_/B _8265_/C gnd _8305_/D vdd OAI21X1
XFILL_4__15589_ gnd vdd FILL
XFILL_1__14429_ gnd vdd FILL
XSFILL79320x76050 gnd vdd FILL
X_7216_ _7202_/B _6960_/B gnd _7216_/Y vdd NAND2X1
XFILL_1__8450_ gnd vdd FILL
XFILL_0__9657_ gnd vdd FILL
XSFILL95080x1050 gnd vdd FILL
X_8196_ _8196_/A _8246_/A _8196_/C gnd _8282_/D vdd OAI21X1
XFILL_2__15719_ gnd vdd FILL
XFILL_0__6869_ gnd vdd FILL
XFILL_3__9366_ gnd vdd FILL
XFILL_0__8608_ gnd vdd FILL
XFILL_1__8381_ gnd vdd FILL
X_7147_ _7093_/A _7147_/CLK _7531_/R vdd _7147_/D gnd vdd DFFSR
XSFILL18760x29050 gnd vdd FILL
XFILL_4__7110_ gnd vdd FILL
XSFILL8600x39050 gnd vdd FILL
XFILL_3__8317_ gnd vdd FILL
XFILL_4__8090_ gnd vdd FILL
XFILL_3__9297_ gnd vdd FILL
XFILL_1__7332_ gnd vdd FILL
XSFILL33800x32050 gnd vdd FILL
XFILL_4__7041_ gnd vdd FILL
X_7078_ _7142_/Q gnd _7078_/Y vdd INVX1
XFILL_3__8248_ gnd vdd FILL
XFILL_5_BUFX2_insert1091 gnd vdd FILL
XFILL_1__9002_ gnd vdd FILL
XFILL_1__7194_ gnd vdd FILL
XFILL_1_BUFX2_insert607 gnd vdd FILL
XFILL111960x42050 gnd vdd FILL
XFILL112440x49050 gnd vdd FILL
XFILL_1_BUFX2_insert618 gnd vdd FILL
XFILL_4__8992_ gnd vdd FILL
XFILL_1_BUFX2_insert629 gnd vdd FILL
XFILL_4__7943_ gnd vdd FILL
X_11650_ _11259_/Y gnd _11650_/Y vdd INVX1
XFILL112040x51050 gnd vdd FILL
X_9719_ _8567_/A _9737_/A gnd _9720_/C vdd NAND2X1
X_10601_ _15837_/A _7664_/CLK _7649_/R vdd _10545_/Y gnd vdd DFFSR
XFILL_4__7874_ gnd vdd FILL
XFILL_1__9904_ gnd vdd FILL
X_11581_ _11623_/A _11623_/B _11402_/Y gnd _11626_/C vdd OAI21X1
XFILL_4__9613_ gnd vdd FILL
X_13320_ _13297_/C _13320_/B gnd _13320_/Y vdd NOR2X1
X_10532_ _10511_/A _8356_/B gnd _10533_/C vdd NAND2X1
XSFILL4280x48050 gnd vdd FILL
XFILL_5_BUFX2_insert540 gnd vdd FILL
XFILL_5_BUFX2_insert551 gnd vdd FILL
XFILL_4__9544_ gnd vdd FILL
XFILL_5_BUFX2_insert562 gnd vdd FILL
X_13251_ _13311_/A _13251_/B _13289_/B gnd _13252_/A vdd AOI21X1
XFILL_5_BUFX2_insert573 gnd vdd FILL
X_10463_ _15437_/A _8815_/CLK _8047_/R vdd _10463_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert584 gnd vdd FILL
XSFILL69080x46050 gnd vdd FILL
XFILL_1__9766_ gnd vdd FILL
XFILL_5_BUFX2_insert595 gnd vdd FILL
XFILL_1__6978_ gnd vdd FILL
XFILL_4__9475_ gnd vdd FILL
X_12202_ _11974_/A gnd _12204_/A vdd INVX1
X_13182_ _13182_/Q _12538_/CLK _12689_/R vdd _13182_/D gnd vdd DFFSR
XFILL_1__8717_ gnd vdd FILL
X_10394_ _15547_/A gnd _10396_/A vdd INVX1
XFILL_2__8490_ gnd vdd FILL
X_12133_ _13097_/A gnd _12135_/A vdd INVX1
XFILL_2__7441_ gnd vdd FILL
XFILL_1__8648_ gnd vdd FILL
XFILL_4__8357_ gnd vdd FILL
XFILL_2_CLKBUF1_insert121 gnd vdd FILL
X_12064_ _12012_/A _12808_/Q _11996_/C gnd _12066_/B vdd NAND3X1
XFILL_2_CLKBUF1_insert132 gnd vdd FILL
XFILL_6__10160_ gnd vdd FILL
XSFILL23800x64050 gnd vdd FILL
XFILL_2_CLKBUF1_insert143 gnd vdd FILL
XFILL_2__7372_ gnd vdd FILL
XFILL_5__10890_ gnd vdd FILL
XFILL_4__7308_ gnd vdd FILL
XFILL_1__8579_ gnd vdd FILL
XSFILL89240x59050 gnd vdd FILL
XFILL_2_CLKBUF1_insert154 gnd vdd FILL
XFILL112120x31050 gnd vdd FILL
XFILL_2_CLKBUF1_insert165 gnd vdd FILL
XFILL_5__7081_ gnd vdd FILL
X_11015_ _11015_/A _11013_/Y _11003_/Y _11015_/D gnd _11015_/Y vdd AOI22X1
XFILL_2_CLKBUF1_insert176 gnd vdd FILL
XFILL_2_CLKBUF1_insert187 gnd vdd FILL
XFILL_2__9111_ gnd vdd FILL
XFILL_2_CLKBUF1_insert198 gnd vdd FILL
XFILL_1__10110_ gnd vdd FILL
XFILL_4__11270_ gnd vdd FILL
XFILL_1__11090_ gnd vdd FILL
XFILL_4__7239_ gnd vdd FILL
X_15823_ _15390_/B _9833_/Q _9577_/Q _15652_/A gnd _15824_/B vdd AOI22X1
XFILL_2__11400_ gnd vdd FILL
XFILL_2__9042_ gnd vdd FILL
XFILL_2_BUFX2_insert430 gnd vdd FILL
XFILL_3__10951_ gnd vdd FILL
XFILL_2__12380_ gnd vdd FILL
XFILL_1__10041_ gnd vdd FILL
XFILL_2_BUFX2_insert441 gnd vdd FILL
XFILL_0__10771_ gnd vdd FILL
XFILL_5__11511_ gnd vdd FILL
XFILL_2_BUFX2_insert452 gnd vdd FILL
XFILL_2_BUFX2_insert463 gnd vdd FILL
XBUFX2_insert9 _13280_/Y gnd _7354_/B vdd BUFX2
X_15754_ _15802_/A _14279_/Y _14268_/D _15774_/C gnd _15757_/B vdd OAI22X1
XFILL_4__10152_ gnd vdd FILL
XFILL_5__12491_ gnd vdd FILL
XFILL_2__11331_ gnd vdd FILL
X_12966_ _6875_/A gnd _12968_/A vdd INVX1
XFILL_2_BUFX2_insert474 gnd vdd FILL
XFILL_3__13670_ gnd vdd FILL
XFILL_0__12510_ gnd vdd FILL
XFILL_2_BUFX2_insert485 gnd vdd FILL
XFILL_3__10882_ gnd vdd FILL
XFILL_2_BUFX2_insert496 gnd vdd FILL
XFILL_5__14230_ gnd vdd FILL
XFILL_0__13490_ gnd vdd FILL
X_14705_ _13868_/B _16117_/D _14705_/C _14496_/A gnd _14705_/Y vdd OAI22X1
XSFILL69160x26050 gnd vdd FILL
X_11917_ _13185_/Q gnd _11919_/A vdd INVX1
XFILL_5__7983_ gnd vdd FILL
XFILL_5__11442_ gnd vdd FILL
XFILL_3__12621_ gnd vdd FILL
X_15685_ _8421_/Q gnd _15686_/A vdd INVX1
XFILL_6__13781_ gnd vdd FILL
XFILL_2__14050_ gnd vdd FILL
XFILL_4__14960_ gnd vdd FILL
XFILL_1__13800_ gnd vdd FILL
X_12897_ _12895_/Y vdd _12897_/C gnd _12943_/D vdd OAI21X1
XFILL_2__11262_ gnd vdd FILL
XFILL_0__12441_ gnd vdd FILL
XSFILL29160x42050 gnd vdd FILL
XFILL_1__14780_ gnd vdd FILL
XFILL_5__9722_ gnd vdd FILL
XFILL_1__11992_ gnd vdd FILL
XFILL_5__6934_ gnd vdd FILL
X_14636_ _13876_/B _14635_/Y _14636_/C _14634_/Y gnd _14636_/Y vdd OAI22X1
XFILL_5__14161_ gnd vdd FILL
XFILL_2__13001_ gnd vdd FILL
XFILL_4__13911_ gnd vdd FILL
XFILL_3__15340_ gnd vdd FILL
X_11848_ _11848_/A _11427_/A _11223_/B _11848_/D gnd _11848_/Y vdd AOI22X1
XFILL_5__11373_ gnd vdd FILL
XSFILL104360x35050 gnd vdd FILL
XFILL_4__14891_ gnd vdd FILL
XFILL_1__10943_ gnd vdd FILL
XFILL_1__13731_ gnd vdd FILL
XFILL_0__15160_ gnd vdd FILL
XFILL_2__11193_ gnd vdd FILL
XFILL_5__9653_ gnd vdd FILL
XFILL_0__12372_ gnd vdd FILL
XFILL_5__13112_ gnd vdd FILL
XSFILL33640x67050 gnd vdd FILL
XFILL_5__6865_ gnd vdd FILL
XSFILL74280x17050 gnd vdd FILL
XFILL_5__10324_ gnd vdd FILL
XFILL_4__13842_ gnd vdd FILL
X_14567_ _14567_/A _14567_/B _14566_/Y _14567_/D gnd _14567_/Y vdd OAI22X1
XFILL_5__14092_ gnd vdd FILL
XFILL_3__11503_ gnd vdd FILL
XFILL_2__10144_ gnd vdd FILL
XFILL_0__14111_ gnd vdd FILL
XFILL_3__15271_ gnd vdd FILL
X_11779_ _11766_/Y _11484_/B _11349_/B _11020_/Y gnd _11779_/Y vdd OAI22X1
XFILL_1__16450_ gnd vdd FILL
XFILL_1__13662_ gnd vdd FILL
XFILL_3__12483_ gnd vdd FILL
XFILL_5__8604_ gnd vdd FILL
XFILL_2__9875_ gnd vdd FILL
XFILL_0__11323_ gnd vdd FILL
XBUFX2_insert440 _15086_/Y gnd _15225_/A vdd BUFX2
XBUFX2_insert451 _13276_/Y gnd _7168_/A vdd BUFX2
XFILL_1__10874_ gnd vdd FILL
X_16306_ _16306_/A _16306_/B _16306_/C _14932_/Y gnd _16306_/Y vdd OAI22X1
XFILL_0__15091_ gnd vdd FILL
XBUFX2_insert462 _15044_/Y gnd _15632_/A vdd BUFX2
X_13518_ _13514_/Y _13518_/B gnd _13518_/Y vdd NOR2X1
XFILL_5__13043_ gnd vdd FILL
XFILL_3__14222_ gnd vdd FILL
XFILL_5__10255_ gnd vdd FILL
XBUFX2_insert473 _15041_/Y gnd _15550_/C vdd BUFX2
XSFILL59080x78050 gnd vdd FILL
XFILL_4__13773_ gnd vdd FILL
XFILL_1__15401_ gnd vdd FILL
X_14498_ _14498_/A _14490_/Y gnd _14499_/A vdd NAND2X1
XFILL_1__12613_ gnd vdd FILL
XFILL_0__8890_ gnd vdd FILL
XFILL_2__8826_ gnd vdd FILL
XFILL_3__11434_ gnd vdd FILL
XFILL112200x11050 gnd vdd FILL
XFILL_0__14042_ gnd vdd FILL
XFILL_2__14952_ gnd vdd FILL
XBUFX2_insert484 _12372_/Y gnd _9362_/B vdd BUFX2
XSFILL99480x83050 gnd vdd FILL
XFILL_1__13593_ gnd vdd FILL
XFILL_1__16381_ gnd vdd FILL
XBUFX2_insert495 BUFX2_insert520/A gnd _8937_/R vdd BUFX2
XFILL_0__11254_ gnd vdd FILL
X_16237_ _9459_/Q _15202_/B _15995_/C gnd _16237_/Y vdd NAND3X1
XFILL_4__15512_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1077 gnd vdd FILL
XSFILL74120x81050 gnd vdd FILL
XFILL_4__12724_ gnd vdd FILL
XFILL_0__7841_ gnd vdd FILL
X_13449_ _13449_/A _14200_/C _14555_/C _13445_/Y gnd _13449_/Y vdd OAI22X1
XFILL_5__10186_ gnd vdd FILL
XFILL_3__14153_ gnd vdd FILL
XFILL_2__13903_ gnd vdd FILL
XFILL_2__8757_ gnd vdd FILL
XFILL_1__15332_ gnd vdd FILL
XFILL_3__7550_ gnd vdd FILL
XFILL_3__11365_ gnd vdd FILL
XFILL_2__14883_ gnd vdd FILL
XFILL_0__11185_ gnd vdd FILL
XFILL_5__8466_ gnd vdd FILL
XFILL_3__13104_ gnd vdd FILL
X_16168_ _15681_/C _16168_/B _15322_/D _14830_/A gnd _16171_/A vdd OAI22X1
XFILL_4__15443_ gnd vdd FILL
XFILL_4__12655_ gnd vdd FILL
XFILL_3__10316_ gnd vdd FILL
XFILL_2__7708_ gnd vdd FILL
XFILL_2__13834_ gnd vdd FILL
XFILL_5__14994_ gnd vdd FILL
XFILL_3__11296_ gnd vdd FILL
XFILL_1__15263_ gnd vdd FILL
XFILL_3__14084_ gnd vdd FILL
XFILL_0__10136_ gnd vdd FILL
XFILL_3__7481_ gnd vdd FILL
XFILL_1__12475_ gnd vdd FILL
XFILL_5__7417_ gnd vdd FILL
XFILL_0__9511_ gnd vdd FILL
X_15119_ _15119_/A _15118_/Y gnd _15119_/Y vdd NOR2X1
XFILL_5__8397_ gnd vdd FILL
XFILL_0__15993_ gnd vdd FILL
X_8050_ _8050_/Q _7411_/CLK _7411_/R vdd _8012_/Y gnd vdd DFFSR
XFILL_4__11606_ gnd vdd FILL
XFILL_4__15374_ gnd vdd FILL
XFILL_1__14214_ gnd vdd FILL
XFILL_3__9220_ gnd vdd FILL
XFILL_3__13035_ gnd vdd FILL
X_16099_ _16099_/A _16099_/B _16099_/C _14725_/B gnd _16100_/A vdd OAI22X1
XFILL_3__10247_ gnd vdd FILL
XFILL_5__13945_ gnd vdd FILL
XFILL_4__12586_ gnd vdd FILL
XFILL_1__11426_ gnd vdd FILL
XFILL_1__15194_ gnd vdd FILL
XFILL_2__13765_ gnd vdd FILL
X_7001_ _6911_/A _8921_/CLK _9049_/R vdd _6913_/Y gnd vdd DFFSR
XFILL_2__10977_ gnd vdd FILL
XFILL_6__13146_ gnd vdd FILL
XFILL_0__10067_ gnd vdd FILL
XFILL_0__14944_ gnd vdd FILL
XFILL_5__7348_ gnd vdd FILL
XFILL_4__14325_ gnd vdd FILL
XFILL_2__15504_ gnd vdd FILL
XFILL_1_BUFX2_insert13 gnd vdd FILL
XFILL_4__11537_ gnd vdd FILL
XFILL_3__9151_ gnd vdd FILL
XFILL_2__12716_ gnd vdd FILL
XFILL_5__13876_ gnd vdd FILL
XFILL_1__14145_ gnd vdd FILL
XFILL_3__10178_ gnd vdd FILL
XFILL_1_BUFX2_insert24 gnd vdd FILL
XFILL_1__11357_ gnd vdd FILL
XFILL_1_BUFX2_insert35 gnd vdd FILL
XFILL_0__14875_ gnd vdd FILL
XFILL_2__13696_ gnd vdd FILL
XSFILL104440x15050 gnd vdd FILL
XFILL_1_BUFX2_insert46 gnd vdd FILL
XFILL_5__15615_ gnd vdd FILL
XFILL_1_BUFX2_insert57 gnd vdd FILL
XFILL_3__8102_ gnd vdd FILL
XFILL_4__14256_ gnd vdd FILL
XFILL_6__10289_ gnd vdd FILL
XFILL_0__9373_ gnd vdd FILL
XFILL_5__12827_ gnd vdd FILL
XFILL_1__10308_ gnd vdd FILL
XFILL_1_BUFX2_insert68 gnd vdd FILL
XFILL_2__15435_ gnd vdd FILL
XSFILL8680x13050 gnd vdd FILL
XFILL_4__11468_ gnd vdd FILL
XFILL_2__12647_ gnd vdd FILL
XFILL_0__13826_ gnd vdd FILL
XFILL_1_BUFX2_insert79 gnd vdd FILL
XSFILL33720x47050 gnd vdd FILL
XFILL_3__14986_ gnd vdd FILL
XFILL_5__9018_ gnd vdd FILL
XFILL_1__14076_ gnd vdd FILL
XFILL_3__9082_ gnd vdd FILL
XFILL_1__11288_ gnd vdd FILL
XFILL_4__13207_ gnd vdd FILL
XFILL_0__8324_ gnd vdd FILL
XFILL_5__12758_ gnd vdd FILL
XFILL_5__15546_ gnd vdd FILL
XFILL_4__10419_ gnd vdd FILL
XFILL_4__14187_ gnd vdd FILL
XFILL_1__13027_ gnd vdd FILL
X_8952_ _8952_/A _8996_/A _8952_/C gnd _9046_/D vdd OAI21X1
XFILL_3__13937_ gnd vdd FILL
XFILL_1__10239_ gnd vdd FILL
XFILL_2__15366_ gnd vdd FILL
XFILL_4__11399_ gnd vdd FILL
XFILL_2__12578_ gnd vdd FILL
XSFILL59160x58050 gnd vdd FILL
XFILL_0__13757_ gnd vdd FILL
XFILL_0__10969_ gnd vdd FILL
XFILL_0__8255_ gnd vdd FILL
XFILL_4__13138_ gnd vdd FILL
XFILL_5__11709_ gnd vdd FILL
X_7903_ _7903_/Q _9194_/CLK _9460_/R vdd _7903_/D gnd vdd DFFSR
XFILL_2__14317_ gnd vdd FILL
X_8883_ _8854_/B _9011_/B gnd _8883_/Y vdd NAND2X1
XFILL_5__15477_ gnd vdd FILL
XFILL_0__12708_ gnd vdd FILL
XFILL_3__13868_ gnd vdd FILL
XFILL_2__11529_ gnd vdd FILL
XSFILL74200x61050 gnd vdd FILL
XFILL_2__15297_ gnd vdd FILL
XFILL_6__9762_ gnd vdd FILL
XFILL_0__7206_ gnd vdd FILL
XFILL_0__13688_ gnd vdd FILL
X_7834_ _7906_/Q gnd _7836_/A vdd INVX1
XFILL_3__15607_ gnd vdd FILL
XFILL_0__8186_ gnd vdd FILL
XFILL_5__14428_ gnd vdd FILL
XFILL_2__14248_ gnd vdd FILL
XFILL_0__15427_ gnd vdd FILL
XFILL_3__13799_ gnd vdd FILL
XFILL_3__9984_ gnd vdd FILL
XFILL_0__12639_ gnd vdd FILL
XFILL_6__8713_ gnd vdd FILL
XFILL_1__14978_ gnd vdd FILL
XSFILL13640x14050 gnd vdd FILL
XFILL_5__14359_ gnd vdd FILL
XFILL_3__15538_ gnd vdd FILL
X_7765_ _7763_/Y _7672_/B _7764_/Y gnd _7797_/D vdd OAI21X1
XFILL_0__15358_ gnd vdd FILL
XFILL_2__14179_ gnd vdd FILL
XFILL_1__13929_ gnd vdd FILL
X_9504_ _9572_/Q gnd _9506_/A vdd INVX1
XFILL_6__15649_ gnd vdd FILL
XFILL_0__7068_ gnd vdd FILL
XFILL_1__7950_ gnd vdd FILL
X_7696_ _7694_/Y _7744_/B _7696_/C gnd _7774_/D vdd OAI21X1
XFILL_0__14309_ gnd vdd FILL
XFILL_3__15469_ gnd vdd FILL
XSFILL38840x80050 gnd vdd FILL
XFILL_3__8866_ gnd vdd FILL
XFILL_0__15289_ gnd vdd FILL
XFILL_5__16029_ gnd vdd FILL
XFILL_1__6901_ gnd vdd FILL
X_9435_ _9435_/Q _9447_/CLK _9447_/R vdd _9351_/Y gnd vdd DFFSR
XFILL_3__7817_ gnd vdd FILL
XFILL_1__7881_ gnd vdd FILL
XFILL_4__7590_ gnd vdd FILL
XFILL_1__9620_ gnd vdd FILL
XSFILL33800x27050 gnd vdd FILL
X_9366_ _9366_/A _9425_/A _9365_/Y gnd _9366_/Y vdd OAI21X1
XFILL_4_BUFX2_insert503 gnd vdd FILL
XFILL_3__7748_ gnd vdd FILL
XSFILL43960x71050 gnd vdd FILL
XFILL_4_BUFX2_insert514 gnd vdd FILL
XFILL_4_BUFX2_insert525 gnd vdd FILL
X_8317_ _8315_/B _9597_/B gnd _8318_/C vdd NAND2X1
XFILL_1__9551_ gnd vdd FILL
XFILL_4_BUFX2_insert536 gnd vdd FILL
XSFILL28760x5050 gnd vdd FILL
XFILL_4_BUFX2_insert547 gnd vdd FILL
X_9297_ _9282_/A _7889_/B gnd _9298_/C vdd NAND2X1
XFILL_4__9260_ gnd vdd FILL
XFILL_3__7679_ gnd vdd FILL
XFILL_4_BUFX2_insert558 gnd vdd FILL
XFILL_1__8502_ gnd vdd FILL
XFILL_4_BUFX2_insert569 gnd vdd FILL
X_8248_ _8248_/A gnd _8250_/A vdd INVX1
XFILL_1__9482_ gnd vdd FILL
XFILL_3__9418_ gnd vdd FILL
XFILL_4__8211_ gnd vdd FILL
XFILL111960x37050 gnd vdd FILL
X_8179_ _8141_/A _7661_/CLK _8819_/R vdd _8143_/Y gnd vdd DFFSR
XSFILL23720x79050 gnd vdd FILL
XFILL_4__8142_ gnd vdd FILL
XFILL_3__9349_ gnd vdd FILL
XFILL112040x46050 gnd vdd FILL
XFILL_1__8364_ gnd vdd FILL
XFILL_4__8073_ gnd vdd FILL
XFILL_6__8009_ gnd vdd FILL
XFILL_3_CLKBUF1_insert205 gnd vdd FILL
XFILL_1__7315_ gnd vdd FILL
XFILL_3_CLKBUF1_insert216 gnd vdd FILL
XSFILL38920x60050 gnd vdd FILL
X_12820_ _12782_/A _12692_/CLK _12692_/R vdd _12820_/D gnd vdd DFFSR
XFILL_1__7246_ gnd vdd FILL
XFILL_1_BUFX2_insert404 gnd vdd FILL
X_12751_ _12751_/A _12777_/A _12751_/C gnd _12751_/Y vdd OAI21X1
XFILL_1_BUFX2_insert415 gnd vdd FILL
XFILL_1__7177_ gnd vdd FILL
XFILL_1_BUFX2_insert426 gnd vdd FILL
XFILL_1_BUFX2_insert437 gnd vdd FILL
XFILL_4__8975_ gnd vdd FILL
X_11702_ _11385_/Y _11379_/Y _11387_/Y gnd _11739_/B vdd AOI21X1
XFILL_1_BUFX2_insert448 gnd vdd FILL
XFILL_1_BUFX2_insert459 gnd vdd FILL
X_15470_ _13959_/A _16099_/B _16099_/C _13956_/A gnd _15471_/A vdd OAI22X1
X_12682_ _12624_/A _12538_/CLK _12689_/R vdd _12682_/D gnd vdd DFFSR
XFILL_2__7990_ gnd vdd FILL
XFILL_4__7926_ gnd vdd FILL
X_14421_ _14417_/Y _14421_/B gnd _14422_/C vdd NOR2X1
X_11633_ _12165_/Y _12282_/Y _11846_/C gnd _11634_/C vdd OAI21X1
XFILL_2__6941_ gnd vdd FILL
XFILL_1_CLKBUF1_insert1083 gnd vdd FILL
XFILL_4__7857_ gnd vdd FILL
X_14352_ _14352_/A _14352_/B gnd _14355_/C vdd NOR2X1
X_11564_ _11553_/B _11559_/Y _11802_/A gnd _11565_/A vdd OAI21X1
XFILL_2__9660_ gnd vdd FILL
XFILL_2__6872_ gnd vdd FILL
X_13303_ _13289_/B _13303_/B _13245_/B gnd _13303_/Y vdd OAI21X1
XFILL112120x26050 gnd vdd FILL
XFILL_5__10040_ gnd vdd FILL
X_10515_ _10515_/A _10548_/B _10514_/Y gnd _10515_/Y vdd OAI21X1
XFILL_5_BUFX2_insert370 gnd vdd FILL
XFILL_2__8611_ gnd vdd FILL
X_11495_ _11175_/Y _11509_/B _11495_/C _11176_/Y gnd _11495_/Y vdd AOI22X1
X_14283_ _9191_/Q _14868_/D _14283_/C _9897_/A gnd _14287_/A vdd AOI22X1
XBUFX2_insert60 _14983_/Y gnd _15842_/A vdd BUFX2
XFILL_4__10770_ gnd vdd FILL
XFILL_4__9527_ gnd vdd FILL
XFILL_5__8320_ gnd vdd FILL
XFILL_5_BUFX2_insert381 gnd vdd FILL
XFILL_2__9591_ gnd vdd FILL
XSFILL64040x11050 gnd vdd FILL
X_16022_ _15187_/A _14610_/Y _15187_/C gnd _16022_/Y vdd NOR3X1
XFILL_5_BUFX2_insert392 gnd vdd FILL
XBUFX2_insert71 _13393_/Y gnd _14697_/C vdd BUFX2
X_10446_ _10443_/A _8910_/B gnd _10447_/C vdd NAND2X1
X_13234_ _13246_/A _13215_/A gnd _13235_/C vdd NOR2X1
XBUFX2_insert82 _13372_/Y gnd _14506_/A vdd BUFX2
XBUFX2_insert93 _12357_/Y gnd _8195_/B vdd BUFX2
XFILL_3__11150_ gnd vdd FILL
XFILL_2__10900_ gnd vdd FILL
XFILL_1__9749_ gnd vdd FILL
XFILL_2__11880_ gnd vdd FILL
XFILL_5__8251_ gnd vdd FILL
XFILL_4__12440_ gnd vdd FILL
X_10377_ _10405_/B _9993_/B gnd _10377_/Y vdd NAND2X1
X_13165_ _13163_/Y _13149_/A _13165_/C gnd _13203_/D vdd OAI21X1
XFILL_5__11991_ gnd vdd FILL
XFILL_3__11081_ gnd vdd FILL
XFILL_2__10831_ gnd vdd FILL
XFILL_2__8473_ gnd vdd FILL
XFILL_5__7202_ gnd vdd FILL
XFILL_1__12260_ gnd vdd FILL
XFILL_5__8182_ gnd vdd FILL
X_12116_ _12823_/A _12150_/B gnd _12117_/C vdd NAND2X1
XFILL_4__9389_ gnd vdd FILL
XFILL_0__12990_ gnd vdd FILL
XFILL_5__10942_ gnd vdd FILL
X_13096_ _13096_/A _13155_/A _13095_/Y gnd _13096_/Y vdd OAI21X1
XFILL_3__10032_ gnd vdd FILL
XFILL_5__13730_ gnd vdd FILL
XFILL_2__7424_ gnd vdd FILL
XFILL_4__12371_ gnd vdd FILL
XFILL_1__11211_ gnd vdd FILL
XFILL_2__10762_ gnd vdd FILL
XFILL_2__13550_ gnd vdd FILL
XFILL_0__11941_ gnd vdd FILL
XFILL_1__12191_ gnd vdd FILL
X_12047_ _12047_/A _12388_/A _12011_/C gnd _12047_/Y vdd NAND3X1
XFILL_4__14110_ gnd vdd FILL
XSFILL84200x24050 gnd vdd FILL
XFILL_5__13661_ gnd vdd FILL
XFILL_4__11322_ gnd vdd FILL
XFILL_3__14840_ gnd vdd FILL
XFILL_2__12501_ gnd vdd FILL
XFILL_4__15090_ gnd vdd FILL
XFILL_5__10873_ gnd vdd FILL
XFILL_2__7355_ gnd vdd FILL
XFILL_1__11142_ gnd vdd FILL
XFILL_2__10693_ gnd vdd FILL
XFILL_0__14660_ gnd vdd FILL
XFILL_2__13481_ gnd vdd FILL
XFILL_0__11872_ gnd vdd FILL
XFILL_5__15400_ gnd vdd FILL
XFILL_5__12612_ gnd vdd FILL
XFILL_5__7064_ gnd vdd FILL
XFILL_4__14041_ gnd vdd FILL
XFILL_5__13592_ gnd vdd FILL
XFILL_2__15220_ gnd vdd FILL
XFILL_5__16380_ gnd vdd FILL
XFILL_4__11253_ gnd vdd FILL
XFILL_2__12432_ gnd vdd FILL
XFILL_0__13611_ gnd vdd FILL
XFILL_3__14771_ gnd vdd FILL
XFILL_3__11983_ gnd vdd FILL
XFILL_2__7286_ gnd vdd FILL
XFILL_1__15950_ gnd vdd FILL
XFILL_1__11073_ gnd vdd FILL
XFILL_0__10823_ gnd vdd FILL
XFILL_0__14591_ gnd vdd FILL
X_15806_ _15806_/A gnd _15806_/Y vdd INVX1
XFILL_5__15331_ gnd vdd FILL
XFILL_2__9025_ gnd vdd FILL
XFILL_2_BUFX2_insert260 gnd vdd FILL
XFILL_3__13722_ gnd vdd FILL
XFILL_3__10934_ gnd vdd FILL
XFILL_2__12363_ gnd vdd FILL
XFILL_0__16330_ gnd vdd FILL
XFILL_1__10024_ gnd vdd FILL
X_13998_ _13997_/Y _13998_/B gnd _14024_/B vdd NOR2X1
XFILL_4__11184_ gnd vdd FILL
XFILL_2__15151_ gnd vdd FILL
XFILL_1__14901_ gnd vdd FILL
XFILL_2_BUFX2_insert271 gnd vdd FILL
XFILL_0__13542_ gnd vdd FILL
XFILL_2_BUFX2_insert282 gnd vdd FILL
XFILL_0__10754_ gnd vdd FILL
XFILL_1__15881_ gnd vdd FILL
XSFILL99480x78050 gnd vdd FILL
XFILL_6__13833_ gnd vdd FILL
X_15737_ _7593_/A _15662_/A gnd _15740_/C vdd NAND2X1
XFILL_5__15262_ gnd vdd FILL
XFILL_2_BUFX2_insert293 gnd vdd FILL
XFILL_5__12474_ gnd vdd FILL
XFILL_4__10135_ gnd vdd FILL
X_12949_ _12949_/Q _8176_/CLK _7408_/R vdd _12949_/D gnd vdd DFFSR
XFILL_2__14102_ gnd vdd FILL
XFILL_2__11314_ gnd vdd FILL
XFILL_3__13653_ gnd vdd FILL
XFILL_4__15992_ gnd vdd FILL
XFILL_1__14832_ gnd vdd FILL
XFILL_2__12294_ gnd vdd FILL
XFILL_0__16261_ gnd vdd FILL
XFILL_2__15082_ gnd vdd FILL
XFILL_5__14213_ gnd vdd FILL
XFILL_0__13473_ gnd vdd FILL
XFILL_0__10685_ gnd vdd FILL
XFILL_5__7966_ gnd vdd FILL
XFILL_5__11425_ gnd vdd FILL
XFILL_3__12604_ gnd vdd FILL
XFILL_5__15193_ gnd vdd FILL
X_15668_ _15667_/Y _15660_/Y gnd _15691_/B vdd NOR2X1
XFILL_6__10976_ gnd vdd FILL
XFILL_0__15212_ gnd vdd FILL
XFILL_2__14033_ gnd vdd FILL
XFILL_4__14943_ gnd vdd FILL
XSFILL13560x29050 gnd vdd FILL
XFILL_3__16372_ gnd vdd FILL
XFILL_1_BUFX2_insert960 gnd vdd FILL
XFILL_4__10066_ gnd vdd FILL
XFILL_2__11245_ gnd vdd FILL
XFILL_1_BUFX2_insert971 gnd vdd FILL
XFILL_0__12424_ gnd vdd FILL
XFILL_3__13584_ gnd vdd FILL
XFILL_1__11975_ gnd vdd FILL
XFILL_0__16192_ gnd vdd FILL
XFILL_1_BUFX2_insert982 gnd vdd FILL
XFILL_3__6981_ gnd vdd FILL
XFILL_3__10796_ gnd vdd FILL
XFILL_5__6917_ gnd vdd FILL
XFILL_1__14763_ gnd vdd FILL
X_14619_ _7662_/Q gnd _14619_/Y vdd INVX1
XFILL_5__14144_ gnd vdd FILL
XFILL_1_BUFX2_insert993 gnd vdd FILL
XFILL_3__15323_ gnd vdd FILL
XFILL_5__11356_ gnd vdd FILL
X_7550_ _7550_/A _7624_/A _7549_/Y gnd _7640_/D vdd OAI21X1
XFILL_3__8720_ gnd vdd FILL
XFILL_4__14874_ gnd vdd FILL
XFILL_0__9991_ gnd vdd FILL
X_15599_ _14104_/A _15940_/B _15802_/D _15599_/D gnd _15602_/B vdd OAI22X1
XFILL_2__9927_ gnd vdd FILL
XFILL_1__10926_ gnd vdd FILL
XFILL_0__15143_ gnd vdd FILL
XFILL_2__11176_ gnd vdd FILL
XFILL_1__13714_ gnd vdd FILL
XFILL_5__9636_ gnd vdd FILL
XFILL_0__12355_ gnd vdd FILL
XFILL_5__6848_ gnd vdd FILL
XFILL_1__14694_ gnd vdd FILL
XFILL_5__10307_ gnd vdd FILL
XFILL_6__15434_ gnd vdd FILL
XFILL_4__13825_ gnd vdd FILL
XFILL_5__14075_ gnd vdd FILL
XSFILL28760x10050 gnd vdd FILL
XFILL_2__10127_ gnd vdd FILL
XFILL_3__15254_ gnd vdd FILL
X_7481_ _7457_/A _9017_/B gnd _7482_/C vdd NAND2X1
XFILL_5__11287_ gnd vdd FILL
XSFILL29240x17050 gnd vdd FILL
XBUFX2_insert270 _13364_/Y gnd _10678_/A vdd BUFX2
XFILL_3__8651_ gnd vdd FILL
XFILL_2__9858_ gnd vdd FILL
XFILL_3__12466_ gnd vdd FILL
XSFILL54040x43050 gnd vdd FILL
XFILL_0__11306_ gnd vdd FILL
XFILL_2__15984_ gnd vdd FILL
XFILL_1__13645_ gnd vdd FILL
XBUFX2_insert281 _15003_/Y gnd _15912_/D vdd BUFX2
XFILL_0__15074_ gnd vdd FILL
XBUFX2_insert292 _13356_/Y gnd _10318_/A vdd BUFX2
X_9220_ _9220_/A _9228_/A _9219_/Y gnd _9220_/Y vdd OAI21X1
XFILL_5__13026_ gnd vdd FILL
XFILL_0__12286_ gnd vdd FILL
XFILL_3__14205_ gnd vdd FILL
XFILL_5__10238_ gnd vdd FILL
XFILL_4__13756_ gnd vdd FILL
XFILL_0__8873_ gnd vdd FILL
XFILL_3__7602_ gnd vdd FILL
XFILL_3__11417_ gnd vdd FILL
XFILL_4__10968_ gnd vdd FILL
XFILL_3__15185_ gnd vdd FILL
XFILL_2__10058_ gnd vdd FILL
XFILL_0__14025_ gnd vdd FILL
XFILL_2__14935_ gnd vdd FILL
XFILL_2__9789_ gnd vdd FILL
XFILL_1__16364_ gnd vdd FILL
XFILL_3__12397_ gnd vdd FILL
XFILL_5__8518_ gnd vdd FILL
XFILL_1__13576_ gnd vdd FILL
XFILL_3__8582_ gnd vdd FILL
XFILL_0__11237_ gnd vdd FILL
XFILL_1__10788_ gnd vdd FILL
XFILL_5_CLKBUF1_insert160 gnd vdd FILL
XFILL_0__7824_ gnd vdd FILL
X_9151_ _9151_/A _7231_/B gnd _9152_/C vdd NAND2X1
XFILL_4__12707_ gnd vdd FILL
XFILL_5__9498_ gnd vdd FILL
XFILL_5_CLKBUF1_insert171 gnd vdd FILL
XFILL_6__11528_ gnd vdd FILL
XFILL_3__14136_ gnd vdd FILL
XFILL_5__10169_ gnd vdd FILL
XFILL_5_CLKBUF1_insert182 gnd vdd FILL
XFILL_6__15296_ gnd vdd FILL
XFILL_1__15315_ gnd vdd FILL
XFILL_1__12527_ gnd vdd FILL
XFILL_4__13687_ gnd vdd FILL
XFILL_3__11348_ gnd vdd FILL
XFILL_5_CLKBUF1_insert193 gnd vdd FILL
XFILL_2__14866_ gnd vdd FILL
XFILL_4__10899_ gnd vdd FILL
XFILL_5__8449_ gnd vdd FILL
X_8102_ _8166_/Q gnd _8102_/Y vdd INVX1
XFILL_1__16295_ gnd vdd FILL
XFILL_0__11168_ gnd vdd FILL
XFILL_6__14247_ gnd vdd FILL
XFILL_4__12638_ gnd vdd FILL
XFILL_0__7755_ gnd vdd FILL
XFILL_4__15426_ gnd vdd FILL
X_9082_ _9116_/B _9082_/B gnd _9082_/Y vdd NAND2X1
XFILL_2__13817_ gnd vdd FILL
XFILL_3__14067_ gnd vdd FILL
XFILL_5__14977_ gnd vdd FILL
XSFILL48920x23050 gnd vdd FILL
XFILL_3__7464_ gnd vdd FILL
XFILL_1__15246_ gnd vdd FILL
XFILL_1__12458_ gnd vdd FILL
XFILL_0__10119_ gnd vdd FILL
XFILL_3__11279_ gnd vdd FILL
XFILL_2__14797_ gnd vdd FILL
XFILL_0__15976_ gnd vdd FILL
X_8033_ _7959_/A _8161_/CLK _8033_/R vdd _8033_/D gnd vdd DFFSR
XFILL_0__11099_ gnd vdd FILL
XFILL_4__15357_ gnd vdd FILL
XFILL_3__13018_ gnd vdd FILL
XFILL_5__13928_ gnd vdd FILL
XFILL_4__12569_ gnd vdd FILL
XFILL_1__11409_ gnd vdd FILL
XFILL_0__7686_ gnd vdd FILL
XFILL_1__15177_ gnd vdd FILL
XFILL_2__13748_ gnd vdd FILL
XFILL_1__12389_ gnd vdd FILL
XFILL_0__14927_ gnd vdd FILL
XSFILL49000x32050 gnd vdd FILL
XFILL_4__14308_ gnd vdd FILL
XFILL_0__9425_ gnd vdd FILL
XFILL_5__13859_ gnd vdd FILL
XFILL_3__9134_ gnd vdd FILL
XFILL_4__15288_ gnd vdd FILL
XFILL_1__14128_ gnd vdd FILL
XFILL_2__13679_ gnd vdd FILL
XFILL_0__14858_ gnd vdd FILL
XFILL_0__9356_ gnd vdd FILL
XFILL_4__14239_ gnd vdd FILL
XSFILL109560x43050 gnd vdd FILL
XFILL_2__15418_ gnd vdd FILL
X_9984_ _9985_/B _9600_/B gnd _9984_/Y vdd NAND2X1
XFILL_1__14059_ gnd vdd FILL
XFILL_3__14969_ gnd vdd FILL
XFILL_0__13809_ gnd vdd FILL
XFILL_2__16398_ gnd vdd FILL
XFILL_1__7100_ gnd vdd FILL
XFILL_0__14789_ gnd vdd FILL
XFILL_1__8080_ gnd vdd FILL
XFILL_5__15529_ gnd vdd FILL
XSFILL54120x23050 gnd vdd FILL
X_8935_ _8873_/A _7400_/CLK _8935_/R vdd _8935_/D gnd vdd DFFSR
XFILL_0__9287_ gnd vdd FILL
XFILL_3__8016_ gnd vdd FILL
XFILL_2__15349_ gnd vdd FILL
XFILL_1__7031_ gnd vdd FILL
XFILL_0__8238_ gnd vdd FILL
X_8866_ _8866_/A _8845_/B _8866_/C gnd _8932_/D vdd OAI21X1
XSFILL43960x66050 gnd vdd FILL
X_7817_ _7824_/B _6921_/B gnd _7818_/C vdd NAND2X1
X_8797_ _8715_/A _7389_/CLK _8285_/R vdd _8717_/Y gnd vdd DFFSR
XFILL_4__8760_ gnd vdd FILL
XSFILL18760x42050 gnd vdd FILL
XSFILL8600x52050 gnd vdd FILL
XFILL_6__6888_ gnd vdd FILL
X_7748_ _7748_/A gnd _7750_/A vdd INVX1
XSFILL44040x75050 gnd vdd FILL
XFILL_1__8982_ gnd vdd FILL
XFILL_4__7711_ gnd vdd FILL
XSFILL98600x74050 gnd vdd FILL
XSFILL59640x54050 gnd vdd FILL
XFILL_3__9898_ gnd vdd FILL
XFILL_1__7933_ gnd vdd FILL
X_7679_ _7769_/Q gnd _7681_/A vdd INVX1
XFILL_3__8849_ gnd vdd FILL
X_9418_ _9418_/A gnd _9418_/Y vdd INVX1
XFILL_1__7864_ gnd vdd FILL
X_10300_ _10318_/A _9532_/B gnd _10301_/C vdd NAND2X1
XFILL_4_BUFX2_insert300 gnd vdd FILL
XFILL_4__7573_ gnd vdd FILL
XFILL_1__9603_ gnd vdd FILL
X_11280_ _11279_/Y gnd _11280_/Y vdd INVX1
XFILL_4_BUFX2_insert311 gnd vdd FILL
XFILL_4_BUFX2_insert322 gnd vdd FILL
XSFILL38920x55050 gnd vdd FILL
X_9349_ _9435_/Q gnd _9351_/A vdd INVX1
XFILL112440x62050 gnd vdd FILL
XFILL_4_BUFX2_insert333 gnd vdd FILL
X_10231_ _8183_/A _10280_/B gnd _10232_/C vdd NAND2X1
XFILL_4_BUFX2_insert344 gnd vdd FILL
XFILL_4_BUFX2_insert355 gnd vdd FILL
XFILL_1__9534_ gnd vdd FILL
XFILL_4_BUFX2_insert366 gnd vdd FILL
XFILL_4__9243_ gnd vdd FILL
XFILL_4_BUFX2_insert377 gnd vdd FILL
XFILL_4_BUFX2_insert388 gnd vdd FILL
XSFILL39000x64050 gnd vdd FILL
X_10162_ _10162_/A gnd _10162_/Y vdd INVX1
XFILL_4_BUFX2_insert399 gnd vdd FILL
XFILL_1__9465_ gnd vdd FILL
X_10093_ _10043_/A _8429_/CLK _9203_/R vdd _10093_/D gnd vdd DFFSR
X_14970_ _7925_/Q gnd _14971_/A vdd INVX1
XFILL_4__8125_ gnd vdd FILL
XFILL_1__9396_ gnd vdd FILL
XSFILL18840x22050 gnd vdd FILL
X_13921_ _13920_/Y _14887_/B _14456_/C _13919_/Y gnd _13921_/Y vdd OAI22X1
XFILL_1__8347_ gnd vdd FILL
XFILL_4__8056_ gnd vdd FILL
X_13852_ _13852_/A _13851_/Y _13852_/C gnd _13863_/A vdd NAND3X1
XSFILL99320x20050 gnd vdd FILL
XFILL_2__7071_ gnd vdd FILL
X_12803_ _11876_/B _7005_/CLK _7133_/R vdd _12733_/Y gnd vdd DFFSR
XSFILL23960x13050 gnd vdd FILL
XSFILL85000x50 gnd vdd FILL
XFILL_1__7229_ gnd vdd FILL
X_13783_ _10332_/Q gnd _13783_/Y vdd INVX1
X_10995_ _10993_/Y _10995_/B gnd _10997_/B vdd NOR2X1
XFILL_5__7820_ gnd vdd FILL
X_15522_ _15522_/A _15521_/Y gnd _15522_/Y vdd NOR2X1
XFILL_1_BUFX2_insert234 gnd vdd FILL
X_12734_ _11879_/B gnd _12736_/A vdd INVX1
XFILL_1_BUFX2_insert245 gnd vdd FILL
XFILL_1_BUFX2_insert256 gnd vdd FILL
XFILL_1_BUFX2_insert267 gnd vdd FILL
XFILL_3__10650_ gnd vdd FILL
XFILL_1_BUFX2_insert278 gnd vdd FILL
XFILL_4__8958_ gnd vdd FILL
XFILL_5__7751_ gnd vdd FILL
XFILL_5__11210_ gnd vdd FILL
XFILL_1_BUFX2_insert289 gnd vdd FILL
X_15453_ _15449_/Y _15453_/B gnd _15454_/B vdd NOR2X1
X_12665_ _12573_/A _7005_/CLK _12799_/R vdd _12665_/D gnd vdd DFFSR
XFILL_4__11940_ gnd vdd FILL
XFILL_2__11030_ gnd vdd FILL
XFILL_5__12190_ gnd vdd FILL
XFILL_0_BUFX2_insert901 gnd vdd FILL
XSFILL89240x72050 gnd vdd FILL
XFILL_0_BUFX2_insert912 gnd vdd FILL
XFILL_2__7973_ gnd vdd FILL
XFILL_0_BUFX2_insert923 gnd vdd FILL
XFILL_3__10581_ gnd vdd FILL
XFILL_1__11760_ gnd vdd FILL
XFILL_6__12500_ gnd vdd FILL
XFILL_0_BUFX2_insert934 gnd vdd FILL
X_14404_ _14358_/B _10802_/A _7658_/Q _14145_/D gnd _14404_/Y vdd AOI22X1
XFILL_5__7682_ gnd vdd FILL
XFILL_4__8889_ gnd vdd FILL
X_11616_ _11431_/Y _11616_/B _11615_/Y gnd _11616_/Y vdd OAI21X1
XFILL_5__11141_ gnd vdd FILL
X_15384_ _15384_/A _13881_/Y _13856_/Y _15384_/D gnd _15387_/B vdd OAI22X1
XFILL_0_BUFX2_insert945 gnd vdd FILL
XFILL_6__10692_ gnd vdd FILL
XFILL_3__12320_ gnd vdd FILL
XFILL_6__13480_ gnd vdd FILL
XFILL_2__6924_ gnd vdd FILL
X_12596_ _12596_/A vdd _12596_/C gnd _12672_/D vdd OAI21X1
XFILL_0_BUFX2_insert956 gnd vdd FILL
XFILL_4__11871_ gnd vdd FILL
XSFILL3720x75050 gnd vdd FILL
XFILL_0_BUFX2_insert967 gnd vdd FILL
XFILL_5__9421_ gnd vdd FILL
XFILL_0__12140_ gnd vdd FILL
XFILL_0_BUFX2_insert978 gnd vdd FILL
XFILL_1__11691_ gnd vdd FILL
XFILL_4__13610_ gnd vdd FILL
XFILL_0_BUFX2_insert989 gnd vdd FILL
X_14335_ _9448_/Q gnd _14335_/Y vdd INVX1
XSFILL84200x19050 gnd vdd FILL
XFILL_4__10822_ gnd vdd FILL
XFILL_5__11072_ gnd vdd FILL
X_11547_ _11521_/C _11437_/A _11537_/Y gnd _11547_/Y vdd NAND3X1
XFILL_4__14590_ gnd vdd FILL
XFILL_1__13430_ gnd vdd FILL
XFILL_3__12251_ gnd vdd FILL
XFILL_2__9643_ gnd vdd FILL
XSFILL94360x63050 gnd vdd FILL
XFILL_2__6855_ gnd vdd FILL
XFILL_1__10642_ gnd vdd FILL
XFILL_0__12071_ gnd vdd FILL
XFILL_5__9352_ gnd vdd FILL
XFILL_2__12981_ gnd vdd FILL
XFILL_6__12362_ gnd vdd FILL
XFILL_5__10023_ gnd vdd FILL
XFILL_5__14900_ gnd vdd FILL
XFILL_4__13541_ gnd vdd FILL
X_14266_ _8423_/Q gnd _14268_/A vdd INVX1
XFILL_3__11202_ gnd vdd FILL
XFILL_4__10753_ gnd vdd FILL
XFILL_2__14720_ gnd vdd FILL
X_11478_ _11360_/C _11478_/B _11477_/Y gnd _11478_/Y vdd NAND3X1
XFILL_5__15880_ gnd vdd FILL
XFILL_1__13361_ gnd vdd FILL
XFILL_2__11932_ gnd vdd FILL
XFILL_3__12182_ gnd vdd FILL
XFILL_0__11022_ gnd vdd FILL
XFILL_1__10573_ gnd vdd FILL
X_16005_ _16004_/Y _16005_/B _16005_/C gnd _16006_/B vdd NOR3X1
X_13217_ _13281_/B gnd _13218_/A vdd INVX1
XFILL_5__9283_ gnd vdd FILL
XFILL_6__11313_ gnd vdd FILL
X_10429_ _10427_/Y _10423_/B _10428_/Y gnd _10477_/D vdd OAI21X1
XFILL_5__14831_ gnd vdd FILL
XFILL_6__15081_ gnd vdd FILL
XFILL_4__16260_ gnd vdd FILL
XFILL_2__8525_ gnd vdd FILL
X_14197_ _9123_/A _14868_/D _14867_/C _9957_/Q gnd _14197_/Y vdd AOI22X1
XFILL_1__15100_ gnd vdd FILL
XFILL_4__13472_ gnd vdd FILL
XFILL_1__12312_ gnd vdd FILL
XFILL_3__11133_ gnd vdd FILL
XFILL_4__10684_ gnd vdd FILL
XFILL_2__14651_ gnd vdd FILL
XFILL_1__16080_ gnd vdd FILL
XFILL_1__13292_ gnd vdd FILL
XFILL_0__15830_ gnd vdd FILL
XFILL_2__11863_ gnd vdd FILL
XSFILL59240x2050 gnd vdd FILL
XFILL_5__8234_ gnd vdd FILL
XFILL_4__15211_ gnd vdd FILL
XFILL_6__14032_ gnd vdd FILL
X_13148_ _12184_/A gnd _13150_/A vdd INVX1
XFILL_4__12423_ gnd vdd FILL
XSFILL64040x9050 gnd vdd FILL
XFILL_2__13602_ gnd vdd FILL
XFILL_5__11974_ gnd vdd FILL
XFILL_4__16191_ gnd vdd FILL
XFILL_1__15031_ gnd vdd FILL
XFILL_3__15941_ gnd vdd FILL
XFILL_3__11064_ gnd vdd FILL
XFILL_5__14762_ gnd vdd FILL
XFILL_2__10814_ gnd vdd FILL
XFILL_2__8456_ gnd vdd FILL
XFILL_1__12243_ gnd vdd FILL
XFILL_2__14582_ gnd vdd FILL
XFILL_0__12973_ gnd vdd FILL
XSFILL74280x30050 gnd vdd FILL
XFILL_2__11794_ gnd vdd FILL
XFILL_0__15761_ gnd vdd FILL
XFILL_5__13713_ gnd vdd FILL
XFILL_4__15142_ gnd vdd FILL
XFILL_6__11175_ gnd vdd FILL
XFILL_4__12354_ gnd vdd FILL
XFILL_5__10925_ gnd vdd FILL
X_13079_ _11887_/A gnd _13081_/A vdd INVX1
XFILL_2__16321_ gnd vdd FILL
XSFILL48440x40050 gnd vdd FILL
XFILL_0__7471_ gnd vdd FILL
XFILL_3__10015_ gnd vdd FILL
XFILL_5__14693_ gnd vdd FILL
XFILL_3__15872_ gnd vdd FILL
XFILL_2__13533_ gnd vdd FILL
XFILL_5__7116_ gnd vdd FILL
XFILL_3__7180_ gnd vdd FILL
XFILL_0__11924_ gnd vdd FILL
XFILL_0__14712_ gnd vdd FILL
XFILL_1__12174_ gnd vdd FILL
XFILL_2__8387_ gnd vdd FILL
XFILL_2__10745_ gnd vdd FILL
XFILL_0__15692_ gnd vdd FILL
XFILL_0__9210_ gnd vdd FILL
XFILL_5__8096_ gnd vdd FILL
XSFILL53960x29050 gnd vdd FILL
XFILL_4__11305_ gnd vdd FILL
XFILL_5__13644_ gnd vdd FILL
XFILL_3__14823_ gnd vdd FILL
XFILL_4__15073_ gnd vdd FILL
XFILL_2__7338_ gnd vdd FILL
XFILL_1__11125_ gnd vdd FILL
XFILL_2__16252_ gnd vdd FILL
XFILL_4__12285_ gnd vdd FILL
XFILL_0__14643_ gnd vdd FILL
XFILL_2__13464_ gnd vdd FILL
XFILL_2__10676_ gnd vdd FILL
XFILL_5__7047_ gnd vdd FILL
XFILL_0__11855_ gnd vdd FILL
XFILL_0__9141_ gnd vdd FILL
XFILL_4__14024_ gnd vdd FILL
XFILL_6__10057_ gnd vdd FILL
XFILL_2__15203_ gnd vdd FILL
XFILL_5__16363_ gnd vdd FILL
XFILL_4__11236_ gnd vdd FILL
XFILL_5__10787_ gnd vdd FILL
XFILL_2__12415_ gnd vdd FILL
X_6981_ _6982_/B _6981_/B gnd _6981_/Y vdd NAND2X1
XSFILL53560x31050 gnd vdd FILL
XFILL_5__13575_ gnd vdd FILL
XFILL_3__14754_ gnd vdd FILL
XFILL_0__10806_ gnd vdd FILL
XFILL_2__16183_ gnd vdd FILL
XFILL_3__11966_ gnd vdd FILL
XFILL_1__15933_ gnd vdd FILL
XFILL_1__11056_ gnd vdd FILL
XFILL_0__14574_ gnd vdd FILL
XFILL_2__13395_ gnd vdd FILL
XFILL_5__15314_ gnd vdd FILL
XFILL_0__11786_ gnd vdd FILL
X_8720_ _8718_/Y _8740_/A _8720_/C gnd _8798_/D vdd OAI21X1
XFILL_5__12526_ gnd vdd FILL
XSFILL94440x43050 gnd vdd FILL
XFILL_2__9008_ gnd vdd FILL
XFILL_3__13705_ gnd vdd FILL
XFILL_3__10917_ gnd vdd FILL
XFILL_1__10007_ gnd vdd FILL
XFILL_2__15134_ gnd vdd FILL
XFILL_4__11167_ gnd vdd FILL
XFILL_5__16294_ gnd vdd FILL
XFILL_2__12346_ gnd vdd FILL
XFILL_0__16313_ gnd vdd FILL
XFILL_3__14685_ gnd vdd FILL
XFILL_0__13525_ gnd vdd FILL
XFILL_3__11897_ gnd vdd FILL
XFILL_1__15864_ gnd vdd FILL
XFILL_5__8998_ gnd vdd FILL
X_8651_ _8655_/B _7499_/B gnd _8652_/C vdd NAND2X1
XFILL_5__12457_ gnd vdd FILL
XFILL_5__15245_ gnd vdd FILL
XFILL_6_BUFX2_insert428 gnd vdd FILL
XFILL_4__10118_ gnd vdd FILL
XFILL_3__13636_ gnd vdd FILL
XFILL_4__15975_ gnd vdd FILL
XFILL_1__14815_ gnd vdd FILL
XFILL_6_BUFX2_insert439 gnd vdd FILL
XFILL_2__15065_ gnd vdd FILL
XFILL_4__11098_ gnd vdd FILL
XFILL_0__16244_ gnd vdd FILL
XFILL_0__13456_ gnd vdd FILL
XFILL_2__12277_ gnd vdd FILL
XFILL_5__7949_ gnd vdd FILL
XFILL_1__15795_ gnd vdd FILL
XFILL_0__10668_ gnd vdd FILL
X_7602_ _7658_/Q gnd _7604_/A vdd INVX1
XFILL_5__11408_ gnd vdd FILL
XFILL_5__15176_ gnd vdd FILL
XFILL_5__12388_ gnd vdd FILL
XFILL_3__16355_ gnd vdd FILL
XFILL_2__14016_ gnd vdd FILL
XFILL_4__10049_ gnd vdd FILL
X_8582_ _8619_/B _8582_/B gnd _8582_/Y vdd NAND2X1
XFILL_1_BUFX2_insert790 gnd vdd FILL
XFILL_4__14926_ gnd vdd FILL
XFILL_0__12407_ gnd vdd FILL
XFILL_3__9752_ gnd vdd FILL
XFILL_3__13567_ gnd vdd FILL
XSFILL48920x18050 gnd vdd FILL
XFILL_2__11228_ gnd vdd FILL
XFILL_0__16175_ gnd vdd FILL
XSFILL18680x57050 gnd vdd FILL
XFILL_3__10779_ gnd vdd FILL
XFILL_3__6964_ gnd vdd FILL
XFILL_1__14746_ gnd vdd FILL
XFILL_1__11958_ gnd vdd FILL
XFILL_0__13387_ gnd vdd FILL
X_7533_ _7533_/Q _8306_/CLK _7533_/R vdd _7485_/Y gnd vdd DFFSR
XFILL_3__15306_ gnd vdd FILL
XFILL_5__14127_ gnd vdd FILL
XFILL_5__11339_ gnd vdd FILL
XFILL_3__8703_ gnd vdd FILL
XFILL_0__9974_ gnd vdd FILL
XFILL_3__12518_ gnd vdd FILL
XFILL_4_BUFX2_insert1007 gnd vdd FILL
XFILL_4__14857_ gnd vdd FILL
XFILL_3__16286_ gnd vdd FILL
XFILL_2__11159_ gnd vdd FILL
XFILL_0__15126_ gnd vdd FILL
XFILL_1__10909_ gnd vdd FILL
XFILL_4_BUFX2_insert1018 gnd vdd FILL
XFILL_3__9683_ gnd vdd FILL
XFILL_0__12338_ gnd vdd FILL
XFILL_3__13498_ gnd vdd FILL
XFILL_4_BUFX2_insert1029 gnd vdd FILL
XFILL_3__6895_ gnd vdd FILL
XFILL_1__14677_ gnd vdd FILL
XFILL_5__9619_ gnd vdd FILL
XSFILL48520x20050 gnd vdd FILL
XFILL_6__12629_ gnd vdd FILL
XFILL_1__11889_ gnd vdd FILL
XFILL_5__14058_ gnd vdd FILL
XFILL_4_BUFX2_insert50 gnd vdd FILL
X_7464_ _7464_/A _7425_/B _7464_/C gnd _7464_/Y vdd OAI21X1
XFILL_4__13808_ gnd vdd FILL
XFILL_3__15237_ gnd vdd FILL
XFILL_4_BUFX2_insert61 gnd vdd FILL
XFILL_4_BUFX2_insert72 gnd vdd FILL
XFILL_3__8634_ gnd vdd FILL
XFILL_3__12449_ gnd vdd FILL
XFILL_1__16416_ gnd vdd FILL
XFILL_1__13628_ gnd vdd FILL
XFILL_4_BUFX2_insert83 gnd vdd FILL
XFILL_0__15057_ gnd vdd FILL
XFILL_2__15967_ gnd vdd FILL
XSFILL89400x32050 gnd vdd FILL
XFILL_4__14788_ gnd vdd FILL
XFILL_0__12269_ gnd vdd FILL
XFILL_5__13009_ gnd vdd FILL
XFILL_4_BUFX2_insert94 gnd vdd FILL
X_9203_ _9203_/Q _8429_/CLK _9203_/R vdd _9203_/D gnd vdd DFFSR
XFILL_0__8856_ gnd vdd FILL
XFILL_3__15168_ gnd vdd FILL
XFILL_0__14008_ gnd vdd FILL
XFILL_2__14918_ gnd vdd FILL
X_7395_ _7325_/A _9077_/CLK _8433_/R vdd _7395_/D gnd vdd DFFSR
XFILL_4__13739_ gnd vdd FILL
XFILL_1__16347_ gnd vdd FILL
XFILL_2__15898_ gnd vdd FILL
XFILL_1__13559_ gnd vdd FILL
XFILL_0__7807_ gnd vdd FILL
X_9134_ _9134_/A _9116_/B _9133_/Y gnd _9134_/Y vdd OAI21X1
XFILL112360x77050 gnd vdd FILL
XFILL_3__14119_ gnd vdd FILL
XSFILL54120x18050 gnd vdd FILL
XFILL_1__7580_ gnd vdd FILL
XFILL_0__8787_ gnd vdd FILL
XFILL_2__14849_ gnd vdd FILL
XFILL_3__15099_ gnd vdd FILL
XFILL_2_BUFX2_insert1000 gnd vdd FILL
XFILL_3__8496_ gnd vdd FILL
XFILL_1__16278_ gnd vdd FILL
XFILL_2_BUFX2_insert1011 gnd vdd FILL
XFILL_3_BUFX2_insert307 gnd vdd FILL
XFILL_4__15409_ gnd vdd FILL
XFILL_3_BUFX2_insert318 gnd vdd FILL
XFILL_0__7738_ gnd vdd FILL
X_9065_ _9065_/Q _7532_/CLK _8816_/R vdd _9009_/Y gnd vdd DFFSR
XFILL_2_BUFX2_insert1022 gnd vdd FILL
XFILL_2_BUFX2_insert1033 gnd vdd FILL
XFILL_4__16389_ gnd vdd FILL
XFILL_1__15229_ gnd vdd FILL
XFILL_3__7447_ gnd vdd FILL
XFILL_3_BUFX2_insert329 gnd vdd FILL
XFILL_2_BUFX2_insert1044 gnd vdd FILL
XFILL_2_BUFX2_insert1055 gnd vdd FILL
XFILL_0__15959_ gnd vdd FILL
X_8016_ _8052_/Q gnd _8018_/A vdd INVX1
XFILL_1__9250_ gnd vdd FILL
XFILL_2_BUFX2_insert1066 gnd vdd FILL
XFILL_2_BUFX2_insert1088 gnd vdd FILL
XFILL_3__7378_ gnd vdd FILL
XFILL_0__9408_ gnd vdd FILL
XFILL_1__8201_ gnd vdd FILL
XSFILL18760x37050 gnd vdd FILL
XFILL_3__9117_ gnd vdd FILL
XSFILL8600x47050 gnd vdd FILL
XSFILL33800x40050 gnd vdd FILL
XFILL_1__8132_ gnd vdd FILL
XFILL_0__9339_ gnd vdd FILL
XFILL_4__9930_ gnd vdd FILL
X_9967_ _9967_/Q _9568_/CLK _8431_/R vdd _9967_/D gnd vdd DFFSR
XFILL_1__8063_ gnd vdd FILL
X_8918_ _8918_/Q _7662_/CLK _8430_/R vdd _8918_/D gnd vdd DFFSR
XSFILL23880x28050 gnd vdd FILL
XFILL_4__9861_ gnd vdd FILL
X_9898_ _9902_/B _9898_/B gnd _9898_/Y vdd NAND2X1
XFILL_0_BUFX2_insert1070 gnd vdd FILL
XFILL_6__7989_ gnd vdd FILL
XFILL_4_CLKBUF1_insert119 gnd vdd FILL
XSFILL108600x54050 gnd vdd FILL
X_10780_ _10778_/Y _10762_/B _10780_/C gnd _10850_/D vdd OAI21X1
XFILL_0_BUFX2_insert1092 gnd vdd FILL
X_8849_ _8927_/Q gnd _8851_/A vdd INVX1
XFILL_4__9792_ gnd vdd FILL
XFILL112440x57050 gnd vdd FILL
XFILL_6_BUFX2_insert940 gnd vdd FILL
XSFILL109240x20050 gnd vdd FILL
XFILL112360x2050 gnd vdd FILL
XFILL_4__8743_ gnd vdd FILL
X_12450_ _12448_/Y vdd _12449_/Y gnd _12450_/Y vdd OAI21X1
XSFILL39000x59050 gnd vdd FILL
XFILL_1__8965_ gnd vdd FILL
X_11401_ _11056_/A _11401_/B _11400_/Y gnd _11623_/B vdd OAI21X1
X_12381_ _12381_/A _12419_/A _12381_/C gnd _12381_/Y vdd OAI21X1
XSFILL114360x11050 gnd vdd FILL
XFILL_1__8896_ gnd vdd FILL
XFILL_4__7625_ gnd vdd FILL
X_14120_ _14120_/A _14112_/Y _14120_/C gnd _14120_/Y vdd NAND3X1
XSFILL18840x17050 gnd vdd FILL
X_11332_ _11201_/Y _11200_/Y gnd _11414_/A vdd NOR2X1
XSFILL114600x73050 gnd vdd FILL
XFILL_1__7847_ gnd vdd FILL
XFILL_4__7556_ gnd vdd FILL
X_14051_ _14050_/Y _14815_/C _14051_/C _14049_/Y gnd _14051_/Y vdd OAI22X1
XSFILL69080x54050 gnd vdd FILL
X_11263_ _11261_/Y _11263_/B gnd _11448_/B vdd NOR2X1
XSFILL85080x9050 gnd vdd FILL
X_13002_ _6887_/A gnd _13002_/Y vdd INVX1
X_10214_ _10214_/Q _8947_/CLK _9069_/R vdd _10152_/Y gnd vdd DFFSR
XFILL_4__7487_ gnd vdd FILL
XFILL_2__8310_ gnd vdd FILL
XFILL_1__9517_ gnd vdd FILL
X_11194_ _12322_/Y _11193_/Y gnd _11194_/Y vdd NOR2X1
XFILL_4__9226_ gnd vdd FILL
XFILL_2__9290_ gnd vdd FILL
X_10145_ _10169_/A _7329_/B gnd _10145_/Y vdd NAND2X1
XFILL_3_BUFX2_insert830 gnd vdd FILL
XSFILL23800x6050 gnd vdd FILL
XFILL_3_BUFX2_insert841 gnd vdd FILL
XFILL_3_BUFX2_insert852 gnd vdd FILL
XFILL_2__8241_ gnd vdd FILL
XFILL_3_BUFX2_insert863 gnd vdd FILL
XFILL_4__9157_ gnd vdd FILL
XFILL_3_BUFX2_insert874 gnd vdd FILL
X_10076_ _9992_/A _7534_/CLK _8156_/R vdd _9994_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert885 gnd vdd FILL
X_14953_ _9043_/A gnd _16314_/B vdd INVX1
XFILL_2__10530_ gnd vdd FILL
XFILL_3_BUFX2_insert896 gnd vdd FILL
XFILL_5__11690_ gnd vdd FILL
XFILL_1__9379_ gnd vdd FILL
XFILL_4__8108_ gnd vdd FILL
XFILL_4__9088_ gnd vdd FILL
X_13904_ _8159_/Q gnd _15429_/C vdd INVX1
XFILL_5__10641_ gnd vdd FILL
XFILL_4__12070_ gnd vdd FILL
XFILL_2__7123_ gnd vdd FILL
XFILL_3__11820_ gnd vdd FILL
X_14884_ _14506_/A _14884_/B _14883_/Y _13630_/B gnd _14888_/A vdd OAI22X1
XFILL_0__11640_ gnd vdd FILL
XFILL_5__13360_ gnd vdd FILL
X_13835_ _8669_/Q gnd _13835_/Y vdd INVX1
XFILL_4__11021_ gnd vdd FILL
XFILL_5__10572_ gnd vdd FILL
XFILL_2__12200_ gnd vdd FILL
XSFILL110280x82050 gnd vdd FILL
XFILL_2__7054_ gnd vdd FILL
XFILL_3__11751_ gnd vdd FILL
XFILL_2__10392_ gnd vdd FILL
XSFILL94360x58050 gnd vdd FILL
XFILL_5__12311_ gnd vdd FILL
XFILL_5__8852_ gnd vdd FILL
XFILL_0__11571_ gnd vdd FILL
XFILL_5__13291_ gnd vdd FILL
XFILL_3__10702_ gnd vdd FILL
X_13766_ _16339_/A gnd _13768_/D vdd INVX1
XFILL_0__13310_ gnd vdd FILL
X_10978_ _10906_/A gnd _10980_/A vdd INVX1
XFILL_3__14470_ gnd vdd FILL
XFILL_2__12131_ gnd vdd FILL
XFILL_0__10522_ gnd vdd FILL
XFILL_5__7803_ gnd vdd FILL
XFILL_3__11682_ gnd vdd FILL
X_15505_ _8801_/Q gnd _15506_/A vdd INVX1
XFILL_1__12861_ gnd vdd FILL
XSFILL69160x34050 gnd vdd FILL
XFILL_0__14290_ gnd vdd FILL
X_12717_ _12777_/A memoryOutData[7] gnd _12718_/C vdd NAND2X1
XFILL_5__8783_ gnd vdd FILL
XFILL_5__15030_ gnd vdd FILL
XFILL_5__12242_ gnd vdd FILL
XFILL_3__13421_ gnd vdd FILL
XFILL_1__14600_ gnd vdd FILL
XFILL_4__12972_ gnd vdd FILL
XFILL_3__10633_ gnd vdd FILL
XFILL_2__12062_ gnd vdd FILL
XFILL_4__15760_ gnd vdd FILL
X_13697_ _13697_/A _13696_/Y gnd _13697_/Y vdd NOR2X1
XFILL_0__13241_ gnd vdd FILL
XFILL_1__11812_ gnd vdd FILL
XFILL_5__7734_ gnd vdd FILL
XFILL_0__10453_ gnd vdd FILL
XFILL_1__15580_ gnd vdd FILL
XFILL_0_BUFX2_insert720 gnd vdd FILL
X_15436_ _15524_/A _13902_/D _15436_/C _15521_/C gnd _15437_/C vdd OAI22X1
X_12648_ _12648_/A gnd _12648_/Y vdd INVX1
XFILL_0_BUFX2_insert731 gnd vdd FILL
XFILL_4__11923_ gnd vdd FILL
XFILL_5__12173_ gnd vdd FILL
XFILL_4__14711_ gnd vdd FILL
XFILL_2__11013_ gnd vdd FILL
XFILL_3__16140_ gnd vdd FILL
XFILL_3__13352_ gnd vdd FILL
XFILL_4__15691_ gnd vdd FILL
XSFILL104360x43050 gnd vdd FILL
XFILL_0_BUFX2_insert742 gnd vdd FILL
XFILL_1__14531_ gnd vdd FILL
XFILL_3__10564_ gnd vdd FILL
XFILL_0_BUFX2_insert753 gnd vdd FILL
XFILL_2__7956_ gnd vdd FILL
XFILL_0__13172_ gnd vdd FILL
XFILL_1__11743_ gnd vdd FILL
XFILL_0_CLKBUF1_insert190 gnd vdd FILL
XFILL_0_BUFX2_insert764 gnd vdd FILL
XFILL_0__10384_ gnd vdd FILL
XFILL_5__11124_ gnd vdd FILL
X_15367_ _15367_/A _15367_/B gnd _15371_/A vdd NOR2X1
XFILL_3__12303_ gnd vdd FILL
XFILL_0_BUFX2_insert775 gnd vdd FILL
XFILL_0__6971_ gnd vdd FILL
X_12579_ _12667_/Q gnd _12579_/Y vdd INVX1
XFILL_4__14642_ gnd vdd FILL
XFILL_0_BUFX2_insert786 gnd vdd FILL
XSFILL48440x35050 gnd vdd FILL
XFILL_2__15821_ gnd vdd FILL
XFILL_2__6907_ gnd vdd FILL
XFILL_3__16071_ gnd vdd FILL
XFILL_4__11854_ gnd vdd FILL
XFILL_3__13283_ gnd vdd FILL
XFILL_5__9404_ gnd vdd FILL
XFILL_0__12123_ gnd vdd FILL
XFILL_0_BUFX2_insert797 gnd vdd FILL
XFILL_2__7887_ gnd vdd FILL
XFILL_3__10495_ gnd vdd FILL
XFILL_1__14462_ gnd vdd FILL
XFILL_1__11674_ gnd vdd FILL
X_14318_ _8168_/Q gnd _14318_/Y vdd INVX1
XFILL_0__8710_ gnd vdd FILL
XFILL_4__10805_ gnd vdd FILL
XFILL_5__15932_ gnd vdd FILL
XFILL_3__15022_ gnd vdd FILL
XFILL_5__7596_ gnd vdd FILL
XFILL_5__11055_ gnd vdd FILL
XFILL_4__14573_ gnd vdd FILL
XFILL_1__16201_ gnd vdd FILL
X_15298_ _10844_/Q _15357_/B _15356_/C _15298_/D gnd _15298_/Y vdd AOI22X1
XFILL_2__9626_ gnd vdd FILL
XFILL_3__12234_ gnd vdd FILL
XFILL_1__10625_ gnd vdd FILL
XFILL_2__6838_ gnd vdd FILL
XFILL_1__13413_ gnd vdd FILL
XFILL_4__11785_ gnd vdd FILL
XFILL_2__15752_ gnd vdd FILL
XFILL_5__9335_ gnd vdd FILL
XFILL_2__12964_ gnd vdd FILL
XFILL_0__12054_ gnd vdd FILL
XFILL_1__14393_ gnd vdd FILL
XFILL_5__10006_ gnd vdd FILL
X_14249_ _15692_/A _13803_/A _13587_/C _14248_/Y gnd _14250_/A vdd OAI22X1
XFILL_4__16312_ gnd vdd FILL
XFILL_0__8641_ gnd vdd FILL
XFILL_4__13524_ gnd vdd FILL
X_7180_ _7181_/B _7180_/B gnd _7180_/Y vdd NAND2X1
XFILL_2__14703_ gnd vdd FILL
XFILL_5__15863_ gnd vdd FILL
XFILL_2__11915_ gnd vdd FILL
XFILL_3__12165_ gnd vdd FILL
XFILL_2__9557_ gnd vdd FILL
XFILL_3__8350_ gnd vdd FILL
XFILL_0__11005_ gnd vdd FILL
XFILL_1__16132_ gnd vdd FILL
XFILL_1__13344_ gnd vdd FILL
XFILL_2__15683_ gnd vdd FILL
XFILL_1__10556_ gnd vdd FILL
XFILL_2__12895_ gnd vdd FILL
XFILL_5__9266_ gnd vdd FILL
XFILL_5__14814_ gnd vdd FILL
XFILL_2__8508_ gnd vdd FILL
XFILL_4__16243_ gnd vdd FILL
XFILL_4__13455_ gnd vdd FILL
XSFILL13560x42050 gnd vdd FILL
XFILL_0__8572_ gnd vdd FILL
XFILL_3__11116_ gnd vdd FILL
XFILL_3__7301_ gnd vdd FILL
XFILL_2__14634_ gnd vdd FILL
XSFILL94440x38050 gnd vdd FILL
XFILL_5__15794_ gnd vdd FILL
XFILL_4__10667_ gnd vdd FILL
XFILL_2__9488_ gnd vdd FILL
XFILL_1__13275_ gnd vdd FILL
XFILL_3__12096_ gnd vdd FILL
XFILL_5__8217_ gnd vdd FILL
XFILL_0__15813_ gnd vdd FILL
XFILL_1__16063_ gnd vdd FILL
XFILL_2__11846_ gnd vdd FILL
XFILL_1__10487_ gnd vdd FILL
XFILL_4__12406_ gnd vdd FILL
XFILL_4__16174_ gnd vdd FILL
XFILL_5__14745_ gnd vdd FILL
XFILL_3__7232_ gnd vdd FILL
XFILL_3__15924_ gnd vdd FILL
XFILL_5__11957_ gnd vdd FILL
XFILL_4__13386_ gnd vdd FILL
XFILL_1__15014_ gnd vdd FILL
XFILL_2__8439_ gnd vdd FILL
XFILL_1__12226_ gnd vdd FILL
XFILL_3__11047_ gnd vdd FILL
XSFILL69240x14050 gnd vdd FILL
XFILL_2__14565_ gnd vdd FILL
XFILL_5__8148_ gnd vdd FILL
XFILL_2__11777_ gnd vdd FILL
XFILL_0__15744_ gnd vdd FILL
XFILL_4__15125_ gnd vdd FILL
XFILL_0__12956_ gnd vdd FILL
XFILL_5__10908_ gnd vdd FILL
XFILL_2__16304_ gnd vdd FILL
XFILL_1_BUFX2_insert9 gnd vdd FILL
XFILL_0__7454_ gnd vdd FILL
XFILL_4__12337_ gnd vdd FILL
XFILL_5__14676_ gnd vdd FILL
XFILL_2__13516_ gnd vdd FILL
XFILL_5__11888_ gnd vdd FILL
XFILL_1__12157_ gnd vdd FILL
XFILL_3__15855_ gnd vdd FILL
XFILL_3__7163_ gnd vdd FILL
XFILL_2__14496_ gnd vdd FILL
XFILL_0__11907_ gnd vdd FILL
XFILL_6__10109_ gnd vdd FILL
XFILL_6__8961_ gnd vdd FILL
XFILL_5__8079_ gnd vdd FILL
XFILL_0__15675_ gnd vdd FILL
XFILL_0__12887_ gnd vdd FILL
XFILL_5__16415_ gnd vdd FILL
XFILL_5__13627_ gnd vdd FILL
X_9821_ _9821_/Q _9707_/CLK _8819_/R vdd _9821_/D gnd vdd DFFSR
XFILL_4__15056_ gnd vdd FILL
XFILL_6__15966_ gnd vdd FILL
XFILL_2__16235_ gnd vdd FILL
XFILL_3__14806_ gnd vdd FILL
XFILL_4__12268_ gnd vdd FILL
XFILL_1__11108_ gnd vdd FILL
XSFILL33720x55050 gnd vdd FILL
XFILL_2__13447_ gnd vdd FILL
XFILL_3__15786_ gnd vdd FILL
XSFILL8680x21050 gnd vdd FILL
XFILL_2__10659_ gnd vdd FILL
XFILL_3__7094_ gnd vdd FILL
XFILL_0__14626_ gnd vdd FILL
XFILL_3__12998_ gnd vdd FILL
XFILL_1__12088_ gnd vdd FILL
XFILL_0__11838_ gnd vdd FILL
XFILL_0__9124_ gnd vdd FILL
XFILL_4__14007_ gnd vdd FILL
XFILL_6__14917_ gnd vdd FILL
XSFILL43080x80050 gnd vdd FILL
XFILL_5__16346_ gnd vdd FILL
XFILL_4__11219_ gnd vdd FILL
X_9752_ _9741_/B _9624_/B gnd _9753_/C vdd NAND2X1
XFILL_3__14737_ gnd vdd FILL
XFILL_5__13558_ gnd vdd FILL
XFILL_1__15916_ gnd vdd FILL
XFILL_2__16166_ gnd vdd FILL
XFILL_3__11949_ gnd vdd FILL
XFILL_4__12199_ gnd vdd FILL
X_6964_ _6962_/Y _6985_/B _6963_/Y gnd _6964_/Y vdd OAI21X1
XSFILL88920x20050 gnd vdd FILL
XFILL_1__11039_ gnd vdd FILL
XFILL_2__13378_ gnd vdd FILL
XSFILL89400x27050 gnd vdd FILL
XFILL_0__14557_ gnd vdd FILL
XSFILL59160x66050 gnd vdd FILL
XFILL_0__11769_ gnd vdd FILL
X_8703_ _8793_/Q gnd _8703_/Y vdd INVX1
XFILL_5__12509_ gnd vdd FILL
XFILL_2__15117_ gnd vdd FILL
XFILL_5__16277_ gnd vdd FILL
X_9683_ _9683_/A gnd _9685_/A vdd INVX1
XFILL_2__12329_ gnd vdd FILL
X_6895_ _6895_/A gnd memoryWriteData[25] vdd BUFX2
XFILL_3__14668_ gnd vdd FILL
XFILL_5__13489_ gnd vdd FILL
XFILL_2__16097_ gnd vdd FILL
XFILL_1__15847_ gnd vdd FILL
XFILL_0__13508_ gnd vdd FILL
XFILL_0__14488_ gnd vdd FILL
XFILL_0__8006_ gnd vdd FILL
XFILL111880x65050 gnd vdd FILL
XFILL_5__15228_ gnd vdd FILL
XFILL_3__13619_ gnd vdd FILL
X_8634_ _8634_/A _8589_/B _8634_/C gnd _8634_/Y vdd OAI21X1
XFILL_3__16407_ gnd vdd FILL
XFILL_6__14779_ gnd vdd FILL
XFILL_3__9804_ gnd vdd FILL
XFILL_2__15048_ gnd vdd FILL
XFILL_4__15958_ gnd vdd FILL
XFILL_3__14599_ gnd vdd FILL
XFILL_0__16227_ gnd vdd FILL
XFILL_0__13439_ gnd vdd FILL
XFILL_3__7996_ gnd vdd FILL
XFILL_1__15778_ gnd vdd FILL
XSFILL94520x18050 gnd vdd FILL
XFILL_6__9513_ gnd vdd FILL
XSFILL13640x22050 gnd vdd FILL
XFILL_5_BUFX2_insert903 gnd vdd FILL
XFILL_5_BUFX2_insert914 gnd vdd FILL
XFILL_3__16338_ gnd vdd FILL
XFILL_5__15159_ gnd vdd FILL
XFILL_4__14909_ gnd vdd FILL
X_8565_ _8531_/A _7010_/CLK _7413_/R vdd _8533_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert925 gnd vdd FILL
XFILL_3__9735_ gnd vdd FILL
XFILL_3__6947_ gnd vdd FILL
XFILL_1__14729_ gnd vdd FILL
XFILL_4__15889_ gnd vdd FILL
XFILL_5_BUFX2_insert936 gnd vdd FILL
XFILL_0__16158_ gnd vdd FILL
XFILL_5_BUFX2_insert947 gnd vdd FILL
X_7516_ _7432_/A _8165_/CLK _9046_/R vdd _7434_/Y gnd vdd DFFSR
XFILL_1__8750_ gnd vdd FILL
XFILL_5_BUFX2_insert958 gnd vdd FILL
XFILL_5_BUFX2_insert969 gnd vdd FILL
X_8496_ _8496_/A _8496_/B gnd _8497_/C vdd NAND2X1
XFILL_3__16269_ gnd vdd FILL
XFILL_3__9666_ gnd vdd FILL
XFILL_0__15109_ gnd vdd FILL
XFILL_0__16089_ gnd vdd FILL
XFILL_3__6878_ gnd vdd FILL
XFILL_0__8908_ gnd vdd FILL
XFILL_1__7701_ gnd vdd FILL
X_7447_ _7447_/A gnd _7449_/A vdd INVX1
XFILL_3__8617_ gnd vdd FILL
XFILL_0__9888_ gnd vdd FILL
XSFILL33800x1050 gnd vdd FILL
XFILL_4__8390_ gnd vdd FILL
XFILL_3__9597_ gnd vdd FILL
XSFILL33800x35050 gnd vdd FILL
XFILL_0__8839_ gnd vdd FILL
XFILL_1__7632_ gnd vdd FILL
X_7378_ _7378_/A _7366_/B _7378_/C gnd _7412_/D vdd OAI21X1
XFILL_4__7341_ gnd vdd FILL
XFILL_6__8257_ gnd vdd FILL
X_9117_ _9117_/A gnd _9117_/Y vdd INVX1
XFILL_1__7563_ gnd vdd FILL
XFILL_3_BUFX2_insert104 gnd vdd FILL
XSFILL84040x72050 gnd vdd FILL
XFILL_6__7208_ gnd vdd FILL
XFILL_3__8479_ gnd vdd FILL
X_9048_ _9048_/Q _8151_/CLK _9048_/R vdd _9048_/D gnd vdd DFFSR
XFILL_4__9011_ gnd vdd FILL
XFILL_1__7494_ gnd vdd FILL
XCLKBUF1_insert1082 clk gnd CLKBUF1_insert220/A vdd CLKBUF1
XFILL_1__9233_ gnd vdd FILL
XFILL_2_BUFX2_insert804 gnd vdd FILL
XFILL_2_BUFX2_insert815 gnd vdd FILL
XFILL_2_BUFX2_insert826 gnd vdd FILL
X_11950_ _13196_/Q gnd _11952_/A vdd INVX1
XFILL_2_BUFX2_insert837 gnd vdd FILL
XFILL_1__9164_ gnd vdd FILL
XFILL112040x54050 gnd vdd FILL
XFILL_2_BUFX2_insert848 gnd vdd FILL
XFILL_2_BUFX2_insert859 gnd vdd FILL
XSFILL79400x59050 gnd vdd FILL
X_10901_ _10898_/Y _10929_/A gnd _16449_/A vdd NOR2X1
XFILL_0_BUFX2_insert70 gnd vdd FILL
XFILL_1__8115_ gnd vdd FILL
X_11881_ _11881_/A gnd _11883_/A vdd INVX1
XFILL_0_BUFX2_insert81 gnd vdd FILL
XFILL_0_BUFX2_insert92 gnd vdd FILL
XFILL_1__9095_ gnd vdd FILL
XFILL_4__9913_ gnd vdd FILL
X_13620_ _13456_/A gnd _13621_/B vdd INVX8
X_10832_ _14883_/A gnd _10834_/A vdd INVX1
XSFILL114600x68050 gnd vdd FILL
X_13551_ _13547_/Y _13551_/B gnd _13559_/A vdd NOR2X1
X_10763_ _10763_/A gnd _10763_/Y vdd INVX1
XBUFX2_insert803 _15091_/Y gnd _15863_/A vdd BUFX2
XBUFX2_insert814 _13329_/Y gnd _9014_/A vdd BUFX2
XBUFX2_insert825 _13287_/Y gnd _7425_/B vdd BUFX2
X_12502_ _12406_/A gnd _12504_/A vdd INVX1
XFILL_4__9775_ gnd vdd FILL
XFILL_4__6987_ gnd vdd FILL
XBUFX2_insert836 _13324_/Y gnd _8567_/B vdd BUFX2
XFILL_6_BUFX2_insert781 gnd vdd FILL
X_16270_ _7248_/A gnd _16270_/Y vdd INVX1
XFILL_2__7810_ gnd vdd FILL
XFILL_6_BUFX2_insert792 gnd vdd FILL
XBUFX2_insert847 _12375_/Y gnd _7445_/B vdd BUFX2
X_13482_ _15095_/A _14934_/B _14320_/C _15110_/C gnd _13482_/Y vdd OAI22X1
X_10694_ _10694_/A _10658_/B _10693_/Y gnd _10694_/Y vdd OAI21X1
XBUFX2_insert858 _13314_/Y gnd _8216_/A vdd BUFX2
XFILL_1__9997_ gnd vdd FILL
XFILL_4__8726_ gnd vdd FILL
X_15221_ _15036_/A _15014_/C _15220_/Y gnd _15382_/B vdd NOR3X1
XBUFX2_insert869 _13379_/Y gnd _14353_/A vdd BUFX2
X_12433_ _12107_/B gnd _12433_/Y vdd INVX1
XFILL_2__7741_ gnd vdd FILL
XFILL_5__7450_ gnd vdd FILL
XFILL_4__8657_ gnd vdd FILL
X_15152_ _13564_/Y _15795_/B _15152_/C gnd _15155_/A vdd OAI21X1
X_12364_ _12364_/A gnd _12364_/Y vdd INVX1
XFILL_4__7608_ gnd vdd FILL
XFILL_3__10280_ gnd vdd FILL
XFILL_2__7672_ gnd vdd FILL
XSFILL38600x27050 gnd vdd FILL
XFILL_1__8879_ gnd vdd FILL
XFILL112120x34050 gnd vdd FILL
X_14103_ _8931_/Q gnd _14104_/A vdd INVX1
XFILL_4__8588_ gnd vdd FILL
XFILL_5__7381_ gnd vdd FILL
X_11315_ _11544_/A _11531_/A _11529_/A gnd _11437_/C vdd AOI21X1
X_15083_ _16199_/C gnd _15696_/A vdd INVX2
XFILL_2__9411_ gnd vdd FILL
XFILL_1__10410_ gnd vdd FILL
X_12295_ _12216_/A gnd _12311_/C gnd _12298_/A vdd NAND3X1
XFILL_4__11570_ gnd vdd FILL
XFILL_5__9120_ gnd vdd FILL
XFILL_1__11390_ gnd vdd FILL
X_14034_ _14033_/Y _14636_/C gnd _14035_/C vdd NOR2X1
XFILL_4__10521_ gnd vdd FILL
X_11246_ _12242_/Y _12135_/Y gnd _11247_/B vdd XOR2X1
XFILL_5__12860_ gnd vdd FILL
XFILL_2__11700_ gnd vdd FILL
XFILL_2__9342_ gnd vdd FILL
XFILL_4__13240_ gnd vdd FILL
XSFILL33960x7050 gnd vdd FILL
XFILL_5__11811_ gnd vdd FILL
XFILL_4__10452_ gnd vdd FILL
X_11177_ _11176_/Y _11175_/Y gnd _11494_/A vdd NOR2X1
XFILL_2__9273_ gnd vdd FILL
XFILL_5__8002_ gnd vdd FILL
XFILL_2__11631_ gnd vdd FILL
XFILL_3__13970_ gnd vdd FILL
XFILL_4__9209_ gnd vdd FILL
XFILL_1__10272_ gnd vdd FILL
XFILL_0__13790_ gnd vdd FILL
XFILL_3_BUFX2_insert660 gnd vdd FILL
X_10128_ _10126_/Y _10127_/A _10128_/C gnd _10206_/D vdd OAI21X1
XFILL_3_BUFX2_insert671 gnd vdd FILL
XFILL_5__14530_ gnd vdd FILL
XSFILL69160x29050 gnd vdd FILL
X_15985_ _15187_/A _14562_/Y _15187_/C gnd _16005_/B vdd NOR3X1
XFILL_2__8224_ gnd vdd FILL
XFILL_1__12011_ gnd vdd FILL
XFILL_4__13171_ gnd vdd FILL
XFILL_3_BUFX2_insert682 gnd vdd FILL
XFILL_5__11742_ gnd vdd FILL
XFILL_4__10383_ gnd vdd FILL
XFILL_2__14350_ gnd vdd FILL
XFILL_0__12741_ gnd vdd FILL
XFILL_3_BUFX2_insert693 gnd vdd FILL
XFILL_2__11562_ gnd vdd FILL
X_10059_ _9985_/B _7243_/B gnd _10059_/Y vdd NAND2X1
X_14936_ _7413_/Q gnd _14937_/A vdd INVX1
XFILL_4__12122_ gnd vdd FILL
XFILL_2__13301_ gnd vdd FILL
XFILL_5__14461_ gnd vdd FILL
XFILL_3__15640_ gnd vdd FILL
XFILL_5__11673_ gnd vdd FILL
XSFILL104360x38050 gnd vdd FILL
XFILL_3__12852_ gnd vdd FILL
XFILL_2__10513_ gnd vdd FILL
XFILL_2__14281_ gnd vdd FILL
XFILL_5__16200_ gnd vdd FILL
XFILL_2__11493_ gnd vdd FILL
XFILL_0__15460_ gnd vdd FILL
XFILL_5__10624_ gnd vdd FILL
XFILL_0__7170_ gnd vdd FILL
XFILL_5__13412_ gnd vdd FILL
XFILL_6__15751_ gnd vdd FILL
X_14867_ _9843_/Q _14470_/B _14867_/C _9933_/A gnd _14867_/Y vdd AOI22X1
XFILL_2__16020_ gnd vdd FILL
XFILL_4__12053_ gnd vdd FILL
XFILL_2__7106_ gnd vdd FILL
XFILL_3__11803_ gnd vdd FILL
XFILL_2__13232_ gnd vdd FILL
XFILL_3__15571_ gnd vdd FILL
XFILL_5__14392_ gnd vdd FILL
XFILL_3__12783_ gnd vdd FILL
XFILL_2__10444_ gnd vdd FILL
XFILL_0__14411_ gnd vdd FILL
XFILL_2__8086_ gnd vdd FILL
XFILL_0__11623_ gnd vdd FILL
XFILL_0__15391_ gnd vdd FILL
XFILL_6__14702_ gnd vdd FILL
XFILL_5__8904_ gnd vdd FILL
XFILL_1__13962_ gnd vdd FILL
X_13818_ _13818_/A _7389_/Q _7901_/Q _13865_/B gnd _13826_/B vdd AOI22X1
XFILL_5__16131_ gnd vdd FILL
XFILL_4__11004_ gnd vdd FILL
XFILL_5__13343_ gnd vdd FILL
XFILL_5__10555_ gnd vdd FILL
XFILL_3__14522_ gnd vdd FILL
XFILL_5__9884_ gnd vdd FILL
XFILL_1__15701_ gnd vdd FILL
X_14798_ _8138_/A gnd _16194_/B vdd INVX1
XFILL_2__7037_ gnd vdd FILL
XFILL_3__11734_ gnd vdd FILL
XFILL112200x14050 gnd vdd FILL
XFILL_2__13163_ gnd vdd FILL
XFILL_0__14342_ gnd vdd FILL
XFILL_1__12913_ gnd vdd FILL
XFILL_2__10375_ gnd vdd FILL
XFILL_0__11554_ gnd vdd FILL
XFILL_5__8835_ gnd vdd FILL
XFILL_1__13893_ gnd vdd FILL
XFILL_5__13274_ gnd vdd FILL
X_13749_ _13749_/A _13749_/B gnd _13750_/C vdd NOR2X1
XFILL_4__15812_ gnd vdd FILL
XFILL_5__16062_ gnd vdd FILL
XFILL_6__11845_ gnd vdd FILL
XFILL_3__14453_ gnd vdd FILL
XFILL_5__10486_ gnd vdd FILL
XFILL_2__12114_ gnd vdd FILL
XFILL_0__10505_ gnd vdd FILL
XFILL_1__15632_ gnd vdd FILL
XFILL_3__7850_ gnd vdd FILL
XFILL_3__11665_ gnd vdd FILL
XFILL_1__12844_ gnd vdd FILL
XFILL_2__13094_ gnd vdd FILL
XFILL_0__14273_ gnd vdd FILL
XFILL_5__8766_ gnd vdd FILL
XFILL_5__15013_ gnd vdd FILL
XFILL_5__12225_ gnd vdd FILL
XFILL_0__11485_ gnd vdd FILL
XFILL_6__14564_ gnd vdd FILL
XFILL_3__13404_ gnd vdd FILL
XFILL_3__10616_ gnd vdd FILL
XFILL_4__15743_ gnd vdd FILL
XFILL_0__13224_ gnd vdd FILL
XFILL_0__16012_ gnd vdd FILL
XFILL_2__12045_ gnd vdd FILL
XFILL_3__14384_ gnd vdd FILL
XFILL_4__12955_ gnd vdd FILL
XFILL_5__7717_ gnd vdd FILL
XFILL_2__8988_ gnd vdd FILL
XFILL_0__10436_ gnd vdd FILL
XFILL_1__15563_ gnd vdd FILL
XFILL_3__11596_ gnd vdd FILL
XFILL_1__12775_ gnd vdd FILL
XFILL_0__9811_ gnd vdd FILL
X_15419_ _9105_/A gnd _15419_/Y vdd INVX1
XFILL_6__13515_ gnd vdd FILL
XFILL_0_BUFX2_insert550 gnd vdd FILL
XFILL_3__16123_ gnd vdd FILL
XFILL_0_BUFX2_insert561 gnd vdd FILL
X_8350_ _8315_/B _7838_/B gnd _8351_/C vdd NAND2X1
XFILL_5__8697_ gnd vdd FILL
XFILL_5__12156_ gnd vdd FILL
XFILL_3__13335_ gnd vdd FILL
XFILL_0_BUFX2_insert572 gnd vdd FILL
XFILL_4__11906_ gnd vdd FILL
X_16399_ _14713_/A gnd _16401_/A vdd INVX1
XFILL_3__9520_ gnd vdd FILL
XFILL_0_BUFX2_insert583 gnd vdd FILL
XSFILL109480x71050 gnd vdd FILL
XFILL_4__15674_ gnd vdd FILL
XFILL_4__12886_ gnd vdd FILL
XFILL_2__7939_ gnd vdd FILL
XFILL_1__14514_ gnd vdd FILL
XFILL_3__10547_ gnd vdd FILL
XFILL_0__13155_ gnd vdd FILL
XFILL_1__11726_ gnd vdd FILL
XFILL_0__10367_ gnd vdd FILL
XFILL_0_BUFX2_insert594 gnd vdd FILL
XFILL_5__11107_ gnd vdd FILL
XFILL_1__15494_ gnd vdd FILL
X_7301_ _7301_/A gnd _7303_/A vdd INVX1
XFILL_0__9742_ gnd vdd FILL
X_8281_ _8191_/A _8025_/CLK _8025_/R vdd _8281_/D gnd vdd DFFSR
XFILL_4__14625_ gnd vdd FILL
XFILL_5__12087_ gnd vdd FILL
XFILL_2__15804_ gnd vdd FILL
XFILL_3__16054_ gnd vdd FILL
XFILL_0__6954_ gnd vdd FILL
XFILL_4__11837_ gnd vdd FILL
XFILL_3__13266_ gnd vdd FILL
XFILL_0__12106_ gnd vdd FILL
XSFILL54040x51050 gnd vdd FILL
XFILL_1__14445_ gnd vdd FILL
XFILL_0__13086_ gnd vdd FILL
XFILL_2__13996_ gnd vdd FILL
XFILL_1__11657_ gnd vdd FILL
X_7232_ _7230_/Y _7184_/B _7232_/C gnd _7278_/D vdd OAI21X1
XFILL_5__15915_ gnd vdd FILL
XFILL_6__16165_ gnd vdd FILL
XFILL_5__7579_ gnd vdd FILL
XFILL_3__15005_ gnd vdd FILL
XFILL_0__10298_ gnd vdd FILL
XSFILL104440x18050 gnd vdd FILL
XFILL_5__11038_ gnd vdd FILL
XFILL_2__9609_ gnd vdd FILL
XFILL_6__13377_ gnd vdd FILL
XFILL_0__9673_ gnd vdd FILL
XFILL_3__12217_ gnd vdd FILL
XFILL_3__8402_ gnd vdd FILL
XFILL_4__14556_ gnd vdd FILL
XFILL_0__6885_ gnd vdd FILL
XFILL_4__11768_ gnd vdd FILL
XFILL_2__15735_ gnd vdd FILL
XFILL_3__9382_ gnd vdd FILL
XFILL_0__12037_ gnd vdd FILL
XSFILL8680x16050 gnd vdd FILL
XFILL_1__14376_ gnd vdd FILL
XFILL_1__11588_ gnd vdd FILL
XFILL_0__8624_ gnd vdd FILL
XFILL_5__15846_ gnd vdd FILL
X_7163_ _7161_/Y _7210_/A _7163_/C gnd _7255_/D vdd OAI21X1
XFILL_4__13507_ gnd vdd FILL
XFILL_3__8333_ gnd vdd FILL
XFILL_4__14487_ gnd vdd FILL
XFILL_3__12148_ gnd vdd FILL
XFILL_1__16115_ gnd vdd FILL
XFILL_1__13327_ gnd vdd FILL
XFILL_2__15666_ gnd vdd FILL
XFILL_1__10539_ gnd vdd FILL
XFILL_4__11699_ gnd vdd FILL
XFILL_5__9249_ gnd vdd FILL
XFILL_2__12878_ gnd vdd FILL
XFILL_4__16226_ gnd vdd FILL
XFILL_6__12259_ gnd vdd FILL
XFILL_4__13438_ gnd vdd FILL
X_7094_ _7095_/B _7094_/B gnd _7094_/Y vdd NAND2X1
XFILL_2__14617_ gnd vdd FILL
XFILL_5__15777_ gnd vdd FILL
XSFILL48920x31050 gnd vdd FILL
XFILL_1__16046_ gnd vdd FILL
XFILL_3__12079_ gnd vdd FILL
XFILL_5__12989_ gnd vdd FILL
XSFILL104440x2050 gnd vdd FILL
XFILL_2__11829_ gnd vdd FILL
XFILL_3__8264_ gnd vdd FILL
XFILL_1__13258_ gnd vdd FILL
XSFILL74200x64050 gnd vdd FILL
XFILL_2__15597_ gnd vdd FILL
XFILL_0__7506_ gnd vdd FILL
XFILL_0__13988_ gnd vdd FILL
XFILL_5__14728_ gnd vdd FILL
XFILL_0__8486_ gnd vdd FILL
XFILL_3__15907_ gnd vdd FILL
XFILL_4__13369_ gnd vdd FILL
XFILL_3__7215_ gnd vdd FILL
XFILL_4__16157_ gnd vdd FILL
XFILL_2__14548_ gnd vdd FILL
XFILL_1__12209_ gnd vdd FILL
XFILL_0__15727_ gnd vdd FILL
XFILL_3__8195_ gnd vdd FILL
XSFILL13640x17050 gnd vdd FILL
XFILL_0__7437_ gnd vdd FILL
XFILL_4__15108_ gnd vdd FILL
XFILL_4__16088_ gnd vdd FILL
XFILL_5__14659_ gnd vdd FILL
XFILL_3__15838_ gnd vdd FILL
XFILL_2__14479_ gnd vdd FILL
XFILL_0__15658_ gnd vdd FILL
X_9804_ _9804_/A _9737_/A _9804_/C gnd _9842_/D vdd OAI21X1
XSFILL109560x51050 gnd vdd FILL
XFILL_2__16218_ gnd vdd FILL
XFILL_4__15039_ gnd vdd FILL
XFILL_0__7368_ gnd vdd FILL
XFILL_3__7077_ gnd vdd FILL
XFILL_0__14609_ gnd vdd FILL
X_7996_ _7997_/B _8764_/B gnd _7997_/C vdd NAND2X1
XFILL_3__15769_ gnd vdd FILL
XSFILL38840x83050 gnd vdd FILL
XFILL_0__9107_ gnd vdd FILL
XFILL_5__16329_ gnd vdd FILL
XFILL_0__15589_ gnd vdd FILL
X_9735_ _9733_/Y _9770_/A _9735_/C gnd _9819_/D vdd OAI21X1
XFILL_0__7299_ gnd vdd FILL
X_6947_ _6947_/A gnd _6947_/Y vdd INVX1
XFILL_2__16149_ gnd vdd FILL
XFILL_4__6910_ gnd vdd FILL
XFILL_4__7890_ gnd vdd FILL
XFILL_0__9038_ gnd vdd FILL
XFILL_1__9920_ gnd vdd FILL
X_9666_ _9597_/A _8642_/B gnd _9666_/Y vdd NAND2X1
XFILL_4__6841_ gnd vdd FILL
X_6878_ _6878_/A gnd memoryWriteData[8] vdd BUFX2
XSFILL43960x74050 gnd vdd FILL
X_8617_ _8617_/A gnd _8619_/A vdd INVX1
XFILL_1__9851_ gnd vdd FILL
XFILL_5_BUFX2_insert700 gnd vdd FILL
XSFILL28760x8050 gnd vdd FILL
XFILL_5_BUFX2_insert711 gnd vdd FILL
X_9597_ _9597_/A _9597_/B gnd _9598_/C vdd NAND2X1
XFILL_5_BUFX2_insert722 gnd vdd FILL
XFILL_3__7979_ gnd vdd FILL
XSFILL18760x50050 gnd vdd FILL
XFILL_5_BUFX2_insert733 gnd vdd FILL
XFILL_5_BUFX2_insert744 gnd vdd FILL
XFILL_1__9782_ gnd vdd FILL
XFILL_4__8511_ gnd vdd FILL
XSFILL8600x60050 gnd vdd FILL
X_8548_ _8548_/Q _8161_/CLK _7140_/R vdd _8548_/D gnd vdd DFFSR
XSFILL44040x83050 gnd vdd FILL
XFILL_3__9718_ gnd vdd FILL
XFILL_5_BUFX2_insert755 gnd vdd FILL
XFILL_1__6994_ gnd vdd FILL
XFILL_5_BUFX2_insert766 gnd vdd FILL
XFILL_4__9491_ gnd vdd FILL
XFILL_5_BUFX2_insert777 gnd vdd FILL
XFILL_5_BUFX2_insert788 gnd vdd FILL
XFILL_1__8733_ gnd vdd FILL
XFILL_5_BUFX2_insert799 gnd vdd FILL
XFILL_3__9649_ gnd vdd FILL
X_8479_ _8479_/A _8469_/A _8479_/C gnd _8547_/D vdd OAI21X1
XFILL_4__8442_ gnd vdd FILL
XSFILL43960x2050 gnd vdd FILL
XFILL112040x49050 gnd vdd FILL
XSFILL23880x41050 gnd vdd FILL
XFILL_4__8373_ gnd vdd FILL
X_11100_ _11099_/Y gnd _11544_/A vdd INVX2
XFILL_1__7615_ gnd vdd FILL
X_12080_ _12072_/A _12812_/Q _12072_/C gnd _12082_/B vdd NAND3X1
XSFILL38920x63050 gnd vdd FILL
XFILL_4__7324_ gnd vdd FILL
XFILL_1__8595_ gnd vdd FILL
XFILL112440x70050 gnd vdd FILL
X_11031_ _12238_/Y _11031_/B gnd _11034_/C vdd NOR2X1
XFILL_1__7546_ gnd vdd FILL
XSFILL39000x72050 gnd vdd FILL
XSFILL89320x1050 gnd vdd FILL
XFILL_1__7477_ gnd vdd FILL
XFILL_2_BUFX2_insert601 gnd vdd FILL
XFILL_2_BUFX2_insert612 gnd vdd FILL
XFILL_4__7186_ gnd vdd FILL
XFILL_1__9216_ gnd vdd FILL
XFILL_2_BUFX2_insert623 gnd vdd FILL
X_15770_ _15770_/A _15769_/Y _15812_/C gnd _12875_/B vdd AOI21X1
XFILL_2_BUFX2_insert634 gnd vdd FILL
X_12982_ vdd _12982_/B gnd _12983_/C vdd NAND2X1
XFILL_2_BUFX2_insert645 gnd vdd FILL
XSFILL18840x30050 gnd vdd FILL
XFILL_2_BUFX2_insert656 gnd vdd FILL
X_14721_ _14721_/A _14719_/Y _14545_/B _14720_/Y gnd _14721_/Y vdd OAI22X1
X_11933_ _11934_/B _12388_/A gnd _11933_/Y vdd NAND2X1
XFILL_2_BUFX2_insert667 gnd vdd FILL
XFILL_1__9147_ gnd vdd FILL
XFILL_2_BUFX2_insert678 gnd vdd FILL
XFILL_2_BUFX2_insert689 gnd vdd FILL
XFILL_5__6950_ gnd vdd FILL
X_14652_ _10177_/A gnd _16069_/C vdd INVX1
X_11864_ _12105_/A _12485_/B gnd _11865_/B vdd NOR2X1
XFILL_1__9078_ gnd vdd FILL
X_13603_ _8153_/Q gnd _13603_/Y vdd INVX1
X_10815_ _10789_/B _8255_/B gnd _10816_/C vdd NAND2X1
XFILL_5_BUFX2_insert16 gnd vdd FILL
XFILL_5__6881_ gnd vdd FILL
XFILL112120x29050 gnd vdd FILL
XFILL_2__8911_ gnd vdd FILL
X_14583_ _14583_/A _14583_/B _13846_/A _14582_/Y gnd _14583_/Y vdd OAI22X1
XFILL_5_BUFX2_insert27 gnd vdd FILL
XFILL_2__10160_ gnd vdd FILL
X_11795_ _11794_/Y _11768_/B _11026_/C gnd _11795_/Y vdd AOI21X1
XFILL_5_BUFX2_insert38 gnd vdd FILL
XFILL_2__9891_ gnd vdd FILL
XFILL_5__8620_ gnd vdd FILL
XBUFX2_insert600 BUFX2_insert600/A gnd _8816_/R vdd BUFX2
XSFILL64040x14050 gnd vdd FILL
X_16322_ gnd gnd gnd _16323_/C vdd NAND2X1
XFILL_5_BUFX2_insert49 gnd vdd FILL
XBUFX2_insert611 _15035_/Y gnd _15550_/A vdd BUFX2
XFILL_1__10890_ gnd vdd FILL
XBUFX2_insert622 _12363_/Y gnd _7177_/B vdd BUFX2
XFILL_6__11630_ gnd vdd FILL
X_13534_ _8408_/Q gnd _13534_/Y vdd INVX1
XFILL_5__10271_ gnd vdd FILL
X_10746_ _10809_/A _8314_/B gnd _10747_/C vdd NAND2X1
XFILL_2__8842_ gnd vdd FILL
XBUFX2_insert633 _12354_/Y gnd _9344_/B vdd BUFX2
XFILL_3__11450_ gnd vdd FILL
XBUFX2_insert644 _13424_/Y gnd _13860_/B vdd BUFX2
XBUFX2_insert655 _12429_/Y gnd _7883_/B vdd BUFX2
XFILL_5__12010_ gnd vdd FILL
XFILL_0__11270_ gnd vdd FILL
XBUFX2_insert666 _12345_/Y gnd _8183_/A vdd BUFX2
XFILL_4__9758_ gnd vdd FILL
X_16253_ _15225_/A _7632_/A _7504_/A _15383_/D gnd _16253_/Y vdd AOI22X1
XFILL_4__12740_ gnd vdd FILL
X_13465_ _13423_/A _13718_/B _13465_/C gnd _13465_/Y vdd NAND3X1
XFILL_3__10401_ gnd vdd FILL
XBUFX2_insert677 _13541_/Y gnd _13864_/C vdd BUFX2
X_10677_ _10677_/A gnd _10677_/Y vdd INVX1
XSFILL89240x80050 gnd vdd FILL
XFILL_5__7502_ gnd vdd FILL
XFILL_2__8773_ gnd vdd FILL
XBUFX2_insert688 _13459_/Y gnd _14545_/B vdd BUFX2
XFILL_3__11381_ gnd vdd FILL
X_15204_ _15204_/A _13607_/Y _13588_/Y _15677_/D gnd _15205_/B vdd OAI22X1
XFILL_4__8709_ gnd vdd FILL
XBUFX2_insert699 _12420_/Y gnd _9794_/B vdd BUFX2
XFILL_6__10512_ gnd vdd FILL
X_12416_ _12380_/A _12639_/A gnd _12417_/C vdd NAND2X1
XFILL_5__8482_ gnd vdd FILL
X_16184_ _16184_/A _16184_/B gnd _16190_/B vdd NOR2X1
XFILL_3__13120_ gnd vdd FILL
X_13396_ _7638_/Q gnd _13399_/D vdd INVX1
XFILL_2__7724_ gnd vdd FILL
XFILL_6__11492_ gnd vdd FILL
XSFILL3720x83050 gnd vdd FILL
XFILL_2__13850_ gnd vdd FILL
XFILL_1__11511_ gnd vdd FILL
XFILL_0__10152_ gnd vdd FILL
XSFILL68920x79050 gnd vdd FILL
XFILL_5__7433_ gnd vdd FILL
XFILL_1__12491_ gnd vdd FILL
XSFILL84200x27050 gnd vdd FILL
X_15135_ _15135_/A _15135_/B gnd _15136_/C vdd NOR2X1
X_12347_ _12359_/A _12570_/A gnd _12348_/C vdd NAND2X1
XFILL_4__14410_ gnd vdd FILL
XFILL_4__11622_ gnd vdd FILL
XFILL_4__15390_ gnd vdd FILL
XFILL_5__13961_ gnd vdd FILL
XFILL_1__14230_ gnd vdd FILL
XFILL_3__10263_ gnd vdd FILL
XFILL_1__11442_ gnd vdd FILL
XSFILL94360x71050 gnd vdd FILL
XFILL_2__13781_ gnd vdd FILL
XFILL_5__15700_ gnd vdd FILL
XFILL_0__14960_ gnd vdd FILL
XFILL_5__7364_ gnd vdd FILL
XFILL_2__10993_ gnd vdd FILL
XFILL_5__12912_ gnd vdd FILL
XFILL_3__12002_ gnd vdd FILL
X_15066_ _16228_/B _15066_/B _15392_/B _13410_/Y gnd _15067_/A vdd OAI22X1
XFILL_4__14341_ gnd vdd FILL
XFILL_2__15520_ gnd vdd FILL
X_12278_ _12278_/A _12278_/B _12278_/C gnd _12278_/Y vdd NAND3X1
XFILL_4__11553_ gnd vdd FILL
XFILL_2__12732_ gnd vdd FILL
XFILL_5__9103_ gnd vdd FILL
XFILL_5__13892_ gnd vdd FILL
XFILL_2__7586_ gnd vdd FILL
XFILL_1__14161_ gnd vdd FILL
XFILL_3__10194_ gnd vdd FILL
XFILL_0__13911_ gnd vdd FILL
XFILL_1__11373_ gnd vdd FILL
X_14017_ _8599_/A gnd _14018_/B vdd INVX1
XFILL_5__7295_ gnd vdd FILL
XFILL_4__10504_ gnd vdd FILL
XFILL_5__15631_ gnd vdd FILL
XFILL_0__14891_ gnd vdd FILL
X_11229_ _10989_/Y _11484_/B _11349_/B _10988_/Y gnd _11229_/Y vdd OAI22X1
XFILL_5__12843_ gnd vdd FILL
XFILL_4__14272_ gnd vdd FILL
XFILL_1__13112_ gnd vdd FILL
XFILL_2__15451_ gnd vdd FILL
XFILL_4__11484_ gnd vdd FILL
XFILL_1__10324_ gnd vdd FILL
XFILL_5__9034_ gnd vdd FILL
XFILL_1__14092_ gnd vdd FILL
XFILL_0__13842_ gnd vdd FILL
XFILL_4__13223_ gnd vdd FILL
XFILL_4__16011_ gnd vdd FILL
XFILL_6__12044_ gnd vdd FILL
XFILL_0__8340_ gnd vdd FILL
XFILL_5__15562_ gnd vdd FILL
XFILL_2__14402_ gnd vdd FILL
XFILL_4__10435_ gnd vdd FILL
XFILL_5__12774_ gnd vdd FILL
XSFILL74120x79050 gnd vdd FILL
XFILL_2__9256_ gnd vdd FILL
XFILL_3__13953_ gnd vdd FILL
XFILL_2__11614_ gnd vdd FILL
XFILL_1__13043_ gnd vdd FILL
XFILL_1__10255_ gnd vdd FILL
XFILL_2__15382_ gnd vdd FILL
XFILL_2__12594_ gnd vdd FILL
XFILL_3_BUFX2_insert490 gnd vdd FILL
XFILL_0__13773_ gnd vdd FILL
XFILL_5__14513_ gnd vdd FILL
XFILL_2__8207_ gnd vdd FILL
XFILL_0__8271_ gnd vdd FILL
XFILL_4__13154_ gnd vdd FILL
XFILL_3__12904_ gnd vdd FILL
XFILL_5__11725_ gnd vdd FILL
X_15968_ _15968_/A _15968_/B _15651_/C gnd _12890_/B vdd AOI21X1
XFILL_2__14333_ gnd vdd FILL
XFILL_4__10366_ gnd vdd FILL
XFILL_5__15493_ gnd vdd FILL
XSFILL49720x74050 gnd vdd FILL
XFILL_3__13884_ gnd vdd FILL
XFILL_0__15512_ gnd vdd FILL
XFILL_2__11545_ gnd vdd FILL
XFILL_0__12724_ gnd vdd FILL
XFILL_1__10186_ gnd vdd FILL
XFILL_0__7222_ gnd vdd FILL
XSFILL89320x60050 gnd vdd FILL
XFILL_4__12105_ gnd vdd FILL
XSFILL53960x37050 gnd vdd FILL
XFILL_5__14444_ gnd vdd FILL
X_14919_ _10192_/A gnd _14919_/Y vdd INVX1
X_15899_ _15899_/A _15899_/B _15899_/C _15899_/D gnd _15901_/A vdd OAI22X1
XFILL_3__15623_ gnd vdd FILL
XFILL_3__12835_ gnd vdd FILL
XFILL_4__13085_ gnd vdd FILL
XFILL_2__8138_ gnd vdd FILL
X_7850_ _7800_/B _9258_/B gnd _7850_/Y vdd NAND2X1
XFILL_5__11656_ gnd vdd FILL
XFILL_2__14264_ gnd vdd FILL
XFILL_4__10297_ gnd vdd FILL
XFILL_0__12655_ gnd vdd FILL
XSFILL89480x7050 gnd vdd FILL
XFILL_2__11476_ gnd vdd FILL
XFILL_0__15443_ gnd vdd FILL
XFILL_1__14994_ gnd vdd FILL
XFILL_5__9936_ gnd vdd FILL
XFILL_2__16003_ gnd vdd FILL
XFILL_4__12036_ gnd vdd FILL
XSFILL28760x13050 gnd vdd FILL
XFILL_2__13215_ gnd vdd FILL
XFILL_3__15554_ gnd vdd FILL
XFILL_5__14375_ gnd vdd FILL
XFILL_5__11587_ gnd vdd FILL
XFILL_3__12766_ gnd vdd FILL
X_7781_ _7781_/Q _7781_/CLK _8025_/R vdd _7781_/D gnd vdd DFFSR
XFILL_2__10427_ gnd vdd FILL
XFILL_3__8951_ gnd vdd FILL
XFILL_2__8069_ gnd vdd FILL
XFILL_2__14195_ gnd vdd FILL
XSFILL54040x46050 gnd vdd FILL
XFILL_0__11606_ gnd vdd FILL
XFILL_1__13945_ gnd vdd FILL
XFILL_0__12586_ gnd vdd FILL
XFILL_0__15374_ gnd vdd FILL
XFILL_5__16114_ gnd vdd FILL
XFILL_6__8660_ gnd vdd FILL
XFILL_5__13326_ gnd vdd FILL
XFILL_5__9867_ gnd vdd FILL
XSFILL94440x51050 gnd vdd FILL
X_9520_ _9529_/A _8496_/B gnd _9521_/C vdd NAND2X1
XFILL_3__14505_ gnd vdd FILL
XFILL_6__12877_ gnd vdd FILL
XFILL_0__7084_ gnd vdd FILL
XFILL_3__11717_ gnd vdd FILL
XFILL_5__10538_ gnd vdd FILL
XFILL_2__13146_ gnd vdd FILL
XFILL_3__15485_ gnd vdd FILL
XFILL_6__7611_ gnd vdd FILL
XFILL_3__12697_ gnd vdd FILL
XFILL_2__10358_ gnd vdd FILL
XFILL_0__14325_ gnd vdd FILL
XFILL_3__8882_ gnd vdd FILL
XFILL_0__11537_ gnd vdd FILL
XFILL_1__13876_ gnd vdd FILL
XFILL_5__16045_ gnd vdd FILL
XFILL_5__13257_ gnd vdd FILL
X_9451_ _9451_/Q _7389_/CLK _7531_/R vdd _9399_/Y gnd vdd DFFSR
XFILL_5__9798_ gnd vdd FILL
XFILL_3__14436_ gnd vdd FILL
XFILL_1__15615_ gnd vdd FILL
XFILL_3__7833_ gnd vdd FILL
XFILL_3__11648_ gnd vdd FILL
XFILL_0__14256_ gnd vdd FILL
XFILL_4__13987_ gnd vdd FILL
XFILL_1__12827_ gnd vdd FILL
XFILL_2__10289_ gnd vdd FILL
XFILL_0__11468_ gnd vdd FILL
XFILL_5__8749_ gnd vdd FILL
XFILL_5__12208_ gnd vdd FILL
X_8402_ _8400_/Y _8345_/B _8401_/Y gnd _8436_/D vdd OAI21X1
XFILL_4__15726_ gnd vdd FILL
X_9382_ _9382_/A gnd _9382_/Y vdd INVX1
XFILL_2__12028_ gnd vdd FILL
XFILL_3__14367_ gnd vdd FILL
XSFILL48920x26050 gnd vdd FILL
XFILL_0__13207_ gnd vdd FILL
XSFILL18680x65050 gnd vdd FILL
XFILL_1__15546_ gnd vdd FILL
XFILL_3__7764_ gnd vdd FILL
XFILL_0__10419_ gnd vdd FILL
XFILL_3__11579_ gnd vdd FILL
XFILL_1__12758_ gnd vdd FILL
XFILL_0__14187_ gnd vdd FILL
XFILL_0_BUFX2_insert380 gnd vdd FILL
XSFILL74200x59050 gnd vdd FILL
XFILL_0_BUFX2_insert391 gnd vdd FILL
XFILL_0__11399_ gnd vdd FILL
X_8333_ _8333_/A _8333_/B _8332_/Y gnd _8333_/Y vdd OAI21X1
XFILL_3__13318_ gnd vdd FILL
XFILL_5__12139_ gnd vdd FILL
XFILL_3__16106_ gnd vdd FILL
XFILL_3__9503_ gnd vdd FILL
XFILL_4__15657_ gnd vdd FILL
XFILL_0__7986_ gnd vdd FILL
XFILL_4__12869_ gnd vdd FILL
XFILL_4_BUFX2_insert707 gnd vdd FILL
XFILL_0__13138_ gnd vdd FILL
XFILL_3__14298_ gnd vdd FILL
XFILL_1__11709_ gnd vdd FILL
XFILL_3__7695_ gnd vdd FILL
XFILL_6__16217_ gnd vdd FILL
XFILL_4_BUFX2_insert718 gnd vdd FILL
XFILL_1__15477_ gnd vdd FILL
XFILL_4_BUFX2_insert729 gnd vdd FILL
XFILL_0__9725_ gnd vdd FILL
XFILL_3__16037_ gnd vdd FILL
XFILL_4__14608_ gnd vdd FILL
XFILL_0__6937_ gnd vdd FILL
X_8264_ _8187_/B _8008_/B gnd _8265_/C vdd NAND2X1
XFILL_3__13249_ gnd vdd FILL
XSFILL89400x40050 gnd vdd FILL
XFILL_4__15588_ gnd vdd FILL
XFILL_1__14428_ gnd vdd FILL
XFILL_2__13979_ gnd vdd FILL
XSFILL109560x46050 gnd vdd FILL
XFILL_0__9656_ gnd vdd FILL
X_7215_ _7273_/Q gnd _7217_/A vdd INVX1
X_8195_ _8246_/A _8195_/B gnd _8196_/C vdd NAND2X1
XFILL_4__14539_ gnd vdd FILL
XFILL_0__6868_ gnd vdd FILL
XFILL_2__15718_ gnd vdd FILL
XFILL_3__9365_ gnd vdd FILL
XFILL_1__14359_ gnd vdd FILL
XFILL_0__8607_ gnd vdd FILL
XFILL_5__15829_ gnd vdd FILL
X_7146_ _7090_/A _7786_/CLK _7153_/R vdd _7146_/D gnd vdd DFFSR
XFILL_1__8380_ gnd vdd FILL
XFILL_3__8316_ gnd vdd FILL
XFILL_2__15649_ gnd vdd FILL
XFILL_3__9296_ gnd vdd FILL
XFILL_4__16209_ gnd vdd FILL
XFILL_1__7331_ gnd vdd FILL
X_7077_ _7075_/Y _7055_/A _7077_/C gnd _7077_/Y vdd OAI21X1
XFILL_4__7040_ gnd vdd FILL
XFILL_3__8247_ gnd vdd FILL
XFILL_1__16029_ gnd vdd FILL
XFILL_5_BUFX2_insert1070 gnd vdd FILL
XSFILL43960x69050 gnd vdd FILL
XFILL_5_BUFX2_insert1092 gnd vdd FILL
XFILL_0__8469_ gnd vdd FILL
XFILL_1__9001_ gnd vdd FILL
XSFILL18760x45050 gnd vdd FILL
XSFILL8600x55050 gnd vdd FILL
XFILL_1__7193_ gnd vdd FILL
XSFILL44040x78050 gnd vdd FILL
XFILL_1_BUFX2_insert608 gnd vdd FILL
XFILL_4__8991_ gnd vdd FILL
XFILL_1_BUFX2_insert619 gnd vdd FILL
XSFILL99240x43050 gnd vdd FILL
XFILL_4__7942_ gnd vdd FILL
X_7979_ _7979_/A _7931_/B _7978_/Y gnd _7979_/Y vdd OAI21X1
X_9718_ _9718_/A gnd _9718_/Y vdd INVX1
XSFILL23880x36050 gnd vdd FILL
X_10600_ _15806_/A _7912_/CLK _7911_/R vdd _10600_/D gnd vdd DFFSR
XFILL_4__7873_ gnd vdd FILL
XSFILL63480x22050 gnd vdd FILL
X_11580_ _11580_/A gnd _12069_/A vdd INVX1
XFILL_1__9903_ gnd vdd FILL
X_9649_ _9647_/Y _9625_/B _9649_/C gnd _9705_/D vdd OAI21X1
XFILL_6__8789_ gnd vdd FILL
XFILL_4__9612_ gnd vdd FILL
XFILL112440x65050 gnd vdd FILL
X_10531_ _10531_/A gnd _10531_/Y vdd INVX1
XFILL_5_BUFX2_insert530 gnd vdd FILL
XSFILL39560x24050 gnd vdd FILL
XFILL_4__9543_ gnd vdd FILL
XFILL_5_BUFX2_insert541 gnd vdd FILL
XSFILL79160x10050 gnd vdd FILL
XFILL_5_BUFX2_insert552 gnd vdd FILL
X_13250_ _13231_/A _13302_/C gnd _13311_/A vdd NAND2X1
XFILL_5_BUFX2_insert563 gnd vdd FILL
X_10462_ _10462_/Q _9817_/CLK _7150_/R vdd _10462_/D gnd vdd DFFSR
XSFILL39000x67050 gnd vdd FILL
XFILL_3_BUFX2_insert0 gnd vdd FILL
XFILL_1__9765_ gnd vdd FILL
XFILL_5_BUFX2_insert574 gnd vdd FILL
XFILL_5_BUFX2_insert585 gnd vdd FILL
XFILL_1__6977_ gnd vdd FILL
XFILL_4__9474_ gnd vdd FILL
XFILL_5_BUFX2_insert596 gnd vdd FILL
X_12201_ _12201_/A _12201_/B _12201_/C gnd _12201_/Y vdd OAI21X1
XFILL_1__8716_ gnd vdd FILL
X_13181_ _13097_/A _9060_/CLK _9060_/R vdd _13181_/D gnd vdd DFFSR
X_10393_ _10393_/A _10372_/B _10393_/C gnd _10465_/D vdd OAI21X1
X_12132_ _12132_/A _12122_/A _12131_/Y gnd _11030_/A vdd OAI21X1
XSFILL114600x81050 gnd vdd FILL
XFILL_2__7440_ gnd vdd FILL
XFILL_1__8647_ gnd vdd FILL
XFILL_4__8356_ gnd vdd FILL
XFILL_2_CLKBUF1_insert111 gnd vdd FILL
XSFILL84520x63050 gnd vdd FILL
XFILL_2_CLKBUF1_insert122 gnd vdd FILL
X_12063_ _11987_/A _12496_/A _12059_/C gnd _12066_/A vdd NAND3X1
XSFILL99320x23050 gnd vdd FILL
XSFILL69080x62050 gnd vdd FILL
XFILL_2_CLKBUF1_insert133 gnd vdd FILL
XFILL_2_CLKBUF1_insert144 gnd vdd FILL
XFILL_2__7371_ gnd vdd FILL
XFILL_4__7307_ gnd vdd FILL
XFILL_1__8578_ gnd vdd FILL
XFILL_2_CLKBUF1_insert155 gnd vdd FILL
XFILL_5__7080_ gnd vdd FILL
XFILL_2_CLKBUF1_insert166 gnd vdd FILL
X_11014_ _12226_/Y _11013_/B gnd _11015_/A vdd OR2X2
XFILL_2__9110_ gnd vdd FILL
XFILL_2_CLKBUF1_insert177 gnd vdd FILL
XFILL_2_CLKBUF1_insert188 gnd vdd FILL
XSFILL99480x2050 gnd vdd FILL
XFILL_2_CLKBUF1_insert199 gnd vdd FILL
XFILL_4__7238_ gnd vdd FILL
X_15822_ _15175_/B _15822_/B _14358_/A _15357_/B gnd _15822_/Y vdd AOI22X1
XFILL_2__9041_ gnd vdd FILL
XFILL_3__10950_ gnd vdd FILL
XFILL_1__10040_ gnd vdd FILL
XFILL_2_BUFX2_insert420 gnd vdd FILL
XFILL_2_BUFX2_insert431 gnd vdd FILL
XFILL_4__7169_ gnd vdd FILL
XFILL_2_BUFX2_insert442 gnd vdd FILL
XFILL_0__10770_ gnd vdd FILL
XSFILL23800x80050 gnd vdd FILL
XFILL_2_BUFX2_insert453 gnd vdd FILL
XFILL_5__11510_ gnd vdd FILL
X_15753_ _15752_/Y _15753_/B gnd _15758_/A vdd NOR2X1
XFILL_4__10151_ gnd vdd FILL
X_12965_ _12963_/Y vdd _12965_/C gnd _13051_/D vdd OAI21X1
XFILL_5__12490_ gnd vdd FILL
XFILL_2_BUFX2_insert464 gnd vdd FILL
XFILL_2__11330_ gnd vdd FILL
XFILL_2_BUFX2_insert475 gnd vdd FILL
XFILL_3__10881_ gnd vdd FILL
XFILL_2_BUFX2_insert486 gnd vdd FILL
X_11916_ _11916_/A _11921_/A _11916_/C gnd _6847_/A vdd OAI21X1
X_14704_ _8304_/Q gnd _16117_/D vdd INVX1
XFILL_5__7982_ gnd vdd FILL
XFILL_2_BUFX2_insert497 gnd vdd FILL
XFILL_5__11441_ gnd vdd FILL
XFILL_3__12620_ gnd vdd FILL
X_15684_ _15684_/A _15684_/B gnd _15689_/A vdd NOR2X1
X_12896_ vdd _12896_/B gnd _12897_/C vdd NAND2X1
XSFILL3720x78050 gnd vdd FILL
XFILL_0__12440_ gnd vdd FILL
XFILL_2__11261_ gnd vdd FILL
XFILL_5__6933_ gnd vdd FILL
XFILL_5__9721_ gnd vdd FILL
X_14635_ _9198_/Q gnd _14635_/Y vdd INVX1
XFILL_1__11991_ gnd vdd FILL
XFILL_2__13000_ gnd vdd FILL
XFILL_5__14160_ gnd vdd FILL
XFILL_4__13910_ gnd vdd FILL
X_11847_ _12218_/Y _12117_/Y gnd _11848_/D vdd NOR2X1
XFILL_5__11372_ gnd vdd FILL
XFILL_1__13730_ gnd vdd FILL
XFILL_2__11192_ gnd vdd FILL
XFILL_4__14890_ gnd vdd FILL
XFILL_1__10942_ gnd vdd FILL
XSFILL94360x66050 gnd vdd FILL
XFILL_0__12371_ gnd vdd FILL
XFILL_5__6864_ gnd vdd FILL
XFILL_5__13111_ gnd vdd FILL
XFILL_5__10323_ gnd vdd FILL
XFILL_5__9652_ gnd vdd FILL
XSFILL68520x76050 gnd vdd FILL
X_14566_ _8173_/Q gnd _14566_/Y vdd INVX1
XFILL_5__14091_ gnd vdd FILL
XFILL_3__11502_ gnd vdd FILL
XFILL_4__13841_ gnd vdd FILL
XFILL_0__14110_ gnd vdd FILL
XFILL_3__15270_ gnd vdd FILL
X_11778_ _11776_/A _11778_/B _11777_/Y gnd _11778_/Y vdd OAI21X1
XFILL_3__12482_ gnd vdd FILL
XFILL_2__9874_ gnd vdd FILL
XFILL_2__10143_ gnd vdd FILL
XBUFX2_insert430 _13326_/Y gnd _8698_/A vdd BUFX2
XFILL_0__11322_ gnd vdd FILL
XFILL_1__13661_ gnd vdd FILL
XFILL_5__8603_ gnd vdd FILL
XFILL_0__15090_ gnd vdd FILL
XBUFX2_insert441 _15086_/Y gnd _15087_/B vdd BUFX2
XSFILL69160x42050 gnd vdd FILL
XFILL_1__10873_ gnd vdd FILL
X_16305_ _16305_/A gnd _16306_/B vdd INVX1
X_13517_ _13517_/A _14317_/C _14768_/D _13517_/D gnd _13518_/B vdd OAI22X1
XFILL_5__10254_ gnd vdd FILL
XFILL_3__14221_ gnd vdd FILL
X_10729_ _10671_/A _7916_/CLK _9964_/R vdd _10729_/D gnd vdd DFFSR
XBUFX2_insert452 _13276_/Y gnd _7166_/B vdd BUFX2
XFILL_5__13042_ gnd vdd FILL
XFILL_6__12593_ gnd vdd FILL
XFILL_1__15400_ gnd vdd FILL
X_14497_ _14496_/Y _14497_/B gnd _14498_/A vdd NOR2X1
XBUFX2_insert463 _15044_/Y gnd _15045_/D vdd BUFX2
XFILL_3__11433_ gnd vdd FILL
XFILL_2__8825_ gnd vdd FILL
XFILL_1__12612_ gnd vdd FILL
XFILL_4__13772_ gnd vdd FILL
XFILL_0__14041_ gnd vdd FILL
XFILL_2__14951_ gnd vdd FILL
XBUFX2_insert474 _15041_/Y gnd _16141_/C vdd BUFX2
XFILL_1__16380_ gnd vdd FILL
XFILL_0__11253_ gnd vdd FILL
XBUFX2_insert485 _12372_/Y gnd _8466_/B vdd BUFX2
XBUFX2_insert496 BUFX2_insert496/A gnd _8424_/R vdd BUFX2
XFILL_1__13592_ gnd vdd FILL
X_16236_ _16236_/A _16236_/B gnd _16242_/A vdd NOR2X1
X_13448_ _13423_/A _13418_/A _13423_/B gnd _14200_/C vdd NAND3X1
XFILL_0__7840_ gnd vdd FILL
XFILL_4__15511_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1078 gnd vdd FILL
XFILL_4__12723_ gnd vdd FILL
XFILL_3__14152_ gnd vdd FILL
XSFILL104360x51050 gnd vdd FILL
XFILL_5__10185_ gnd vdd FILL
XFILL_2__13902_ gnd vdd FILL
XFILL_1__15331_ gnd vdd FILL
XFILL_2__8756_ gnd vdd FILL
XFILL_3__11364_ gnd vdd FILL
XFILL_2__14882_ gnd vdd FILL
XFILL_0__11184_ gnd vdd FILL
XFILL_5__8465_ gnd vdd FILL
XFILL_3__13103_ gnd vdd FILL
X_16167_ _7114_/A gnd _16168_/B vdd INVX1
XSFILL74280x33050 gnd vdd FILL
XFILL_3__10315_ gnd vdd FILL
XFILL_2__7707_ gnd vdd FILL
X_13379_ _13843_/C gnd _13379_/Y vdd INVX8
XFILL_4__15442_ gnd vdd FILL
XFILL_4__12654_ gnd vdd FILL
XFILL_2__13833_ gnd vdd FILL
XFILL_5__14993_ gnd vdd FILL
XFILL_3__14083_ gnd vdd FILL
XFILL_6__16002_ gnd vdd FILL
XFILL_5__7416_ gnd vdd FILL
XFILL_0__10135_ gnd vdd FILL
XFILL_3__7480_ gnd vdd FILL
XFILL_3__11295_ gnd vdd FILL
XFILL_1__15262_ gnd vdd FILL
XFILL_6__13214_ gnd vdd FILL
XFILL_0__9510_ gnd vdd FILL
XFILL_1__12474_ gnd vdd FILL
X_15118_ _16301_/A _15116_/Y _15117_/Y _15761_/D gnd _15118_/Y vdd OAI22X1
XFILL_0__15992_ gnd vdd FILL
XFILL_5__8396_ gnd vdd FILL
X_16098_ _15351_/A _14720_/Y _16098_/C _15351_/D gnd _16100_/B vdd OAI22X1
XFILL_3__13034_ gnd vdd FILL
XFILL_4__11605_ gnd vdd FILL
XFILL_5__13944_ gnd vdd FILL
XFILL_4__12585_ gnd vdd FILL
XFILL_1__14213_ gnd vdd FILL
XFILL_4__15373_ gnd vdd FILL
XFILL_3__10246_ gnd vdd FILL
XFILL_2__13764_ gnd vdd FILL
XFILL_1__11425_ gnd vdd FILL
XFILL_2__10976_ gnd vdd FILL
XFILL_1__15193_ gnd vdd FILL
XFILL_0__14943_ gnd vdd FILL
X_7000_ _6908_/A _7640_/CLK _7000_/R vdd _6910_/Y gnd vdd DFFSR
XFILL_0__10066_ gnd vdd FILL
XFILL_5__7347_ gnd vdd FILL
X_15049_ _15045_/Y _15048_/Y gnd _15058_/B vdd NOR2X1
XFILL_2__15503_ gnd vdd FILL
XFILL_4__14324_ gnd vdd FILL
XFILL_4__11536_ gnd vdd FILL
XFILL_2__12715_ gnd vdd FILL
XFILL_5__13875_ gnd vdd FILL
XFILL_3__9150_ gnd vdd FILL
XFILL_1__14144_ gnd vdd FILL
XFILL_1_BUFX2_insert14 gnd vdd FILL
XFILL_3__10177_ gnd vdd FILL
XFILL_2__7569_ gnd vdd FILL
XFILL_1__11356_ gnd vdd FILL
XFILL_2__13695_ gnd vdd FILL
XFILL_1_BUFX2_insert25 gnd vdd FILL
XFILL_0__14874_ gnd vdd FILL
XFILL_5__15614_ gnd vdd FILL
XFILL_1_BUFX2_insert36 gnd vdd FILL
XFILL_6_BUFX2_insert4 gnd vdd FILL
XFILL_0__9372_ gnd vdd FILL
XFILL_1_BUFX2_insert47 gnd vdd FILL
XFILL_3__8101_ gnd vdd FILL
XFILL_5__12826_ gnd vdd FILL
XFILL_4__14255_ gnd vdd FILL
XSFILL94440x46050 gnd vdd FILL
XFILL_2__15434_ gnd vdd FILL
XFILL_4__11467_ gnd vdd FILL
XFILL_2__12646_ gnd vdd FILL
XFILL_5__9017_ gnd vdd FILL
XFILL_1__10307_ gnd vdd FILL
XFILL_1_BUFX2_insert58 gnd vdd FILL
XFILL_3__9081_ gnd vdd FILL
XFILL_0__13825_ gnd vdd FILL
XFILL_3__14985_ gnd vdd FILL
XFILL_1_BUFX2_insert69 gnd vdd FILL
XFILL_1__14075_ gnd vdd FILL
XFILL_1__11287_ gnd vdd FILL
XFILL_0__8323_ gnd vdd FILL
XFILL_5__15545_ gnd vdd FILL
XFILL_4__10418_ gnd vdd FILL
XFILL_4__14186_ gnd vdd FILL
XFILL_5__12757_ gnd vdd FILL
X_8951_ _8951_/A _8996_/A gnd _8952_/C vdd NAND2X1
XFILL_2__9239_ gnd vdd FILL
XFILL_2__15365_ gnd vdd FILL
XFILL_1__13026_ gnd vdd FILL
XFILL_4__11398_ gnd vdd FILL
XFILL_3__13936_ gnd vdd FILL
XFILL_1__10238_ gnd vdd FILL
XFILL_2__12577_ gnd vdd FILL
XFILL_0__13756_ gnd vdd FILL
XFILL_0__10968_ gnd vdd FILL
XFILL_0__8254_ gnd vdd FILL
X_7902_ _7902_/Q _7902_/CLK _9566_/R vdd _7824_/Y gnd vdd DFFSR
XFILL_4__13137_ gnd vdd FILL
XFILL_5__11708_ gnd vdd FILL
XFILL_2__14316_ gnd vdd FILL
XFILL_5__15476_ gnd vdd FILL
XFILL_2__11528_ gnd vdd FILL
X_8882_ _8938_/Q gnd _8884_/A vdd INVX1
XFILL_3__13867_ gnd vdd FILL
XFILL_0__12707_ gnd vdd FILL
XFILL_1__10169_ gnd vdd FILL
XFILL_2__15296_ gnd vdd FILL
XFILL_0__7205_ gnd vdd FILL
XSFILL104440x31050 gnd vdd FILL
XFILL_0__10899_ gnd vdd FILL
XFILL_0__13687_ gnd vdd FILL
XFILL_5__14427_ gnd vdd FILL
X_7833_ _7833_/A _7821_/B _7833_/C gnd _7833_/Y vdd OAI21X1
XFILL_5__11639_ gnd vdd FILL
XFILL_3__15606_ gnd vdd FILL
XFILL_0__8185_ gnd vdd FILL
XFILL_2__14247_ gnd vdd FILL
XFILL_3__13798_ gnd vdd FILL
XFILL_2__11459_ gnd vdd FILL
XFILL_0__15426_ gnd vdd FILL
XFILL_0__12638_ gnd vdd FILL
XFILL_3__9983_ gnd vdd FILL
XFILL_5__9919_ gnd vdd FILL
XFILL_1__14977_ gnd vdd FILL
XFILL_4__12019_ gnd vdd FILL
XSFILL8120x72050 gnd vdd FILL
XFILL_5__14358_ gnd vdd FILL
XFILL_3__12749_ gnd vdd FILL
XFILL_3__15537_ gnd vdd FILL
X_7764_ _7672_/B _9556_/B gnd _7764_/Y vdd NAND2X1
XFILL_2__14178_ gnd vdd FILL
XSFILL89400x35050 gnd vdd FILL
XFILL_1__13928_ gnd vdd FILL
XFILL_0__15357_ gnd vdd FILL
XFILL_5__13309_ gnd vdd FILL
XFILL_0__12569_ gnd vdd FILL
X_9503_ _9501_/Y _9514_/A _9503_/C gnd _9503_/Y vdd OAI21X1
XFILL_0__7067_ gnd vdd FILL
XFILL_2__13129_ gnd vdd FILL
XFILL_5__14289_ gnd vdd FILL
X_7695_ _7690_/B _9487_/B gnd _7696_/C vdd NAND2X1
XFILL_3__8865_ gnd vdd FILL
XFILL_0__14308_ gnd vdd FILL
XFILL_3__15468_ gnd vdd FILL
XFILL_1__13859_ gnd vdd FILL
XFILL111880x73050 gnd vdd FILL
XFILL_5__16028_ gnd vdd FILL
XFILL_0__15288_ gnd vdd FILL
XFILL_1__6900_ gnd vdd FILL
X_9434_ _9434_/Q _7389_/CLK _8285_/R vdd _9348_/Y gnd vdd DFFSR
XFILL_3__14419_ gnd vdd FILL
XFILL_1__7880_ gnd vdd FILL
XFILL_3__15399_ gnd vdd FILL
XFILL_3__7816_ gnd vdd FILL
XFILL_0__14239_ gnd vdd FILL
XSFILL13640x30050 gnd vdd FILL
XFILL_4__15709_ gnd vdd FILL
X_9365_ _9425_/A _6933_/B gnd _9365_/Y vdd NAND2X1
XFILL_1__15529_ gnd vdd FILL
XFILL_3__7747_ gnd vdd FILL
XFILL_4_BUFX2_insert504 gnd vdd FILL
XFILL_4_BUFX2_insert515 gnd vdd FILL
XFILL_6__7456_ gnd vdd FILL
XFILL_1__9550_ gnd vdd FILL
X_8316_ _8408_/Q gnd _8318_/A vdd INVX1
XFILL_0__7969_ gnd vdd FILL
XFILL_4_BUFX2_insert526 gnd vdd FILL
X_9296_ _9332_/Q gnd _9296_/Y vdd INVX1
XFILL_4_BUFX2_insert537 gnd vdd FILL
XFILL_4_BUFX2_insert548 gnd vdd FILL
XFILL_3__7678_ gnd vdd FILL
XFILL_4_BUFX2_insert559 gnd vdd FILL
XFILL_1__8501_ gnd vdd FILL
X_8247_ _8245_/Y _8246_/A _8247_/C gnd _8299_/D vdd OAI21X1
XFILL_1__9481_ gnd vdd FILL
XFILL_4__8210_ gnd vdd FILL
XFILL_3__9417_ gnd vdd FILL
XSFILL104520x11050 gnd vdd FILL
XFILL_6__9126_ gnd vdd FILL
XFILL_0__9639_ gnd vdd FILL
XSFILL83960x71050 gnd vdd FILL
XSFILL33800x43050 gnd vdd FILL
XFILL_4__8141_ gnd vdd FILL
XFILL_3__9348_ gnd vdd FILL
X_8178_ _8138_/A _8818_/CLK _8278_/R vdd _8178_/D gnd vdd DFFSR
X_7129_ _7039_/A _7129_/CLK _9049_/R vdd _7129_/D gnd vdd DFFSR
XFILL_1__8363_ gnd vdd FILL
XFILL_3__9279_ gnd vdd FILL
XFILL_4__8072_ gnd vdd FILL
XFILL_1__7314_ gnd vdd FILL
XFILL_3_CLKBUF1_insert206 gnd vdd FILL
XFILL_3_CLKBUF1_insert217 gnd vdd FILL
XFILL111960x53050 gnd vdd FILL
XSFILL23480x33050 gnd vdd FILL
XFILL_1__7245_ gnd vdd FILL
XSFILL13720x10050 gnd vdd FILL
XFILL112360x5050 gnd vdd FILL
X_12750_ _12777_/A memoryOutData[18] gnd _12751_/C vdd NAND2X1
XFILL_1_BUFX2_insert405 gnd vdd FILL
XFILL112040x62050 gnd vdd FILL
XFILL_1__7176_ gnd vdd FILL
XFILL_1_BUFX2_insert416 gnd vdd FILL
XFILL_1_BUFX2_insert427 gnd vdd FILL
XFILL_1_BUFX2_insert438 gnd vdd FILL
X_11701_ _11720_/A gnd _11703_/C vdd INVX1
XFILL_4__8974_ gnd vdd FILL
XFILL_1_BUFX2_insert449 gnd vdd FILL
X_12681_ _12621_/A _12809_/CLK _12809_/R vdd _12681_/D gnd vdd DFFSR
X_14420_ _14418_/Y _14160_/B _13876_/C _14419_/Y gnd _14421_/B vdd OAI22X1
XSFILL4280x59050 gnd vdd FILL
X_11632_ _11138_/Y _11748_/A _11366_/B _11137_/Y gnd _11632_/Y vdd OAI22X1
XSFILL114600x76050 gnd vdd FILL
XSFILL43640x46050 gnd vdd FILL
XFILL_2__6940_ gnd vdd FILL
X_14351_ _14351_/A _14045_/A _13456_/A _14349_/Y gnd _14352_/A vdd OAI22X1
XFILL_4__7856_ gnd vdd FILL
X_11563_ _11553_/B _11559_/Y _11563_/C gnd _11563_/Y vdd NAND3X1
XSFILL69080x57050 gnd vdd FILL
XSFILL99320x18050 gnd vdd FILL
XFILL_2__6871_ gnd vdd FILL
X_13302_ _13209_/Y _13222_/B _13302_/C gnd _13303_/B vdd OAI21X1
X_10514_ _10548_/B _7314_/B gnd _10514_/Y vdd NAND2X1
XSFILL84120x60050 gnd vdd FILL
XFILL_2__8610_ gnd vdd FILL
X_14282_ _14278_/Y _14282_/B gnd _14287_/C vdd NOR2X1
XFILL_5_BUFX2_insert360 gnd vdd FILL
X_11494_ _11494_/A _11764_/A gnd _11494_/Y vdd NAND2X1
XFILL_2__9590_ gnd vdd FILL
XBUFX2_insert50 _13381_/Y gnd _14071_/B vdd BUFX2
XFILL_5_BUFX2_insert371 gnd vdd FILL
XFILL_4__9526_ gnd vdd FILL
X_16021_ _16021_/A _16012_/Y gnd _16046_/A vdd NOR2X1
XBUFX2_insert61 _14983_/Y gnd _15369_/A vdd BUFX2
XFILL_5_BUFX2_insert382 gnd vdd FILL
X_13233_ _13231_/A gnd _13236_/B vdd INVX2
XBUFX2_insert72 _12366_/Y gnd _6924_/B vdd BUFX2
XFILL_5_BUFX2_insert393 gnd vdd FILL
XSFILL23800x9050 gnd vdd FILL
X_10445_ _10483_/Q gnd _10445_/Y vdd INVX1
XBUFX2_insert83 _13372_/Y gnd _13871_/A vdd BUFX2
XFILL_1__9748_ gnd vdd FILL
XBUFX2_insert94 _15068_/Y gnd _15581_/C vdd BUFX2
XFILL_5__8250_ gnd vdd FILL
X_13164_ _13149_/A _13164_/B gnd _13165_/C vdd NAND2X1
XSFILL23800x75050 gnd vdd FILL
X_10376_ _15300_/A gnd _10378_/A vdd INVX1
XFILL_2__10830_ gnd vdd FILL
XFILL_1__9679_ gnd vdd FILL
XFILL_2__8472_ gnd vdd FILL
XFILL_5__11990_ gnd vdd FILL
XFILL_5__7201_ gnd vdd FILL
XFILL_3__11080_ gnd vdd FILL
X_12115_ _11887_/A gnd _12117_/A vdd INVX1
XFILL112120x42050 gnd vdd FILL
XFILL_4__9388_ gnd vdd FILL
XFILL_5__10941_ gnd vdd FILL
XFILL_2__7423_ gnd vdd FILL
XFILL_4__12370_ gnd vdd FILL
X_13095_ _13155_/A _13095_/B gnd _13095_/Y vdd NAND2X1
XFILL_3__10031_ gnd vdd FILL
XFILL_1__11210_ gnd vdd FILL
XFILL_2__10761_ gnd vdd FILL
XFILL_4__8339_ gnd vdd FILL
XSFILL114600x50 gnd vdd FILL
XFILL_1__12190_ gnd vdd FILL
XFILL_0__11940_ gnd vdd FILL
X_12046_ _12046_/A _12046_/B _12046_/C gnd _13122_/B vdd NAND3X1
XFILL_4__11321_ gnd vdd FILL
XFILL_5__13660_ gnd vdd FILL
XFILL_2__12500_ gnd vdd FILL
XFILL_2__7354_ gnd vdd FILL
XFILL_5__10872_ gnd vdd FILL
XFILL_1__11141_ gnd vdd FILL
XFILL_2__13480_ gnd vdd FILL
XFILL_5__7063_ gnd vdd FILL
XFILL_2__10692_ gnd vdd FILL
XFILL_0__11871_ gnd vdd FILL
XSFILL43720x26050 gnd vdd FILL
XFILL_5__12611_ gnd vdd FILL
XFILL_4__14040_ gnd vdd FILL
XFILL_4__11252_ gnd vdd FILL
XFILL_2__12431_ gnd vdd FILL
XFILL_5__13591_ gnd vdd FILL
XSFILL53880x70050 gnd vdd FILL
XFILL_0__13610_ gnd vdd FILL
XFILL_3__11982_ gnd vdd FILL
XFILL_3__14770_ gnd vdd FILL
XFILL_1__11072_ gnd vdd FILL
XFILL_0__10822_ gnd vdd FILL
XFILL_0__14590_ gnd vdd FILL
XFILL_5__15330_ gnd vdd FILL
X_15805_ _15804_/Y _15328_/B _15376_/B _15805_/D gnd _15809_/A vdd OAI22X1
XSFILL69160x37050 gnd vdd FILL
XFILL_6__14881_ gnd vdd FILL
XSFILL3640x2050 gnd vdd FILL
XFILL_2__9024_ gnd vdd FILL
XFILL_3__10933_ gnd vdd FILL
XFILL_1__10023_ gnd vdd FILL
X_13997_ _13988_/Y _13997_/B _13997_/C gnd _13997_/Y vdd NAND3X1
XFILL_4__11183_ gnd vdd FILL
XFILL_1__14900_ gnd vdd FILL
XFILL_2__15150_ gnd vdd FILL
XFILL_3__13721_ gnd vdd FILL
XFILL_2_BUFX2_insert250 gnd vdd FILL
XFILL_2__12362_ gnd vdd FILL
XFILL_2_BUFX2_insert261 gnd vdd FILL
XFILL_0__10753_ gnd vdd FILL
XFILL_0__13541_ gnd vdd FILL
XSFILL84200x40050 gnd vdd FILL
XFILL_1__15880_ gnd vdd FILL
XFILL_2_BUFX2_insert272 gnd vdd FILL
XFILL_2_BUFX2_insert283 gnd vdd FILL
X_12948_ _12910_/A _9050_/CLK _9050_/R vdd _12948_/D gnd vdd DFFSR
XFILL_4__10134_ gnd vdd FILL
XFILL_5__15261_ gnd vdd FILL
XFILL_2__14101_ gnd vdd FILL
X_15736_ _15736_/A _15736_/B _15733_/Y gnd _15736_/Y vdd NAND3X1
XFILL_3__13652_ gnd vdd FILL
XFILL_5__12473_ gnd vdd FILL
XFILL_2_BUFX2_insert294 gnd vdd FILL
XFILL_2__11313_ gnd vdd FILL
XFILL_4__15991_ gnd vdd FILL
XFILL_1__14831_ gnd vdd FILL
XFILL_2__15081_ gnd vdd FILL
XFILL_2__12293_ gnd vdd FILL
XFILL_0__16260_ gnd vdd FILL
XFILL_0__10684_ gnd vdd FILL
XFILL_5__14212_ gnd vdd FILL
XFILL_0__13472_ gnd vdd FILL
XFILL_3__12603_ gnd vdd FILL
XSFILL74280x28050 gnd vdd FILL
XFILL_5__7965_ gnd vdd FILL
XFILL_5__11424_ gnd vdd FILL
XFILL_5__15192_ gnd vdd FILL
X_15667_ _15667_/A _15662_/Y _15667_/C gnd _15667_/Y vdd NAND3X1
XFILL_2__14032_ gnd vdd FILL
XFILL_4__14942_ gnd vdd FILL
X_12879_ _12877_/Y vdd _12879_/C gnd _12937_/D vdd OAI21X1
XFILL_1_BUFX2_insert950 gnd vdd FILL
XFILL_4__10065_ gnd vdd FILL
XFILL_3__16371_ gnd vdd FILL
XFILL_0__15211_ gnd vdd FILL
XFILL_3__13583_ gnd vdd FILL
XFILL_2__11244_ gnd vdd FILL
XFILL_0__12423_ gnd vdd FILL
XFILL_3__6980_ gnd vdd FILL
XFILL_1_BUFX2_insert961 gnd vdd FILL
XFILL_3__10795_ gnd vdd FILL
XFILL_1__14762_ gnd vdd FILL
XFILL_1__11974_ gnd vdd FILL
XFILL_5__6916_ gnd vdd FILL
XFILL_1_BUFX2_insert972 gnd vdd FILL
XFILL_0__16191_ gnd vdd FILL
XFILL_1_BUFX2_insert983 gnd vdd FILL
X_14618_ _14618_/A _14617_/Y gnd _14647_/A vdd NOR2X1
XFILL_5__14143_ gnd vdd FILL
XFILL_1_BUFX2_insert994 gnd vdd FILL
XFILL_3__15322_ gnd vdd FILL
XFILL_3__12534_ gnd vdd FILL
XFILL_0__9990_ gnd vdd FILL
XFILL_6__13694_ gnd vdd FILL
X_15598_ _15598_/A _15598_/B gnd _15609_/A vdd NAND2X1
XFILL_5__11355_ gnd vdd FILL
XFILL_4__14873_ gnd vdd FILL
XFILL_2__9926_ gnd vdd FILL
XFILL_1__13713_ gnd vdd FILL
XFILL112200x22050 gnd vdd FILL
XFILL_0__12354_ gnd vdd FILL
XFILL_1__10925_ gnd vdd FILL
XFILL_0__15142_ gnd vdd FILL
XFILL_2__11175_ gnd vdd FILL
XFILL_5__9635_ gnd vdd FILL
XFILL_1__14693_ gnd vdd FILL
X_14549_ _14527_/Y _14549_/B _15651_/C gnd _13018_/B vdd AOI21X1
XFILL_5__6847_ gnd vdd FILL
XFILL_5__10306_ gnd vdd FILL
XFILL_4__13824_ gnd vdd FILL
XFILL_3__15253_ gnd vdd FILL
X_7480_ _7480_/A gnd _7482_/A vdd INVX1
XFILL_5__14074_ gnd vdd FILL
XFILL_5__11286_ gnd vdd FILL
XFILL_2__10126_ gnd vdd FILL
XFILL_3__8650_ gnd vdd FILL
XFILL_3__12465_ gnd vdd FILL
XFILL_0__11305_ gnd vdd FILL
XBUFX2_insert260 _11225_/Y gnd _11778_/B vdd BUFX2
XFILL_2__9857_ gnd vdd FILL
XFILL_1__13644_ gnd vdd FILL
XFILL_2__15983_ gnd vdd FILL
XFILL_0__15073_ gnd vdd FILL
XBUFX2_insert271 _13364_/Y gnd _10658_/B vdd BUFX2
XFILL_0__12285_ gnd vdd FILL
XFILL_3__14204_ gnd vdd FILL
XBUFX2_insert282 _15003_/Y gnd _15677_/D vdd BUFX2
XFILL_5__13025_ gnd vdd FILL
XFILL_5__10237_ gnd vdd FILL
XFILL_0__8872_ gnd vdd FILL
XSFILL18680x2050 gnd vdd FILL
XBUFX2_insert293 _13356_/Y gnd _10264_/A vdd BUFX2
XFILL_3__11416_ gnd vdd FILL
XFILL_3__7601_ gnd vdd FILL
XFILL_3__15184_ gnd vdd FILL
XFILL_4__13755_ gnd vdd FILL
XFILL_4__10967_ gnd vdd FILL
XFILL_1__16363_ gnd vdd FILL
XFILL_0__14024_ gnd vdd FILL
XFILL_3__12396_ gnd vdd FILL
XFILL_2__14934_ gnd vdd FILL
XFILL_3__8581_ gnd vdd FILL
XFILL_2__10057_ gnd vdd FILL
XFILL_0__11236_ gnd vdd FILL
XFILL_2__9788_ gnd vdd FILL
XFILL_5__8517_ gnd vdd FILL
XFILL_5_CLKBUF1_insert150 gnd vdd FILL
XFILL_1__13575_ gnd vdd FILL
XFILL_0__7823_ gnd vdd FILL
XFILL_1__10787_ gnd vdd FILL
X_16219_ _16219_/A _16219_/B _16219_/C gnd _16220_/A vdd NAND3X1
XSFILL53960x50050 gnd vdd FILL
XFILL_4__12706_ gnd vdd FILL
X_9150_ _9198_/Q gnd _9150_/Y vdd INVX1
XFILL_5__9497_ gnd vdd FILL
XSFILL54440x57050 gnd vdd FILL
XFILL_3__14135_ gnd vdd FILL
XFILL_5__10168_ gnd vdd FILL
XFILL_5_CLKBUF1_insert161 gnd vdd FILL
XFILL_1__15314_ gnd vdd FILL
XFILL_5_CLKBUF1_insert172 gnd vdd FILL
XFILL_3__11347_ gnd vdd FILL
XFILL_2__8739_ gnd vdd FILL
XFILL_4__10898_ gnd vdd FILL
XFILL_2__14865_ gnd vdd FILL
XFILL_4__13686_ gnd vdd FILL
XFILL_1__12526_ gnd vdd FILL
XFILL_5_CLKBUF1_insert183 gnd vdd FILL
XSFILL69240x17050 gnd vdd FILL
XFILL_5_CLKBUF1_insert194 gnd vdd FILL
XFILL_0__11167_ gnd vdd FILL
XFILL_1__16294_ gnd vdd FILL
XFILL_5__8448_ gnd vdd FILL
X_8101_ _8101_/A _8100_/A _8101_/C gnd _8101_/Y vdd OAI21X1
XFILL_0__7754_ gnd vdd FILL
XFILL_4__15425_ gnd vdd FILL
XFILL_4__12637_ gnd vdd FILL
XFILL_2__13816_ gnd vdd FILL
XFILL_3__14066_ gnd vdd FILL
XFILL_5__14976_ gnd vdd FILL
X_9081_ _9175_/Q gnd _9081_/Y vdd INVX1
XFILL_3__7463_ gnd vdd FILL
XFILL_1__15245_ gnd vdd FILL
XFILL_0__10118_ gnd vdd FILL
XFILL_3__11278_ gnd vdd FILL
XFILL_1__12457_ gnd vdd FILL
XFILL_2__14796_ gnd vdd FILL
XFILL_5__8379_ gnd vdd FILL
XFILL_0__15975_ gnd vdd FILL
XFILL_6__7172_ gnd vdd FILL
XSFILL104440x26050 gnd vdd FILL
XFILL_0__11098_ gnd vdd FILL
XFILL_3__13017_ gnd vdd FILL
X_8032_ _7956_/A _7274_/CLK _7274_/R vdd _8032_/D gnd vdd DFFSR
XFILL_5__13927_ gnd vdd FILL
XFILL_4__15356_ gnd vdd FILL
XFILL_0__7685_ gnd vdd FILL
XFILL_4__12568_ gnd vdd FILL
XFILL_2__13747_ gnd vdd FILL
XFILL_1__11408_ gnd vdd FILL
XSFILL8680x24050 gnd vdd FILL
XFILL_2__10959_ gnd vdd FILL
XFILL_1__15176_ gnd vdd FILL
XFILL_0__10049_ gnd vdd FILL
XFILL_0__14926_ gnd vdd FILL
XFILL_1__12388_ gnd vdd FILL
XFILL_0__9424_ gnd vdd FILL
XFILL_4__14307_ gnd vdd FILL
XFILL_5__13858_ gnd vdd FILL
XFILL_3__9133_ gnd vdd FILL
XFILL_4__11519_ gnd vdd FILL
XFILL_1__14127_ gnd vdd FILL
XFILL_4__12499_ gnd vdd FILL
XFILL_4__15287_ gnd vdd FILL
XFILL_2__13678_ gnd vdd FILL
XFILL_1__11339_ gnd vdd FILL
XSFILL59160x69050 gnd vdd FILL
XFILL_0__14857_ gnd vdd FILL
XFILL_0__9355_ gnd vdd FILL
XFILL_4__14238_ gnd vdd FILL
XFILL_2__15417_ gnd vdd FILL
X_9983_ _9983_/A gnd _9983_/Y vdd INVX1
XFILL_2__12629_ gnd vdd FILL
XFILL_5__13789_ gnd vdd FILL
XFILL_0__13808_ gnd vdd FILL
XFILL_1__14058_ gnd vdd FILL
XFILL_3__14968_ gnd vdd FILL
XFILL_2__16397_ gnd vdd FILL
XSFILL74200x72050 gnd vdd FILL
XFILL_5__15528_ gnd vdd FILL
XFILL_0__14788_ gnd vdd FILL
XFILL_3__8015_ gnd vdd FILL
X_8934_ _8870_/A _8921_/CLK _9049_/R vdd _8934_/D gnd vdd DFFSR
XFILL_0__9286_ gnd vdd FILL
XFILL_2__15348_ gnd vdd FILL
XFILL_4__14169_ gnd vdd FILL
XFILL_1__13009_ gnd vdd FILL
XFILL_3__13919_ gnd vdd FILL
XSFILL109160x38050 gnd vdd FILL
XFILL_6__9813_ gnd vdd FILL
XFILL_3__14899_ gnd vdd FILL
XFILL_0__13739_ gnd vdd FILL
XFILL_1__7030_ gnd vdd FILL
XFILL_0__8237_ gnd vdd FILL
XSFILL13640x25050 gnd vdd FILL
XFILL_5__15459_ gnd vdd FILL
X_8865_ _8845_/B _9889_/B gnd _8866_/C vdd NAND2X1
XSFILL79880x39050 gnd vdd FILL
XFILL_2__15279_ gnd vdd FILL
X_7816_ _7900_/Q gnd _7816_/Y vdd INVX1
XFILL_0__15409_ gnd vdd FILL
X_8796_ _8796_/Q _7662_/CLK _9454_/R vdd _8714_/Y gnd vdd DFFSR
XSFILL114280x29050 gnd vdd FILL
XFILL_0__7119_ gnd vdd FILL
XFILL_0__16389_ gnd vdd FILL
XFILL_0__8099_ gnd vdd FILL
X_7747_ _7747_/A _7753_/B _7747_/C gnd _7791_/D vdd OAI21X1
XFILL_1__8981_ gnd vdd FILL
XFILL_4__7710_ gnd vdd FILL
XFILL_3__8917_ gnd vdd FILL
XFILL_3__9897_ gnd vdd FILL
XFILL_1__7932_ gnd vdd FILL
XSFILL33800x38050 gnd vdd FILL
X_7678_ _7676_/Y _7723_/B _7678_/C gnd _7768_/D vdd OAI21X1
XFILL_3__8848_ gnd vdd FILL
XSFILL43960x82050 gnd vdd FILL
X_9417_ _9417_/A _9401_/A _9416_/Y gnd _9457_/D vdd OAI21X1
XFILL_1__7863_ gnd vdd FILL
XFILL_4__7572_ gnd vdd FILL
XFILL_3__8779_ gnd vdd FILL
XFILL_6__7508_ gnd vdd FILL
XFILL_4_BUFX2_insert301 gnd vdd FILL
XFILL_1__9602_ gnd vdd FILL
X_9348_ _9348_/A _9398_/A _9347_/Y gnd _9348_/Y vdd OAI21X1
XFILL_4_BUFX2_insert312 gnd vdd FILL
XFILL_4_BUFX2_insert323 gnd vdd FILL
XFILL111960x48050 gnd vdd FILL
XFILL_4_BUFX2_insert334 gnd vdd FILL
X_10230_ _13452_/A gnd _10232_/A vdd INVX1
XFILL_1__9533_ gnd vdd FILL
XFILL_4_BUFX2_insert345 gnd vdd FILL
XFILL_4_BUFX2_insert356 gnd vdd FILL
X_9279_ _9232_/B _8255_/B gnd _9279_/Y vdd NAND2X1
XFILL_4__9242_ gnd vdd FILL
XFILL_4_BUFX2_insert367 gnd vdd FILL
XFILL_4_BUFX2_insert378 gnd vdd FILL
XFILL_4_BUFX2_insert389 gnd vdd FILL
X_10161_ _10161_/A _10160_/A _10161_/C gnd _10217_/D vdd OAI21X1
XFILL112040x57050 gnd vdd FILL
XFILL_1__9464_ gnd vdd FILL
XFILL_4__9173_ gnd vdd FILL
X_10092_ _15962_/A _7020_/CLK _9580_/R vdd _10042_/Y gnd vdd DFFSR
XFILL_4__8124_ gnd vdd FILL
XSFILL38920x71050 gnd vdd FILL
XFILL_1__9395_ gnd vdd FILL
X_13920_ _13920_/A gnd _13920_/Y vdd INVX1
XFILL_1__8346_ gnd vdd FILL
XFILL_4__8055_ gnd vdd FILL
X_13851_ _10462_/Q _14389_/B _13850_/Y gnd _13851_/Y vdd AOI21X1
XFILL_1__8277_ gnd vdd FILL
XFILL_2__7070_ gnd vdd FILL
X_12802_ _12802_/Q _12685_/CLK _12685_/R vdd _12802_/D gnd vdd DFFSR
XFILL_1__7228_ gnd vdd FILL
X_13782_ _13780_/Y _14830_/B _14203_/C _13781_/Y gnd _13782_/Y vdd OAI22X1
X_10994_ _12338_/Y gnd _10995_/B vdd INVX1
X_12733_ _12731_/Y _12768_/A _12733_/C gnd _12733_/Y vdd OAI21X1
X_15521_ _15915_/C _13985_/D _15521_/C _13995_/D gnd _15521_/Y vdd OAI22X1
XFILL_1_BUFX2_insert235 gnd vdd FILL
XFILL_1_BUFX2_insert246 gnd vdd FILL
XFILL_1__7159_ gnd vdd FILL
XFILL_1_BUFX2_insert257 gnd vdd FILL
XFILL_1_BUFX2_insert268 gnd vdd FILL
XFILL_4__8957_ gnd vdd FILL
X_15452_ _15842_/A _15451_/Y _15452_/C _16137_/C gnd _15453_/B vdd OAI22X1
XFILL_1_BUFX2_insert279 gnd vdd FILL
XFILL_5__7750_ gnd vdd FILL
X_12664_ _12570_/A _12667_/CLK _12795_/R vdd _12664_/D gnd vdd DFFSR
XFILL_6__10760_ gnd vdd FILL
XFILL_0_BUFX2_insert902 gnd vdd FILL
XFILL_2__7972_ gnd vdd FILL
XFILL_3__10580_ gnd vdd FILL
XFILL_0_BUFX2_insert913 gnd vdd FILL
X_14403_ _8626_/A _13864_/B _14403_/C _8498_/A gnd _14403_/Y vdd AOI22X1
XFILL_5__7681_ gnd vdd FILL
XFILL112120x37050 gnd vdd FILL
XFILL_0_BUFX2_insert924 gnd vdd FILL
XFILL_5__11140_ gnd vdd FILL
X_11615_ _11138_/Y gnd _11615_/Y vdd INVX2
X_15383_ _15383_/A _7646_/Q _7518_/Q _15383_/D gnd _15388_/B vdd AOI22X1
XFILL_0_BUFX2_insert935 gnd vdd FILL
XFILL_4__8888_ gnd vdd FILL
XFILL_2__6923_ gnd vdd FILL
X_12595_ vdd memoryOutData[9] gnd _12596_/C vdd NAND2X1
XFILL_0_BUFX2_insert946 gnd vdd FILL
XFILL_4__11870_ gnd vdd FILL
XFILL_0_BUFX2_insert957 gnd vdd FILL
XSFILL23400x72050 gnd vdd FILL
XFILL_5__9420_ gnd vdd FILL
XFILL_0_BUFX2_insert968 gnd vdd FILL
X_14334_ _9644_/A gnd _14336_/A vdd INVX1
XFILL_1__11690_ gnd vdd FILL
XSFILL38200x32050 gnd vdd FILL
XFILL_4__7839_ gnd vdd FILL
XFILL_0_BUFX2_insert979 gnd vdd FILL
X_11546_ _11546_/A _11846_/C _11545_/Y gnd _11546_/Y vdd AOI21X1
XFILL_5__11071_ gnd vdd FILL
XFILL_3__12250_ gnd vdd FILL
XFILL_4__10821_ gnd vdd FILL
XFILL_2__6854_ gnd vdd FILL
XFILL_2__9642_ gnd vdd FILL
XFILL_0__12070_ gnd vdd FILL
XFILL_2__12980_ gnd vdd FILL
XFILL_1__10641_ gnd vdd FILL
XFILL_5__10022_ gnd vdd FILL
XFILL_5__9351_ gnd vdd FILL
X_14265_ _14265_/A _14265_/B _14265_/C gnd _13000_/B vdd AOI21X1
XFILL_3__11201_ gnd vdd FILL
XFILL_4__10752_ gnd vdd FILL
X_11477_ _11476_/Y _11477_/B _11461_/A gnd _11477_/Y vdd OAI21X1
XFILL_4__13540_ gnd vdd FILL
XFILL_2__11931_ gnd vdd FILL
XFILL_3__12181_ gnd vdd FILL
XFILL_0__11021_ gnd vdd FILL
XFILL_4__9509_ gnd vdd FILL
XFILL_1__13360_ gnd vdd FILL
X_16004_ _15998_/Y _16004_/B gnd _16004_/Y vdd NAND2X1
X_13216_ _13220_/A _13305_/A gnd _13281_/B vdd NAND2X1
XFILL_1__10572_ gnd vdd FILL
XFILL_5__9282_ gnd vdd FILL
X_10428_ _10423_/B _9788_/B gnd _10428_/Y vdd NAND2X1
XFILL_5__14830_ gnd vdd FILL
X_14196_ _14626_/A _7397_/Q _7909_/Q _13865_/B gnd _14196_/Y vdd AOI22X1
XFILL_2__8524_ gnd vdd FILL
XFILL_3__11132_ gnd vdd FILL
XFILL_4__10683_ gnd vdd FILL
XFILL_4__13471_ gnd vdd FILL
XFILL_1__12311_ gnd vdd FILL
XFILL_2__14650_ gnd vdd FILL
XSFILL28680x41050 gnd vdd FILL
XFILL_5__8233_ gnd vdd FILL
XFILL_2__11862_ gnd vdd FILL
XFILL_1__13291_ gnd vdd FILL
XFILL_4__15210_ gnd vdd FILL
X_13147_ _13145_/Y _13149_/A _13147_/C gnd _13197_/D vdd OAI21X1
XFILL_4_BUFX2_insert890 gnd vdd FILL
XFILL_2__13601_ gnd vdd FILL
XFILL_4__12422_ gnd vdd FILL
X_10359_ _8823_/A _10405_/B gnd _10360_/C vdd NAND2X1
XFILL_5__14761_ gnd vdd FILL
XFILL_2__10813_ gnd vdd FILL
XFILL_5__11973_ gnd vdd FILL
XFILL_4__16190_ gnd vdd FILL
XFILL_1__15030_ gnd vdd FILL
XFILL_3__15940_ gnd vdd FILL
XFILL_3__11063_ gnd vdd FILL
XFILL_2__8455_ gnd vdd FILL
XFILL_2__14581_ gnd vdd FILL
XFILL_1__12242_ gnd vdd FILL
XFILL_0__15760_ gnd vdd FILL
XFILL_2__11793_ gnd vdd FILL
XFILL_0__12972_ gnd vdd FILL
XFILL_5__13712_ gnd vdd FILL
XFILL_4__12353_ gnd vdd FILL
XFILL_5__10924_ gnd vdd FILL
XFILL_2__16320_ gnd vdd FILL
X_13078_ _6901_/A _8176_/CLK _7408_/R vdd _13078_/D gnd vdd DFFSR
XFILL_0__7470_ gnd vdd FILL
XFILL_3__10014_ gnd vdd FILL
XFILL_4__15141_ gnd vdd FILL
XFILL_5__14692_ gnd vdd FILL
XFILL_2__13532_ gnd vdd FILL
XFILL_5__7115_ gnd vdd FILL
XFILL_2__10744_ gnd vdd FILL
XFILL_0__14711_ gnd vdd FILL
XFILL_2__8386_ gnd vdd FILL
XFILL_3__15871_ gnd vdd FILL
XFILL_0__11923_ gnd vdd FILL
XFILL_1__12173_ gnd vdd FILL
XFILL_0__15691_ gnd vdd FILL
X_12029_ _12029_/A _12025_/B _12025_/C gnd gnd _12029_/Y vdd AOI22X1
XFILL_5__8095_ gnd vdd FILL
XFILL_4__11304_ gnd vdd FILL
XFILL_5__13643_ gnd vdd FILL
XFILL_3__14822_ gnd vdd FILL
XFILL_4__15072_ gnd vdd FILL
XFILL_2__7337_ gnd vdd FILL
XFILL_4__12284_ gnd vdd FILL
XFILL_2__16251_ gnd vdd FILL
XFILL_2__13463_ gnd vdd FILL
XFILL_1__11124_ gnd vdd FILL
XFILL_0__14642_ gnd vdd FILL
XFILL_5__7046_ gnd vdd FILL
XFILL_2__10675_ gnd vdd FILL
XFILL_0__9140_ gnd vdd FILL
XFILL_0__11854_ gnd vdd FILL
XFILL_2__15202_ gnd vdd FILL
XFILL_4__14023_ gnd vdd FILL
XFILL_5__16362_ gnd vdd FILL
XFILL_4__11235_ gnd vdd FILL
XFILL_6__14933_ gnd vdd FILL
XFILL_2__12414_ gnd vdd FILL
XFILL_5__13574_ gnd vdd FILL
XFILL_2__16182_ gnd vdd FILL
XFILL_3__11965_ gnd vdd FILL
XFILL_1__15932_ gnd vdd FILL
XFILL_5__10786_ gnd vdd FILL
X_6980_ _6980_/A gnd _6982_/A vdd INVX1
XFILL_3__14753_ gnd vdd FILL
XFILL_1__11055_ gnd vdd FILL
XFILL_0__10805_ gnd vdd FILL
XFILL_2__13394_ gnd vdd FILL
XFILL_0__14573_ gnd vdd FILL
XFILL_5__15313_ gnd vdd FILL
XFILL_5__12525_ gnd vdd FILL
XFILL_2__9007_ gnd vdd FILL
XFILL_0__11785_ gnd vdd FILL
XFILL_3__10916_ gnd vdd FILL
XFILL_5__16293_ gnd vdd FILL
XFILL_1__10006_ gnd vdd FILL
XFILL_2__15133_ gnd vdd FILL
XFILL_3__13704_ gnd vdd FILL
XFILL_4__11166_ gnd vdd FILL
XFILL_2__12345_ gnd vdd FILL
XFILL_0__16312_ gnd vdd FILL
XFILL_3__11896_ gnd vdd FILL
XFILL_3__14684_ gnd vdd FILL
XFILL_2__7199_ gnd vdd FILL
XFILL_0__13524_ gnd vdd FILL
XFILL_1__15863_ gnd vdd FILL
X_15719_ _15719_/A _15719_/B _15719_/C gnd _15720_/A vdd NOR3X1
XFILL_5__15244_ gnd vdd FILL
XSFILL53960x45050 gnd vdd FILL
XFILL_4__10117_ gnd vdd FILL
XFILL_5__8997_ gnd vdd FILL
X_8650_ _8690_/Q gnd _8650_/Y vdd INVX1
XFILL_5__12456_ gnd vdd FILL
XFILL_6_BUFX2_insert418 gnd vdd FILL
XSFILL109480x74050 gnd vdd FILL
XFILL_3__13635_ gnd vdd FILL
XFILL_4__15974_ gnd vdd FILL
XFILL_1__14814_ gnd vdd FILL
XFILL_2__15064_ gnd vdd FILL
XFILL_4__11097_ gnd vdd FILL
XFILL_0__16243_ gnd vdd FILL
XFILL_2__12276_ gnd vdd FILL
XFILL_0__13455_ gnd vdd FILL
XFILL_1__15794_ gnd vdd FILL
XFILL_0__10667_ gnd vdd FILL
XFILL_5__7948_ gnd vdd FILL
XFILL_6__13746_ gnd vdd FILL
XFILL_5__11407_ gnd vdd FILL
X_7601_ _7601_/A _7577_/B _7600_/Y gnd _7601_/Y vdd OAI21X1
XFILL_5__15175_ gnd vdd FILL
XFILL_4__10048_ gnd vdd FILL
XFILL_2__14015_ gnd vdd FILL
XFILL_1_BUFX2_insert780 gnd vdd FILL
XFILL_4__14925_ gnd vdd FILL
XSFILL28760x21050 gnd vdd FILL
XFILL_5__12387_ gnd vdd FILL
XFILL_3__16354_ gnd vdd FILL
XFILL_3__13566_ gnd vdd FILL
X_8581_ _8667_/Q gnd _8583_/A vdd INVX1
XFILL_2__11227_ gnd vdd FILL
XFILL_0__12406_ gnd vdd FILL
XSFILL54040x54050 gnd vdd FILL
XFILL_3__9751_ gnd vdd FILL
XFILL_3__10778_ gnd vdd FILL
XFILL_3__6963_ gnd vdd FILL
XFILL_1_BUFX2_insert791 gnd vdd FILL
XFILL_1__14745_ gnd vdd FILL
XFILL_0__16174_ gnd vdd FILL
XFILL_1__11957_ gnd vdd FILL
XFILL_5__14126_ gnd vdd FILL
XFILL_0__13386_ gnd vdd FILL
XFILL_3__15305_ gnd vdd FILL
X_7532_ _7480_/A _7532_/CLK _9313_/R vdd _7532_/D gnd vdd DFFSR
XFILL_5__7879_ gnd vdd FILL
XFILL_5__11338_ gnd vdd FILL
XFILL_2__9909_ gnd vdd FILL
XFILL_4__14856_ gnd vdd FILL
XFILL_3__12517_ gnd vdd FILL
XFILL_6__10889_ gnd vdd FILL
XFILL_3__8702_ gnd vdd FILL
XFILL_1__10908_ gnd vdd FILL
XFILL_3__16285_ gnd vdd FILL
XFILL_4_BUFX2_insert1008 gnd vdd FILL
XFILL_3__13497_ gnd vdd FILL
XFILL_2__11158_ gnd vdd FILL
XFILL_0__15125_ gnd vdd FILL
XSFILL8680x19050 gnd vdd FILL
XFILL_3__6894_ gnd vdd FILL
XFILL_4_BUFX2_insert1019 gnd vdd FILL
XFILL_1__14676_ gnd vdd FILL
XFILL_5__9618_ gnd vdd FILL
XFILL_3__9682_ gnd vdd FILL
XFILL_0__12337_ gnd vdd FILL
XFILL_4_BUFX2_insert40 gnd vdd FILL
XFILL_1__11888_ gnd vdd FILL
XFILL_4_BUFX2_insert51 gnd vdd FILL
XFILL_4__13807_ gnd vdd FILL
XFILL_5__14057_ gnd vdd FILL
XFILL_6__16396_ gnd vdd FILL
X_7463_ _7425_/B _9383_/B gnd _7464_/C vdd NAND2X1
XFILL_3__12448_ gnd vdd FILL
XFILL_3__15236_ gnd vdd FILL
XFILL_4_BUFX2_insert62 gnd vdd FILL
XFILL_1__16415_ gnd vdd FILL
XFILL_2__10109_ gnd vdd FILL
XSFILL33880x12050 gnd vdd FILL
XFILL_5__11269_ gnd vdd FILL
XFILL_1__13627_ gnd vdd FILL
XFILL_3__8633_ gnd vdd FILL
XFILL_4__14787_ gnd vdd FILL
XFILL_4_BUFX2_insert73 gnd vdd FILL
XFILL_4__11999_ gnd vdd FILL
XFILL_0__15056_ gnd vdd FILL
XFILL_2__15966_ gnd vdd FILL
XFILL_0__12268_ gnd vdd FILL
XFILL_2__11089_ gnd vdd FILL
XFILL_5__9549_ gnd vdd FILL
XFILL_6__15347_ gnd vdd FILL
X_9202_ _9162_/A _7282_/CLK _7411_/R vdd _9202_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert84 gnd vdd FILL
XFILL_5__13008_ gnd vdd FILL
XFILL_4_BUFX2_insert95 gnd vdd FILL
XFILL_0__8855_ gnd vdd FILL
XFILL_3__15167_ gnd vdd FILL
XFILL_4__13738_ gnd vdd FILL
XSFILL18680x73050 gnd vdd FILL
XFILL_1__16346_ gnd vdd FILL
XFILL_0__14007_ gnd vdd FILL
XFILL_3__12379_ gnd vdd FILL
X_7394_ _7394_/Q _7382_/CLK _8674_/R vdd _7324_/Y gnd vdd DFFSR
XSFILL48920x34050 gnd vdd FILL
XFILL_2__14917_ gnd vdd FILL
XSFILL104440x5050 gnd vdd FILL
XFILL_1__13558_ gnd vdd FILL
XFILL_0__11219_ gnd vdd FILL
XFILL_2__15897_ gnd vdd FILL
XSFILL74200x67050 gnd vdd FILL
XFILL_0__12199_ gnd vdd FILL
XFILL_0__7806_ gnd vdd FILL
XFILL_6__8273_ gnd vdd FILL
X_9133_ _9116_/B _6957_/B gnd _9133_/Y vdd NAND2X1
XFILL_0__8786_ gnd vdd FILL
XFILL_3__14118_ gnd vdd FILL
XFILL_4__13669_ gnd vdd FILL
XFILL_1__12509_ gnd vdd FILL
XFILL_3__15098_ gnd vdd FILL
XSFILL108680x26050 gnd vdd FILL
XFILL_2__14848_ gnd vdd FILL
XFILL_6__7224_ gnd vdd FILL
XFILL_3__8495_ gnd vdd FILL
XFILL_1__16277_ gnd vdd FILL
XFILL_1__13489_ gnd vdd FILL
XFILL_4__15408_ gnd vdd FILL
XSFILL49000x43050 gnd vdd FILL
XFILL_2_BUFX2_insert1001 gnd vdd FILL
XFILL_0__7737_ gnd vdd FILL
XFILL_2_BUFX2_insert1012 gnd vdd FILL
XFILL_3_BUFX2_insert308 gnd vdd FILL
XFILL_3__14049_ gnd vdd FILL
XFILL_5__14959_ gnd vdd FILL
X_9064_ _9004_/A _7400_/CLK _9064_/R vdd _9064_/D gnd vdd DFFSR
XFILL_4__16388_ gnd vdd FILL
XFILL_1__15228_ gnd vdd FILL
XFILL_3_BUFX2_insert319 gnd vdd FILL
XFILL_3__7446_ gnd vdd FILL
XFILL_2_BUFX2_insert1023 gnd vdd FILL
XFILL_2_BUFX2_insert1034 gnd vdd FILL
XFILL_2__14779_ gnd vdd FILL
XFILL_0__15958_ gnd vdd FILL
X_8015_ _8015_/A _7948_/A _8014_/Y gnd _8051_/D vdd OAI21X1
XFILL_2_BUFX2_insert1045 gnd vdd FILL
XFILL_4__15339_ gnd vdd FILL
XFILL_2_BUFX2_insert1056 gnd vdd FILL
XFILL_2_BUFX2_insert1067 gnd vdd FILL
XFILL_1__15159_ gnd vdd FILL
XFILL_0__14909_ gnd vdd FILL
XFILL_3__7377_ gnd vdd FILL
XFILL_2_BUFX2_insert1089 gnd vdd FILL
XFILL_0__9407_ gnd vdd FILL
XFILL_1__8200_ gnd vdd FILL
XFILL_0__15889_ gnd vdd FILL
XFILL_3__9116_ gnd vdd FILL
XSFILL54120x34050 gnd vdd FILL
XFILL_0__7599_ gnd vdd FILL
XFILL_2__16449_ gnd vdd FILL
XFILL_1__8131_ gnd vdd FILL
XFILL_0__9338_ gnd vdd FILL
X_9966_ _9918_/A _7662_/CLK _9454_/R vdd _9966_/D gnd vdd DFFSR
XSFILL43960x77050 gnd vdd FILL
XFILL_0__9269_ gnd vdd FILL
XFILL_1__8062_ gnd vdd FILL
X_8917_ _8915_/Y _8916_/A _8917_/C gnd _8949_/D vdd OAI21X1
X_9897_ _9897_/A gnd _9897_/Y vdd INVX1
XFILL_4__9860_ gnd vdd FILL
XFILL_0_BUFX2_insert1060 gnd vdd FILL
XFILL_0_BUFX2_insert1071 gnd vdd FILL
XSFILL18760x53050 gnd vdd FILL
X_8848_ _8846_/Y _8823_/B _8847_/Y gnd _8848_/Y vdd OAI21X1
XSFILL8600x63050 gnd vdd FILL
XFILL_0_BUFX2_insert1093 gnd vdd FILL
XFILL_6_BUFX2_insert930 gnd vdd FILL
XFILL_4__9791_ gnd vdd FILL
X_8779_ _8714_/B _9803_/B gnd _8779_/Y vdd NAND2X1
XFILL_4__8742_ gnd vdd FILL
XSFILL43960x5050 gnd vdd FILL
XFILL_6_BUFX2_insert996 gnd vdd FILL
XFILL_6__9658_ gnd vdd FILL
XFILL_1__8964_ gnd vdd FILL
X_11400_ _11048_/A _11400_/B _11400_/C gnd _11400_/Y vdd AOI21X1
XFILL_6__8609_ gnd vdd FILL
X_12380_ _12380_/A _12675_/Q gnd _12381_/C vdd NAND2X1
XFILL_1__8895_ gnd vdd FILL
XSFILL38920x66050 gnd vdd FILL
XFILL112440x73050 gnd vdd FILL
XFILL_4__7624_ gnd vdd FILL
X_11331_ _11513_/A _11331_/B _11440_/A gnd _11358_/B vdd OAI21X1
XFILL_1__7846_ gnd vdd FILL
XFILL_4__7555_ gnd vdd FILL
X_14050_ _9570_/Q gnd _14050_/Y vdd INVX1
XSFILL39000x75050 gnd vdd FILL
X_11262_ _11054_/A _11720_/A gnd _11263_/B vdd NAND2X1
X_13001_ _12999_/Y vdd _13001_/C gnd _13063_/D vdd OAI21X1
X_10213_ _10213_/Q _7269_/CLK _9061_/R vdd _10149_/Y gnd vdd DFFSR
XFILL_4__7486_ gnd vdd FILL
XFILL_1__9516_ gnd vdd FILL
X_11193_ _12195_/Y gnd _11193_/Y vdd INVX1
XFILL_4__9225_ gnd vdd FILL
XSFILL69480x68050 gnd vdd FILL
XSFILL18840x33050 gnd vdd FILL
XFILL_3_BUFX2_insert820 gnd vdd FILL
X_10144_ _14123_/A gnd _10146_/A vdd INVX1
XFILL_3_BUFX2_insert831 gnd vdd FILL
XFILL_2__8240_ gnd vdd FILL
XFILL_3_BUFX2_insert842 gnd vdd FILL
XFILL_3_BUFX2_insert853 gnd vdd FILL
XFILL_4__9156_ gnd vdd FILL
XSFILL49640x5050 gnd vdd FILL
XFILL_3_BUFX2_insert864 gnd vdd FILL
XFILL_3_BUFX2_insert875 gnd vdd FILL
X_10075_ _9989_/A _8663_/CLK _8664_/R vdd _9991_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert886 gnd vdd FILL
XSFILL99320x31050 gnd vdd FILL
X_14952_ _14952_/A _14952_/B gnd _14978_/B vdd NOR2X1
XSFILL104680x77050 gnd vdd FILL
XFILL_1__9378_ gnd vdd FILL
XFILL_3_BUFX2_insert897 gnd vdd FILL
XFILL_4__8107_ gnd vdd FILL
XFILL_4__9087_ gnd vdd FILL
X_13903_ _8927_/Q gnd _13905_/A vdd INVX1
XFILL_5__10640_ gnd vdd FILL
XFILL_1__8329_ gnd vdd FILL
XFILL_2__7122_ gnd vdd FILL
X_14883_ _14883_/A gnd _14883_/Y vdd INVX1
XSFILL64040x17050 gnd vdd FILL
XFILL_4__11020_ gnd vdd FILL
X_13834_ _8971_/A gnd _15341_/A vdd INVX1
XFILL_2__7053_ gnd vdd FILL
XFILL_5__10571_ gnd vdd FILL
XFILL_3__11750_ gnd vdd FILL
XFILL_2__10391_ gnd vdd FILL
XFILL_0__11570_ gnd vdd FILL
XFILL_5__12310_ gnd vdd FILL
XFILL_5__8851_ gnd vdd FILL
XFILL_3__10701_ gnd vdd FILL
X_13765_ _13764_/Y _13617_/D gnd _13769_/A vdd NOR2X1
XFILL_5__13290_ gnd vdd FILL
X_10977_ _10977_/A vdd _10977_/C gnd _10985_/D vdd OAI21X1
XFILL_2__12130_ gnd vdd FILL
XSFILL89240x83050 gnd vdd FILL
XFILL_0__10521_ gnd vdd FILL
XFILL_3__11681_ gnd vdd FILL
XFILL_1__12860_ gnd vdd FILL
XFILL_5__7802_ gnd vdd FILL
XSFILL3480x24050 gnd vdd FILL
X_15504_ _15504_/A _15503_/Y _15504_/C gnd _15504_/Y vdd NAND3X1
XFILL_6__14580_ gnd vdd FILL
X_12716_ _12716_/A gnd _12718_/A vdd INVX1
XFILL_5__8782_ gnd vdd FILL
XFILL_3__13420_ gnd vdd FILL
XFILL_5__12241_ gnd vdd FILL
XFILL_4__9989_ gnd vdd FILL
XSFILL13880x76050 gnd vdd FILL
XFILL_3__10632_ gnd vdd FILL
X_13696_ _13694_/Y _14071_/B _14030_/C _13696_/D gnd _13696_/Y vdd OAI22X1
XFILL_2__12061_ gnd vdd FILL
XFILL_4__12971_ gnd vdd FILL
XFILL_1__11811_ gnd vdd FILL
XFILL_0__13240_ gnd vdd FILL
XFILL_0__10452_ gnd vdd FILL
XFILL_5__7733_ gnd vdd FILL
XFILL_0_BUFX2_insert710 gnd vdd FILL
XFILL_6__13531_ gnd vdd FILL
X_12647_ _12647_/A vdd _12647_/C gnd _12689_/D vdd OAI21X1
XFILL_0_BUFX2_insert721 gnd vdd FILL
XFILL_4__14710_ gnd vdd FILL
X_15435_ _13920_/A _15863_/A gnd _15440_/A vdd NAND2X1
XFILL_3__13351_ gnd vdd FILL
XFILL_0_BUFX2_insert732 gnd vdd FILL
XFILL_4__11922_ gnd vdd FILL
XFILL_5__12172_ gnd vdd FILL
XFILL_2__11012_ gnd vdd FILL
XFILL_4__15690_ gnd vdd FILL
XFILL_1__14530_ gnd vdd FILL
XFILL_3__10563_ gnd vdd FILL
XSFILL94360x74050 gnd vdd FILL
XFILL_0__13171_ gnd vdd FILL
XFILL_0_BUFX2_insert743 gnd vdd FILL
XFILL_2__7955_ gnd vdd FILL
XFILL_1__11742_ gnd vdd FILL
XFILL_0_CLKBUF1_insert180 gnd vdd FILL
XFILL_0__10383_ gnd vdd FILL
XFILL_0_BUFX2_insert754 gnd vdd FILL
XFILL_0_CLKBUF1_insert191 gnd vdd FILL
X_15366_ _15364_/Y _15981_/B _15922_/C _15366_/D gnd _15367_/A vdd OAI22X1
XFILL_0_BUFX2_insert765 gnd vdd FILL
XFILL_3__12302_ gnd vdd FILL
XFILL_5__11123_ gnd vdd FILL
XFILL_4__14641_ gnd vdd FILL
X_12578_ _12578_/A vdd _12577_/Y gnd _12666_/D vdd OAI21X1
XFILL_0_BUFX2_insert776 gnd vdd FILL
XFILL_0__6970_ gnd vdd FILL
XFILL_3__16070_ gnd vdd FILL
XFILL_3__13282_ gnd vdd FILL
XFILL_2__15820_ gnd vdd FILL
XFILL_2__6906_ gnd vdd FILL
XFILL_0__12122_ gnd vdd FILL
XFILL_4__11853_ gnd vdd FILL
XFILL_2__7886_ gnd vdd FILL
XFILL_1__14461_ gnd vdd FILL
XFILL_5__9403_ gnd vdd FILL
XFILL_0_BUFX2_insert787 gnd vdd FILL
XFILL_3__10494_ gnd vdd FILL
XSFILL99400x11050 gnd vdd FILL
XFILL_6__12413_ gnd vdd FILL
XSFILL69160x50050 gnd vdd FILL
XFILL_0_BUFX2_insert798 gnd vdd FILL
XFILL_1__11673_ gnd vdd FILL
XFILL_6__16181_ gnd vdd FILL
XFILL_3__15021_ gnd vdd FILL
XFILL_5__15931_ gnd vdd FILL
X_14317_ _14316_/Y _13775_/B _14317_/C _15795_/A gnd _14317_/Y vdd OAI22X1
XFILL_5__7595_ gnd vdd FILL
X_11529_ _11529_/A _11509_/B _11495_/C _11105_/Y gnd _11529_/Y vdd AOI22X1
X_15297_ _10716_/Q _15916_/B gnd _15297_/Y vdd NAND2X1
XFILL_1__16200_ gnd vdd FILL
XFILL_6__13393_ gnd vdd FILL
XFILL_3__12233_ gnd vdd FILL
XFILL_5__11054_ gnd vdd FILL
XFILL_4__10804_ gnd vdd FILL
XFILL_2__6837_ gnd vdd FILL
XFILL_4__14572_ gnd vdd FILL
XFILL_1__13412_ gnd vdd FILL
XFILL_2__9625_ gnd vdd FILL
XFILL_1__10624_ gnd vdd FILL
XFILL_2__12963_ gnd vdd FILL
XFILL_0__12053_ gnd vdd FILL
XFILL_2__15751_ gnd vdd FILL
XFILL_4__11784_ gnd vdd FILL
XFILL_5__9334_ gnd vdd FILL
XFILL_1__14392_ gnd vdd FILL
XFILL_6__15132_ gnd vdd FILL
X_14248_ _7590_/A gnd _14248_/Y vdd INVX1
XFILL_0__8640_ gnd vdd FILL
XSFILL48840x49050 gnd vdd FILL
XFILL_4__16311_ gnd vdd FILL
XFILL_5__10005_ gnd vdd FILL
XFILL_4__13523_ gnd vdd FILL
XFILL_5__15862_ gnd vdd FILL
XFILL_2__11914_ gnd vdd FILL
XFILL_3__12164_ gnd vdd FILL
XFILL_2__14702_ gnd vdd FILL
XFILL_1__16131_ gnd vdd FILL
XFILL_0__11004_ gnd vdd FILL
XFILL_1__13343_ gnd vdd FILL
XFILL_2__15682_ gnd vdd FILL
XFILL_2__9556_ gnd vdd FILL
XFILL_2__12894_ gnd vdd FILL
XFILL_1__10555_ gnd vdd FILL
XFILL_5__14813_ gnd vdd FILL
XFILL_5__9265_ gnd vdd FILL
X_14179_ _14179_/A _14179_/B _14178_/Y gnd _14179_/Y vdd NOR3X1
XFILL_4__16242_ gnd vdd FILL
XFILL_3__7300_ gnd vdd FILL
XFILL_6__12275_ gnd vdd FILL
XFILL_0__8571_ gnd vdd FILL
XFILL_3__11115_ gnd vdd FILL
XFILL_2__8507_ gnd vdd FILL
XFILL_2__14633_ gnd vdd FILL
XFILL_4__13454_ gnd vdd FILL
XFILL_5__15793_ gnd vdd FILL
XFILL_2__9487_ gnd vdd FILL
XFILL_3__12095_ gnd vdd FILL
XFILL_0__15812_ gnd vdd FILL
XFILL_4__10666_ gnd vdd FILL
XFILL_1__16062_ gnd vdd FILL
XFILL_2__11845_ gnd vdd FILL
XFILL_1__13274_ gnd vdd FILL
XFILL_5__8216_ gnd vdd FILL
XFILL_1__10486_ gnd vdd FILL
XFILL_6__11226_ gnd vdd FILL
XSFILL89320x63050 gnd vdd FILL
XFILL_4__12405_ gnd vdd FILL
XFILL_5__14744_ gnd vdd FILL
XFILL_3__7231_ gnd vdd FILL
XFILL_3__15923_ gnd vdd FILL
XFILL_4__16173_ gnd vdd FILL
XFILL_5__11956_ gnd vdd FILL
XFILL_1__15013_ gnd vdd FILL
XFILL_2__8438_ gnd vdd FILL
XFILL_3__11046_ gnd vdd FILL
XFILL_2__14564_ gnd vdd FILL
XFILL_4__13385_ gnd vdd FILL
XFILL_1__12225_ gnd vdd FILL
XSFILL109480x69050 gnd vdd FILL
XFILL_2__11776_ gnd vdd FILL
XFILL_0__15743_ gnd vdd FILL
XFILL_5__8147_ gnd vdd FILL
XFILL_0__12955_ gnd vdd FILL
XFILL_5__10907_ gnd vdd FILL
XSFILL3800x66050 gnd vdd FILL
XFILL_0__7453_ gnd vdd FILL
XFILL_4__15124_ gnd vdd FILL
XFILL_2__16303_ gnd vdd FILL
XFILL_4__12336_ gnd vdd FILL
XFILL_5__14675_ gnd vdd FILL
XFILL_2__13515_ gnd vdd FILL
XFILL_5__11887_ gnd vdd FILL
XFILL_3__15854_ gnd vdd FILL
XFILL_2__8369_ gnd vdd FILL
XFILL_3__7162_ gnd vdd FILL
XFILL_2__14495_ gnd vdd FILL
XFILL_0__11906_ gnd vdd FILL
XSFILL54040x49050 gnd vdd FILL
XFILL_1__12156_ gnd vdd FILL
XFILL_5__8078_ gnd vdd FILL
XFILL_0__15674_ gnd vdd FILL
XFILL_5__16414_ gnd vdd FILL
XFILL_5__13626_ gnd vdd FILL
XFILL_0__12886_ gnd vdd FILL
X_9820_ _9820_/Q _9436_/CLK _8156_/R vdd _9738_/Y gnd vdd DFFSR
XFILL_3__14805_ gnd vdd FILL
XSFILL94440x54050 gnd vdd FILL
XFILL_4__15055_ gnd vdd FILL
XFILL_6__11088_ gnd vdd FILL
XFILL_2__16234_ gnd vdd FILL
XFILL_2__13446_ gnd vdd FILL
XFILL_4__12267_ gnd vdd FILL
XFILL_1__11107_ gnd vdd FILL
XFILL_3__7093_ gnd vdd FILL
XFILL_0__14625_ gnd vdd FILL
XFILL_2__10658_ gnd vdd FILL
XFILL_3__15785_ gnd vdd FILL
XFILL_0__9123_ gnd vdd FILL
XFILL_3__12997_ gnd vdd FILL
XFILL_1__12087_ gnd vdd FILL
XFILL_0__11837_ gnd vdd FILL
XFILL_5__16345_ gnd vdd FILL
XFILL_4__14006_ gnd vdd FILL
X_9751_ _9751_/A gnd _9751_/Y vdd INVX1
XFILL_5__13557_ gnd vdd FILL
XFILL_4__11218_ gnd vdd FILL
XFILL_2__16165_ gnd vdd FILL
XFILL_3__14736_ gnd vdd FILL
XSFILL69240x30050 gnd vdd FILL
XFILL_4__12198_ gnd vdd FILL
XFILL_5__10769_ gnd vdd FILL
X_6963_ _6985_/B _8243_/B gnd _6963_/Y vdd NAND2X1
XFILL_1__15915_ gnd vdd FILL
XFILL_2__13377_ gnd vdd FILL
XFILL_3__11948_ gnd vdd FILL
XFILL_1__11038_ gnd vdd FILL
XFILL_0__14556_ gnd vdd FILL
XFILL_5__12508_ gnd vdd FILL
X_8702_ _8702_/A _8698_/A _8701_/Y gnd _8792_/D vdd OAI21X1
XFILL_0__11768_ gnd vdd FILL
XFILL_4__11149_ gnd vdd FILL
XFILL_2__15116_ gnd vdd FILL
XFILL_5__16276_ gnd vdd FILL
XFILL_2__12328_ gnd vdd FILL
XFILL_5__13488_ gnd vdd FILL
X_9682_ _9680_/Y _9652_/B _9682_/C gnd _9682_/Y vdd OAI21X1
X_6894_ _6894_/A gnd memoryWriteData[24] vdd BUFX2
XFILL_2__16096_ gnd vdd FILL
XSFILL48920x29050 gnd vdd FILL
XFILL_3__14667_ gnd vdd FILL
XFILL_0__13507_ gnd vdd FILL
XFILL_3__11879_ gnd vdd FILL
XFILL_0__8005_ gnd vdd FILL
XFILL_1__15846_ gnd vdd FILL
XFILL_0__14487_ gnd vdd FILL
XFILL_5__15227_ gnd vdd FILL
X_8633_ _8589_/B _8377_/B gnd _8634_/C vdd NAND2X1
XFILL_5__12439_ gnd vdd FILL
XFILL_3__16406_ gnd vdd FILL
XFILL_0__11699_ gnd vdd FILL
XFILL_3__13618_ gnd vdd FILL
XFILL_3__9803_ gnd vdd FILL
XFILL_4__15957_ gnd vdd FILL
XFILL_2__15047_ gnd vdd FILL
XFILL_0__16226_ gnd vdd FILL
XFILL_2__12259_ gnd vdd FILL
XFILL_3__14598_ gnd vdd FILL
XFILL_1__15777_ gnd vdd FILL
XFILL_0__13438_ gnd vdd FILL
XFILL_3__7995_ gnd vdd FILL
XFILL_1__12989_ gnd vdd FILL
XSFILL49000x38050 gnd vdd FILL
XFILL_5__15158_ gnd vdd FILL
XFILL_4__14908_ gnd vdd FILL
XFILL_5_BUFX2_insert904 gnd vdd FILL
XFILL_3__16337_ gnd vdd FILL
X_8564_ _8564_/Q _9578_/CLK _9460_/R vdd _8564_/D gnd vdd DFFSR
XFILL_1__14728_ gnd vdd FILL
XFILL_5_BUFX2_insert915 gnd vdd FILL
XFILL_3__13549_ gnd vdd FILL
XFILL_3__9734_ gnd vdd FILL
XFILL_4__15888_ gnd vdd FILL
XSFILL59160x82050 gnd vdd FILL
XFILL_3__6946_ gnd vdd FILL
XFILL_5_BUFX2_insert926 gnd vdd FILL
XFILL_0__16157_ gnd vdd FILL
XFILL_0__13369_ gnd vdd FILL
XFILL_5_BUFX2_insert937 gnd vdd FILL
XFILL_5__14109_ gnd vdd FILL
XFILL_5_BUFX2_insert948 gnd vdd FILL
X_7515_ _7515_/Q _7515_/CLK _7515_/R vdd _7515_/D gnd vdd DFFSR
XFILL_4__14839_ gnd vdd FILL
XSFILL109560x49050 gnd vdd FILL
XFILL_5__15089_ gnd vdd FILL
X_8495_ _8495_/A gnd _8495_/Y vdd INVX1
XFILL_5_BUFX2_insert959 gnd vdd FILL
XFILL_3__16268_ gnd vdd FILL
XFILL_0__15108_ gnd vdd FILL
XFILL_3__6877_ gnd vdd FILL
XFILL_3__9665_ gnd vdd FILL
XFILL_1__14659_ gnd vdd FILL
XFILL_0__16088_ gnd vdd FILL
XFILL_1__7700_ gnd vdd FILL
XFILL_0__8907_ gnd vdd FILL
XFILL_6__9374_ gnd vdd FILL
XFILL_3__15219_ gnd vdd FILL
XSFILL54120x29050 gnd vdd FILL
X_7446_ _7446_/A _7472_/A _7445_/Y gnd _7520_/D vdd OAI21X1
XFILL_3__8616_ gnd vdd FILL
XFILL_0__9887_ gnd vdd FILL
XFILL_3__16199_ gnd vdd FILL
XFILL_0__15039_ gnd vdd FILL
XFILL_2__15949_ gnd vdd FILL
XFILL_3__9596_ gnd vdd FILL
XFILL_6__8325_ gnd vdd FILL
XFILL_1__7631_ gnd vdd FILL
XSFILL79080x33050 gnd vdd FILL
XFILL_0__8838_ gnd vdd FILL
XFILL_4__7340_ gnd vdd FILL
XFILL_1__16329_ gnd vdd FILL
X_7377_ _7366_/B _9041_/B gnd _7378_/C vdd NAND2X1
XSFILL13720x3050 gnd vdd FILL
X_9116_ _9114_/Y _9116_/B _9116_/C gnd _9116_/Y vdd OAI21X1
XFILL_1__7562_ gnd vdd FILL
XFILL_0__8769_ gnd vdd FILL
XFILL_3_BUFX2_insert105 gnd vdd FILL
XFILL_3__8478_ gnd vdd FILL
XFILL_1__9301_ gnd vdd FILL
X_9047_ _9047_/Q _6999_/CLK _7000_/R vdd _9047_/D gnd vdd DFFSR
XFILL_4__9010_ gnd vdd FILL
XSFILL8600x58050 gnd vdd FILL
XFILL_1__7493_ gnd vdd FILL
XFILL_3__7429_ gnd vdd FILL
XSFILL58360x34050 gnd vdd FILL
XFILL_1__9232_ gnd vdd FILL
XCLKBUF1_insert1083 clk gnd CLKBUF1_insert187/A vdd CLKBUF1
XFILL_2_BUFX2_insert805 gnd vdd FILL
XFILL_2_BUFX2_insert816 gnd vdd FILL
XFILL_2_BUFX2_insert827 gnd vdd FILL
XFILL_6__7069_ gnd vdd FILL
XFILL_2_BUFX2_insert838 gnd vdd FILL
XFILL_1__9163_ gnd vdd FILL
XFILL_2_BUFX2_insert849 gnd vdd FILL
X_10900_ _10984_/Q _10903_/A gnd _10929_/A vdd NAND2X1
XFILL_0_BUFX2_insert60 gnd vdd FILL
XFILL_1__8114_ gnd vdd FILL
X_11880_ _11880_/A _11874_/B _11879_/Y gnd _13215_/A vdd OAI21X1
X_9949_ _9949_/Q _9707_/CLK _8819_/R vdd _9869_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert71 gnd vdd FILL
XFILL_1__9094_ gnd vdd FILL
XFILL111960x61050 gnd vdd FILL
XFILL_0_BUFX2_insert82 gnd vdd FILL
XFILL_4__9912_ gnd vdd FILL
XFILL112440x68050 gnd vdd FILL
XFILL_0_BUFX2_insert93 gnd vdd FILL
X_10831_ _10831_/A _10831_/B _10830_/Y gnd _10831_/Y vdd OAI21X1
XSFILL109240x31050 gnd vdd FILL
X_13550_ _15145_/B _14778_/B _14342_/B _15157_/B gnd _13551_/B vdd OAI22X1
XSFILL79160x13050 gnd vdd FILL
X_10762_ _10760_/Y _10762_/B _10762_/C gnd _10844_/D vdd OAI21X1
XBUFX2_insert804 _15091_/Y gnd _16294_/C vdd BUFX2
X_12501_ _12499_/Y vdd _12500_/Y gnd _12555_/D vdd OAI21X1
XBUFX2_insert815 _13329_/Y gnd _9017_/A vdd BUFX2
XFILL_4__9774_ gnd vdd FILL
XBUFX2_insert826 _13287_/Y gnd _7430_/A vdd BUFX2
XFILL_4__6986_ gnd vdd FILL
XFILL_6_BUFX2_insert771 gnd vdd FILL
X_13481_ _8057_/A gnd _15110_/C vdd INVX1
X_10693_ _10658_/B _7877_/B gnd _10693_/Y vdd NAND2X1
XBUFX2_insert837 _13324_/Y gnd _8619_/B vdd BUFX2
XBUFX2_insert848 _13269_/Y gnd _7061_/A vdd BUFX2
XFILL_1__9996_ gnd vdd FILL
X_15220_ _12812_/Q _15220_/B gnd _15220_/Y vdd NAND2X1
XBUFX2_insert859 _13314_/Y gnd _8237_/A vdd BUFX2
XFILL_4__8725_ gnd vdd FILL
X_12432_ _12430_/Y _12407_/A _12432_/C gnd _12432_/Y vdd OAI21X1
XSFILL18840x28050 gnd vdd FILL
XFILL_2__7740_ gnd vdd FILL
X_15151_ _9340_/A _15114_/C _15764_/C gnd _15152_/C vdd NAND3X1
XFILL_4__8656_ gnd vdd FILL
X_12363_ _12361_/Y _12380_/A _12363_/C gnd _12363_/Y vdd OAI21X1
XSFILL69080x65050 gnd vdd FILL
XFILL_1_CLKBUF1_insert220 gnd vdd FILL
XSFILL99320x26050 gnd vdd FILL
XFILL_2__7671_ gnd vdd FILL
XFILL_4__7607_ gnd vdd FILL
XFILL_1__8878_ gnd vdd FILL
X_14102_ _9245_/A gnd _15595_/A vdd INVX1
XFILL_5__7380_ gnd vdd FILL
X_11314_ _11105_/Y gnd _11531_/A vdd INVX1
XFILL_4__8587_ gnd vdd FILL
X_15082_ _8023_/Q _15081_/Y gnd _15085_/A vdd NAND2X1
X_12294_ _12294_/A _12292_/Y _12293_/Y gnd _12294_/Y vdd NAND3X1
XFILL_2__9410_ gnd vdd FILL
XFILL_1__7829_ gnd vdd FILL
X_14033_ _10138_/A gnd _14033_/Y vdd INVX1
X_11245_ _11384_/A _12138_/Y gnd _11245_/Y vdd XOR2X1
XFILL_4__10520_ gnd vdd FILL
XFILL_2__9341_ gnd vdd FILL
XSFILL109320x11050 gnd vdd FILL
XFILL_6__12060_ gnd vdd FILL
XFILL_4__7469_ gnd vdd FILL
XFILL_5__11810_ gnd vdd FILL
XSFILL23800x83050 gnd vdd FILL
XFILL_4__10451_ gnd vdd FILL
X_11176_ _12192_/Y _12318_/Y gnd _11176_/Y vdd NOR2X1
XFILL_5__12790_ gnd vdd FILL
XFILL_2__9272_ gnd vdd FILL
XFILL_2__11630_ gnd vdd FILL
XSFILL89240x78050 gnd vdd FILL
XFILL_4__9208_ gnd vdd FILL
XFILL_1__10271_ gnd vdd FILL
XFILL_5__8001_ gnd vdd FILL
XFILL112120x50050 gnd vdd FILL
XFILL_3_BUFX2_insert650 gnd vdd FILL
XFILL_6__11011_ gnd vdd FILL
X_10127_ _10127_/A _9615_/B gnd _10128_/C vdd NAND2X1
XFILL_3_BUFX2_insert661 gnd vdd FILL
XFILL_4__13170_ gnd vdd FILL
XFILL_2__8223_ gnd vdd FILL
XFILL_5__11741_ gnd vdd FILL
XFILL_4__10382_ gnd vdd FILL
X_15984_ _15984_/A _15984_/B gnd _16006_/A vdd NOR2X1
XFILL_3_BUFX2_insert672 gnd vdd FILL
XFILL_1__12010_ gnd vdd FILL
XFILL_2__11561_ gnd vdd FILL
XFILL_3_BUFX2_insert683 gnd vdd FILL
XFILL_0__12740_ gnd vdd FILL
XFILL_3_BUFX2_insert694 gnd vdd FILL
XFILL_4__9139_ gnd vdd FILL
XFILL_2__13300_ gnd vdd FILL
XFILL_5__14460_ gnd vdd FILL
X_10058_ _10098_/Q gnd _10058_/Y vdd INVX1
XFILL_4__12121_ gnd vdd FILL
X_14935_ _9555_/A gnd _14937_/D vdd INVX1
XFILL_2__10512_ gnd vdd FILL
XFILL_5__11672_ gnd vdd FILL
XFILL_3__12851_ gnd vdd FILL
XFILL_2__14280_ gnd vdd FILL
XSFILL94360x69050 gnd vdd FILL
XFILL_2__11492_ gnd vdd FILL
XFILL_5__13411_ gnd vdd FILL
XFILL_5__10623_ gnd vdd FILL
XFILL_4__12052_ gnd vdd FILL
XFILL_2__7105_ gnd vdd FILL
XFILL_2__13231_ gnd vdd FILL
X_14866_ _14866_/A _14866_/B gnd _14869_/C vdd NOR2X1
XFILL_5__14391_ gnd vdd FILL
XFILL_3__11802_ gnd vdd FILL
XFILL_3__12782_ gnd vdd FILL
XFILL_2__10443_ gnd vdd FILL
XFILL_3__15570_ gnd vdd FILL
XFILL_0__14410_ gnd vdd FILL
XFILL_2__8085_ gnd vdd FILL
XFILL_5__8903_ gnd vdd FILL
XFILL_0__11622_ gnd vdd FILL
XFILL_1__13961_ gnd vdd FILL
XFILL_0__15390_ gnd vdd FILL
XSFILL69160x45050 gnd vdd FILL
XFILL_5__16130_ gnd vdd FILL
XFILL_4__11003_ gnd vdd FILL
XFILL_5__13342_ gnd vdd FILL
X_13817_ _13865_/C _7773_/Q _7645_/Q _13848_/C gnd _13826_/A vdd AOI22X1
XFILL_5__9883_ gnd vdd FILL
XFILL_3__14521_ gnd vdd FILL
XFILL_5__10554_ gnd vdd FILL
XFILL_2__7036_ gnd vdd FILL
XFILL_1__15700_ gnd vdd FILL
XFILL_1__12912_ gnd vdd FILL
X_14797_ _10186_/A gnd _14797_/Y vdd INVX1
XFILL_2__13162_ gnd vdd FILL
XFILL_3__11733_ gnd vdd FILL
XFILL_0__14341_ gnd vdd FILL
XFILL_2__10374_ gnd vdd FILL
XFILL_5__8834_ gnd vdd FILL
XFILL_1__13892_ gnd vdd FILL
XFILL_0__11553_ gnd vdd FILL
XFILL_4__15811_ gnd vdd FILL
XFILL_5__16061_ gnd vdd FILL
XFILL_5__13273_ gnd vdd FILL
X_13748_ _15307_/D _14615_/B _13857_/C _15299_/B gnd _13749_/B vdd OAI22X1
XFILL_2__12113_ gnd vdd FILL
XFILL_3__14452_ gnd vdd FILL
XFILL_1__15631_ gnd vdd FILL
XFILL_3__11664_ gnd vdd FILL
XFILL_0__10504_ gnd vdd FILL
XFILL_1__12843_ gnd vdd FILL
XFILL_2__13093_ gnd vdd FILL
XFILL_5__15012_ gnd vdd FILL
XFILL_0__11484_ gnd vdd FILL
XFILL_0__14272_ gnd vdd FILL
XFILL_5__8765_ gnd vdd FILL
XFILL_5__12224_ gnd vdd FILL
XFILL_3__13403_ gnd vdd FILL
XFILL_3__10615_ gnd vdd FILL
XFILL_4__15742_ gnd vdd FILL
XFILL_0__16011_ gnd vdd FILL
X_13679_ _13679_/A gnd _13679_/Y vdd INVX1
XFILL_2__12044_ gnd vdd FILL
XFILL_4__12954_ gnd vdd FILL
XFILL_0__13223_ gnd vdd FILL
XFILL_1__15562_ gnd vdd FILL
XFILL_3__14383_ gnd vdd FILL
XFILL_3__11595_ gnd vdd FILL
XFILL_1__12774_ gnd vdd FILL
XFILL_5__7716_ gnd vdd FILL
XFILL_2__8987_ gnd vdd FILL
XFILL_0__10435_ gnd vdd FILL
XFILL_0_BUFX2_insert540 gnd vdd FILL
XFILL_0_BUFX2_insert551 gnd vdd FILL
X_15418_ _15417_/Y _15656_/B _15656_/C gnd _15421_/B vdd NOR3X1
XFILL_0__9810_ gnd vdd FILL
XSFILL89320x58050 gnd vdd FILL
XFILL_4__11905_ gnd vdd FILL
XFILL_5__8696_ gnd vdd FILL
XFILL_3__16122_ gnd vdd FILL
XFILL_5__12155_ gnd vdd FILL
XFILL_3__13334_ gnd vdd FILL
XFILL_4__15673_ gnd vdd FILL
XFILL_0_BUFX2_insert562 gnd vdd FILL
XFILL_1__14513_ gnd vdd FILL
XFILL112200x30050 gnd vdd FILL
X_16398_ _16396_/Y gnd _16398_/C gnd _16398_/Y vdd OAI21X1
XFILL_3__10546_ gnd vdd FILL
XFILL_2__7938_ gnd vdd FILL
XFILL_0_BUFX2_insert573 gnd vdd FILL
XFILL_1__11725_ gnd vdd FILL
XFILL_4__12885_ gnd vdd FILL
XFILL_0_BUFX2_insert584 gnd vdd FILL
XFILL_0__13154_ gnd vdd FILL
XFILL_0__10366_ gnd vdd FILL
XFILL_1__15493_ gnd vdd FILL
XFILL_0_BUFX2_insert595 gnd vdd FILL
X_7300_ _7300_/A _7308_/A _7299_/Y gnd _7386_/D vdd OAI21X1
XFILL_5__11106_ gnd vdd FILL
X_15349_ _7005_/Q _15382_/B _16096_/C _7389_/Q gnd _15354_/A vdd AOI22X1
XFILL_0__9741_ gnd vdd FILL
XFILL_4__14624_ gnd vdd FILL
XFILL_6__10657_ gnd vdd FILL
XFILL_0__6953_ gnd vdd FILL
XFILL_3__13265_ gnd vdd FILL
XFILL_5__12086_ gnd vdd FILL
XFILL_2__15803_ gnd vdd FILL
X_8280_ _8280_/Q _6999_/CLK _7000_/R vdd _8280_/D gnd vdd DFFSR
XFILL_3__16053_ gnd vdd FILL
XFILL_4__11836_ gnd vdd FILL
XFILL_0__12105_ gnd vdd FILL
XFILL_1__14444_ gnd vdd FILL
XFILL_2__7869_ gnd vdd FILL
XFILL_1__11656_ gnd vdd FILL
XFILL_0__13085_ gnd vdd FILL
XFILL_2__13995_ gnd vdd FILL
XFILL_0__10297_ gnd vdd FILL
X_7231_ _7184_/B _7231_/B gnd _7232_/C vdd NAND2X1
XFILL_5__15914_ gnd vdd FILL
XFILL_5__7578_ gnd vdd FILL
XFILL_0__9672_ gnd vdd FILL
XFILL_3__12216_ gnd vdd FILL
XFILL_5__11037_ gnd vdd FILL
XFILL_3__15004_ gnd vdd FILL
XFILL_2__9608_ gnd vdd FILL
XFILL_4__14555_ gnd vdd FILL
XSFILL94440x49050 gnd vdd FILL
XFILL_0__6884_ gnd vdd FILL
XSFILL43800x14050 gnd vdd FILL
XFILL_3__8401_ gnd vdd FILL
XFILL_3__9381_ gnd vdd FILL
XFILL_4__11767_ gnd vdd FILL
XFILL_2__15734_ gnd vdd FILL
XFILL_0__12036_ gnd vdd FILL
XFILL_1__14375_ gnd vdd FILL
XFILL_6__9090_ gnd vdd FILL
XFILL_0__8623_ gnd vdd FILL
XFILL_1__11587_ gnd vdd FILL
XFILL_4__13506_ gnd vdd FILL
XFILL_3__8332_ gnd vdd FILL
XFILL_5__15845_ gnd vdd FILL
XFILL_1__16114_ gnd vdd FILL
XFILL_3__12147_ gnd vdd FILL
X_7162_ _7210_/A _9466_/B gnd _7163_/C vdd NAND2X1
XFILL_1__13326_ gnd vdd FILL
XFILL_4__14486_ gnd vdd FILL
XFILL_2__9539_ gnd vdd FILL
XSFILL69240x25050 gnd vdd FILL
XFILL_2__15665_ gnd vdd FILL
XFILL_2__12877_ gnd vdd FILL
XFILL_4__11698_ gnd vdd FILL
XFILL_1__10538_ gnd vdd FILL
XFILL_5__9248_ gnd vdd FILL
XFILL_4__16225_ gnd vdd FILL
X_7093_ _7093_/A gnd _7095_/A vdd INVX1
XFILL_4__13437_ gnd vdd FILL
XFILL_5__15776_ gnd vdd FILL
XFILL_1__16045_ gnd vdd FILL
XFILL_2__14616_ gnd vdd FILL
XFILL_3__12078_ gnd vdd FILL
XFILL_4__10649_ gnd vdd FILL
XFILL_5__12988_ gnd vdd FILL
XFILL_2__11828_ gnd vdd FILL
XFILL_3__8263_ gnd vdd FILL
XFILL_1__13257_ gnd vdd FILL
XSFILL104440x34050 gnd vdd FILL
XFILL_2__15596_ gnd vdd FILL
XFILL_0__7505_ gnd vdd FILL
XFILL_0__13987_ gnd vdd FILL
XFILL_5__14727_ gnd vdd FILL
XFILL_3__15906_ gnd vdd FILL
XFILL_0__8485_ gnd vdd FILL
XFILL_3__7214_ gnd vdd FILL
XFILL_5__11939_ gnd vdd FILL
XFILL_3__11029_ gnd vdd FILL
XFILL_4__16156_ gnd vdd FILL
XFILL_4__13368_ gnd vdd FILL
XFILL_1__12208_ gnd vdd FILL
XSFILL8680x32050 gnd vdd FILL
XFILL_0__15726_ gnd vdd FILL
XFILL_3__8194_ gnd vdd FILL
XFILL_2__14547_ gnd vdd FILL
XFILL_2__11759_ gnd vdd FILL
XFILL_0__7436_ gnd vdd FILL
XFILL_4__15107_ gnd vdd FILL
XFILL_4__12319_ gnd vdd FILL
XFILL_5__14658_ gnd vdd FILL
XFILL_3__15837_ gnd vdd FILL
XFILL_4__16087_ gnd vdd FILL
XFILL_4__13299_ gnd vdd FILL
XFILL_2__14478_ gnd vdd FILL
XFILL_1__12139_ gnd vdd FILL
XFILL_0__15657_ gnd vdd FILL
XSFILL89400x38050 gnd vdd FILL
XFILL_5__13609_ gnd vdd FILL
XFILL_0__12869_ gnd vdd FILL
X_9803_ _9737_/A _9803_/B gnd _9804_/C vdd NAND2X1
XFILL_4__15038_ gnd vdd FILL
XFILL_0__7367_ gnd vdd FILL
XFILL_5__14589_ gnd vdd FILL
XFILL_2__16217_ gnd vdd FILL
XFILL_2__13429_ gnd vdd FILL
XFILL_3__7076_ gnd vdd FILL
XFILL_0__14608_ gnd vdd FILL
X_7995_ _8045_/Q gnd _7995_/Y vdd INVX1
XFILL_3__15768_ gnd vdd FILL
XFILL_0__9106_ gnd vdd FILL
XFILL111880x76050 gnd vdd FILL
XFILL_5__16328_ gnd vdd FILL
XFILL_0__15588_ gnd vdd FILL
X_9734_ _9770_/A _8582_/B gnd _9735_/C vdd NAND2X1
XFILL_0__7298_ gnd vdd FILL
X_6946_ _6946_/A _6967_/B _6946_/C gnd _7012_/D vdd OAI21X1
XFILL_3__14719_ gnd vdd FILL
XFILL_6__15879_ gnd vdd FILL
XFILL_2__16148_ gnd vdd FILL
XFILL_3__15699_ gnd vdd FILL
XFILL_0__14539_ gnd vdd FILL
XFILL_0__9037_ gnd vdd FILL
XSFILL13640x33050 gnd vdd FILL
XFILL_5__16259_ gnd vdd FILL
X_9665_ _9711_/Q gnd _9665_/Y vdd INVX1
X_6877_ _6877_/A gnd memoryWriteData[7] vdd BUFX2
XFILL_2__16079_ gnd vdd FILL
XFILL_4__6840_ gnd vdd FILL
XFILL_1__15829_ gnd vdd FILL
X_8616_ _8614_/Y _8655_/B _8615_/Y gnd _8678_/D vdd OAI21X1
XFILL_6__7756_ gnd vdd FILL
XFILL_1__9850_ gnd vdd FILL
XFILL_0__16209_ gnd vdd FILL
X_9596_ _9596_/A gnd _9596_/Y vdd INVX1
XFILL_5_BUFX2_insert701 gnd vdd FILL
XFILL_5_BUFX2_insert712 gnd vdd FILL
XFILL_3__7978_ gnd vdd FILL
XFILL_5_BUFX2_insert723 gnd vdd FILL
XFILL_5_BUFX2_insert734 gnd vdd FILL
X_8547_ _8477_/A _7651_/CLK _7011_/R vdd _8547_/D gnd vdd DFFSR
XFILL_1__9781_ gnd vdd FILL
XFILL_4__8510_ gnd vdd FILL
XFILL_5_BUFX2_insert745 gnd vdd FILL
XSFILL104520x14050 gnd vdd FILL
XFILL_1__6993_ gnd vdd FILL
XFILL_5_BUFX2_insert756 gnd vdd FILL
XFILL_3__6929_ gnd vdd FILL
XFILL_5_BUFX2_insert767 gnd vdd FILL
XFILL_4__9490_ gnd vdd FILL
XSFILL8760x12050 gnd vdd FILL
XFILL_5_BUFX2_insert778 gnd vdd FILL
XSFILL33800x46050 gnd vdd FILL
XFILL_1__8732_ gnd vdd FILL
XFILL_0__9939_ gnd vdd FILL
XFILL_5_BUFX2_insert789 gnd vdd FILL
X_8478_ _8469_/A _8606_/B gnd _8479_/C vdd NAND2X1
XFILL_3__9648_ gnd vdd FILL
XFILL_4__8441_ gnd vdd FILL
X_7429_ _7515_/Q gnd _7429_/Y vdd INVX1
XFILL_4__8372_ gnd vdd FILL
XSFILL23880x4050 gnd vdd FILL
XFILL_1__7614_ gnd vdd FILL
XFILL_1__8594_ gnd vdd FILL
XFILL111960x56050 gnd vdd FILL
XFILL_4__7323_ gnd vdd FILL
X_11030_ _11030_/A gnd _11031_/B vdd INVX1
XFILL_1__7545_ gnd vdd FILL
XSFILL63880x41050 gnd vdd FILL
XSFILL13720x13050 gnd vdd FILL
XFILL112040x65050 gnd vdd FILL
XFILL_1__7476_ gnd vdd FILL
XFILL_2_BUFX2_insert602 gnd vdd FILL
XFILL_4__7185_ gnd vdd FILL
XFILL_2_BUFX2_insert613 gnd vdd FILL
XFILL_1__9215_ gnd vdd FILL
X_12981_ _6880_/A gnd _12983_/A vdd INVX1
XFILL_2_BUFX2_insert624 gnd vdd FILL
XFILL_2_BUFX2_insert635 gnd vdd FILL
XFILL_2_BUFX2_insert646 gnd vdd FILL
XFILL_2_BUFX2_insert657 gnd vdd FILL
X_14720_ _8048_/Q gnd _14720_/Y vdd INVX1
X_11932_ _13190_/Q gnd _11934_/A vdd INVX1
XFILL_1__9146_ gnd vdd FILL
XSFILL114600x79050 gnd vdd FILL
XFILL_2_BUFX2_insert668 gnd vdd FILL
XFILL_2_BUFX2_insert679 gnd vdd FILL
X_11863_ _11863_/A _11862_/Y _11860_/Y gnd _11865_/A vdd NOR3X1
X_14651_ _16070_/A gnd _14651_/Y vdd INVX1
X_10814_ _10862_/Q gnd _10814_/Y vdd INVX1
X_13602_ _13602_/A _13602_/B gnd _13602_/Y vdd NOR2X1
XFILL_5_BUFX2_insert17 gnd vdd FILL
XFILL_5__6880_ gnd vdd FILL
XFILL_2__8910_ gnd vdd FILL
X_14582_ _10171_/A gnd _14582_/Y vdd INVX1
X_11794_ _11025_/Y gnd _11794_/Y vdd INVX1
XFILL_5_BUFX2_insert28 gnd vdd FILL
XFILL_2__9890_ gnd vdd FILL
XFILL_5_BUFX2_insert39 gnd vdd FILL
X_16321_ _16417_/Q gnd _16321_/Y vdd INVX1
XBUFX2_insert601 BUFX2_insert494/A gnd _9460_/R vdd BUFX2
XBUFX2_insert612 _10926_/Y gnd _12111_/A vdd BUFX2
X_10745_ _13485_/A gnd _10745_/Y vdd INVX1
X_13533_ _13533_/A _13504_/Y _15812_/C gnd _12955_/B vdd AOI21X1
XBUFX2_insert623 _12363_/Y gnd _9993_/B vdd BUFX2
XFILL_5__10270_ gnd vdd FILL
XBUFX2_insert634 _12354_/Y gnd _8832_/B vdd BUFX2
XFILL_2__8841_ gnd vdd FILL
XBUFX2_insert645 _13424_/Y gnd _14697_/B vdd BUFX2
XFILL_4__9757_ gnd vdd FILL
XBUFX2_insert656 _12429_/Y gnd _7243_/B vdd BUFX2
XFILL_3__10400_ gnd vdd FILL
X_13464_ _7510_/Q gnd _13464_/Y vdd INVX1
XFILL_4__6969_ gnd vdd FILL
X_16252_ _6992_/A _15382_/B _16096_/C _7376_/A gnd _16252_/Y vdd AOI22X1
XSFILL23800x78050 gnd vdd FILL
XSFILL23000x59050 gnd vdd FILL
XBUFX2_insert667 _12345_/Y gnd _8823_/A vdd BUFX2
X_10676_ _10676_/A _10676_/B _10675_/Y gnd _10730_/D vdd OAI21X1
XFILL_3__11380_ gnd vdd FILL
XBUFX2_insert678 _13541_/Y gnd _14273_/C vdd BUFX2
XBUFX2_insert689 _13362_/Y gnd _10535_/A vdd BUFX2
XFILL_5__7501_ gnd vdd FILL
XFILL_4__8708_ gnd vdd FILL
XFILL_2__8772_ gnd vdd FILL
XFILL_1__9979_ gnd vdd FILL
X_12415_ _12083_/B gnd _12415_/Y vdd INVX1
X_15203_ _13599_/Y _15203_/B _15203_/C gnd _15203_/Y vdd OAI21X1
XFILL_5__8481_ gnd vdd FILL
X_16183_ _15394_/C _14809_/B _16183_/C _16026_/D gnd _16184_/A vdd OAI22X1
X_13395_ _8310_/A gnd _13395_/Y vdd INVX1
XFILL_1__11510_ gnd vdd FILL
XFILL_2__7723_ gnd vdd FILL
XFILL_0__10151_ gnd vdd FILL
XSFILL64040x30050 gnd vdd FILL
XFILL_4__8639_ gnd vdd FILL
XFILL_5__7432_ gnd vdd FILL
XFILL_1__12490_ gnd vdd FILL
X_12346_ _11991_/B gnd _12346_/Y vdd INVX1
X_15134_ _13574_/A _15565_/B _15801_/A _15133_/Y gnd _15135_/A vdd OAI22X1
XFILL_4__11621_ gnd vdd FILL
XFILL_5__13960_ gnd vdd FILL
XFILL_3__10262_ gnd vdd FILL
XFILL_2__13780_ gnd vdd FILL
XFILL_1__11441_ gnd vdd FILL
XFILL_2__10992_ gnd vdd FILL
XFILL_5__12911_ gnd vdd FILL
XFILL_3__12001_ gnd vdd FILL
X_15065_ _14986_/A _14982_/Y _15061_/C gnd _15065_/Y vdd NAND3X1
XFILL_6__13161_ gnd vdd FILL
XFILL_5__7363_ gnd vdd FILL
X_12277_ _6885_/A _12277_/B _12309_/C _11879_/B gnd _12278_/C vdd AOI22X1
XFILL_4__14340_ gnd vdd FILL
XFILL_6__10373_ gnd vdd FILL
XFILL_2__12731_ gnd vdd FILL
XFILL_5__13891_ gnd vdd FILL
XFILL_4__11552_ gnd vdd FILL
XFILL_5__9102_ gnd vdd FILL
XFILL_2__7585_ gnd vdd FILL
XFILL_1__14160_ gnd vdd FILL
XFILL_3__10193_ gnd vdd FILL
XFILL_0__13910_ gnd vdd FILL
X_14016_ _14016_/A gnd _14018_/D vdd INVX1
XFILL_1__11372_ gnd vdd FILL
XFILL_5__15630_ gnd vdd FILL
XFILL_5__7294_ gnd vdd FILL
X_11228_ _11214_/Y _10882_/Y _11224_/Y gnd _11228_/Y vdd NAND3X1
XFILL_0__14890_ gnd vdd FILL
XFILL_5__12842_ gnd vdd FILL
XFILL_4__10503_ gnd vdd FILL
XFILL_1__13111_ gnd vdd FILL
XSFILL3640x5050 gnd vdd FILL
XFILL_4__14271_ gnd vdd FILL
XFILL_2__12662_ gnd vdd FILL
XFILL_2__15450_ gnd vdd FILL
XFILL_4__11483_ gnd vdd FILL
XFILL_1__10323_ gnd vdd FILL
XFILL_0__13841_ gnd vdd FILL
XSFILL29160x56050 gnd vdd FILL
XFILL_1__14091_ gnd vdd FILL
XFILL_5__9033_ gnd vdd FILL
XFILL_4__16010_ gnd vdd FILL
XSFILL84200x43050 gnd vdd FILL
XFILL_4__13222_ gnd vdd FILL
XFILL_5__15561_ gnd vdd FILL
X_11159_ _11108_/Y _12302_/Y _11159_/C gnd _11159_/Y vdd OAI21X1
XFILL_5__12773_ gnd vdd FILL
XFILL_2__11613_ gnd vdd FILL
XFILL_2__14401_ gnd vdd FILL
XFILL_4__10434_ gnd vdd FILL
XFILL_2__15381_ gnd vdd FILL
XFILL_2__9255_ gnd vdd FILL
XSFILL104360x49050 gnd vdd FILL
XFILL_3__13952_ gnd vdd FILL
XFILL_1__13042_ gnd vdd FILL
XFILL_2__12593_ gnd vdd FILL
XFILL_1__10254_ gnd vdd FILL
XFILL_3_BUFX2_insert480 gnd vdd FILL
XFILL_0__13772_ gnd vdd FILL
XFILL_5__14512_ gnd vdd FILL
XFILL_0__8270_ gnd vdd FILL
XFILL_5__11724_ gnd vdd FILL
XFILL_3_BUFX2_insert491 gnd vdd FILL
XFILL_2__8206_ gnd vdd FILL
XFILL_4__13153_ gnd vdd FILL
X_15967_ _15955_/Y _15967_/B _15967_/C gnd _15968_/B vdd NOR3X1
XFILL_3__12903_ gnd vdd FILL
XFILL_2__14332_ gnd vdd FILL
XFILL_4__10365_ gnd vdd FILL
XFILL_5__15492_ gnd vdd FILL
XFILL_0__15511_ gnd vdd FILL
XFILL_2__11544_ gnd vdd FILL
XFILL_0__12723_ gnd vdd FILL
XFILL_3__13883_ gnd vdd FILL
XFILL_0__7221_ gnd vdd FILL
XFILL_6__15802_ gnd vdd FILL
XFILL_1__10185_ gnd vdd FILL
XFILL_4__12104_ gnd vdd FILL
X_14918_ _14918_/A gnd _16247_/A vdd INVX1
XFILL_5__14443_ gnd vdd FILL
XFILL_3__15622_ gnd vdd FILL
XFILL_2__8137_ gnd vdd FILL
XFILL_5__11655_ gnd vdd FILL
X_15898_ _9835_/Q gnd _15899_/B vdd INVX1
XFILL_2__14263_ gnd vdd FILL
XFILL_3__12834_ gnd vdd FILL
XFILL_4__10296_ gnd vdd FILL
XFILL_4__13084_ gnd vdd FILL
XFILL112200x25050 gnd vdd FILL
XFILL_2__11475_ gnd vdd FILL
XFILL_0__15442_ gnd vdd FILL
XFILL_0__12654_ gnd vdd FILL
XFILL_5__9935_ gnd vdd FILL
XFILL_1__14993_ gnd vdd FILL
XFILL_2__13214_ gnd vdd FILL
XFILL_2__16002_ gnd vdd FILL
X_14849_ _14849_/A _14849_/B gnd _14850_/C vdd NOR2X1
XFILL_4__12035_ gnd vdd FILL
XFILL_5__14374_ gnd vdd FILL
XSFILL64120x10050 gnd vdd FILL
XFILL_2__8068_ gnd vdd FILL
X_7780_ _7780_/Q _9818_/CLK _9441_/R vdd _7714_/Y gnd vdd DFFSR
XFILL_3__15553_ gnd vdd FILL
XFILL_2__10426_ gnd vdd FILL
XFILL_5__11586_ gnd vdd FILL
XFILL_3__8950_ gnd vdd FILL
XFILL_3__12765_ gnd vdd FILL
XFILL_2__14194_ gnd vdd FILL
XFILL_0__11605_ gnd vdd FILL
XFILL_1__13944_ gnd vdd FILL
XFILL_0__15373_ gnd vdd FILL
XFILL_5__16113_ gnd vdd FILL
XFILL_5__13325_ gnd vdd FILL
XFILL_0__12585_ gnd vdd FILL
XFILL_5__9866_ gnd vdd FILL
XFILL_6__15664_ gnd vdd FILL
XFILL_3__14504_ gnd vdd FILL
XFILL_0__7083_ gnd vdd FILL
XFILL_5__10537_ gnd vdd FILL
XFILL_2__13145_ gnd vdd FILL
XSFILL18680x5050 gnd vdd FILL
XFILL_3__11716_ gnd vdd FILL
XSFILL3400x58050 gnd vdd FILL
XFILL_0__14324_ gnd vdd FILL
XFILL_3__15484_ gnd vdd FILL
XFILL_3__12696_ gnd vdd FILL
XFILL_1__13875_ gnd vdd FILL
XFILL_0__11536_ gnd vdd FILL
XFILL_3__8881_ gnd vdd FILL
XFILL_5__16044_ gnd vdd FILL
XFILL_6__14615_ gnd vdd FILL
XFILL_5__13256_ gnd vdd FILL
XFILL_5__9797_ gnd vdd FILL
X_9450_ _9394_/A _7786_/CLK _7153_/R vdd _9450_/D gnd vdd DFFSR
XFILL_3__14435_ gnd vdd FILL
XFILL_1__15614_ gnd vdd FILL
XFILL_3__7832_ gnd vdd FILL
XFILL_4__13986_ gnd vdd FILL
XFILL_3__11647_ gnd vdd FILL
XFILL_1__12826_ gnd vdd FILL
XFILL_0__14255_ gnd vdd FILL
XFILL_2__10288_ gnd vdd FILL
XFILL_5__8748_ gnd vdd FILL
XFILL_5__12207_ gnd vdd FILL
XFILL_0__11467_ gnd vdd FILL
X_8401_ _8345_/B _8401_/B gnd _8401_/Y vdd NAND2X1
XFILL_4__15725_ gnd vdd FILL
XFILL_6__11758_ gnd vdd FILL
X_9381_ _9381_/A _9359_/A _9380_/Y gnd _9445_/D vdd OAI21X1
XFILL_2__12027_ gnd vdd FILL
XSFILL54040x62050 gnd vdd FILL
XFILL_1__15545_ gnd vdd FILL
XFILL_3__14366_ gnd vdd FILL
XFILL_5__10399_ gnd vdd FILL
XFILL_3__11578_ gnd vdd FILL
XFILL_1__12757_ gnd vdd FILL
XFILL_3__7763_ gnd vdd FILL
XFILL_0_BUFX2_insert370 gnd vdd FILL
XFILL_0__10418_ gnd vdd FILL
XFILL_0__14186_ gnd vdd FILL
X_8332_ _8333_/B _7948_/B gnd _8332_/Y vdd NAND2X1
XFILL_0_BUFX2_insert381 gnd vdd FILL
XFILL_6__14477_ gnd vdd FILL
XFILL_5__12138_ gnd vdd FILL
XFILL_3__16105_ gnd vdd FILL
XFILL_6__7472_ gnd vdd FILL
XFILL_0__11398_ gnd vdd FILL
XFILL_3__13317_ gnd vdd FILL
XFILL_4__15656_ gnd vdd FILL
XFILL_3__10529_ gnd vdd FILL
XFILL_0_BUFX2_insert392 gnd vdd FILL
XFILL_0__7985_ gnd vdd FILL
XFILL_3__9502_ gnd vdd FILL
XFILL_4__12868_ gnd vdd FILL
XFILL_1__11708_ gnd vdd FILL
XFILL_4_BUFX2_insert708 gnd vdd FILL
XFILL_0__13137_ gnd vdd FILL
XSFILL8680x27050 gnd vdd FILL
XFILL_1__15476_ gnd vdd FILL
XFILL_3__14297_ gnd vdd FILL
XFILL_3__7694_ gnd vdd FILL
XFILL_4_BUFX2_insert719 gnd vdd FILL
XFILL_4__14607_ gnd vdd FILL
XFILL_6__13428_ gnd vdd FILL
XFILL_0__9724_ gnd vdd FILL
XFILL_3__16036_ gnd vdd FILL
XFILL_5__12069_ gnd vdd FILL
XFILL_0__6936_ gnd vdd FILL
XFILL_4__11819_ gnd vdd FILL
X_8263_ _8305_/Q gnd _8263_/Y vdd INVX1
XFILL_3__13248_ gnd vdd FILL
XFILL_4__15587_ gnd vdd FILL
XFILL_1__14427_ gnd vdd FILL
XFILL_1__11639_ gnd vdd FILL
XFILL_2__13978_ gnd vdd FILL
X_7214_ _7214_/A _7207_/A _7213_/Y gnd _7272_/D vdd OAI21X1
XFILL_0__6867_ gnd vdd FILL
XFILL_0__9655_ gnd vdd FILL
XFILL_4__14538_ gnd vdd FILL
XSFILL18680x81050 gnd vdd FILL
X_8194_ _8282_/Q gnd _8196_/A vdd INVX1
XFILL_2__15717_ gnd vdd FILL
XFILL_0__12019_ gnd vdd FILL
XFILL_1__14358_ gnd vdd FILL
XFILL_3__9364_ gnd vdd FILL
XSFILL74200x75050 gnd vdd FILL
XFILL_0__8606_ gnd vdd FILL
XFILL_6__16078_ gnd vdd FILL
XFILL_5__15828_ gnd vdd FILL
X_7145_ _7145_/Q _9705_/CLK _9964_/R vdd _7089_/Y gnd vdd DFFSR
XFILL_1__13309_ gnd vdd FILL
XFILL_4__14469_ gnd vdd FILL
XFILL_3__8315_ gnd vdd FILL
XFILL_2__15648_ gnd vdd FILL
XFILL_3__9295_ gnd vdd FILL
XFILL_1__14289_ gnd vdd FILL
XFILL_4__16208_ gnd vdd FILL
XFILL_1__7330_ gnd vdd FILL
XSFILL13640x28050 gnd vdd FILL
X_7076_ _7055_/A _8868_/B gnd _7077_/C vdd NAND2X1
XFILL_1__16028_ gnd vdd FILL
XFILL_5__15759_ gnd vdd FILL
XFILL_3__8246_ gnd vdd FILL
XFILL_5_BUFX2_insert1060 gnd vdd FILL
XFILL_5_BUFX2_insert1071 gnd vdd FILL
XFILL_2__15579_ gnd vdd FILL
XFILL_5_BUFX2_insert1093 gnd vdd FILL
XFILL_0__8468_ gnd vdd FILL
XFILL_4__16139_ gnd vdd FILL
XFILL_1__9000_ gnd vdd FILL
XFILL_0__15709_ gnd vdd FILL
XFILL_0__7419_ gnd vdd FILL
XSFILL54120x42050 gnd vdd FILL
XFILL_0__8399_ gnd vdd FILL
XFILL_1__7192_ gnd vdd FILL
XSFILL33800x7050 gnd vdd FILL
XFILL_4__8990_ gnd vdd FILL
XFILL_1_BUFX2_insert609 gnd vdd FILL
XFILL_3__7059_ gnd vdd FILL
X_7978_ _7931_/B _9898_/B gnd _7978_/Y vdd NAND2X1
XFILL_4__7941_ gnd vdd FILL
XFILL_6__8857_ gnd vdd FILL
X_9717_ _9683_/A _7010_/CLK _7413_/R vdd _9717_/D gnd vdd DFFSR
X_6929_ _7007_/Q gnd _6931_/A vdd INVX1
XFILL_4__7872_ gnd vdd FILL
XFILL_6__7808_ gnd vdd FILL
XSFILL18760x61050 gnd vdd FILL
XFILL_1__9902_ gnd vdd FILL
XSFILL8600x71050 gnd vdd FILL
XSFILL19240x68050 gnd vdd FILL
X_9648_ _9625_/B _6960_/B gnd _9649_/C vdd NAND2X1
XFILL_4__9611_ gnd vdd FILL
X_10530_ _10528_/Y _10557_/B _10529_/Y gnd _10530_/Y vdd OAI21X1
XFILL_5_BUFX2_insert520 gnd vdd FILL
X_9579_ _9579_/Q _9195_/CLK _8051_/R vdd _9579_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert531 gnd vdd FILL
XFILL_5_BUFX2_insert542 gnd vdd FILL
XFILL_4__9542_ gnd vdd FILL
XFILL_5_BUFX2_insert553 gnd vdd FILL
X_10461_ _10379_/A _9195_/CLK _7915_/R vdd _10461_/D gnd vdd DFFSR
XSFILL23880x52050 gnd vdd FILL
XFILL_5_BUFX2_insert564 gnd vdd FILL
XFILL_1__9764_ gnd vdd FILL
XFILL_5_BUFX2_insert575 gnd vdd FILL
XFILL_3_BUFX2_insert1 gnd vdd FILL
XFILL_1__6976_ gnd vdd FILL
XSFILL109640x42050 gnd vdd FILL
X_12200_ _12150_/B _12907_/A gnd _12201_/C vdd NAND2X1
XFILL_5_BUFX2_insert586 gnd vdd FILL
XFILL_4__9473_ gnd vdd FILL
X_13180_ _13180_/Q _13180_/CLK _13180_/R vdd _13096_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert597 gnd vdd FILL
XFILL_1__8715_ gnd vdd FILL
X_10392_ _10372_/B _8088_/B gnd _10393_/C vdd NAND2X1
XSFILL38920x74050 gnd vdd FILL
XFILL112440x81050 gnd vdd FILL
X_12131_ _12122_/A _12131_/B gnd _12131_/Y vdd NAND2X1
XSFILL78520x60050 gnd vdd FILL
XFILL_1__8646_ gnd vdd FILL
XFILL_4__8355_ gnd vdd FILL
XSFILL69080x50 gnd vdd FILL
XSFILL39000x83050 gnd vdd FILL
XFILL_2_CLKBUF1_insert112 gnd vdd FILL
X_12062_ _12062_/A _12062_/B _12061_/Y gnd _13134_/B vdd NAND3X1
XFILL_2_CLKBUF1_insert123 gnd vdd FILL
XFILL_2__7370_ gnd vdd FILL
XFILL_2_CLKBUF1_insert134 gnd vdd FILL
XFILL_1__8577_ gnd vdd FILL
XFILL_4__7306_ gnd vdd FILL
XFILL_2_CLKBUF1_insert145 gnd vdd FILL
X_11013_ _12226_/Y _11013_/B gnd _11013_/Y vdd NAND2X1
XFILL_2_CLKBUF1_insert156 gnd vdd FILL
XFILL_2_CLKBUF1_insert167 gnd vdd FILL
XFILL_2_CLKBUF1_insert178 gnd vdd FILL
XFILL_2_CLKBUF1_insert189 gnd vdd FILL
XFILL_4__7237_ gnd vdd FILL
XSFILL18840x41050 gnd vdd FILL
X_15821_ _8809_/Q _15821_/B _15821_/C gnd _15824_/C vdd AOI21X1
XFILL_2__9040_ gnd vdd FILL
XFILL_1__7459_ gnd vdd FILL
XFILL_2_BUFX2_insert410 gnd vdd FILL
XFILL_2_BUFX2_insert421 gnd vdd FILL
XFILL_4__7168_ gnd vdd FILL
XFILL_2_BUFX2_insert432 gnd vdd FILL
XFILL_4__10150_ gnd vdd FILL
XFILL_2_BUFX2_insert443 gnd vdd FILL
XSFILL63960x16050 gnd vdd FILL
X_15752_ _15563_/A _15751_/Y _15563_/C _14284_/Y gnd _15752_/Y vdd OAI22X1
XFILL_2_BUFX2_insert454 gnd vdd FILL
X_12964_ vdd _12964_/B gnd _12965_/C vdd NAND2X1
XFILL_3__10880_ gnd vdd FILL
XFILL_2_BUFX2_insert465 gnd vdd FILL
XFILL_2_BUFX2_insert476 gnd vdd FILL
XFILL_4__7099_ gnd vdd FILL
X_14703_ _14703_/A gnd _14705_/C vdd INVX1
X_11915_ _11921_/A _12023_/B gnd _11916_/C vdd NAND2X1
XFILL_5__7981_ gnd vdd FILL
XFILL_2_BUFX2_insert487 gnd vdd FILL
XFILL_5__11440_ gnd vdd FILL
X_15683_ _15683_/A _15683_/B _15683_/C _14210_/Y gnd _15684_/A vdd OAI22X1
XFILL_6__10991_ gnd vdd FILL
XFILL_2_BUFX2_insert498 gnd vdd FILL
XFILL_1__9129_ gnd vdd FILL
X_12895_ _12895_/A gnd _12895_/Y vdd INVX1
XFILL_2__11260_ gnd vdd FILL
XFILL_5__9720_ gnd vdd FILL
XSFILL64040x25050 gnd vdd FILL
XFILL_1__11990_ gnd vdd FILL
XFILL_5__6932_ gnd vdd FILL
X_14634_ _10222_/Q gnd _14634_/Y vdd INVX1
XFILL_5__11371_ gnd vdd FILL
X_11846_ _12218_/Y _12117_/Y _11846_/C gnd _11849_/A vdd OAI21X1
XFILL_1__10941_ gnd vdd FILL
XFILL_2__11191_ gnd vdd FILL
XFILL_0__12370_ gnd vdd FILL
XFILL_5__13110_ gnd vdd FILL
XFILL_5__9651_ gnd vdd FILL
XFILL_5__6863_ gnd vdd FILL
XFILL_5__10322_ gnd vdd FILL
X_14565_ _8813_/Q gnd _14567_/B vdd INVX1
XFILL_4__13840_ gnd vdd FILL
XFILL_5__14090_ gnd vdd FILL
XSFILL115320x7050 gnd vdd FILL
XFILL_3__11501_ gnd vdd FILL
X_11777_ _11020_/Y _11764_/D gnd _11777_/Y vdd NAND2X1
XFILL_3__12481_ gnd vdd FILL
XFILL_2__10142_ gnd vdd FILL
XFILL_1__13660_ gnd vdd FILL
XFILL_5__8602_ gnd vdd FILL
XBUFX2_insert420 _14991_/Y gnd _15794_/B vdd BUFX2
XFILL_2__9873_ gnd vdd FILL
XFILL_0__11321_ gnd vdd FILL
XFILL_4__9809_ gnd vdd FILL
XBUFX2_insert431 _13326_/Y gnd _8714_/B vdd BUFX2
X_16304_ _14960_/Y _15595_/B _16304_/C gnd _16307_/A vdd OAI21X1
XFILL_1__10872_ gnd vdd FILL
XFILL_6__14400_ gnd vdd FILL
XBUFX2_insert442 _12378_/Y gnd _8088_/B vdd BUFX2
X_10728_ _10668_/A _7912_/CLK _8424_/R vdd _10728_/D gnd vdd DFFSR
X_13516_ _9303_/Q gnd _13517_/A vdd INVX1
XFILL_5__13041_ gnd vdd FILL
XBUFX2_insert453 _13276_/Y gnd _7184_/B vdd BUFX2
XFILL_5__10253_ gnd vdd FILL
XSFILL13080x65050 gnd vdd FILL
XFILL_3__14220_ gnd vdd FILL
XFILL_3__11432_ gnd vdd FILL
X_14496_ _14496_/A _14496_/B _14495_/Y _13795_/B gnd _14496_/Y vdd OAI22X1
XFILL_1__12611_ gnd vdd FILL
XFILL_2__8824_ gnd vdd FILL
XFILL_4__13771_ gnd vdd FILL
XBUFX2_insert464 _13318_/Y gnd _8315_/B vdd BUFX2
XFILL_4__10983_ gnd vdd FILL
XFILL_0__14040_ gnd vdd FILL
XFILL_2__14950_ gnd vdd FILL
XFILL_1__13591_ gnd vdd FILL
XBUFX2_insert475 _15041_/Y gnd _15187_/C vdd BUFX2
XFILL_5__8533_ gnd vdd FILL
XFILL_0__11252_ gnd vdd FILL
X_16235_ _16235_/A _16234_/Y _14843_/Y _16026_/D gnd _16236_/B vdd OAI22X1
XFILL_4__15510_ gnd vdd FILL
XFILL_6__11543_ gnd vdd FILL
XBUFX2_insert486 _12372_/Y gnd _7314_/B vdd BUFX2
X_10659_ _10659_/A gnd _10661_/A vdd INVX1
XFILL_4__12722_ gnd vdd FILL
X_13447_ _13423_/A _13418_/A _13465_/C gnd _14555_/C vdd NAND3X1
XBUFX2_insert497 BUFX2_insert494/A gnd _9711_/R vdd BUFX2
XFILL_1__15330_ gnd vdd FILL
XFILL_3__14151_ gnd vdd FILL
XFILL_5__10184_ gnd vdd FILL
XFILL_2__13901_ gnd vdd FILL
XFILL_3__11363_ gnd vdd FILL
XSFILL94360x82050 gnd vdd FILL
XFILL_2__8755_ gnd vdd FILL
XFILL_2_CLKBUF1_insert1079 gnd vdd FILL
XFILL_2__14881_ gnd vdd FILL
XFILL_0__11183_ gnd vdd FILL
XFILL_5__8464_ gnd vdd FILL
XFILL_6__14262_ gnd vdd FILL
XFILL_3__10314_ gnd vdd FILL
XFILL_3__13102_ gnd vdd FILL
X_13378_ _13377_/Y _13718_/B gnd _13843_/C vdd NAND2X1
X_16166_ _16166_/A _10354_/Q _7626_/A _15383_/A gnd _16172_/B vdd AOI22X1
XFILL_4__15441_ gnd vdd FILL
XSFILL59000x14050 gnd vdd FILL
XFILL_4__12653_ gnd vdd FILL
XFILL_2__7706_ gnd vdd FILL
XFILL_5__14992_ gnd vdd FILL
XFILL_3__14082_ gnd vdd FILL
XFILL_2__13832_ gnd vdd FILL
XFILL_0__10134_ gnd vdd FILL
XFILL_3__11294_ gnd vdd FILL
XFILL_1__15261_ gnd vdd FILL
XFILL_5__7415_ gnd vdd FILL
XFILL_1__12473_ gnd vdd FILL
XFILL_0__15991_ gnd vdd FILL
X_15117_ _6999_/Q gnd _15117_/Y vdd INVX1
XFILL_5__8395_ gnd vdd FILL
X_12329_ _6898_/A _12301_/B _12301_/C _12313_/D gnd _12330_/C vdd AOI22X1
XFILL_4__11604_ gnd vdd FILL
XFILL_5__13943_ gnd vdd FILL
XFILL_3__13033_ gnd vdd FILL
XFILL_4__15372_ gnd vdd FILL
XFILL_1__14212_ gnd vdd FILL
X_16097_ _15225_/A _7620_/A _7536_/Q _15383_/D gnd _16097_/Y vdd AOI22X1
XFILL_3__10245_ gnd vdd FILL
XFILL_4__12584_ gnd vdd FILL
XFILL_2__7637_ gnd vdd FILL
XFILL_1__11424_ gnd vdd FILL
XFILL_2__10975_ gnd vdd FILL
XFILL_1__15192_ gnd vdd FILL
XFILL_2__13763_ gnd vdd FILL
XFILL_0__14942_ gnd vdd FILL
XFILL_0__10065_ gnd vdd FILL
XFILL_5__7346_ gnd vdd FILL
X_15048_ _15384_/A _15048_/B _13422_/Y _15384_/D gnd _15048_/Y vdd OAI22X1
XFILL_4__14323_ gnd vdd FILL
XFILL_5__13874_ gnd vdd FILL
XFILL_4__11535_ gnd vdd FILL
XFILL_2__15502_ gnd vdd FILL
XFILL_2__12714_ gnd vdd FILL
XFILL_3__10176_ gnd vdd FILL
XFILL_1__14143_ gnd vdd FILL
XFILL_2__7568_ gnd vdd FILL
XFILL_1_BUFX2_insert15 gnd vdd FILL
XFILL_2__13694_ gnd vdd FILL
XFILL_1__11355_ gnd vdd FILL
XFILL_0__14873_ gnd vdd FILL
XFILL_1_BUFX2_insert26 gnd vdd FILL
XFILL_5__15613_ gnd vdd FILL
XFILL_5__12825_ gnd vdd FILL
XFILL_0__9371_ gnd vdd FILL
XFILL_3__8100_ gnd vdd FILL
XFILL_4__14254_ gnd vdd FILL
XFILL_1_BUFX2_insert37 gnd vdd FILL
XFILL_2__12645_ gnd vdd FILL
XFILL_1_BUFX2_insert48 gnd vdd FILL
XFILL_3__9080_ gnd vdd FILL
XFILL_1__10306_ gnd vdd FILL
XFILL_2__15433_ gnd vdd FILL
XFILL_4__11466_ gnd vdd FILL
XFILL_0__13824_ gnd vdd FILL
XFILL_2__7499_ gnd vdd FILL
XFILL_1_BUFX2_insert59 gnd vdd FILL
XFILL_3__14984_ gnd vdd FILL
XFILL_1__14074_ gnd vdd FILL
XFILL_5__9016_ gnd vdd FILL
XFILL_0__8322_ gnd vdd FILL
XFILL_1__11286_ gnd vdd FILL
XSFILL89320x71050 gnd vdd FILL
XSFILL53960x48050 gnd vdd FILL
XFILL_5__15544_ gnd vdd FILL
X_8950_ _8950_/A gnd _8952_/A vdd INVX1
XFILL_5__12756_ gnd vdd FILL
XFILL_4__10417_ gnd vdd FILL
XSFILL3560x12050 gnd vdd FILL
XFILL_4__14185_ gnd vdd FILL
XFILL_1__13025_ gnd vdd FILL
XFILL_3__13935_ gnd vdd FILL
XFILL_2__9238_ gnd vdd FILL
XFILL_2__12576_ gnd vdd FILL
XFILL_2__15364_ gnd vdd FILL
XFILL_4__11397_ gnd vdd FILL
XFILL_1__10237_ gnd vdd FILL
XFILL_0__13755_ gnd vdd FILL
XFILL_0__10967_ gnd vdd FILL
X_7901_ _7901_/Q _7915_/CLK _7915_/R vdd _7821_/Y gnd vdd DFFSR
XFILL_0__8253_ gnd vdd FILL
XFILL_5__11707_ gnd vdd FILL
XFILL_4__13136_ gnd vdd FILL
XFILL_5__15475_ gnd vdd FILL
XFILL_2__14315_ gnd vdd FILL
XFILL_2__11527_ gnd vdd FILL
X_8881_ _8881_/A _8902_/B _8881_/C gnd _8881_/Y vdd OAI21X1
XFILL_0__12706_ gnd vdd FILL
XFILL_3__13866_ gnd vdd FILL
XFILL_2__15295_ gnd vdd FILL
XFILL_2__9169_ gnd vdd FILL
XFILL_0__7204_ gnd vdd FILL
XFILL_1__10168_ gnd vdd FILL
XFILL_0__13686_ gnd vdd FILL
XFILL_5__14426_ gnd vdd FILL
XFILL_0__10898_ gnd vdd FILL
XSFILL94440x62050 gnd vdd FILL
X_7832_ _7821_/B _9624_/B gnd _7833_/C vdd NAND2X1
XFILL_0__8184_ gnd vdd FILL
XFILL_5__11638_ gnd vdd FILL
XFILL_3__15605_ gnd vdd FILL
XSFILL68600x72050 gnd vdd FILL
XFILL_2__14246_ gnd vdd FILL
XFILL_4__10279_ gnd vdd FILL
XFILL_2__11458_ gnd vdd FILL
XFILL_0__15425_ gnd vdd FILL
XFILL_0__12637_ gnd vdd FILL
XFILL_3__13797_ gnd vdd FILL
XFILL_5__9918_ gnd vdd FILL
XFILL_3__9982_ gnd vdd FILL
XFILL_1__14976_ gnd vdd FILL
XFILL_4__12018_ gnd vdd FILL
XFILL_5__14357_ gnd vdd FILL
XFILL_3__15536_ gnd vdd FILL
X_7763_ _7763_/A gnd _7763_/Y vdd INVX1
XFILL_2__10409_ gnd vdd FILL
XFILL_5__11569_ gnd vdd FILL
XSFILL33880x15050 gnd vdd FILL
XFILL_3__12748_ gnd vdd FILL
XFILL_2__14177_ gnd vdd FILL
XFILL_0__15356_ gnd vdd FILL
XFILL_2__11389_ gnd vdd FILL
XFILL_1__13927_ gnd vdd FILL
XFILL_5__13308_ gnd vdd FILL
XFILL_0__12568_ gnd vdd FILL
XFILL_5__9849_ gnd vdd FILL
X_9502_ _9514_/A _7838_/B gnd _9503_/C vdd NAND2X1
XFILL_0__7066_ gnd vdd FILL
XSFILL13720x50 gnd vdd FILL
XFILL_2__13128_ gnd vdd FILL
XFILL_5__14288_ gnd vdd FILL
X_7694_ _7694_/A gnd _7694_/Y vdd INVX1
XSFILL18680x76050 gnd vdd FILL
XSFILL48920x37050 gnd vdd FILL
XFILL_0__14307_ gnd vdd FILL
XFILL_3__15467_ gnd vdd FILL
XFILL_1__13858_ gnd vdd FILL
XFILL_3__8864_ gnd vdd FILL
XFILL_0__11519_ gnd vdd FILL
XSFILL104440x8050 gnd vdd FILL
XFILL_5__16027_ gnd vdd FILL
XFILL_0__15287_ gnd vdd FILL
XFILL_5__13239_ gnd vdd FILL
X_9433_ _9343_/A _7129_/CLK _8542_/R vdd _9433_/D gnd vdd DFFSR
XFILL_0__12499_ gnd vdd FILL
XFILL_6__8573_ gnd vdd FILL
XSFILL88520x23050 gnd vdd FILL
XFILL_3__14418_ gnd vdd FILL
XFILL_3__7815_ gnd vdd FILL
XFILL_4__13969_ gnd vdd FILL
XFILL_3__15398_ gnd vdd FILL
XFILL_0__14238_ gnd vdd FILL
XFILL_1__13789_ gnd vdd FILL
XSFILL49000x46050 gnd vdd FILL
XFILL_4__15708_ gnd vdd FILL
X_9364_ _9440_/Q gnd _9366_/A vdd INVX1
XFILL_3__14349_ gnd vdd FILL
XSFILL89400x51050 gnd vdd FILL
XFILL_1__15528_ gnd vdd FILL
XFILL_3__7746_ gnd vdd FILL
XFILL_0__14169_ gnd vdd FILL
XFILL_4_BUFX2_insert505 gnd vdd FILL
X_8315_ _8315_/A _8315_/B _8314_/Y gnd _8315_/Y vdd OAI21X1
XSFILL109560x57050 gnd vdd FILL
XFILL_4__15639_ gnd vdd FILL
XFILL_4_BUFX2_insert516 gnd vdd FILL
X_9295_ _9293_/Y _9232_/B _9295_/C gnd _9331_/D vdd OAI21X1
XFILL_0__7968_ gnd vdd FILL
XFILL_4_BUFX2_insert527 gnd vdd FILL
XFILL_4_BUFX2_insert538 gnd vdd FILL
XFILL_3__7677_ gnd vdd FILL
XFILL_1__15459_ gnd vdd FILL
XFILL_4_BUFX2_insert549 gnd vdd FILL
XFILL_1__8500_ gnd vdd FILL
X_8246_ _8246_/A _7094_/B gnd _8247_/C vdd NAND2X1
XFILL_3__16019_ gnd vdd FILL
XFILL_0__6919_ gnd vdd FILL
XFILL_1__9480_ gnd vdd FILL
XFILL_3__9416_ gnd vdd FILL
XSFILL94520x42050 gnd vdd FILL
XFILL_0__9638_ gnd vdd FILL
X_8177_ _8177_/Q _7537_/CLK _8053_/R vdd _8137_/Y gnd vdd DFFSR
XFILL_3__9347_ gnd vdd FILL
XFILL_4__8140_ gnd vdd FILL
XFILL_1__8362_ gnd vdd FILL
X_7128_ _7128_/Q _7640_/CLK _7896_/R vdd _7038_/Y gnd vdd DFFSR
XFILL_4__8071_ gnd vdd FILL
XFILL_3__9278_ gnd vdd FILL
XFILL_1__7313_ gnd vdd FILL
XSFILL18760x56050 gnd vdd FILL
X_7059_ _7059_/A _7064_/A _7058_/Y gnd _7059_/Y vdd OAI21X1
XFILL_3__8229_ gnd vdd FILL
XFILL_3_CLKBUF1_insert207 gnd vdd FILL
XFILL_3_CLKBUF1_insert218 gnd vdd FILL
XFILL_1__7244_ gnd vdd FILL
XSFILL43960x8050 gnd vdd FILL
XFILL_1_BUFX2_insert406 gnd vdd FILL
XSFILL23880x47050 gnd vdd FILL
XFILL_1__7175_ gnd vdd FILL
XFILL_1_BUFX2_insert417 gnd vdd FILL
XFILL_1_BUFX2_insert428 gnd vdd FILL
XFILL_4__8973_ gnd vdd FILL
X_11700_ _11700_/A gnd _12476_/B vdd INVX1
X_12680_ _12618_/A _12685_/CLK _12685_/R vdd _12680_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert439 gnd vdd FILL
XSFILL64760x59050 gnd vdd FILL
XSFILL38920x69050 gnd vdd FILL
XSFILL79560x19050 gnd vdd FILL
XFILL112440x76050 gnd vdd FILL
X_11631_ _11802_/A _11624_/C _11630_/Y gnd _11631_/Y vdd NAND3X1
XFILL_1_CLKBUF1_insert1074 gnd vdd FILL
XFILL_4__7855_ gnd vdd FILL
XSFILL79160x21050 gnd vdd FILL
X_14350_ _7212_/A gnd _14351_/A vdd INVX1
X_11562_ _11562_/A _11562_/B _11577_/B gnd _11563_/C vdd OAI21X1
XSFILL89320x7050 gnd vdd FILL
XSFILL79400x83050 gnd vdd FILL
XFILL_2__6870_ gnd vdd FILL
X_13301_ _13297_/C _13300_/Y gnd _13301_/Y vdd NOR2X1
X_10513_ _13919_/A gnd _10515_/A vdd INVX1
X_14281_ _14555_/C _15761_/C _14342_/B _14279_/Y gnd _14282_/B vdd OAI22X1
XFILL_5_BUFX2_insert350 gnd vdd FILL
X_11493_ _11492_/A _11492_/B _11553_/C gnd _11493_/Y vdd OAI21X1
XBUFX2_insert40 _13265_/Y gnd _6951_/A vdd BUFX2
XFILL_5_BUFX2_insert361 gnd vdd FILL
XFILL_4__9525_ gnd vdd FILL
XBUFX2_insert51 _13309_/Y gnd _8142_/A vdd BUFX2
XFILL_5_BUFX2_insert372 gnd vdd FILL
X_13232_ _13230_/Y _13231_/A _13294_/A gnd _13260_/B vdd OAI21X1
X_16020_ _16013_/Y _16020_/B _16020_/C gnd _16021_/A vdd NAND3X1
XSFILL18840x36050 gnd vdd FILL
X_10444_ _10444_/A _10443_/A _10443_/Y gnd _10482_/D vdd OAI21X1
XBUFX2_insert62 _14983_/Y gnd _15687_/A vdd BUFX2
XSFILL84280x12050 gnd vdd FILL
XFILL_5_BUFX2_insert383 gnd vdd FILL
XBUFX2_insert73 _12366_/Y gnd _7180_/B vdd BUFX2
XFILL_5_BUFX2_insert394 gnd vdd FILL
XBUFX2_insert84 _13372_/Y gnd _14555_/B vdd BUFX2
XFILL_1__9747_ gnd vdd FILL
XBUFX2_insert95 _15068_/Y gnd _15981_/B vdd BUFX2
XFILL_1__6959_ gnd vdd FILL
XSFILL84520x74050 gnd vdd FILL
X_13163_ _11971_/A gnd _13163_/Y vdd INVX1
XSFILL99320x34050 gnd vdd FILL
X_10375_ _10373_/Y _10363_/B _10375_/C gnd _10375_/Y vdd OAI21X1
XFILL_1__9678_ gnd vdd FILL
XFILL_2__8471_ gnd vdd FILL
XFILL_5__7200_ gnd vdd FILL
X_12114_ _12114_/A _12114_/B _12113_/Y gnd _13173_/B vdd NAND3X1
XFILL_4__9387_ gnd vdd FILL
XFILL_5__10940_ gnd vdd FILL
X_13094_ _13180_/Q gnd _13096_/A vdd INVX1
XFILL_3__10030_ gnd vdd FILL
XFILL_6__11190_ gnd vdd FILL
XFILL_1__8629_ gnd vdd FILL
XFILL_2__7422_ gnd vdd FILL
XFILL_2__10760_ gnd vdd FILL
XFILL_4__8338_ gnd vdd FILL
X_12045_ _12482_/B _12025_/B _12025_/C gnd gnd _12046_/C vdd AOI22X1
XFILL_4__11320_ gnd vdd FILL
XFILL_2__7353_ gnd vdd FILL
XFILL_5__10871_ gnd vdd FILL
XFILL_1__11140_ gnd vdd FILL
XFILL_2__10691_ gnd vdd FILL
XFILL_5__7062_ gnd vdd FILL
XFILL_4__8269_ gnd vdd FILL
XFILL_5__12610_ gnd vdd FILL
XFILL_0__11870_ gnd vdd FILL
XFILL_2__12430_ gnd vdd FILL
XFILL_5__13590_ gnd vdd FILL
XFILL_4__11251_ gnd vdd FILL
XSFILL38600x51050 gnd vdd FILL
XFILL_3__11981_ gnd vdd FILL
XFILL_0__10821_ gnd vdd FILL
XFILL_1__11071_ gnd vdd FILL
X_15804_ _7852_/A gnd _15804_/Y vdd INVX1
XSFILL113800x44050 gnd vdd FILL
XFILL_2__9023_ gnd vdd FILL
XFILL_2_BUFX2_insert240 gnd vdd FILL
XFILL_3__13720_ gnd vdd FILL
XFILL_4__11182_ gnd vdd FILL
XFILL_3__10932_ gnd vdd FILL
XFILL_1__10022_ gnd vdd FILL
XFILL_2__12361_ gnd vdd FILL
X_13996_ _13995_/Y _13996_/B gnd _13997_/C vdd NOR2X1
XFILL_2_BUFX2_insert251 gnd vdd FILL
XFILL_0__13540_ gnd vdd FILL
XFILL_0__10752_ gnd vdd FILL
XSFILL114440x10050 gnd vdd FILL
XFILL_2_BUFX2_insert262 gnd vdd FILL
XFILL_2_BUFX2_insert273 gnd vdd FILL
XFILL_5__15260_ gnd vdd FILL
X_15735_ _10087_/Q _15696_/A gnd _15736_/B vdd NAND2X1
XFILL_5__12472_ gnd vdd FILL
XFILL_2_BUFX2_insert284 gnd vdd FILL
X_12947_ _12907_/A _7532_/CLK _8816_/R vdd _12947_/D gnd vdd DFFSR
XFILL_4__10133_ gnd vdd FILL
XFILL_2__14100_ gnd vdd FILL
XFILL_2__11312_ gnd vdd FILL
XFILL_2_BUFX2_insert295 gnd vdd FILL
XFILL_4__15990_ gnd vdd FILL
XFILL_3__13651_ gnd vdd FILL
XSFILL114440x3050 gnd vdd FILL
XFILL_2__15080_ gnd vdd FILL
XSFILL94360x77050 gnd vdd FILL
XFILL_1__14830_ gnd vdd FILL
XFILL_2__12292_ gnd vdd FILL
XFILL_5__14211_ gnd vdd FILL
XFILL_0__13471_ gnd vdd FILL
XFILL_0__10683_ gnd vdd FILL
XFILL_5__7964_ gnd vdd FILL
XFILL_5__11423_ gnd vdd FILL
XFILL_3__12602_ gnd vdd FILL
XFILL_5__15191_ gnd vdd FILL
X_15666_ _15666_/A _15663_/Y gnd _15667_/C vdd NOR2X1
XFILL_2__14031_ gnd vdd FILL
XFILL_4__14941_ gnd vdd FILL
XFILL_4__10064_ gnd vdd FILL
XFILL_0__15210_ gnd vdd FILL
XFILL_3__16370_ gnd vdd FILL
X_12878_ vdd _15812_/Y gnd _12879_/C vdd NAND2X1
XFILL_1_BUFX2_insert940 gnd vdd FILL
XFILL_2__11243_ gnd vdd FILL
XFILL_0__12422_ gnd vdd FILL
XFILL_1_BUFX2_insert951 gnd vdd FILL
XFILL_3__13582_ gnd vdd FILL
XFILL_1__14761_ gnd vdd FILL
XFILL_3__10794_ gnd vdd FILL
XFILL_1_BUFX2_insert962 gnd vdd FILL
XFILL_5__6915_ gnd vdd FILL
XFILL_1__11973_ gnd vdd FILL
XFILL_0__16190_ gnd vdd FILL
XSFILL69160x53050 gnd vdd FILL
XSFILL99400x14050 gnd vdd FILL
X_14617_ _14608_/Y _14617_/B _14617_/C gnd _14617_/Y vdd NAND3X1
XFILL_5__14142_ gnd vdd FILL
XFILL_1_BUFX2_insert973 gnd vdd FILL
XFILL_3__15321_ gnd vdd FILL
X_11829_ _11829_/A _11828_/Y gnd _11830_/A vdd NOR2X1
XFILL_5__11354_ gnd vdd FILL
XFILL_4__14872_ gnd vdd FILL
XFILL_2__9925_ gnd vdd FILL
XFILL_3__12533_ gnd vdd FILL
X_15597_ _15597_/A _15596_/Y gnd _15598_/B vdd NOR2X1
XFILL_1__13712_ gnd vdd FILL
XFILL_1_BUFX2_insert984 gnd vdd FILL
XFILL_1_BUFX2_insert995 gnd vdd FILL
XFILL_1__10924_ gnd vdd FILL
XFILL_0__15141_ gnd vdd FILL
XFILL_2__11174_ gnd vdd FILL
XFILL_0__12353_ gnd vdd FILL
XFILL_5__9634_ gnd vdd FILL
XFILL_1__14692_ gnd vdd FILL
XFILL_5__6846_ gnd vdd FILL
XFILL_5__10305_ gnd vdd FILL
XFILL_4__13823_ gnd vdd FILL
XSFILL73640x78050 gnd vdd FILL
XFILL_6__12644_ gnd vdd FILL
X_14548_ _14537_/Y _14548_/B gnd _14549_/B vdd NOR2X1
XFILL_5__14073_ gnd vdd FILL
XFILL_2__10125_ gnd vdd FILL
XFILL_3__15252_ gnd vdd FILL
XFILL_5__11285_ gnd vdd FILL
XFILL_2__9856_ gnd vdd FILL
XFILL_1__13643_ gnd vdd FILL
XFILL_3__12464_ gnd vdd FILL
XFILL_0__11304_ gnd vdd FILL
XBUFX2_insert250 _10922_/Y gnd _14791_/C vdd BUFX2
XFILL_2__15982_ gnd vdd FILL
XFILL_0__15072_ gnd vdd FILL
XBUFX2_insert261 _11225_/Y gnd _11574_/B vdd BUFX2
XFILL_5__13024_ gnd vdd FILL
XSFILL74280x44050 gnd vdd FILL
XFILL_0__12284_ gnd vdd FILL
XBUFX2_insert272 _13364_/Y gnd _10681_/A vdd BUFX2
XFILL_3__14203_ gnd vdd FILL
XBUFX2_insert283 _15003_/Y gnd _15521_/C vdd BUFX2
XFILL_5__10236_ gnd vdd FILL
XFILL_0__8871_ gnd vdd FILL
X_14479_ _14478_/Y _14479_/B _14862_/C _14477_/Y gnd _14480_/B vdd OAI22X1
XFILL_4__13754_ gnd vdd FILL
XFILL_3__11415_ gnd vdd FILL
XFILL_3__7600_ gnd vdd FILL
XFILL_4__10966_ gnd vdd FILL
XFILL_3__15183_ gnd vdd FILL
XFILL_0__14023_ gnd vdd FILL
XBUFX2_insert294 _13356_/Y gnd _10280_/B vdd BUFX2
XFILL_3__12395_ gnd vdd FILL
XFILL_1__16362_ gnd vdd FILL
XFILL_2__10056_ gnd vdd FILL
XFILL_2__14933_ gnd vdd FILL
XFILL_2__9787_ gnd vdd FILL
XFILL_3__8580_ gnd vdd FILL
XFILL_5__8516_ gnd vdd FILL
XFILL_1__13574_ gnd vdd FILL
XFILL_0__11235_ gnd vdd FILL
X_16218_ _16218_/A _16217_/Y _16218_/C gnd _16219_/C vdd NOR3X1
XFILL_5_CLKBUF1_insert140 gnd vdd FILL
XFILL_1__10786_ gnd vdd FILL
XFILL_6__14314_ gnd vdd FILL
XFILL_0__7822_ gnd vdd FILL
XFILL_4__12705_ gnd vdd FILL
XSFILL89320x66050 gnd vdd FILL
XFILL_5__9496_ gnd vdd FILL
XFILL_5_CLKBUF1_insert151 gnd vdd FILL
XFILL_5__10167_ gnd vdd FILL
XFILL_3__14134_ gnd vdd FILL
XFILL_5_CLKBUF1_insert162 gnd vdd FILL
XFILL_5_CLKBUF1_insert173 gnd vdd FILL
XFILL_4__13685_ gnd vdd FILL
XFILL_1__12525_ gnd vdd FILL
XFILL_1__15313_ gnd vdd FILL
XFILL_2__8738_ gnd vdd FILL
XFILL_3__11346_ gnd vdd FILL
XFILL_2__14864_ gnd vdd FILL
XFILL_4__10897_ gnd vdd FILL
XFILL_1__16293_ gnd vdd FILL
X_8100_ _8100_/A _7972_/B gnd _8101_/C vdd NAND2X1
XFILL_5__8447_ gnd vdd FILL
XFILL_5_CLKBUF1_insert184 gnd vdd FILL
XFILL_0__11166_ gnd vdd FILL
XFILL_5_CLKBUF1_insert195 gnd vdd FILL
X_16149_ _14747_/Y _15595_/B _16148_/Y gnd _16152_/A vdd OAI21X1
XSFILL38760x9050 gnd vdd FILL
XFILL_4__15424_ gnd vdd FILL
XFILL_4__12636_ gnd vdd FILL
X_9080_ _9078_/Y _9151_/A _9080_/C gnd _9174_/D vdd OAI21X1
XFILL_0__7753_ gnd vdd FILL
XSFILL28760x19050 gnd vdd FILL
XFILL_2__13815_ gnd vdd FILL
XFILL_1__15244_ gnd vdd FILL
XFILL_3__14065_ gnd vdd FILL
XFILL_5__14975_ gnd vdd FILL
XFILL_3__11277_ gnd vdd FILL
XFILL_3__7462_ gnd vdd FILL
XFILL_1__12456_ gnd vdd FILL
XFILL_0__10117_ gnd vdd FILL
XFILL_6__10408_ gnd vdd FILL
XFILL_0__15974_ gnd vdd FILL
XFILL_2__14795_ gnd vdd FILL
XFILL_5__8378_ gnd vdd FILL
XFILL_0__11097_ gnd vdd FILL
X_8031_ _7953_/A _7647_/CLK _9823_/R vdd _8031_/D gnd vdd DFFSR
XFILL_3__13016_ gnd vdd FILL
XFILL_4__15355_ gnd vdd FILL
XSFILL94440x57050 gnd vdd FILL
XFILL_0__7684_ gnd vdd FILL
XFILL_5__13926_ gnd vdd FILL
XFILL_4__12567_ gnd vdd FILL
XFILL_1__11407_ gnd vdd FILL
XFILL_1__15175_ gnd vdd FILL
XFILL_2__13746_ gnd vdd FILL
XFILL_2__10958_ gnd vdd FILL
XFILL_0__10048_ gnd vdd FILL
XFILL_1__12387_ gnd vdd FILL
XFILL_5__7329_ gnd vdd FILL
XFILL_0__14925_ gnd vdd FILL
XFILL_0__9423_ gnd vdd FILL
XFILL_4__14306_ gnd vdd FILL
XFILL_4__11518_ gnd vdd FILL
XFILL_5__13857_ gnd vdd FILL
XFILL_1__14126_ gnd vdd FILL
XFILL_3__9132_ gnd vdd FILL
XFILL_3__10159_ gnd vdd FILL
XFILL_4__15286_ gnd vdd FILL
XFILL_4__12498_ gnd vdd FILL
XSFILL53960x3050 gnd vdd FILL
XFILL_1__11338_ gnd vdd FILL
XFILL_0__14856_ gnd vdd FILL
XFILL_2__13677_ gnd vdd FILL
XFILL_2__10889_ gnd vdd FILL
XFILL_0__9354_ gnd vdd FILL
XFILL_4__14237_ gnd vdd FILL
XFILL_5__13788_ gnd vdd FILL
XFILL_4__11449_ gnd vdd FILL
X_9982_ _9980_/Y _9979_/B _9982_/C gnd _9982_/Y vdd OAI21X1
XFILL_2__15416_ gnd vdd FILL
XFILL_0__13807_ gnd vdd FILL
XFILL_2__12628_ gnd vdd FILL
XFILL_1__14057_ gnd vdd FILL
XFILL_3__14967_ gnd vdd FILL
XSFILL73720x58050 gnd vdd FILL
XFILL_6__12009_ gnd vdd FILL
XFILL_2__16396_ gnd vdd FILL
XFILL_1__11269_ gnd vdd FILL
XFILL_0__14787_ gnd vdd FILL
X_8933_ _8933_/Q _8926_/CLK _7262_/R vdd _8933_/D gnd vdd DFFSR
XFILL_5__12739_ gnd vdd FILL
XFILL_0__11999_ gnd vdd FILL
XSFILL58280x57050 gnd vdd FILL
XFILL_5__15527_ gnd vdd FILL
XFILL_0__9285_ gnd vdd FILL
XFILL_3__8014_ gnd vdd FILL
XFILL_4__14168_ gnd vdd FILL
XFILL_1__13008_ gnd vdd FILL
XFILL_3__13918_ gnd vdd FILL
XFILL_2__15347_ gnd vdd FILL
XSFILL8680x40050 gnd vdd FILL
XFILL_0__13738_ gnd vdd FILL
XFILL_3__14898_ gnd vdd FILL
XFILL_0__8236_ gnd vdd FILL
XFILL_4__13119_ gnd vdd FILL
X_8864_ _8864_/A gnd _8866_/A vdd INVX1
XFILL_5__15458_ gnd vdd FILL
XFILL_3__13849_ gnd vdd FILL
XFILL_4__14099_ gnd vdd FILL
XSFILL89400x46050 gnd vdd FILL
XFILL_2__15278_ gnd vdd FILL
XFILL_0__13669_ gnd vdd FILL
XFILL_5__14409_ gnd vdd FILL
X_7815_ _7815_/A _7814_/A _7815_/C gnd _7815_/Y vdd OAI21X1
XFILL_6__6955_ gnd vdd FILL
XFILL_5__15389_ gnd vdd FILL
XFILL_2__14229_ gnd vdd FILL
XFILL_0__15408_ gnd vdd FILL
X_8795_ _8795_/Q _8151_/CLK _9048_/R vdd _8795_/D gnd vdd DFFSR
XFILL_0_CLKBUF1_insert1080 gnd vdd FILL
XFILL_0__7118_ gnd vdd FILL
XFILL_0__16388_ gnd vdd FILL
XFILL_1__14959_ gnd vdd FILL
XFILL_3__15519_ gnd vdd FILL
XFILL_0__8098_ gnd vdd FILL
X_7746_ _7753_/B _7490_/B gnd _7747_/C vdd NAND2X1
XFILL_1__8980_ gnd vdd FILL
XFILL_3__8916_ gnd vdd FILL
XFILL_0__15339_ gnd vdd FILL
XFILL_3__9896_ gnd vdd FILL
XFILL_0__7049_ gnd vdd FILL
XFILL_1__7931_ gnd vdd FILL
X_7677_ _7723_/B _7293_/B gnd _7678_/C vdd NAND2X1
XFILL_3__8847_ gnd vdd FILL
XSFILL39080x52050 gnd vdd FILL
X_9416_ _9401_/A _8136_/B gnd _9416_/Y vdd NAND2X1
XSFILL13720x6050 gnd vdd FILL
XSFILL69320x13050 gnd vdd FILL
XFILL_1__7862_ gnd vdd FILL
XFILL_3__8778_ gnd vdd FILL
XFILL_4__7571_ gnd vdd FILL
XFILL_1__9601_ gnd vdd FILL
XFILL_4_BUFX2_insert302 gnd vdd FILL
X_9347_ _9398_/A _9347_/B gnd _9347_/Y vdd NAND2X1
XFILL_4_BUFX2_insert313 gnd vdd FILL
XFILL_3__7729_ gnd vdd FILL
XFILL_4_BUFX2_insert324 gnd vdd FILL
XSFILL8760x20050 gnd vdd FILL
XFILL_4_BUFX2_insert335 gnd vdd FILL
XFILL_1__9532_ gnd vdd FILL
XSFILL33800x54050 gnd vdd FILL
XFILL_4_BUFX2_insert346 gnd vdd FILL
X_9278_ _9326_/Q gnd _9278_/Y vdd INVX1
XFILL_4_BUFX2_insert357 gnd vdd FILL
XFILL_4__9241_ gnd vdd FILL
XFILL_4_BUFX2_insert368 gnd vdd FILL
XSFILL109240x4050 gnd vdd FILL
X_10160_ _10160_/A _8496_/B gnd _10161_/C vdd NAND2X1
XFILL_4_BUFX2_insert379 gnd vdd FILL
XSFILL34440x20050 gnd vdd FILL
X_8229_ _8227_/Y _8208_/B _8229_/C gnd _8229_/Y vdd OAI21X1
XFILL_1__9463_ gnd vdd FILL
XFILL_4__9172_ gnd vdd FILL
X_10091_ _10091_/Q _7915_/CLK _8669_/R vdd _10091_/D gnd vdd DFFSR
XFILL_4__8123_ gnd vdd FILL
XFILL111960x64050 gnd vdd FILL
XFILL_1__9394_ gnd vdd FILL
XFILL_1__8345_ gnd vdd FILL
XSFILL13720x21050 gnd vdd FILL
XFILL_4__8054_ gnd vdd FILL
XSFILL79160x16050 gnd vdd FILL
XFILL112040x73050 gnd vdd FILL
X_13850_ _13850_/A _13850_/B gnd _13850_/Y vdd NOR2X1
XFILL_1__8276_ gnd vdd FILL
X_12801_ _12801_/Q _12685_/CLK _12799_/R vdd _12727_/Y gnd vdd DFFSR
XFILL_1__7227_ gnd vdd FILL
X_13781_ _9564_/Q gnd _13781_/Y vdd INVX1
X_10993_ _12207_/Y gnd _10993_/Y vdd INVX1
X_15520_ _14010_/A _15342_/B _15520_/C gnd _15522_/A vdd OAI21X1
XFILL_1_BUFX2_insert225 gnd vdd FILL
X_12732_ _12768_/A memoryOutData[12] gnd _12733_/C vdd NAND2X1
XFILL_1__7158_ gnd vdd FILL
XFILL_1_BUFX2_insert236 gnd vdd FILL
XFILL_1_BUFX2_insert247 gnd vdd FILL
XFILL_1_BUFX2_insert258 gnd vdd FILL
XFILL_4__8956_ gnd vdd FILL
X_15451_ _8465_/A gnd _15451_/Y vdd INVX1
XFILL_1_BUFX2_insert269 gnd vdd FILL
X_12663_ _12663_/Q _12667_/CLK _12809_/R vdd _12663_/D gnd vdd DFFSR
XSFILL99320x29050 gnd vdd FILL
XFILL_1__7089_ gnd vdd FILL
XFILL_0_BUFX2_insert903 gnd vdd FILL
XFILL_2__7971_ gnd vdd FILL
X_14402_ _14402_/A _14402_/B _14402_/C gnd _13009_/B vdd AOI21X1
XFILL_0_BUFX2_insert914 gnd vdd FILL
XFILL_5__7680_ gnd vdd FILL
XFILL_4__8887_ gnd vdd FILL
XFILL_0_BUFX2_insert925 gnd vdd FILL
X_11614_ _11614_/A gnd _11618_/B vdd INVX1
X_15382_ _6926_/A _15382_/B _16096_/C _7390_/Q gnd _15388_/A vdd AOI22X1
X_12594_ _12594_/A gnd _12596_/A vdd INVX1
XFILL_2__6922_ gnd vdd FILL
XFILL_0_BUFX2_insert936 gnd vdd FILL
XFILL_0_BUFX2_insert947 gnd vdd FILL
XFILL_0_BUFX2_insert958 gnd vdd FILL
XFILL_4__7838_ gnd vdd FILL
XFILL_0_BUFX2_insert969 gnd vdd FILL
X_14333_ _14333_/A _14332_/Y gnd _14357_/A vdd NOR2X1
XFILL_4__10820_ gnd vdd FILL
X_11545_ _11521_/C _11574_/B _11544_/Y gnd _11545_/Y vdd OAI21X1
XFILL_5__11070_ gnd vdd FILL
XFILL_2__9641_ gnd vdd FILL
XFILL_1__10640_ gnd vdd FILL
XFILL_2__6853_ gnd vdd FILL
XSFILL109320x14050 gnd vdd FILL
XFILL_5__9350_ gnd vdd FILL
XFILL_5__10021_ gnd vdd FILL
X_14264_ _14253_/Y _14264_/B gnd _14265_/B vdd NOR2X1
X_11476_ _11327_/Y _11486_/C _11174_/C gnd _11476_/Y vdd AOI21X1
XFILL_3__11200_ gnd vdd FILL
XFILL_4__10751_ gnd vdd FILL
XSFILL88760x74050 gnd vdd FILL
XFILL_3__12180_ gnd vdd FILL
XFILL_4__9508_ gnd vdd FILL
XFILL_2__11930_ gnd vdd FILL
XFILL_0__11020_ gnd vdd FILL
X_16003_ _16003_/A _16003_/B gnd _16004_/B vdd NOR2X1
XFILL112120x53050 gnd vdd FILL
XFILL_1__10571_ gnd vdd FILL
X_13215_ _13215_/A _13215_/B gnd _13231_/B vdd NOR2X1
X_10427_ _10427_/A gnd _10427_/Y vdd INVX1
XFILL_5__9281_ gnd vdd FILL
XFILL_3__11131_ gnd vdd FILL
X_14195_ _14194_/Y _14195_/B gnd _14217_/B vdd NOR2X1
XFILL_4__13470_ gnd vdd FILL
XFILL_2__8523_ gnd vdd FILL
XFILL_1__12310_ gnd vdd FILL
XFILL_4__10682_ gnd vdd FILL
XFILL_2__11861_ gnd vdd FILL
XFILL_1__13290_ gnd vdd FILL
XFILL_5__8232_ gnd vdd FILL
XFILL_6_CLKBUF1_insert224 gnd vdd FILL
X_10358_ _10358_/A gnd _10360_/A vdd INVX1
XFILL_4__12421_ gnd vdd FILL
X_13146_ _13149_/A _13146_/B gnd _13147_/C vdd NAND2X1
XFILL_2__13600_ gnd vdd FILL
XFILL_5__11972_ gnd vdd FILL
XFILL_4_BUFX2_insert880 gnd vdd FILL
XFILL_3__11062_ gnd vdd FILL
XFILL_5__14760_ gnd vdd FILL
XFILL_4_BUFX2_insert891 gnd vdd FILL
XFILL_2__10812_ gnd vdd FILL
XFILL_1__12241_ gnd vdd FILL
XFILL_2__8454_ gnd vdd FILL
XFILL_2__14580_ gnd vdd FILL
XFILL_2__11792_ gnd vdd FILL
XFILL_0__12971_ gnd vdd FILL
XFILL_5__10923_ gnd vdd FILL
XFILL_3__10013_ gnd vdd FILL
XFILL_4__15140_ gnd vdd FILL
XFILL_5__13711_ gnd vdd FILL
X_13077_ _6900_/A _8169_/CLK _8937_/R vdd _13077_/D gnd vdd DFFSR
XFILL_4__12352_ gnd vdd FILL
X_10289_ _10287_/Y _10264_/A _10289_/C gnd _10345_/D vdd OAI21X1
XFILL_5__14691_ gnd vdd FILL
XFILL_2__10743_ gnd vdd FILL
XFILL_0__14710_ gnd vdd FILL
XFILL_2__13531_ gnd vdd FILL
XFILL_3__15870_ gnd vdd FILL
XFILL_5__7114_ gnd vdd FILL
XFILL_0__11922_ gnd vdd FILL
XFILL_1__12172_ gnd vdd FILL
XFILL_2__8385_ gnd vdd FILL
XFILL_6__10124_ gnd vdd FILL
XFILL_0__15690_ gnd vdd FILL
XSFILL69160x48050 gnd vdd FILL
X_12028_ _12028_/A _12719_/A _12024_/C gnd _12030_/B vdd NAND3X1
XFILL_5__13642_ gnd vdd FILL
XFILL_4__11303_ gnd vdd FILL
XFILL_5__8094_ gnd vdd FILL
XFILL_6__15981_ gnd vdd FILL
XFILL_3__14821_ gnd vdd FILL
XFILL_4__15071_ gnd vdd FILL
XFILL_2__7336_ gnd vdd FILL
XFILL_1__11123_ gnd vdd FILL
XFILL_2__16250_ gnd vdd FILL
XFILL_4__12283_ gnd vdd FILL
XFILL_0__14641_ gnd vdd FILL
XFILL_2__13462_ gnd vdd FILL
XFILL_2__10674_ gnd vdd FILL
XSFILL84200x51050 gnd vdd FILL
XFILL_5__7045_ gnd vdd FILL
XFILL_0__11853_ gnd vdd FILL
XFILL_4__14022_ gnd vdd FILL
XFILL_2__15201_ gnd vdd FILL
XFILL_5__16361_ gnd vdd FILL
XFILL_5__13573_ gnd vdd FILL
XFILL_4__11234_ gnd vdd FILL
XFILL_2__12413_ gnd vdd FILL
XFILL_5__10785_ gnd vdd FILL
XFILL_3__14752_ gnd vdd FILL
XFILL_2__16181_ gnd vdd FILL
XFILL_2__13393_ gnd vdd FILL
XFILL_1__15931_ gnd vdd FILL
XFILL_3__11964_ gnd vdd FILL
XFILL_1__11054_ gnd vdd FILL
XFILL_0__10804_ gnd vdd FILL
XFILL_0__14572_ gnd vdd FILL
XFILL_5__15312_ gnd vdd FILL
XFILL_5__12524_ gnd vdd FILL
XFILL_0__11784_ gnd vdd FILL
XFILL_5__16292_ gnd vdd FILL
XFILL_2__9006_ gnd vdd FILL
XFILL_3__13703_ gnd vdd FILL
XFILL_3__10915_ gnd vdd FILL
XFILL_2__12344_ gnd vdd FILL
X_13979_ _8801_/Q _13853_/B _13978_/Y gnd _13987_/B vdd AOI21X1
XFILL_0__16311_ gnd vdd FILL
XFILL_4__11165_ gnd vdd FILL
XFILL_1__10005_ gnd vdd FILL
XFILL_2__15132_ gnd vdd FILL
XFILL_0__13523_ gnd vdd FILL
XFILL_2__7198_ gnd vdd FILL
XFILL_3__14683_ gnd vdd FILL
XFILL_3__11895_ gnd vdd FILL
XFILL_0__8021_ gnd vdd FILL
XFILL_1__15862_ gnd vdd FILL
X_15718_ _14222_/Y _15386_/B _15386_/C _15718_/D gnd _15719_/A vdd OAI22X1
XFILL_5__15243_ gnd vdd FILL
XFILL_6_BUFX2_insert408 gnd vdd FILL
XFILL_5__8996_ gnd vdd FILL
XFILL_4__10116_ gnd vdd FILL
XFILL_5__12455_ gnd vdd FILL
XSFILL49080x15050 gnd vdd FILL
XFILL_3__13634_ gnd vdd FILL
XFILL_6__14794_ gnd vdd FILL
XFILL112200x33050 gnd vdd FILL
XFILL_4__15973_ gnd vdd FILL
XFILL_0__16242_ gnd vdd FILL
XFILL_1__14813_ gnd vdd FILL
XFILL_2__15063_ gnd vdd FILL
XFILL_2__12275_ gnd vdd FILL
XFILL_4__11096_ gnd vdd FILL
XFILL_0__13454_ gnd vdd FILL
XSFILL23720x1050 gnd vdd FILL
XFILL_5__7947_ gnd vdd FILL
XFILL_1__15793_ gnd vdd FILL
XFILL_0__10666_ gnd vdd FILL
XFILL_5__11406_ gnd vdd FILL
X_7600_ _7577_/B _8624_/B gnd _7600_/Y vdd NAND2X1
XFILL_5__15174_ gnd vdd FILL
X_15649_ _15645_/Y _15649_/B gnd _15650_/C vdd NAND2X1
XFILL_4__10047_ gnd vdd FILL
X_8580_ _8580_/A _8589_/B _8579_/Y gnd _8666_/D vdd OAI21X1
XFILL_5__12386_ gnd vdd FILL
XFILL_2__14014_ gnd vdd FILL
XFILL_3__16353_ gnd vdd FILL
XFILL_1_BUFX2_insert770 gnd vdd FILL
XFILL_4__14924_ gnd vdd FILL
XFILL_2__11226_ gnd vdd FILL
XFILL_0__12405_ gnd vdd FILL
XFILL_3__9750_ gnd vdd FILL
XFILL_3__13565_ gnd vdd FILL
XFILL_1_BUFX2_insert781 gnd vdd FILL
XFILL_0__16173_ gnd vdd FILL
XFILL_1__11956_ gnd vdd FILL
XFILL_3__10777_ gnd vdd FILL
XFILL_1_BUFX2_insert792 gnd vdd FILL
XFILL_3__6962_ gnd vdd FILL
XFILL_1__14744_ gnd vdd FILL
XFILL_5__14125_ gnd vdd FILL
XFILL_0__13385_ gnd vdd FILL
X_7531_ _7531_/Q _7261_/CLK _7531_/R vdd _7479_/Y gnd vdd DFFSR
XFILL_3__15304_ gnd vdd FILL
XFILL_5__7878_ gnd vdd FILL
XFILL_5__11337_ gnd vdd FILL
XFILL_4__14855_ gnd vdd FILL
XFILL_3__12516_ gnd vdd FILL
XFILL_2__9908_ gnd vdd FILL
XFILL112200x5050 gnd vdd FILL
XFILL_3__8701_ gnd vdd FILL
XFILL_1__10907_ gnd vdd FILL
XFILL_3__16284_ gnd vdd FILL
XFILL_2__11157_ gnd vdd FILL
XFILL_0__15124_ gnd vdd FILL
XFILL_0__12336_ gnd vdd FILL
XFILL_3__13496_ gnd vdd FILL
XSFILL28360x16050 gnd vdd FILL
XFILL_5__9617_ gnd vdd FILL
XFILL_3__9681_ gnd vdd FILL
XFILL_3__6893_ gnd vdd FILL
XSFILL53960x61050 gnd vdd FILL
XFILL_1__11887_ gnd vdd FILL
XFILL_4_BUFX2_insert30 gnd vdd FILL
XFILL_4_BUFX2_insert1009 gnd vdd FILL
XFILL_1__14675_ gnd vdd FILL
XFILL_4__13806_ gnd vdd FILL
XFILL_5__14056_ gnd vdd FILL
X_7462_ _7526_/Q gnd _7464_/A vdd INVX1
XFILL_3__15235_ gnd vdd FILL
XFILL_4_BUFX2_insert41 gnd vdd FILL
XFILL_2__10108_ gnd vdd FILL
XFILL_5__11268_ gnd vdd FILL
XFILL_3__8632_ gnd vdd FILL
XFILL_3__12447_ gnd vdd FILL
XFILL_1__16414_ gnd vdd FILL
XFILL_4__14786_ gnd vdd FILL
XSFILL69240x28050 gnd vdd FILL
XFILL_4_BUFX2_insert52 gnd vdd FILL
XFILL_1__13626_ gnd vdd FILL
XFILL_4__11998_ gnd vdd FILL
XFILL_0__15055_ gnd vdd FILL
XFILL_2__15965_ gnd vdd FILL
XFILL_4_BUFX2_insert63 gnd vdd FILL
XFILL_2__11088_ gnd vdd FILL
XFILL_5__9548_ gnd vdd FILL
XFILL_4_BUFX2_insert74 gnd vdd FILL
XFILL_5__13007_ gnd vdd FILL
XFILL_0__12267_ gnd vdd FILL
X_9201_ _9159_/A _9077_/CLK _8433_/R vdd _9161_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert85 gnd vdd FILL
XFILL_0__8854_ gnd vdd FILL
XFILL_4__13737_ gnd vdd FILL
XFILL_4__10949_ gnd vdd FILL
XFILL_2__10039_ gnd vdd FILL
XFILL_4_BUFX2_insert96 gnd vdd FILL
XFILL_0__14006_ gnd vdd FILL
X_7393_ _7319_/A _9188_/CLK _8929_/R vdd _7393_/D gnd vdd DFFSR
XFILL_3__15166_ gnd vdd FILL
XFILL_2__14916_ gnd vdd FILL
XFILL_5__11199_ gnd vdd FILL
XFILL_1__16345_ gnd vdd FILL
XFILL_3__12378_ gnd vdd FILL
XFILL_1__13557_ gnd vdd FILL
XFILL_0__11218_ gnd vdd FILL
XFILL_2__15896_ gnd vdd FILL
XFILL_1__10769_ gnd vdd FILL
XSFILL104440x37050 gnd vdd FILL
X_9132_ _9192_/Q gnd _9134_/A vdd INVX1
XFILL_0__12198_ gnd vdd FILL
XFILL_5__9479_ gnd vdd FILL
XFILL_0__7805_ gnd vdd FILL
XFILL_3__14117_ gnd vdd FILL
XFILL_4__13668_ gnd vdd FILL
XFILL_1__12508_ gnd vdd FILL
XFILL_0__8785_ gnd vdd FILL
XFILL_3__11329_ gnd vdd FILL
XFILL_2__14847_ gnd vdd FILL
XFILL_3__15097_ gnd vdd FILL
XSFILL8680x35050 gnd vdd FILL
XFILL_3__8494_ gnd vdd FILL
XFILL_0__11149_ gnd vdd FILL
XFILL_1__13488_ gnd vdd FILL
XFILL_1__16276_ gnd vdd FILL
XFILL_4__15407_ gnd vdd FILL
XFILL_4__12619_ gnd vdd FILL
XFILL_0__7736_ gnd vdd FILL
XFILL_2_BUFX2_insert1002 gnd vdd FILL
X_9063_ _9063_/Q _8551_/CLK _9064_/R vdd _9063_/D gnd vdd DFFSR
XFILL_4__16387_ gnd vdd FILL
XFILL_3__14048_ gnd vdd FILL
XFILL_5__14958_ gnd vdd FILL
XFILL_3_BUFX2_insert309 gnd vdd FILL
XFILL_4__13599_ gnd vdd FILL
XFILL_1__15227_ gnd vdd FILL
XFILL_1__12439_ gnd vdd FILL
XFILL_2_BUFX2_insert1013 gnd vdd FILL
XFILL_3__7445_ gnd vdd FILL
XFILL_2_BUFX2_insert1024 gnd vdd FILL
XFILL_2__14778_ gnd vdd FILL
X_8014_ _7948_/A _8014_/B gnd _8014_/Y vdd NAND2X1
XFILL_2_BUFX2_insert1035 gnd vdd FILL
XFILL_0__15957_ gnd vdd FILL
XFILL_4__15338_ gnd vdd FILL
XFILL_5__13909_ gnd vdd FILL
XFILL_2_BUFX2_insert1046 gnd vdd FILL
XFILL_2_BUFX2_insert1057 gnd vdd FILL
XFILL_1__15158_ gnd vdd FILL
XFILL_2__13729_ gnd vdd FILL
XFILL_5__14889_ gnd vdd FILL
XFILL_2_BUFX2_insert1068 gnd vdd FILL
XFILL_3__7376_ gnd vdd FILL
XFILL_0__14908_ gnd vdd FILL
XFILL_0__9406_ gnd vdd FILL
XFILL_0__15888_ gnd vdd FILL
XFILL_3__9115_ gnd vdd FILL
XFILL_0__7598_ gnd vdd FILL
XFILL_1__14109_ gnd vdd FILL
XFILL_4__15269_ gnd vdd FILL
XFILL_3__15999_ gnd vdd FILL
XFILL_1__15089_ gnd vdd FILL
XFILL_0__14839_ gnd vdd FILL
XSFILL13640x36050 gnd vdd FILL
XFILL_1__8130_ gnd vdd FILL
XFILL_0__9337_ gnd vdd FILL
X_9965_ _9965_/Q _8947_/CLK _9069_/R vdd _9917_/Y gnd vdd DFFSR
XFILL_2__16379_ gnd vdd FILL
XFILL_1__8061_ gnd vdd FILL
XFILL_0__9268_ gnd vdd FILL
X_8916_ _8916_/A _9172_/B gnd _8917_/C vdd NAND2X1
X_9896_ _9896_/A _9896_/B _9896_/C gnd _9958_/D vdd OAI21X1
XFILL_0_BUFX2_insert1050 gnd vdd FILL
XFILL_0_BUFX2_insert1061 gnd vdd FILL
XFILL_0__8219_ gnd vdd FILL
XFILL_0_BUFX2_insert1072 gnd vdd FILL
X_8847_ _8823_/B _9615_/B gnd _8847_/Y vdd NAND2X1
XSFILL104520x17050 gnd vdd FILL
XFILL_4__9790_ gnd vdd FILL
XFILL_6_BUFX2_insert920 gnd vdd FILL
XFILL_6__9726_ gnd vdd FILL
XSFILL33800x49050 gnd vdd FILL
XSFILL8760x15050 gnd vdd FILL
X_8778_ _8778_/A gnd _8778_/Y vdd INVX1
XFILL_4__8741_ gnd vdd FILL
XFILL_6_BUFX2_insert986 gnd vdd FILL
X_7729_ _7729_/A _7729_/B _7728_/Y gnd _7785_/D vdd OAI21X1
XFILL_1__8963_ gnd vdd FILL
XFILL_3__9879_ gnd vdd FILL
XSFILL23880x7050 gnd vdd FILL
XFILL_1__8894_ gnd vdd FILL
XFILL_4__7623_ gnd vdd FILL
XFILL111960x59050 gnd vdd FILL
X_11330_ _11472_/B _11321_/Y _11330_/C gnd _11440_/A vdd AOI21X1
XFILL_1__7845_ gnd vdd FILL
XSFILL13720x16050 gnd vdd FILL
XFILL_4__7554_ gnd vdd FILL
XFILL_4_BUFX2_insert110 gnd vdd FILL
X_11261_ _11731_/B _11050_/Y gnd _11261_/Y vdd NAND2X1
XFILL112040x68050 gnd vdd FILL
X_13000_ vdd _13000_/B gnd _13001_/C vdd NAND2X1
X_10212_ _14123_/A _7642_/CLK _8676_/R vdd _10146_/Y gnd vdd DFFSR
XFILL_4__7485_ gnd vdd FILL
XSFILL94200x14050 gnd vdd FILL
X_11192_ _12198_/Y gnd _11196_/A vdd INVX1
XFILL_1__9515_ gnd vdd FILL
XSFILL38920x82050 gnd vdd FILL
XFILL_4__9224_ gnd vdd FILL
XFILL_3_BUFX2_insert810 gnd vdd FILL
X_10143_ _10143_/A _10106_/A _10143_/C gnd _10211_/D vdd OAI21X1
XFILL_3_BUFX2_insert821 gnd vdd FILL
XFILL_3_BUFX2_insert832 gnd vdd FILL
XFILL_3_BUFX2_insert843 gnd vdd FILL
XFILL_3_BUFX2_insert854 gnd vdd FILL
XFILL_4__9155_ gnd vdd FILL
X_10074_ _9986_/A _9306_/CLK _9306_/R vdd _9988_/Y gnd vdd DFFSR
X_14951_ _14951_/A _14951_/B _14950_/Y gnd _14952_/A vdd NAND3X1
XFILL_3_BUFX2_insert865 gnd vdd FILL
XFILL_3_BUFX2_insert876 gnd vdd FILL
XFILL_1__9377_ gnd vdd FILL
XFILL_3_BUFX2_insert887 gnd vdd FILL
XFILL_4__8106_ gnd vdd FILL
XFILL_3_BUFX2_insert898 gnd vdd FILL
X_13902_ _13901_/Y _14901_/B _14894_/B _13902_/D gnd _13906_/B vdd OAI22X1
XFILL_4__9086_ gnd vdd FILL
XFILL_1__8328_ gnd vdd FILL
XFILL_2__7121_ gnd vdd FILL
X_14882_ _14882_/A gnd _14884_/B vdd INVX1
X_13833_ _13467_/A _13833_/B _14865_/C _13833_/D gnd _13833_/Y vdd OAI22X1
XFILL_2__7052_ gnd vdd FILL
XFILL_5__10570_ gnd vdd FILL
XFILL_1__8259_ gnd vdd FILL
XSFILL23560x19050 gnd vdd FILL
XFILL_2__10390_ gnd vdd FILL
XFILL_5__8850_ gnd vdd FILL
XFILL_3__10700_ gnd vdd FILL
X_13764_ _7900_/Q gnd _13764_/Y vdd INVX1
XFILL_6__11860_ gnd vdd FILL
X_10976_ vdd _10976_/B gnd _10977_/C vdd NAND2X1
XFILL_0__10520_ gnd vdd FILL
XFILL_5__7801_ gnd vdd FILL
XFILL_3__11680_ gnd vdd FILL
X_15503_ _7831_/A _16204_/B _16212_/A _8599_/A gnd _15503_/Y vdd AOI22X1
XFILL_6__10811_ gnd vdd FILL
X_12715_ _12713_/Y _12768_/A _12715_/C gnd _12797_/D vdd OAI21X1
XFILL_5__8781_ gnd vdd FILL
XFILL_4__9988_ gnd vdd FILL
XFILL112120x48050 gnd vdd FILL
XFILL_5__12240_ gnd vdd FILL
XFILL_2__12060_ gnd vdd FILL
XFILL_4__12970_ gnd vdd FILL
XFILL_3__10631_ gnd vdd FILL
X_13695_ _9989_/A gnd _13696_/D vdd INVX1
XFILL_1__11810_ gnd vdd FILL
XSFILL64040x33050 gnd vdd FILL
XFILL_1__12790_ gnd vdd FILL
XFILL_5__7732_ gnd vdd FILL
XFILL_0__10451_ gnd vdd FILL
XFILL_0_BUFX2_insert700 gnd vdd FILL
X_15434_ _15433_/Y _15434_/B gnd _15456_/B vdd NOR2X1
X_12646_ vdd memoryOutData[26] gnd _12647_/C vdd NAND2X1
XFILL_4__11921_ gnd vdd FILL
XFILL_0_BUFX2_insert711 gnd vdd FILL
XFILL_5__12171_ gnd vdd FILL
XFILL_2__11011_ gnd vdd FILL
XFILL_3__13350_ gnd vdd FILL
XFILL_0_BUFX2_insert722 gnd vdd FILL
XFILL_0_BUFX2_insert733 gnd vdd FILL
XFILL_1__11741_ gnd vdd FILL
XFILL_2__7954_ gnd vdd FILL
XFILL_3__10562_ gnd vdd FILL
XFILL_0_BUFX2_insert744 gnd vdd FILL
XFILL_0__13170_ gnd vdd FILL
XFILL_0__10382_ gnd vdd FILL
XFILL_0_CLKBUF1_insert170 gnd vdd FILL
XFILL_5__11122_ gnd vdd FILL
XFILL_0_CLKBUF1_insert181 gnd vdd FILL
X_15365_ _7773_/Q gnd _15366_/D vdd INVX1
XFILL_4__14640_ gnd vdd FILL
XFILL_3__12301_ gnd vdd FILL
XFILL_0_BUFX2_insert755 gnd vdd FILL
XFILL_0_CLKBUF1_insert192 gnd vdd FILL
X_12577_ vdd memoryOutData[3] gnd _12577_/Y vdd NAND2X1
XFILL_0_BUFX2_insert766 gnd vdd FILL
XFILL_2__6905_ gnd vdd FILL
XFILL_4__11852_ gnd vdd FILL
XFILL_3__13281_ gnd vdd FILL
XSFILL53880x76050 gnd vdd FILL
XFILL_1__14460_ gnd vdd FILL
XFILL_0_BUFX2_insert777 gnd vdd FILL
XFILL_0__12121_ gnd vdd FILL
XFILL_5__9402_ gnd vdd FILL
XFILL_3__10493_ gnd vdd FILL
XFILL_2__7885_ gnd vdd FILL
XFILL_0_BUFX2_insert788 gnd vdd FILL
XFILL_1__11672_ gnd vdd FILL
XFILL_0_BUFX2_insert799 gnd vdd FILL
X_14316_ _8936_/Q gnd _14316_/Y vdd INVX1
XFILL_5__15930_ gnd vdd FILL
XFILL_3__15020_ gnd vdd FILL
XFILL_5__7594_ gnd vdd FILL
X_11528_ _11571_/A _11522_/Y _11527_/Y gnd _11541_/A vdd NAND3X1
XFILL_5__11053_ gnd vdd FILL
XFILL_4__10803_ gnd vdd FILL
XFILL_4__14571_ gnd vdd FILL
XFILL_2__9624_ gnd vdd FILL
XFILL_1__13411_ gnd vdd FILL
XFILL_3__12232_ gnd vdd FILL
XSFILL3640x8050 gnd vdd FILL
X_15296_ _15296_/A _15296_/B _14791_/C gnd _12839_/B vdd AOI21X1
XFILL_2__6836_ gnd vdd FILL
XFILL_1__10623_ gnd vdd FILL
XFILL_4__11783_ gnd vdd FILL
XFILL_2__15750_ gnd vdd FILL
XFILL_2__12962_ gnd vdd FILL
XFILL_0__12052_ gnd vdd FILL
XFILL_1__14391_ gnd vdd FILL
XFILL_4__16310_ gnd vdd FILL
XFILL_5__10004_ gnd vdd FILL
X_14247_ _9318_/Q gnd _15692_/A vdd INVX1
XFILL_4__13522_ gnd vdd FILL
XFILL_2__14701_ gnd vdd FILL
X_11459_ _11411_/A _11411_/B _11184_/A gnd _11502_/B vdd AOI21X1
XFILL_5__15861_ gnd vdd FILL
XFILL_1__13342_ gnd vdd FILL
XFILL_2__11913_ gnd vdd FILL
XFILL_3__12163_ gnd vdd FILL
XFILL_2__9555_ gnd vdd FILL
XFILL_1__16130_ gnd vdd FILL
XFILL_0__11003_ gnd vdd FILL
XFILL_2__15681_ gnd vdd FILL
XFILL_1__10554_ gnd vdd FILL
XFILL_2__12893_ gnd vdd FILL
XFILL_5__9264_ gnd vdd FILL
XFILL_4__16241_ gnd vdd FILL
XFILL_5__14812_ gnd vdd FILL
XSFILL59000x22050 gnd vdd FILL
X_14178_ _14177_/Y _14593_/C gnd _14178_/Y vdd NOR2X1
XFILL_2__8506_ gnd vdd FILL
XFILL_4__13453_ gnd vdd FILL
XSFILL64200x50 gnd vdd FILL
XFILL_0__8570_ gnd vdd FILL
XFILL_3__11114_ gnd vdd FILL
XFILL_2__14632_ gnd vdd FILL
XFILL_3__12094_ gnd vdd FILL
XFILL_5__15792_ gnd vdd FILL
XFILL_4__10665_ gnd vdd FILL
XFILL_1__16061_ gnd vdd FILL
XFILL_2__9486_ gnd vdd FILL
XFILL_1__13273_ gnd vdd FILL
XFILL_5__8215_ gnd vdd FILL
XFILL_0__15811_ gnd vdd FILL
XFILL_2__11844_ gnd vdd FILL
XFILL_4__12404_ gnd vdd FILL
X_13129_ _13129_/A _13099_/B _13128_/Y gnd _13191_/D vdd OAI21X1
XFILL_3__15922_ gnd vdd FILL
XFILL_4__16172_ gnd vdd FILL
XFILL_5__11955_ gnd vdd FILL
XFILL_1__15012_ gnd vdd FILL
XFILL_5__14743_ gnd vdd FILL
XFILL_3__11045_ gnd vdd FILL
XFILL111720x21050 gnd vdd FILL
XFILL_3__7230_ gnd vdd FILL
XFILL_4__13384_ gnd vdd FILL
XFILL_1__12224_ gnd vdd FILL
XFILL112200x28050 gnd vdd FILL
XFILL_2__14563_ gnd vdd FILL
XFILL_0__12954_ gnd vdd FILL
XFILL_5__8146_ gnd vdd FILL
XFILL_0__15742_ gnd vdd FILL
XFILL_2__11775_ gnd vdd FILL
XFILL_5__10906_ gnd vdd FILL
XFILL_0__7452_ gnd vdd FILL
XFILL_4__15123_ gnd vdd FILL
XFILL_2__16302_ gnd vdd FILL
XFILL_4__12335_ gnd vdd FILL
XSFILL64120x13050 gnd vdd FILL
XFILL_5__11886_ gnd vdd FILL
XFILL_3__15853_ gnd vdd FILL
XFILL_5__14674_ gnd vdd FILL
XFILL_2__13514_ gnd vdd FILL
XFILL_0__11905_ gnd vdd FILL
XFILL_2__8368_ gnd vdd FILL
XFILL_1__12155_ gnd vdd FILL
XFILL_3__7161_ gnd vdd FILL
XSFILL89720x77050 gnd vdd FILL
XFILL_2__14494_ gnd vdd FILL
XFILL_0__15673_ gnd vdd FILL
XFILL_5__8077_ gnd vdd FILL
XFILL_5__16413_ gnd vdd FILL
XFILL_0__12885_ gnd vdd FILL
XFILL_5__13625_ gnd vdd FILL
XFILL_3__14804_ gnd vdd FILL
XFILL_4__15054_ gnd vdd FILL
XFILL_5__10837_ gnd vdd FILL
XFILL_2__16233_ gnd vdd FILL
XFILL_2__7319_ gnd vdd FILL
XFILL_4__12266_ gnd vdd FILL
XFILL_1__11106_ gnd vdd FILL
XSFILL18680x8050 gnd vdd FILL
XFILL_0__14624_ gnd vdd FILL
XFILL_2__10657_ gnd vdd FILL
XFILL_2__13445_ gnd vdd FILL
XFILL_3__15784_ gnd vdd FILL
XFILL_3__7092_ gnd vdd FILL
XFILL_3__12996_ gnd vdd FILL
XFILL_1__12086_ gnd vdd FILL
XFILL_0__11836_ gnd vdd FILL
XFILL_0__9122_ gnd vdd FILL
XFILL_4__14005_ gnd vdd FILL
XFILL_5__16344_ gnd vdd FILL
XSFILL53960x56050 gnd vdd FILL
XFILL_5__13556_ gnd vdd FILL
XFILL_4__11217_ gnd vdd FILL
XFILL_5__10768_ gnd vdd FILL
XFILL_3__14735_ gnd vdd FILL
X_9750_ _9750_/A _9813_/B _9750_/C gnd _9750_/Y vdd OAI21X1
X_6962_ _6962_/A gnd _6962_/Y vdd INVX1
XSFILL3560x20050 gnd vdd FILL
XFILL_1__15914_ gnd vdd FILL
XFILL_3__11947_ gnd vdd FILL
XFILL_4__12197_ gnd vdd FILL
XFILL_1__11037_ gnd vdd FILL
XFILL_2__16164_ gnd vdd FILL
XFILL_0__14555_ gnd vdd FILL
XFILL_2__13376_ gnd vdd FILL
XFILL_0__11767_ gnd vdd FILL
XFILL_6__14846_ gnd vdd FILL
XFILL_5__12507_ gnd vdd FILL
XSFILL28760x32050 gnd vdd FILL
X_8701_ _8698_/A _8701_/B gnd _8701_/Y vdd NAND2X1
XFILL_5__13487_ gnd vdd FILL
XFILL_4__11148_ gnd vdd FILL
XFILL_2__15115_ gnd vdd FILL
X_9681_ _9652_/B _8529_/B gnd _9682_/C vdd NAND2X1
XFILL_5__16275_ gnd vdd FILL
X_6893_ _6893_/A gnd memoryWriteData[23] vdd BUFX2
XFILL_5__10699_ gnd vdd FILL
XFILL_2__12327_ gnd vdd FILL
XFILL_3__14666_ gnd vdd FILL
XFILL_0__13506_ gnd vdd FILL
XFILL_3__11878_ gnd vdd FILL
XSFILL54040x65050 gnd vdd FILL
XFILL_2__16095_ gnd vdd FILL
XFILL_1__15845_ gnd vdd FILL
XFILL_0__14486_ gnd vdd FILL
XFILL_0__8004_ gnd vdd FILL
XSFILL33880x2050 gnd vdd FILL
XSFILL94440x70050 gnd vdd FILL
X_8632_ _8632_/A gnd _8634_/A vdd INVX1
XFILL_5__15226_ gnd vdd FILL
XFILL_3__16405_ gnd vdd FILL
XFILL_5__12438_ gnd vdd FILL
XFILL_0__11698_ gnd vdd FILL
XFILL_5__8979_ gnd vdd FILL
XFILL_3__13617_ gnd vdd FILL
XFILL_3__9802_ gnd vdd FILL
XFILL_3__10829_ gnd vdd FILL
XFILL_0__16225_ gnd vdd FILL
XFILL_4__15956_ gnd vdd FILL
XFILL_2__15046_ gnd vdd FILL
XFILL_2__12258_ gnd vdd FILL
XFILL_4__11079_ gnd vdd FILL
XFILL_6_BUFX2_insert249 gnd vdd FILL
XFILL_3__14597_ gnd vdd FILL
XFILL_0__13437_ gnd vdd FILL
XFILL_0__10649_ gnd vdd FILL
XFILL_3__7994_ gnd vdd FILL
XFILL_1__15776_ gnd vdd FILL
XFILL_1__12988_ gnd vdd FILL
XFILL_5__12369_ gnd vdd FILL
X_8563_ _8525_/A _9707_/CLK _8819_/R vdd _8563_/D gnd vdd DFFSR
XFILL_3__16336_ gnd vdd FILL
XFILL_5__15157_ gnd vdd FILL
XFILL_4__14907_ gnd vdd FILL
XSFILL33880x23050 gnd vdd FILL
XFILL_5_BUFX2_insert905 gnd vdd FILL
XSFILL104840x53050 gnd vdd FILL
XFILL_3__13548_ gnd vdd FILL
XFILL_3__9733_ gnd vdd FILL
XFILL_2__11209_ gnd vdd FILL
XFILL_2__12189_ gnd vdd FILL
XFILL_5_BUFX2_insert916 gnd vdd FILL
XFILL_3__6945_ gnd vdd FILL
XFILL_1__14727_ gnd vdd FILL
XFILL_0__16156_ gnd vdd FILL
XFILL_4__15887_ gnd vdd FILL
XFILL_0__13368_ gnd vdd FILL
XFILL_1__11939_ gnd vdd FILL
X_7514_ _7514_/Q _9306_/CLK _9306_/R vdd _7428_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert927 gnd vdd FILL
XFILL_5__14108_ gnd vdd FILL
XFILL_6__13659_ gnd vdd FILL
XFILL_5__15088_ gnd vdd FILL
XFILL_5_BUFX2_insert938 gnd vdd FILL
XFILL_4__14838_ gnd vdd FILL
XFILL_5_BUFX2_insert949 gnd vdd FILL
X_8494_ _8494_/A _8494_/B _8493_/Y gnd _8494_/Y vdd OAI21X1
XFILL_0__15107_ gnd vdd FILL
XFILL_3__16267_ gnd vdd FILL
XFILL_3__9664_ gnd vdd FILL
XFILL_0__12319_ gnd vdd FILL
XFILL_3__13479_ gnd vdd FILL
XFILL_3__6876_ gnd vdd FILL
XFILL_1__14658_ gnd vdd FILL
XFILL_0__16087_ gnd vdd FILL
XFILL_0__13299_ gnd vdd FILL
XFILL_0__8906_ gnd vdd FILL
XFILL_5__14039_ gnd vdd FILL
XFILL_3__15218_ gnd vdd FILL
X_7445_ _7472_/A _7445_/B gnd _7445_/Y vdd NAND2X1
XFILL_3__8615_ gnd vdd FILL
XFILL_0__9886_ gnd vdd FILL
XSFILL79240x1050 gnd vdd FILL
XFILL_4__14769_ gnd vdd FILL
XFILL_1__13609_ gnd vdd FILL
XFILL_3__16198_ gnd vdd FILL
XFILL_0__15038_ gnd vdd FILL
XFILL_2__15948_ gnd vdd FILL
XFILL_3__9595_ gnd vdd FILL
XFILL_1__14589_ gnd vdd FILL
XSFILL49000x54050 gnd vdd FILL
XFILL_1__7630_ gnd vdd FILL
XFILL_0__8837_ gnd vdd FILL
XFILL_3__15149_ gnd vdd FILL
X_7376_ _7376_/A gnd _7378_/A vdd INVX1
XFILL_1__16328_ gnd vdd FILL
XFILL_2__15879_ gnd vdd FILL
X_9115_ _9151_/A _8987_/B gnd _9116_/C vdd NAND2X1
XFILL_0__8768_ gnd vdd FILL
XFILL_1__7561_ gnd vdd FILL
XFILL_3_BUFX2_insert106 gnd vdd FILL
XFILL_3__8477_ gnd vdd FILL
XFILL_1__16259_ gnd vdd FILL
XFILL_1__9300_ gnd vdd FILL
XFILL_0__7719_ gnd vdd FILL
XSFILL54120x45050 gnd vdd FILL
X_9046_ _8950_/A _8022_/CLK _9046_/R vdd _9046_/D gnd vdd DFFSR
XFILL_6__8186_ gnd vdd FILL
XFILL_1__7492_ gnd vdd FILL
XFILL_3__7428_ gnd vdd FILL
XFILL_0__8699_ gnd vdd FILL
XFILL_1__9231_ gnd vdd FILL
XSFILL114680x56050 gnd vdd FILL
XFILL_3__7359_ gnd vdd FILL
XFILL_2_BUFX2_insert806 gnd vdd FILL
XFILL_2_BUFX2_insert817 gnd vdd FILL
XFILL_2_BUFX2_insert828 gnd vdd FILL
XFILL_1__9162_ gnd vdd FILL
XFILL_2_BUFX2_insert839 gnd vdd FILL
XSFILL94920x1050 gnd vdd FILL
XFILL_0_BUFX2_insert50 gnd vdd FILL
XFILL_1__8113_ gnd vdd FILL
XSFILL18760x64050 gnd vdd FILL
XFILL_0_BUFX2_insert61 gnd vdd FILL
XFILL_4__9911_ gnd vdd FILL
XSFILL8600x74050 gnd vdd FILL
XFILL_0_BUFX2_insert72 gnd vdd FILL
X_9948_ _9864_/A _9436_/CLK _7644_/R vdd _9948_/D gnd vdd DFFSR
XFILL_3__9029_ gnd vdd FILL
XFILL_1__9093_ gnd vdd FILL
XFILL_0_BUFX2_insert83 gnd vdd FILL
XSFILL39000x4050 gnd vdd FILL
X_10830_ _10831_/B _7502_/B gnd _10830_/Y vdd NAND2X1
XFILL_0_BUFX2_insert94 gnd vdd FILL
X_9879_ _9879_/A gnd _9881_/A vdd INVX1
X_10761_ _10762_/B _9737_/B gnd _10762_/C vdd NAND2X1
XSFILL23880x55050 gnd vdd FILL
X_12500_ vdd _12069_/A gnd _12500_/Y vdd NAND2X1
XBUFX2_insert805 _13490_/Y gnd _14145_/D vdd BUFX2
XFILL_4__9773_ gnd vdd FILL
XBUFX2_insert816 _13329_/Y gnd _8961_/B vdd BUFX2
XFILL_6_BUFX2_insert761 gnd vdd FILL
XFILL_4__6985_ gnd vdd FILL
XBUFX2_insert827 _13287_/Y gnd _7503_/B vdd BUFX2
X_10692_ _10736_/Q gnd _10694_/A vdd INVX1
X_13480_ _8919_/Q gnd _15095_/A vdd INVX1
XBUFX2_insert838 _13324_/Y gnd _8577_/B vdd BUFX2
XFILL_1__9995_ gnd vdd FILL
XFILL_4__8724_ gnd vdd FILL
XBUFX2_insert849 _13269_/Y gnd _7067_/A vdd BUFX2
X_12431_ _12407_/A _12654_/A gnd _12432_/C vdd NAND2X1
XFILL_4__8655_ gnd vdd FILL
X_15150_ _15150_/A _15149_/Y gnd _15156_/A vdd NOR2X1
X_12362_ _12380_/A _12362_/B gnd _12363_/C vdd NAND2X1
XFILL_1_CLKBUF1_insert210 gnd vdd FILL
XFILL_1_CLKBUF1_insert221 gnd vdd FILL
XFILL_4__7606_ gnd vdd FILL
XFILL_2__7670_ gnd vdd FILL
XFILL_1__8877_ gnd vdd FILL
X_14101_ _14101_/A _14778_/B _13420_/C _14101_/D gnd _14105_/B vdd OAI22X1
XFILL_4__8586_ gnd vdd FILL
X_11313_ _11312_/Y _11313_/B gnd _11313_/Y vdd NAND2X1
X_15081_ _15384_/A gnd _15081_/Y vdd INVX2
X_12293_ _6889_/A _12289_/B _12289_/C _12297_/D gnd _12293_/Y vdd AOI22X1
XFILL_1__7828_ gnd vdd FILL
X_14032_ _7906_/Q _13865_/B _13865_/C _7706_/A gnd _14032_/Y vdd AOI22X1
X_11244_ _11447_/B _11241_/Y gnd _11768_/B vdd NAND2X1
XSFILL84280x20050 gnd vdd FILL
XFILL_2__9340_ gnd vdd FILL
XFILL_1__7759_ gnd vdd FILL
XFILL_4__7468_ gnd vdd FILL
XSFILL99320x42050 gnd vdd FILL
X_11175_ _12192_/Y _12318_/Y gnd _11175_/Y vdd AND2X2
XFILL_4__10450_ gnd vdd FILL
XFILL_5__8000_ gnd vdd FILL
XFILL_2__9271_ gnd vdd FILL
XFILL_4__9207_ gnd vdd FILL
XFILL_1__10270_ gnd vdd FILL
X_10126_ _10206_/Q gnd _10126_/Y vdd INVX1
XFILL_3_BUFX2_insert640 gnd vdd FILL
XFILL_3_BUFX2_insert651 gnd vdd FILL
XFILL_5__11740_ gnd vdd FILL
X_15983_ _15983_/A _15978_/Y _15983_/C gnd _15984_/A vdd NAND3X1
XFILL_1__9429_ gnd vdd FILL
XFILL_2__8222_ gnd vdd FILL
XFILL_3_BUFX2_insert662 gnd vdd FILL
XFILL_4__10381_ gnd vdd FILL
XFILL_3_BUFX2_insert673 gnd vdd FILL
XFILL_2__11560_ gnd vdd FILL
XFILL_4__9138_ gnd vdd FILL
XFILL_3_BUFX2_insert684 gnd vdd FILL
XSFILL64040x28050 gnd vdd FILL
XFILL_3_BUFX2_insert695 gnd vdd FILL
X_14934_ _14934_/A _14934_/B _13574_/C _14932_/Y gnd _14934_/Y vdd OAI22X1
X_10057_ _10057_/A _10066_/B _10056_/Y gnd _10057_/Y vdd OAI21X1
XFILL_4__12120_ gnd vdd FILL
XSFILL63800x83050 gnd vdd FILL
XFILL_2__10511_ gnd vdd FILL
XFILL_5__11671_ gnd vdd FILL
XFILL_3__12850_ gnd vdd FILL
XFILL_2__11491_ gnd vdd FILL
XFILL_5__13410_ gnd vdd FILL
XFILL_5__10622_ gnd vdd FILL
XFILL_2__7104_ gnd vdd FILL
X_14865_ _14863_/Y _14865_/B _14865_/C _14864_/Y gnd _14866_/B vdd OAI22X1
XFILL_4__12051_ gnd vdd FILL
XFILL_5__14390_ gnd vdd FILL
XFILL_3__11801_ gnd vdd FILL
XFILL_2__13230_ gnd vdd FILL
XFILL_2__10442_ gnd vdd FILL
XFILL_3__12781_ gnd vdd FILL
XFILL_5__8902_ gnd vdd FILL
XFILL_2__8084_ gnd vdd FILL
XFILL_0__11621_ gnd vdd FILL
XFILL_1__13960_ gnd vdd FILL
XFILL_5__13341_ gnd vdd FILL
X_13816_ _13816_/A _13805_/Y gnd _13840_/A vdd NOR2X1
XFILL_5__9882_ gnd vdd FILL
XFILL_4__11002_ gnd vdd FILL
XFILL_3__14520_ gnd vdd FILL
XFILL_5__10553_ gnd vdd FILL
XFILL_6__12892_ gnd vdd FILL
X_14796_ _14795_/Y _13775_/B _13601_/B _14796_/D gnd _14796_/Y vdd OAI22X1
XFILL_2__13161_ gnd vdd FILL
XFILL_2__7035_ gnd vdd FILL
XFILL_3__11732_ gnd vdd FILL
XFILL_1__12911_ gnd vdd FILL
XFILL_0__14340_ gnd vdd FILL
XFILL_2__10373_ gnd vdd FILL
XFILL_5__8833_ gnd vdd FILL
XFILL_0__11552_ gnd vdd FILL
XFILL_6__14631_ gnd vdd FILL
XFILL_1__13891_ gnd vdd FILL
XFILL_5__16060_ gnd vdd FILL
XFILL_5__13272_ gnd vdd FILL
X_13747_ _8796_/Q gnd _15307_/D vdd INVX1
XFILL_2__12112_ gnd vdd FILL
XFILL_4__15810_ gnd vdd FILL
X_10959_ _10955_/A _10959_/B _10943_/C gnd _10964_/A vdd NAND3X1
XFILL_3__14451_ gnd vdd FILL
XFILL_1__15630_ gnd vdd FILL
XFILL_2__13092_ gnd vdd FILL
XFILL_3__11663_ gnd vdd FILL
XFILL_0__10503_ gnd vdd FILL
XFILL_1__12842_ gnd vdd FILL
XFILL_0__14271_ gnd vdd FILL
XFILL_5__8764_ gnd vdd FILL
XFILL_5__15011_ gnd vdd FILL
XFILL_5__12223_ gnd vdd FILL
XFILL_0__11483_ gnd vdd FILL
XFILL_3__13402_ gnd vdd FILL
XSFILL59000x17050 gnd vdd FILL
XFILL_0__16010_ gnd vdd FILL
X_13678_ _15234_/A gnd _13678_/Y vdd INVX1
XFILL_3__10614_ gnd vdd FILL
XFILL_2__12043_ gnd vdd FILL
XFILL_4__12953_ gnd vdd FILL
XFILL_4__15741_ gnd vdd FILL
XFILL_0__13222_ gnd vdd FILL
XFILL_3__14382_ gnd vdd FILL
XFILL_1__12773_ gnd vdd FILL
XFILL_5__7715_ gnd vdd FILL
XSFILL69160x61050 gnd vdd FILL
XFILL_2__8986_ gnd vdd FILL
XFILL_1__15561_ gnd vdd FILL
XFILL_0__10434_ gnd vdd FILL
XFILL_3__11594_ gnd vdd FILL
XSFILL99400x22050 gnd vdd FILL
XFILL_0_BUFX2_insert530 gnd vdd FILL
X_15417_ _9361_/A gnd _15417_/Y vdd INVX1
X_12629_ _12627_/Y vdd _12629_/C gnd _12683_/D vdd OAI21X1
XFILL_5__8695_ gnd vdd FILL
XFILL_3__16121_ gnd vdd FILL
XFILL_4__11904_ gnd vdd FILL
XFILL_5__12154_ gnd vdd FILL
XFILL_0_BUFX2_insert541 gnd vdd FILL
XFILL_3__13333_ gnd vdd FILL
XFILL_6__14493_ gnd vdd FILL
XFILL_4__15672_ gnd vdd FILL
X_16397_ gnd gnd gnd _16398_/C vdd NAND2X1
XFILL_0_BUFX2_insert552 gnd vdd FILL
XFILL_2__7937_ gnd vdd FILL
XFILL_0_BUFX2_insert563 gnd vdd FILL
XFILL_1__14512_ gnd vdd FILL
XFILL_3__10545_ gnd vdd FILL
XFILL_1__11724_ gnd vdd FILL
XFILL_4__12884_ gnd vdd FILL
XFILL_0__13153_ gnd vdd FILL
XFILL_0_BUFX2_insert574 gnd vdd FILL
XFILL_6__16232_ gnd vdd FILL
XFILL_5__11105_ gnd vdd FILL
XFILL_0__10365_ gnd vdd FILL
XFILL_1__15492_ gnd vdd FILL
XFILL_0__9740_ gnd vdd FILL
X_15348_ _15348_/A _15348_/B _15343_/Y gnd _15355_/B vdd NAND3X1
XFILL_6__13444_ gnd vdd FILL
XFILL_0_BUFX2_insert585 gnd vdd FILL
XFILL_0__6952_ gnd vdd FILL
XFILL_4__14623_ gnd vdd FILL
XSFILL104360x70050 gnd vdd FILL
XFILL_5__12085_ gnd vdd FILL
XFILL_0_BUFX2_insert596 gnd vdd FILL
XFILL_2__15802_ gnd vdd FILL
XFILL_3__16052_ gnd vdd FILL
XFILL_4__11835_ gnd vdd FILL
XFILL_3__13264_ gnd vdd FILL
XFILL_0__12104_ gnd vdd FILL
XFILL_2__7868_ gnd vdd FILL
XFILL_1__11655_ gnd vdd FILL
XFILL_1__14443_ gnd vdd FILL
XFILL_2__13994_ gnd vdd FILL
XFILL_0__13084_ gnd vdd FILL
X_7230_ _7230_/A gnd _7230_/Y vdd INVX1
XFILL_5__15913_ gnd vdd FILL
XFILL_3__15003_ gnd vdd FILL
XFILL_0__10296_ gnd vdd FILL
XFILL_5__7577_ gnd vdd FILL
XFILL_5__11036_ gnd vdd FILL
XFILL_4__14554_ gnd vdd FILL
XFILL_0__9671_ gnd vdd FILL
XFILL_3__12215_ gnd vdd FILL
XFILL_2__9607_ gnd vdd FILL
X_15279_ _16301_/A _13704_/B _15279_/C _15761_/D gnd _15280_/B vdd OAI22X1
XFILL_3__8400_ gnd vdd FILL
XFILL_0__6883_ gnd vdd FILL
XFILL_2__15733_ gnd vdd FILL
XFILL_4__11766_ gnd vdd FILL
XFILL_3__9380_ gnd vdd FILL
XFILL_0__12035_ gnd vdd FILL
XFILL_1__14374_ gnd vdd FILL
XFILL_2__7799_ gnd vdd FILL
XFILL_1__11586_ gnd vdd FILL
XFILL_0__8622_ gnd vdd FILL
XFILL_4__13505_ gnd vdd FILL
XFILL_6__12326_ gnd vdd FILL
XFILL_6__16094_ gnd vdd FILL
XFILL_5__15844_ gnd vdd FILL
X_7161_ _7161_/A gnd _7161_/Y vdd INVX1
XFILL_3__8331_ gnd vdd FILL
XFILL_4__14485_ gnd vdd FILL
XFILL_1__16113_ gnd vdd FILL
XFILL_2__9538_ gnd vdd FILL
XFILL_3__12146_ gnd vdd FILL
XSFILL3560x15050 gnd vdd FILL
XFILL_1__13325_ gnd vdd FILL
XFILL_2__15664_ gnd vdd FILL
XFILL_4__11697_ gnd vdd FILL
XFILL_1__10537_ gnd vdd FILL
XFILL_2__12876_ gnd vdd FILL
XFILL_5__9247_ gnd vdd FILL
XCLKBUF1_insert220 CLKBUF1_insert220/A gnd _7382_/CLK vdd CLKBUF1
XFILL_6__15045_ gnd vdd FILL
XFILL_4__16224_ gnd vdd FILL
XFILL_4__13436_ gnd vdd FILL
XFILL_2__14615_ gnd vdd FILL
XFILL_4__10648_ gnd vdd FILL
XFILL_5__15775_ gnd vdd FILL
X_7092_ _7092_/A _7124_/A _7091_/Y gnd _7146_/D vdd OAI21X1
XSFILL28760x27050 gnd vdd FILL
XFILL_1__13256_ gnd vdd FILL
XFILL_1__16044_ gnd vdd FILL
XFILL_3__12077_ gnd vdd FILL
XFILL_3__8262_ gnd vdd FILL
XFILL_5__12987_ gnd vdd FILL
XFILL_2__9469_ gnd vdd FILL
XFILL_2__11827_ gnd vdd FILL
XFILL_2__15595_ gnd vdd FILL
XFILL_0__13986_ gnd vdd FILL
XFILL_0__7504_ gnd vdd FILL
XFILL_6__12188_ gnd vdd FILL
XFILL_5__14726_ gnd vdd FILL
XFILL_4__16155_ gnd vdd FILL
XSFILL94440x65050 gnd vdd FILL
XFILL_3__15905_ gnd vdd FILL
XFILL_0__8484_ gnd vdd FILL
XFILL_4__13367_ gnd vdd FILL
XFILL_3__7213_ gnd vdd FILL
XFILL_5__11938_ gnd vdd FILL
XFILL_1__12207_ gnd vdd FILL
XFILL_3__11028_ gnd vdd FILL
XFILL_2__14546_ gnd vdd FILL
XFILL_4__10579_ gnd vdd FILL
XFILL_3__8193_ gnd vdd FILL
XFILL_0__15725_ gnd vdd FILL
XFILL_5__8129_ gnd vdd FILL
XFILL_2__11758_ gnd vdd FILL
XFILL_1__10399_ gnd vdd FILL
XFILL_6__11139_ gnd vdd FILL
XFILL_4__15106_ gnd vdd FILL
XFILL_0__7435_ gnd vdd FILL
XFILL_4__12318_ gnd vdd FILL
XFILL_5__14657_ gnd vdd FILL
XFILL_4__16086_ gnd vdd FILL
XFILL_4__13298_ gnd vdd FILL
XFILL_1__12138_ gnd vdd FILL
XFILL_5__11869_ gnd vdd FILL
XFILL_3__15836_ gnd vdd FILL
XFILL_2__10709_ gnd vdd FILL
XSFILL33880x18050 gnd vdd FILL
XFILL_2__14477_ gnd vdd FILL
XFILL_0__15656_ gnd vdd FILL
XFILL_0__12868_ gnd vdd FILL
XFILL_2__11689_ gnd vdd FILL
XFILL_5__13608_ gnd vdd FILL
X_9802_ _9802_/A gnd _9804_/A vdd INVX1
XFILL_4__15037_ gnd vdd FILL
XFILL_2__16216_ gnd vdd FILL
XFILL_4__12249_ gnd vdd FILL
XFILL_0__7366_ gnd vdd FILL
XFILL_5__14588_ gnd vdd FILL
XFILL_2__13428_ gnd vdd FILL
X_7994_ _7994_/A _7970_/B _7994_/C gnd _8044_/D vdd OAI21X1
XFILL_3__15767_ gnd vdd FILL
XSFILL18680x79050 gnd vdd FILL
XFILL_3__7075_ gnd vdd FILL
XFILL_0__14607_ gnd vdd FILL
XFILL_1__12069_ gnd vdd FILL
XFILL_3__12979_ gnd vdd FILL
XFILL_0__11819_ gnd vdd FILL
XSFILL104440x50050 gnd vdd FILL
XFILL_0__9105_ gnd vdd FILL
XFILL_0__15587_ gnd vdd FILL
XFILL_5__16327_ gnd vdd FILL
XFILL_0__7297_ gnd vdd FILL
X_6945_ _6967_/B _8225_/B gnd _6946_/C vdd NAND2X1
XFILL_3__14718_ gnd vdd FILL
X_9733_ _9733_/A gnd _9733_/Y vdd INVX1
XFILL_5__13539_ gnd vdd FILL
XFILL_2__16147_ gnd vdd FILL
XFILL_2__13359_ gnd vdd FILL
XFILL_3__15698_ gnd vdd FILL
XFILL_6__7824_ gnd vdd FILL
XFILL_0__14538_ gnd vdd FILL
XFILL_0__9036_ gnd vdd FILL
XFILL_5__16258_ gnd vdd FILL
X_9664_ _9664_/A _9615_/A _9664_/C gnd _9710_/D vdd OAI21X1
X_6876_ _6876_/A gnd memoryWriteData[6] vdd BUFX2
XFILL_3__14649_ gnd vdd FILL
XFILL_1__15828_ gnd vdd FILL
XFILL_2__16078_ gnd vdd FILL
XFILL_0__14469_ gnd vdd FILL
XFILL_5__15209_ gnd vdd FILL
X_8615_ _8655_/B _9383_/B gnd _8615_/Y vdd NAND2X1
XFILL_5__16189_ gnd vdd FILL
XFILL_2__15029_ gnd vdd FILL
XFILL_4__15939_ gnd vdd FILL
X_9595_ _9595_/A _9628_/B _9595_/C gnd _9687_/D vdd OAI21X1
XFILL_0__16208_ gnd vdd FILL
XFILL_5_BUFX2_insert702 gnd vdd FILL
XFILL_1__15759_ gnd vdd FILL
XFILL_3__7977_ gnd vdd FILL
XFILL_5_BUFX2_insert713 gnd vdd FILL
XFILL_5_BUFX2_insert724 gnd vdd FILL
XFILL_3__16319_ gnd vdd FILL
X_8546_ _8474_/A _6998_/CLK _8418_/R vdd _8546_/D gnd vdd DFFSR
XFILL_1__9780_ gnd vdd FILL
XFILL_5_BUFX2_insert735 gnd vdd FILL
XFILL_3__6928_ gnd vdd FILL
XFILL_1__6992_ gnd vdd FILL
XFILL_5_BUFX2_insert746 gnd vdd FILL
XFILL_6__9425_ gnd vdd FILL
XFILL_0__16139_ gnd vdd FILL
XFILL_5_BUFX2_insert757 gnd vdd FILL
XFILL_5_BUFX2_insert768 gnd vdd FILL
XFILL_1__8731_ gnd vdd FILL
XFILL_0__9938_ gnd vdd FILL
XFILL_5_BUFX2_insert779 gnd vdd FILL
X_8477_ _8477_/A gnd _8479_/A vdd INVX1
XFILL_4__8440_ gnd vdd FILL
XFILL_3__9647_ gnd vdd FILL
XFILL_3__6859_ gnd vdd FILL
XSFILL69320x21050 gnd vdd FILL
X_7428_ _7428_/A _7503_/B _7428_/C gnd _7428_/Y vdd OAI21X1
XFILL_0__9869_ gnd vdd FILL
XFILL_4__8371_ gnd vdd FILL
XFILL_1__7613_ gnd vdd FILL
X_7359_ _7359_/A _7359_/B gnd _7360_/C vdd NAND2X1
XSFILL18760x59050 gnd vdd FILL
XFILL_4__7322_ gnd vdd FILL
XSFILL104520x30050 gnd vdd FILL
XFILL_1__8593_ gnd vdd FILL
XFILL_3__8529_ gnd vdd FILL
XSFILL33800x62050 gnd vdd FILL
XFILL_1__7544_ gnd vdd FILL
XFILL_4__7253_ gnd vdd FILL
X_9029_ _9017_/A _8005_/B gnd _9030_/C vdd NAND2X1
XFILL_1__7475_ gnd vdd FILL
XFILL_4__7184_ gnd vdd FILL
XFILL_2_BUFX2_insert603 gnd vdd FILL
XFILL_1__9214_ gnd vdd FILL
XFILL_2_BUFX2_insert614 gnd vdd FILL
X_12980_ _12978_/Y vdd _12980_/C gnd _13056_/D vdd OAI21X1
XFILL_2_BUFX2_insert625 gnd vdd FILL
XFILL_2_BUFX2_insert636 gnd vdd FILL
X_11931_ _11931_/A _11921_/A _11930_/Y gnd _6852_/A vdd OAI21X1
XFILL_2_BUFX2_insert647 gnd vdd FILL
XFILL_2_BUFX2_insert658 gnd vdd FILL
XFILL_1__9145_ gnd vdd FILL
XFILL_2_BUFX2_insert669 gnd vdd FILL
XSFILL79160x24050 gnd vdd FILL
X_14650_ _14650_/A _13843_/C _14200_/C _14650_/D gnd _14654_/A vdd OAI22X1
X_11862_ _11516_/A _11862_/B gnd _11862_/Y vdd NAND2X1
X_13601_ _13599_/Y _13601_/B _13850_/B _13600_/Y gnd _13602_/A vdd OAI22X1
X_10813_ _10813_/A _10831_/B _10812_/Y gnd _10813_/Y vdd OAI21X1
X_14581_ _10427_/A gnd _14583_/A vdd INVX1
XFILL_5_BUFX2_insert18 gnd vdd FILL
XSFILL83640x49050 gnd vdd FILL
X_11793_ _11253_/B _11846_/C _11792_/Y gnd _11798_/C vdd AOI21X1
XFILL_5_BUFX2_insert29 gnd vdd FILL
X_16320_ _16320_/A _16319_/Y _15812_/C gnd _12917_/B vdd AOI21X1
XBUFX2_insert602 BUFX2_insert520/A gnd _9332_/R vdd BUFX2
X_13532_ _13532_/A _13532_/B gnd _13533_/A vdd NOR2X1
X_10744_ _10742_/Y _10762_/B _10743_/Y gnd _10838_/D vdd OAI21X1
XBUFX2_insert613 _10926_/Y gnd _12031_/A vdd BUFX2
XSFILL84280x15050 gnd vdd FILL
XFILL_2__8840_ gnd vdd FILL
XBUFX2_insert624 _12363_/Y gnd _6921_/B vdd BUFX2
XBUFX2_insert635 _12354_/Y gnd _7424_/B vdd BUFX2
XFILL_4__9756_ gnd vdd FILL
XBUFX2_insert646 _13424_/Y gnd _13813_/B vdd BUFX2
XFILL_4__6968_ gnd vdd FILL
X_16251_ _16245_/Y _16251_/B _16251_/C gnd _16259_/A vdd NAND3X1
X_13463_ _8438_/A gnd _14987_/B vdd INVX1
XBUFX2_insert657 _11988_/Y gnd _12025_/C vdd BUFX2
XSFILL99320x37050 gnd vdd FILL
XBUFX2_insert668 _12345_/Y gnd _8951_/A vdd BUFX2
X_10675_ _10676_/B _9011_/B gnd _10675_/Y vdd NAND2X1
XFILL_5__7500_ gnd vdd FILL
XFILL_4__8707_ gnd vdd FILL
XFILL_2__8771_ gnd vdd FILL
XFILL_1__9978_ gnd vdd FILL
X_15202_ _9343_/A _15202_/B _16037_/C gnd _15203_/C vdd NAND3X1
XBUFX2_insert679 _15005_/Y gnd _15392_/C vdd BUFX2
X_12414_ _12412_/Y _12368_/A _12414_/C gnd _12414_/Y vdd OAI21X1
XFILL_5__8480_ gnd vdd FILL
X_16182_ _6986_/A gnd _16183_/C vdd INVX1
XFILL_4__6899_ gnd vdd FILL
X_13394_ _13601_/B _15056_/A _14615_/B _14993_/A gnd _13394_/Y vdd OAI22X1
XFILL_2__7722_ gnd vdd FILL
XFILL_0__10150_ gnd vdd FILL
XFILL_4__8638_ gnd vdd FILL
XFILL_5__7431_ gnd vdd FILL
X_15133_ _9816_/Q gnd _15133_/Y vdd INVX1
X_12345_ _12343_/Y _12422_/A _12345_/C gnd _12345_/Y vdd OAI21X1
XFILL_4__11620_ gnd vdd FILL
XFILL_3__10261_ gnd vdd FILL
XFILL_1__11440_ gnd vdd FILL
XFILL_2__10991_ gnd vdd FILL
XFILL_5__7362_ gnd vdd FILL
XFILL_4__8569_ gnd vdd FILL
XFILL_5__12910_ gnd vdd FILL
XFILL_3__12000_ gnd vdd FILL
X_15064_ _15064_/A _15212_/B _14982_/Y gnd _15064_/Y vdd NAND3X1
X_12276_ _12272_/A _11885_/B _12272_/C gnd _12278_/B vdd NAND3X1
XFILL_4__11551_ gnd vdd FILL
XFILL_5__9101_ gnd vdd FILL
XFILL_2__12730_ gnd vdd FILL
XFILL_5__13890_ gnd vdd FILL
XFILL_3__10192_ gnd vdd FILL
XFILL_2__7584_ gnd vdd FILL
XFILL_1__11371_ gnd vdd FILL
XFILL112120x61050 gnd vdd FILL
X_14015_ _14014_/Y _13868_/B _13467_/A _14013_/Y gnd _14019_/A vdd OAI22X1
XFILL_6__12111_ gnd vdd FILL
XSFILL24440x60050 gnd vdd FILL
XFILL_4__10502_ gnd vdd FILL
XFILL_5__7293_ gnd vdd FILL
X_11227_ _11227_/A _11224_/Y gnd _11484_/B vdd NAND2X1
XFILL_5__12841_ gnd vdd FILL
XSFILL113800x47050 gnd vdd FILL
XFILL_1__13110_ gnd vdd FILL
XFILL_4__14270_ gnd vdd FILL
XFILL_1__10322_ gnd vdd FILL
XFILL_4__11482_ gnd vdd FILL
XFILL_2__12661_ gnd vdd FILL
XFILL_0__13840_ gnd vdd FILL
XFILL_1__14090_ gnd vdd FILL
XFILL_5__9032_ gnd vdd FILL
XFILL_4__13221_ gnd vdd FILL
XSFILL114440x13050 gnd vdd FILL
XFILL_5__12772_ gnd vdd FILL
XFILL_5__15560_ gnd vdd FILL
XFILL_2__14400_ gnd vdd FILL
XFILL_4__10433_ gnd vdd FILL
X_11158_ _11110_/Y _11111_/Y _11157_/Y gnd _11159_/C vdd OAI21X1
XFILL_2__9254_ gnd vdd FILL
XFILL_2__11612_ gnd vdd FILL
XFILL_3__13951_ gnd vdd FILL
XFILL_1__13041_ gnd vdd FILL
XFILL_1__10253_ gnd vdd FILL
XFILL_2__15380_ gnd vdd FILL
XSFILL114440x6050 gnd vdd FILL
XFILL_2__12592_ gnd vdd FILL
XFILL_0__13771_ gnd vdd FILL
XFILL_3_BUFX2_insert470 gnd vdd FILL
XFILL_0__10983_ gnd vdd FILL
XFILL_5__14511_ gnd vdd FILL
XFILL_3_BUFX2_insert481 gnd vdd FILL
X_10109_ _10106_/A _9597_/B gnd _10110_/C vdd NAND2X1
XFILL_2__8205_ gnd vdd FILL
XFILL_4__13152_ gnd vdd FILL
X_15966_ _15959_/Y _15965_/Y gnd _15967_/C vdd NAND2X1
XFILL_3__12902_ gnd vdd FILL
XFILL_5__11723_ gnd vdd FILL
X_11089_ _12266_/Y _11064_/Y gnd _11089_/Y vdd NOR2X1
XFILL_3_BUFX2_insert492 gnd vdd FILL
XFILL_2__14331_ gnd vdd FILL
XFILL_4__10364_ gnd vdd FILL
XFILL_5__15491_ gnd vdd FILL
XFILL_3__13882_ gnd vdd FILL
XFILL_0__12722_ gnd vdd FILL
XFILL_0__15510_ gnd vdd FILL
XFILL_2__11543_ gnd vdd FILL
XFILL_1__10184_ gnd vdd FILL
XSFILL99400x17050 gnd vdd FILL
XFILL_4__12103_ gnd vdd FILL
XFILL_0__7220_ gnd vdd FILL
X_14917_ _14908_/Y _14909_/Y _14916_/Y gnd _14917_/Y vdd NAND3X1
XFILL_3__15621_ gnd vdd FILL
XFILL_5__11654_ gnd vdd FILL
XFILL_5__14442_ gnd vdd FILL
X_15897_ _9963_/Q gnd _15899_/D vdd INVX1
XFILL_3__12833_ gnd vdd FILL
XFILL_4__13083_ gnd vdd FILL
XFILL_2__8136_ gnd vdd FILL
XFILL_4__10295_ gnd vdd FILL
XFILL_2__14262_ gnd vdd FILL
XFILL_0__15441_ gnd vdd FILL
XFILL_0__12653_ gnd vdd FILL
XFILL_2__11474_ gnd vdd FILL
XFILL_5__9934_ gnd vdd FILL
XFILL_1__14992_ gnd vdd FILL
X_14848_ _8013_/A gnd _14849_/A vdd INVX1
XFILL_2__16001_ gnd vdd FILL
XFILL_4__12034_ gnd vdd FILL
XFILL_2__13213_ gnd vdd FILL
XSFILL104360x65050 gnd vdd FILL
XFILL_3__15552_ gnd vdd FILL
XFILL_5__14373_ gnd vdd FILL
XFILL_5__11585_ gnd vdd FILL
XFILL_3__12764_ gnd vdd FILL
XFILL_2__8067_ gnd vdd FILL
XFILL_2__10425_ gnd vdd FILL
XFILL_0__11604_ gnd vdd FILL
XFILL_0__15372_ gnd vdd FILL
XFILL_2__14193_ gnd vdd FILL
XFILL_1__13943_ gnd vdd FILL
XFILL_0__12584_ gnd vdd FILL
XFILL_5__16112_ gnd vdd FILL
XFILL_5__10536_ gnd vdd FILL
XFILL_5__13324_ gnd vdd FILL
XFILL_5__9865_ gnd vdd FILL
XSFILL74280x47050 gnd vdd FILL
XFILL_3__14503_ gnd vdd FILL
XFILL_0__7082_ gnd vdd FILL
XFILL_3__11715_ gnd vdd FILL
X_14779_ _10225_/Q gnd _14779_/Y vdd INVX1
XFILL_2__13144_ gnd vdd FILL
XFILL_0__14323_ gnd vdd FILL
XFILL_3__15483_ gnd vdd FILL
XFILL_3__12695_ gnd vdd FILL
XFILL_3__8880_ gnd vdd FILL
XFILL_0__11535_ gnd vdd FILL
XFILL_1__13874_ gnd vdd FILL
XFILL_5__13255_ gnd vdd FILL
XFILL_5__16043_ gnd vdd FILL
XFILL_5__9796_ gnd vdd FILL
XSFILL89320x69050 gnd vdd FILL
XFILL112200x41050 gnd vdd FILL
XSFILL49080x23050 gnd vdd FILL
XFILL_3__14434_ gnd vdd FILL
XFILL_1__15613_ gnd vdd FILL
XFILL_3__7831_ gnd vdd FILL
XFILL_3__11646_ gnd vdd FILL
XFILL_0__14254_ gnd vdd FILL
XFILL_4__13985_ gnd vdd FILL
XFILL_1__12825_ gnd vdd FILL
XFILL_2__10287_ gnd vdd FILL
XFILL_5__12206_ gnd vdd FILL
XFILL_5__8747_ gnd vdd FILL
XFILL_0__11466_ gnd vdd FILL
X_16449_ _16449_/A gnd _16451_/A vdd INVX1
X_8400_ _8436_/Q gnd _8400_/Y vdd INVX1
X_9380_ _9359_/A _9380_/B gnd _9380_/Y vdd NAND2X1
XFILL_4__15724_ gnd vdd FILL
XFILL_2__12026_ gnd vdd FILL
XFILL_3__14365_ gnd vdd FILL
XFILL_5__10398_ gnd vdd FILL
XFILL_2__8969_ gnd vdd FILL
XFILL_1__15544_ gnd vdd FILL
XFILL_0__10417_ gnd vdd FILL
XFILL_3__11577_ gnd vdd FILL
XFILL_3__7762_ gnd vdd FILL
XFILL_1__12756_ gnd vdd FILL
XFILL_0__14185_ gnd vdd FILL
XFILL_0_BUFX2_insert360 gnd vdd FILL
X_8331_ _8413_/Q gnd _8333_/A vdd INVX1
XFILL_5__12137_ gnd vdd FILL
XFILL_3__16104_ gnd vdd FILL
XFILL_6__10708_ gnd vdd FILL
XFILL_0__11397_ gnd vdd FILL
XFILL_0_BUFX2_insert371 gnd vdd FILL
XFILL_3__13316_ gnd vdd FILL
XFILL_3__9501_ gnd vdd FILL
XFILL_0_BUFX2_insert382 gnd vdd FILL
XFILL_4__15655_ gnd vdd FILL
XFILL_0_BUFX2_insert393 gnd vdd FILL
XFILL_3__10528_ gnd vdd FILL
XFILL_4__12867_ gnd vdd FILL
XFILL_0__7984_ gnd vdd FILL
XFILL_0__13136_ gnd vdd FILL
XFILL_1__11707_ gnd vdd FILL
XFILL_3__14296_ gnd vdd FILL
XFILL_5__7629_ gnd vdd FILL
XFILL_3__7693_ gnd vdd FILL
XFILL_1__15475_ gnd vdd FILL
XFILL_4_BUFX2_insert709 gnd vdd FILL
XFILL_0__9723_ gnd vdd FILL
XFILL_4__14606_ gnd vdd FILL
XFILL_3__16035_ gnd vdd FILL
XFILL_5__12068_ gnd vdd FILL
XFILL_0__6935_ gnd vdd FILL
X_8262_ _8262_/A _8216_/A _8262_/C gnd _8304_/D vdd OAI21X1
XFILL_4__11818_ gnd vdd FILL
XFILL_3__13247_ gnd vdd FILL
XSFILL69240x36050 gnd vdd FILL
XSFILL53960x6050 gnd vdd FILL
XFILL_4__15586_ gnd vdd FILL
XFILL_1__14426_ gnd vdd FILL
XFILL_6__9141_ gnd vdd FILL
XFILL_2__13977_ gnd vdd FILL
XFILL_1__11638_ gnd vdd FILL
XFILL_0__10279_ gnd vdd FILL
X_7213_ _7207_/A _6957_/B gnd _7213_/Y vdd NAND2X1
XFILL_5__11019_ gnd vdd FILL
XFILL_0__9654_ gnd vdd FILL
X_8193_ _8191_/Y _8208_/B _8193_/C gnd _8281_/D vdd OAI21X1
XFILL_2__15716_ gnd vdd FILL
XFILL_0__6866_ gnd vdd FILL
XFILL_4__14537_ gnd vdd FILL
XFILL_4__11749_ gnd vdd FILL
XFILL_0__12018_ gnd vdd FILL
XFILL_3__9363_ gnd vdd FILL
XFILL_1__14357_ gnd vdd FILL
XFILL_1__11569_ gnd vdd FILL
XSFILL104440x45050 gnd vdd FILL
XFILL_0__8605_ gnd vdd FILL
XFILL_5__15827_ gnd vdd FILL
X_7144_ _7084_/A _7400_/CLK _9704_/R vdd _7144_/D gnd vdd DFFSR
XFILL_4__14468_ gnd vdd FILL
XFILL_3__12129_ gnd vdd FILL
XFILL_3__8314_ gnd vdd FILL
XFILL_1__13308_ gnd vdd FILL
XFILL_2__15647_ gnd vdd FILL
XSFILL8680x43050 gnd vdd FILL
XFILL_3__9294_ gnd vdd FILL
XFILL_2__12859_ gnd vdd FILL
XFILL_1__14288_ gnd vdd FILL
XFILL_4__16207_ gnd vdd FILL
XFILL_4__13419_ gnd vdd FILL
X_7075_ _7141_/Q gnd _7075_/Y vdd INVX1
XFILL_5__15758_ gnd vdd FILL
XFILL_3__8245_ gnd vdd FILL
XFILL_1__16027_ gnd vdd FILL
XFILL_4__14399_ gnd vdd FILL
XFILL_5_BUFX2_insert1050 gnd vdd FILL
XFILL_1__13239_ gnd vdd FILL
XFILL_5_BUFX2_insert1061 gnd vdd FILL
XFILL_2__15578_ gnd vdd FILL
XSFILL89400x49050 gnd vdd FILL
XFILL_5_BUFX2_insert1072 gnd vdd FILL
XFILL_5__14709_ gnd vdd FILL
XFILL_0__13969_ gnd vdd FILL
XFILL_0__8467_ gnd vdd FILL
XFILL_4__16138_ gnd vdd FILL
XFILL_5__15689_ gnd vdd FILL
XFILL_2__14529_ gnd vdd FILL
XFILL_0__15708_ gnd vdd FILL
XFILL_0__7418_ gnd vdd FILL
XFILL_6__9974_ gnd vdd FILL
XFILL_1__7191_ gnd vdd FILL
XFILL_4__16069_ gnd vdd FILL
XFILL_0__8398_ gnd vdd FILL
XFILL_3__15819_ gnd vdd FILL
XFILL_0__15639_ gnd vdd FILL
XSFILL13640x44050 gnd vdd FILL
XFILL_0__7349_ gnd vdd FILL
XFILL_4__7940_ gnd vdd FILL
XFILL_3__7058_ gnd vdd FILL
X_7977_ _8039_/Q gnd _7979_/A vdd INVX1
XSFILL13720x9050 gnd vdd FILL
X_9716_ _9680_/A _9716_/CLK _9460_/R vdd _9682_/Y gnd vdd DFFSR
X_6928_ _6926_/Y _6988_/B _6928_/C gnd _7006_/D vdd OAI21X1
XFILL_4__7871_ gnd vdd FILL
XFILL_0__9019_ gnd vdd FILL
XFILL_1__9901_ gnd vdd FILL
XFILL_4__9610_ gnd vdd FILL
X_9647_ _9647_/A gnd _9647_/Y vdd INVX1
X_6859_ _6859_/A gnd memoryAddress[21] vdd BUFX2
XFILL_5_BUFX2_insert510 gnd vdd FILL
XSFILL8760x23050 gnd vdd FILL
XFILL_5_BUFX2_insert521 gnd vdd FILL
XFILL_4__9541_ gnd vdd FILL
X_9578_ _9578_/Q _9578_/CLK _7153_/R vdd _9578_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert532 gnd vdd FILL
X_10460_ _15300_/A _7534_/CLK _8156_/R vdd _10378_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert543 gnd vdd FILL
XFILL_5_BUFX2_insert554 gnd vdd FILL
XFILL_1__9763_ gnd vdd FILL
X_8529_ _8496_/A _8529_/B gnd _8530_/C vdd NAND2X1
XFILL_1__6975_ gnd vdd FILL
XFILL_5_BUFX2_insert565 gnd vdd FILL
XFILL_3_BUFX2_insert2 gnd vdd FILL
XFILL_4__9472_ gnd vdd FILL
XFILL_5_BUFX2_insert576 gnd vdd FILL
XFILL_5_BUFX2_insert587 gnd vdd FILL
XFILL_1__8714_ gnd vdd FILL
XFILL_5_BUFX2_insert598 gnd vdd FILL
X_10391_ _10465_/Q gnd _10393_/A vdd INVX1
XFILL111960x67050 gnd vdd FILL
X_12130_ _13180_/Q gnd _12132_/A vdd INVX1
XSFILL108760x30050 gnd vdd FILL
XFILL_1__8645_ gnd vdd FILL
XSFILL13720x24050 gnd vdd FILL
XFILL_4__8354_ gnd vdd FILL
X_12061_ _12494_/B _12093_/B _12061_/C gnd gnd _12061_/Y vdd AOI22X1
XFILL112040x76050 gnd vdd FILL
XFILL_2_CLKBUF1_insert113 gnd vdd FILL
XFILL_1__8576_ gnd vdd FILL
XFILL_4__7305_ gnd vdd FILL
XFILL_2_CLKBUF1_insert124 gnd vdd FILL
XFILL_2_CLKBUF1_insert135 gnd vdd FILL
XFILL_2_CLKBUF1_insert146 gnd vdd FILL
X_11012_ _12218_/Y _11009_/Y _11011_/Y _11010_/Y gnd _11012_/Y vdd AOI22X1
XFILL_2_CLKBUF1_insert157 gnd vdd FILL
XFILL_2_CLKBUF1_insert168 gnd vdd FILL
XSFILL114360x28050 gnd vdd FILL
XFILL_2_CLKBUF1_insert179 gnd vdd FILL
XFILL_4__7236_ gnd vdd FILL
X_15820_ _15820_/A _16099_/B _15980_/C _14360_/Y gnd _15821_/C vdd OAI22X1
XFILL_2_BUFX2_insert400 gnd vdd FILL
XFILL_1__7458_ gnd vdd FILL
XFILL_2_BUFX2_insert411 gnd vdd FILL
XFILL_4__7167_ gnd vdd FILL
XFILL_2_BUFX2_insert422 gnd vdd FILL
XFILL_2_BUFX2_insert433 gnd vdd FILL
X_15751_ _7081_/A gnd _15751_/Y vdd INVX1
XFILL_2_BUFX2_insert444 gnd vdd FILL
X_12963_ _6874_/A gnd _12963_/Y vdd INVX1
XFILL_2_BUFX2_insert455 gnd vdd FILL
XFILL_2_BUFX2_insert466 gnd vdd FILL
X_14702_ _14702_/A _14694_/Y _14701_/Y gnd _14702_/Y vdd NAND3X1
XFILL_4__7098_ gnd vdd FILL
X_11914_ _11914_/A gnd _11916_/A vdd INVX1
XFILL_2_BUFX2_insert477 gnd vdd FILL
XFILL_5__7980_ gnd vdd FILL
X_15682_ _7909_/Q gnd _15683_/A vdd INVX1
XFILL_1__9128_ gnd vdd FILL
XFILL_2_BUFX2_insert488 gnd vdd FILL
X_12894_ _12892_/Y vdd _12894_/C gnd _12894_/Y vdd OAI21X1
XFILL_2_BUFX2_insert499 gnd vdd FILL
XFILL_5__6931_ gnd vdd FILL
X_14633_ _13871_/D _14631_/Y _13857_/C _14632_/Y gnd _14637_/B vdd OAI22X1
XFILL_5__11370_ gnd vdd FILL
X_11845_ _11837_/Y _11845_/B _11844_/Y gnd _11849_/B vdd OAI21X1
XFILL_2__9941_ gnd vdd FILL
XFILL_2__11190_ gnd vdd FILL
XFILL_1__10940_ gnd vdd FILL
XFILL_5__9650_ gnd vdd FILL
XFILL_5__6862_ gnd vdd FILL
XFILL_5__10321_ gnd vdd FILL
XFILL_6__12660_ gnd vdd FILL
X_14564_ _14562_/Y _14174_/C _13617_/D _14563_/Y gnd _14568_/A vdd OAI22X1
XSFILL63960x32050 gnd vdd FILL
XFILL_3__11500_ gnd vdd FILL
XFILL_2__10141_ gnd vdd FILL
X_11776_ _11776_/A _11776_/B _11776_/C gnd _11784_/C vdd OAI21X1
XFILL_2__9872_ gnd vdd FILL
XFILL_5__8601_ gnd vdd FILL
XBUFX2_insert410 _13484_/Y gnd _13884_/C vdd BUFX2
XFILL_3__12480_ gnd vdd FILL
XFILL_0__11320_ gnd vdd FILL
XBUFX2_insert421 _14991_/Y gnd _15636_/B vdd BUFX2
X_16303_ _9461_/Q _15044_/C _15071_/C gnd _16304_/C vdd NAND3X1
XFILL_1__10871_ gnd vdd FILL
XFILL_4__9808_ gnd vdd FILL
XFILL112120x56050 gnd vdd FILL
XFILL_5__13040_ gnd vdd FILL
XBUFX2_insert432 _13326_/Y gnd _8788_/A vdd BUFX2
X_13515_ _9593_/A gnd _13517_/D vdd INVX1
XFILL_5__10252_ gnd vdd FILL
X_10727_ _10727_/Q _7400_/CLK _9704_/R vdd _10667_/Y gnd vdd DFFSR
X_14495_ _9195_/Q gnd _14495_/Y vdd INVX1
XFILL_2__8823_ gnd vdd FILL
XFILL_4__13770_ gnd vdd FILL
XBUFX2_insert443 _12378_/Y gnd _8600_/B vdd BUFX2
XFILL_3__11431_ gnd vdd FILL
XBUFX2_insert454 _13276_/Y gnd _7181_/B vdd BUFX2
XFILL_4__10982_ gnd vdd FILL
XFILL_1__12610_ gnd vdd FILL
XSFILL64040x41050 gnd vdd FILL
XFILL_1__13590_ gnd vdd FILL
XSFILL64840x60050 gnd vdd FILL
XFILL_5__8532_ gnd vdd FILL
XFILL_0__11251_ gnd vdd FILL
XBUFX2_insert465 _13318_/Y gnd _8372_/B vdd BUFX2
X_16234_ _10739_/Q gnd _16234_/Y vdd INVX1
XFILL_4__9739_ gnd vdd FILL
XBUFX2_insert476 _15038_/Y gnd _15527_/A vdd BUFX2
XFILL_4__12721_ gnd vdd FILL
X_13446_ _7030_/A gnd _13449_/A vdd INVX1
XBUFX2_insert487 _12372_/Y gnd _7954_/B vdd BUFX2
XFILL_3__14150_ gnd vdd FILL
X_10658_ _10656_/Y _10658_/B _10657_/Y gnd _10724_/D vdd OAI21X1
XFILL_5__10183_ gnd vdd FILL
XFILL_2__13900_ gnd vdd FILL
XBUFX2_insert498 BUFX2_insert524/A gnd _7665_/R vdd BUFX2
XFILL_2__8754_ gnd vdd FILL
XFILL_3__11362_ gnd vdd FILL
XFILL_2__14880_ gnd vdd FILL
XSFILL2840x82050 gnd vdd FILL
XFILL_5__8463_ gnd vdd FILL
XFILL_0__11182_ gnd vdd FILL
XFILL_3__13101_ gnd vdd FILL
X_16165_ _8778_/A _15821_/B _15978_/C _8522_/A gnd _16172_/A vdd AOI22X1
XFILL_4__12652_ gnd vdd FILL
X_13377_ _11884_/A _12808_/Q _12807_/Q gnd _13377_/Y vdd NOR3X1
XFILL_2__7705_ gnd vdd FILL
XFILL_3__10313_ gnd vdd FILL
XFILL_4__15440_ gnd vdd FILL
X_10589_ _10589_/Q _9963_/CLK _9963_/R vdd _10509_/Y gnd vdd DFFSR
XFILL_2__13831_ gnd vdd FILL
XFILL_5__14991_ gnd vdd FILL
XFILL_3__14081_ gnd vdd FILL
XFILL_5__7414_ gnd vdd FILL
XFILL_1__12472_ gnd vdd FILL
XFILL_3__11293_ gnd vdd FILL
XFILL_0__10133_ gnd vdd FILL
XFILL_1__15260_ gnd vdd FILL
X_15116_ _13530_/A gnd _15116_/Y vdd INVX1
XFILL_5__8394_ gnd vdd FILL
XFILL_0__15990_ gnd vdd FILL
XFILL_6__10424_ gnd vdd FILL
X_12328_ _12312_/A _12340_/B _12312_/C gnd _12328_/Y vdd NAND3X1
XFILL_4__11603_ gnd vdd FILL
XFILL_4__15371_ gnd vdd FILL
X_16096_ _6980_/A _15382_/B _16096_/C _7364_/A gnd _16096_/Y vdd AOI22X1
XFILL_3__13032_ gnd vdd FILL
XFILL_5__13942_ gnd vdd FILL
XFILL_1__14211_ gnd vdd FILL
XFILL_4__12583_ gnd vdd FILL
XFILL_3__10244_ gnd vdd FILL
XFILL_2__7636_ gnd vdd FILL
XFILL_1__11423_ gnd vdd FILL
XFILL_2__13762_ gnd vdd FILL
XFILL_2__10974_ gnd vdd FILL
XFILL_1__15191_ gnd vdd FILL
XFILL_0__14941_ gnd vdd FILL
XFILL_5__7345_ gnd vdd FILL
XFILL_0__10064_ gnd vdd FILL
X_15047_ _14983_/A _16035_/B _15024_/C gnd _15047_/Y vdd NAND3X1
XFILL_4__14322_ gnd vdd FILL
XFILL_2__15501_ gnd vdd FILL
X_12259_ _12255_/A gnd _12255_/C gnd _12259_/Y vdd NAND3X1
XFILL_4__11534_ gnd vdd FILL
XFILL_5__13873_ gnd vdd FILL
XFILL_2__12713_ gnd vdd FILL
XFILL_2__7567_ gnd vdd FILL
XFILL_3__10175_ gnd vdd FILL
XFILL_1__14142_ gnd vdd FILL
XFILL_1__11354_ gnd vdd FILL
XFILL_2__13693_ gnd vdd FILL
XFILL_0__14872_ gnd vdd FILL
XFILL_5__15612_ gnd vdd FILL
XFILL_1_BUFX2_insert16 gnd vdd FILL
XSFILL59000x30050 gnd vdd FILL
XFILL_4__14253_ gnd vdd FILL
XFILL_5__12824_ gnd vdd FILL
XFILL_0__9370_ gnd vdd FILL
XFILL_1_BUFX2_insert27 gnd vdd FILL
XFILL_1__10305_ gnd vdd FILL
XFILL_2__15432_ gnd vdd FILL
XFILL_4__11465_ gnd vdd FILL
XFILL_1_BUFX2_insert38 gnd vdd FILL
XFILL_5__9015_ gnd vdd FILL
XFILL_2__12644_ gnd vdd FILL
XFILL_3__14983_ gnd vdd FILL
XFILL_1__14073_ gnd vdd FILL
XFILL_0__13823_ gnd vdd FILL
XFILL_2__7498_ gnd vdd FILL
XFILL_1_BUFX2_insert49 gnd vdd FILL
XFILL_1__11285_ gnd vdd FILL
XFILL_0__8321_ gnd vdd FILL
XFILL_5__15543_ gnd vdd FILL
XFILL_4__10416_ gnd vdd FILL
XFILL_5__12755_ gnd vdd FILL
XFILL_4__14184_ gnd vdd FILL
XFILL_1__13024_ gnd vdd FILL
XFILL_3__13934_ gnd vdd FILL
XFILL_2__9237_ gnd vdd FILL
XSFILL49080x18050 gnd vdd FILL
XFILL_2__15363_ gnd vdd FILL
XFILL112200x36050 gnd vdd FILL
XFILL_4__11396_ gnd vdd FILL
XFILL_1__10236_ gnd vdd FILL
XFILL_2__12575_ gnd vdd FILL
XFILL_0__10966_ gnd vdd FILL
XFILL_0__13754_ gnd vdd FILL
XFILL_0__8252_ gnd vdd FILL
X_7900_ _7900_/Q _7534_/CLK _8156_/R vdd _7900_/D gnd vdd DFFSR
XFILL_4__13135_ gnd vdd FILL
XFILL_5__11706_ gnd vdd FILL
XSFILL64120x21050 gnd vdd FILL
X_15949_ _15946_/Y _15948_/Y gnd _15949_/Y vdd NOR2X1
XFILL_2__14314_ gnd vdd FILL
XFILL_5__15474_ gnd vdd FILL
XFILL_3__13865_ gnd vdd FILL
X_8880_ _8902_/B _9008_/B gnd _8881_/C vdd NAND2X1
XFILL_2__11526_ gnd vdd FILL
XFILL_2__9168_ gnd vdd FILL
XFILL_0__12705_ gnd vdd FILL
XFILL_1__10167_ gnd vdd FILL
XFILL_2__15294_ gnd vdd FILL
XFILL_0__7203_ gnd vdd FILL
XFILL_0__13685_ gnd vdd FILL
XFILL_0__10897_ gnd vdd FILL
XFILL_5__14425_ gnd vdd FILL
XFILL_2__8119_ gnd vdd FILL
X_7831_ _7831_/A gnd _7833_/A vdd INVX1
XFILL_6__13976_ gnd vdd FILL
XFILL_0__8183_ gnd vdd FILL
XFILL_5__11637_ gnd vdd FILL
XFILL_3__15604_ gnd vdd FILL
XFILL_2__14245_ gnd vdd FILL
XFILL_4__10278_ gnd vdd FILL
XSFILL27880x12050 gnd vdd FILL
XFILL_2__9099_ gnd vdd FILL
XFILL_0__12636_ gnd vdd FILL
XFILL_3__13796_ gnd vdd FILL
XFILL_3__9981_ gnd vdd FILL
XFILL_0__15424_ gnd vdd FILL
XFILL_2__11457_ gnd vdd FILL
XFILL_5__9917_ gnd vdd FILL
XFILL_6__15715_ gnd vdd FILL
XFILL_1__14975_ gnd vdd FILL
XSFILL53960x64050 gnd vdd FILL
XFILL_4__12017_ gnd vdd FILL
XFILL_3__15535_ gnd vdd FILL
XFILL_5__14356_ gnd vdd FILL
XFILL_5__11568_ gnd vdd FILL
XFILL_3__12747_ gnd vdd FILL
XFILL_2__10408_ gnd vdd FILL
X_7762_ _7762_/A _7729_/B _7761_/Y gnd _7796_/D vdd OAI21X1
XFILL_2__14176_ gnd vdd FILL
XFILL_1__13926_ gnd vdd FILL
XSFILL13960x80050 gnd vdd FILL
XFILL_0__12567_ gnd vdd FILL
XFILL_0__15355_ gnd vdd FILL
XFILL_2__11388_ gnd vdd FILL
XFILL_5__13307_ gnd vdd FILL
XFILL_5__9848_ gnd vdd FILL
XSFILL28760x40050 gnd vdd FILL
X_9501_ _9501_/A gnd _9501_/Y vdd INVX1
XFILL_5__10519_ gnd vdd FILL
XFILL_0__7065_ gnd vdd FILL
X_7693_ _7691_/Y _7759_/B _7693_/C gnd _7773_/D vdd OAI21X1
XFILL_2__13127_ gnd vdd FILL
XFILL_5__11499_ gnd vdd FILL
XFILL_3__15466_ gnd vdd FILL
XFILL_5__14287_ gnd vdd FILL
XSFILL54040x73050 gnd vdd FILL
XFILL_3__8863_ gnd vdd FILL
XFILL_0__11518_ gnd vdd FILL
XFILL_0__14306_ gnd vdd FILL
XFILL_1__13857_ gnd vdd FILL
XFILL_0__15286_ gnd vdd FILL
XFILL_5__16026_ gnd vdd FILL
XFILL_0__12498_ gnd vdd FILL
XFILL_6__11809_ gnd vdd FILL
XFILL_5__13238_ gnd vdd FILL
X_9432_ _9340_/A _7640_/CLK _7000_/R vdd _9432_/D gnd vdd DFFSR
XFILL_6__15577_ gnd vdd FILL
XFILL_5__9779_ gnd vdd FILL
XFILL_3__14417_ gnd vdd FILL
XFILL_6__12789_ gnd vdd FILL
XFILL_3__11629_ gnd vdd FILL
XFILL_3__7814_ gnd vdd FILL
XFILL_3__15397_ gnd vdd FILL
XFILL_0__14237_ gnd vdd FILL
XFILL_4__13968_ gnd vdd FILL
XFILL_0__11449_ gnd vdd FILL
XFILL_1__13788_ gnd vdd FILL
XFILL_6__14528_ gnd vdd FILL
XFILL_4__15707_ gnd vdd FILL
XFILL_5__13169_ gnd vdd FILL
XFILL_2__12009_ gnd vdd FILL
XFILL_3__14348_ gnd vdd FILL
X_9363_ _9363_/A _9425_/A _9362_/Y gnd _9439_/D vdd OAI21X1
XFILL_1__15527_ gnd vdd FILL
XFILL_3__7745_ gnd vdd FILL
XFILL_1__12739_ gnd vdd FILL
XFILL_0__14168_ gnd vdd FILL
XFILL_4__13899_ gnd vdd FILL
XFILL_4_BUFX2_insert506 gnd vdd FILL
X_8314_ _8315_/B _8314_/B gnd _8314_/Y vdd NAND2X1
X_9294_ _9232_/B _8910_/B gnd _9295_/C vdd NAND2X1
XFILL_4__15638_ gnd vdd FILL
XFILL_0__7967_ gnd vdd FILL
XFILL_0__13119_ gnd vdd FILL
XFILL_4_BUFX2_insert517 gnd vdd FILL
XFILL_3__14279_ gnd vdd FILL
XFILL_4_BUFX2_insert528 gnd vdd FILL
XFILL_3__7676_ gnd vdd FILL
XFILL_1__15458_ gnd vdd FILL
XFILL_4_BUFX2_insert539 gnd vdd FILL
XFILL_0__14099_ gnd vdd FILL
X_8245_ _8299_/Q gnd _8245_/Y vdd INVX1
XFILL_3__16018_ gnd vdd FILL
XFILL_0__6918_ gnd vdd FILL
XFILL_3__9415_ gnd vdd FILL
XFILL_4__15569_ gnd vdd FILL
XFILL_1__14409_ gnd vdd FILL
XFILL_1__15389_ gnd vdd FILL
XSFILL49000x62050 gnd vdd FILL
XFILL_0__9637_ gnd vdd FILL
XSFILL13640x39050 gnd vdd FILL
XFILL_0__6849_ gnd vdd FILL
X_8176_ _8132_/A _8176_/CLK _8176_/R vdd _8176_/D gnd vdd DFFSR
XFILL_3__9346_ gnd vdd FILL
XSFILL109560x73050 gnd vdd FILL
X_7127_ _7127_/Q _7515_/CLK _7000_/R vdd _7127_/D gnd vdd DFFSR
XSFILL13240x41050 gnd vdd FILL
XFILL_1__8361_ gnd vdd FILL
XFILL_3__9277_ gnd vdd FILL
XFILL_4__8070_ gnd vdd FILL
XFILL_1__7312_ gnd vdd FILL
XFILL_0__8519_ gnd vdd FILL
XSFILL54120x53050 gnd vdd FILL
XSFILL23880x50 gnd vdd FILL
X_7058_ _7064_/A _7314_/B gnd _7058_/Y vdd NAND2X1
XFILL_3__8228_ gnd vdd FILL
XFILL_0__9499_ gnd vdd FILL
XFILL_3_CLKBUF1_insert208 gnd vdd FILL
XFILL_3_CLKBUF1_insert219 gnd vdd FILL
XFILL_1__7243_ gnd vdd FILL
XSFILL33960x11050 gnd vdd FILL
XFILL_1__7174_ gnd vdd FILL
XFILL_1_BUFX2_insert407 gnd vdd FILL
XFILL_4__8972_ gnd vdd FILL
XFILL_1_BUFX2_insert418 gnd vdd FILL
XFILL_6__8908_ gnd vdd FILL
XFILL_1_BUFX2_insert429 gnd vdd FILL
XSFILL18760x72050 gnd vdd FILL
X_11630_ _11615_/Y _11630_/B gnd _11630_/Y vdd NAND2X1
XFILL_4__7854_ gnd vdd FILL
XFILL_1_CLKBUF1_insert1075 gnd vdd FILL
X_11561_ _11561_/A _11311_/Y gnd _11577_/B vdd NAND2X1
XSFILL23080x44050 gnd vdd FILL
X_13300_ _13297_/A _13300_/B gnd _13300_/Y vdd OR2X2
XSFILL109640x53050 gnd vdd FILL
X_10512_ _10510_/Y _10511_/A _10512_/C gnd _10590_/D vdd OAI21X1
X_14280_ _7015_/Q gnd _15761_/C vdd INVX1
XFILL_5_BUFX2_insert340 gnd vdd FILL
X_11492_ _11492_/A _11492_/B gnd _11492_/Y vdd AND2X2
XBUFX2_insert30 _13320_/Y gnd _8484_/A vdd BUFX2
XFILL_5_BUFX2_insert351 gnd vdd FILL
XFILL_4__9524_ gnd vdd FILL
XBUFX2_insert41 _13265_/Y gnd _6937_/B vdd BUFX2
XSFILL54200x33050 gnd vdd FILL
XFILL_5_BUFX2_insert362 gnd vdd FILL
XSFILL69240x9050 gnd vdd FILL
X_13231_ _13231_/A _13231_/B gnd _13294_/A vdd NAND2X1
XFILL_5_BUFX2_insert373 gnd vdd FILL
XBUFX2_insert52 _13309_/Y gnd _8082_/A vdd BUFX2
X_10443_ _10443_/A _7499_/B gnd _10443_/Y vdd NAND2X1
XFILL_5_BUFX2_insert384 gnd vdd FILL
XBUFX2_insert63 _12215_/Y gnd _12249_/B vdd BUFX2
XBUFX2_insert74 _12366_/Y gnd _9100_/B vdd BUFX2
XFILL_1__9746_ gnd vdd FILL
XFILL_1__6958_ gnd vdd FILL
XFILL_5_BUFX2_insert395 gnd vdd FILL
XBUFX2_insert85 _13390_/Y gnd _14725_/A vdd BUFX2
XBUFX2_insert96 _15068_/Y gnd _15328_/B vdd BUFX2
X_13162_ _13160_/Y _13173_/A _13162_/C gnd _13202_/D vdd OAI21X1
X_10374_ _10363_/B _9478_/B gnd _10375_/C vdd NAND2X1
XFILL_1__9677_ gnd vdd FILL
XFILL_2__8470_ gnd vdd FILL
XFILL_1__6889_ gnd vdd FILL
X_12113_ _12113_/A _12113_/B _12113_/C gnd gnd _12113_/Y vdd AOI22X1
XFILL_4__9386_ gnd vdd FILL
X_13093_ _13093_/A _13099_/B _13093_/C gnd _13179_/D vdd OAI21X1
XFILL_2__7421_ gnd vdd FILL
XFILL_1__8628_ gnd vdd FILL
XSFILL84120x69050 gnd vdd FILL
XFILL_4__8337_ gnd vdd FILL
XFILL_6__10140_ gnd vdd FILL
X_12044_ _12028_/A _11876_/B _12024_/C gnd _12046_/B vdd NAND3X1
XFILL_5__10870_ gnd vdd FILL
XFILL_2__7352_ gnd vdd FILL
XFILL_4__8268_ gnd vdd FILL
XFILL_2__10690_ gnd vdd FILL
XFILL_5__7061_ gnd vdd FILL
XSFILL99320x50050 gnd vdd FILL
XFILL_4__11250_ gnd vdd FILL
XFILL_3__11980_ gnd vdd FILL
XFILL_0__10820_ gnd vdd FILL
XFILL_1__11070_ gnd vdd FILL
XFILL_4__7219_ gnd vdd FILL
XSFILL84920x9050 gnd vdd FILL
X_15803_ _15801_/Y _15803_/B gnd _15803_/Y vdd NOR2X1
XFILL_4__8199_ gnd vdd FILL
XFILL_2__9022_ gnd vdd FILL
XFILL_3__10931_ gnd vdd FILL
XFILL_1__10021_ gnd vdd FILL
X_13995_ _13995_/A _13680_/B _14466_/C _13995_/D gnd _13995_/Y vdd OAI22X1
XFILL_2_BUFX2_insert230 gnd vdd FILL
XFILL_4__11181_ gnd vdd FILL
XFILL_2_BUFX2_insert241 gnd vdd FILL
XFILL_2__12360_ gnd vdd FILL
XFILL112280x10050 gnd vdd FILL
XFILL_0__10751_ gnd vdd FILL
XFILL_2_BUFX2_insert252 gnd vdd FILL
XSFILL64040x36050 gnd vdd FILL
XFILL_2_BUFX2_insert263 gnd vdd FILL
X_15734_ _8039_/Q _15081_/Y gnd _15736_/A vdd NAND2X1
XFILL_2_BUFX2_insert274 gnd vdd FILL
XFILL_5__12471_ gnd vdd FILL
X_12946_ _12946_/Q _9328_/CLK _7920_/R vdd _12906_/Y gnd vdd DFFSR
XFILL_4__10132_ gnd vdd FILL
XFILL_3__13650_ gnd vdd FILL
XFILL_2__11311_ gnd vdd FILL
XFILL_2_BUFX2_insert285 gnd vdd FILL
XFILL_2_BUFX2_insert296 gnd vdd FILL
XFILL_0__13470_ gnd vdd FILL
XFILL_2__12291_ gnd vdd FILL
XFILL_5__14210_ gnd vdd FILL
XFILL_5__7963_ gnd vdd FILL
XFILL_0__10682_ gnd vdd FILL
XFILL_5__11422_ gnd vdd FILL
XFILL_3__12601_ gnd vdd FILL
X_15665_ _14190_/Y _15386_/B _15386_/C _15665_/D gnd _15666_/A vdd OAI22X1
XFILL_6__13761_ gnd vdd FILL
XFILL_4__10063_ gnd vdd FILL
XFILL_5__15190_ gnd vdd FILL
XFILL_2__14030_ gnd vdd FILL
XFILL_4__14940_ gnd vdd FILL
X_12877_ _12170_/B gnd _12877_/Y vdd INVX1
XFILL_1_BUFX2_insert930 gnd vdd FILL
XSFILL53880x79050 gnd vdd FILL
XFILL_0__12421_ gnd vdd FILL
XFILL_3__13581_ gnd vdd FILL
XFILL_2__11242_ gnd vdd FILL
XFILL_1_BUFX2_insert941 gnd vdd FILL
XFILL_5__6914_ gnd vdd FILL
XFILL_6__15500_ gnd vdd FILL
XFILL_3__10793_ gnd vdd FILL
XFILL_1__14760_ gnd vdd FILL
XFILL_6__12712_ gnd vdd FILL
X_14616_ _14616_/A _14615_/Y gnd _14617_/C vdd NOR2X1
XFILL_1__11972_ gnd vdd FILL
XFILL_1_BUFX2_insert952 gnd vdd FILL
XFILL_1_BUFX2_insert963 gnd vdd FILL
XFILL_3__15320_ gnd vdd FILL
XFILL_5__14141_ gnd vdd FILL
X_11828_ _11828_/A _11828_/B _11827_/Y gnd _11828_/Y vdd NAND3X1
XFILL_5__11353_ gnd vdd FILL
XFILL_1_BUFX2_insert974 gnd vdd FILL
XFILL_3__12532_ gnd vdd FILL
X_15596_ _16306_/A _14089_/Y _16306_/C _14083_/D gnd _15596_/Y vdd OAI22X1
XFILL_4__14871_ gnd vdd FILL
XFILL_2__9924_ gnd vdd FILL
XFILL_0__15140_ gnd vdd FILL
XFILL_1__13711_ gnd vdd FILL
XFILL_2__11173_ gnd vdd FILL
XFILL_1_BUFX2_insert985 gnd vdd FILL
XFILL_0__12352_ gnd vdd FILL
XFILL_1__10923_ gnd vdd FILL
XFILL_1_BUFX2_insert996 gnd vdd FILL
XFILL_5__10304_ gnd vdd FILL
XFILL_5__6845_ gnd vdd FILL
XFILL_5__9633_ gnd vdd FILL
XFILL_1__14691_ gnd vdd FILL
X_14547_ _14547_/A _14547_/B _14546_/Y gnd _14548_/B vdd NAND3X1
XFILL_5__14072_ gnd vdd FILL
XFILL_2__10124_ gnd vdd FILL
XFILL_4__13822_ gnd vdd FILL
XFILL_3__15251_ gnd vdd FILL
XFILL_5__11284_ gnd vdd FILL
X_11759_ _11037_/Y gnd _11761_/A vdd INVX1
XFILL_2__9855_ gnd vdd FILL
XFILL_3__12463_ gnd vdd FILL
XBUFX2_insert240 _15065_/Y gnd _15239_/B vdd BUFX2
XFILL_0__11303_ gnd vdd FILL
XFILL_2__15981_ gnd vdd FILL
XFILL_1__13642_ gnd vdd FILL
XFILL_0__15071_ gnd vdd FILL
XBUFX2_insert251 _10922_/Y gnd _15812_/C vdd BUFX2
XFILL_5__13023_ gnd vdd FILL
XFILL_0__12283_ gnd vdd FILL
XFILL_3__14202_ gnd vdd FILL
XFILL_6__15362_ gnd vdd FILL
XFILL_5__10235_ gnd vdd FILL
XBUFX2_insert262 _11225_/Y gnd _11748_/A vdd BUFX2
XSFILL59000x25050 gnd vdd FILL
XFILL_0__8870_ gnd vdd FILL
XBUFX2_insert273 _13364_/Y gnd _10661_/B vdd BUFX2
X_14478_ _7915_/Q gnd _14478_/Y vdd INVX1
XFILL_3__11414_ gnd vdd FILL
XFILL_4__10965_ gnd vdd FILL
XFILL_3__15182_ gnd vdd FILL
XFILL_4__13753_ gnd vdd FILL
XFILL_0__14022_ gnd vdd FILL
XBUFX2_insert284 _15003_/Y gnd _15558_/D vdd BUFX2
XFILL_2__14932_ gnd vdd FILL
XFILL_2__10055_ gnd vdd FILL
XBUFX2_insert295 _13356_/Y gnd _10294_/A vdd BUFX2
XFILL_3__12394_ gnd vdd FILL
XFILL_2__9786_ gnd vdd FILL
XSFILL99400x30050 gnd vdd FILL
XFILL_1__16361_ gnd vdd FILL
XFILL_5__8515_ gnd vdd FILL
XFILL_0__11234_ gnd vdd FILL
X_16217_ _16217_/A _16216_/Y _15656_/C gnd _16217_/Y vdd NOR3X1
XFILL_1__10785_ gnd vdd FILL
XFILL_1__13573_ gnd vdd FILL
XFILL_5_CLKBUF1_insert130 gnd vdd FILL
XFILL_0__7821_ gnd vdd FILL
XFILL_5_CLKBUF1_insert141 gnd vdd FILL
XFILL_5__9495_ gnd vdd FILL
X_13429_ _13423_/A _13418_/A _13404_/B gnd _14045_/A vdd NAND3X1
XFILL_4__12704_ gnd vdd FILL
XFILL_5__10166_ gnd vdd FILL
XFILL_3__14133_ gnd vdd FILL
XFILL_1__15312_ gnd vdd FILL
XFILL_4__13684_ gnd vdd FILL
XFILL_2__8737_ gnd vdd FILL
XFILL_5_CLKBUF1_insert152 gnd vdd FILL
XFILL_3__11345_ gnd vdd FILL
XFILL_2__14863_ gnd vdd FILL
XFILL_1__12524_ gnd vdd FILL
XFILL_4__10896_ gnd vdd FILL
XFILL_5_CLKBUF1_insert163 gnd vdd FILL
XFILL_1__16292_ gnd vdd FILL
XFILL_0__11165_ gnd vdd FILL
XFILL_5__8446_ gnd vdd FILL
XFILL_5_CLKBUF1_insert174 gnd vdd FILL
XFILL_5_CLKBUF1_insert185 gnd vdd FILL
X_16148_ _9457_/Q _15945_/C _16148_/C gnd _16148_/Y vdd NAND3X1
XFILL_4__12635_ gnd vdd FILL
XFILL_5_CLKBUF1_insert196 gnd vdd FILL
XFILL_6__11456_ gnd vdd FILL
XFILL_4__15423_ gnd vdd FILL
XFILL_0__7752_ gnd vdd FILL
XFILL_2__13814_ gnd vdd FILL
XFILL_3__14064_ gnd vdd FILL
XFILL_5__14974_ gnd vdd FILL
XFILL_3__7461_ gnd vdd FILL
XFILL_0__10116_ gnd vdd FILL
XFILL_1__15243_ gnd vdd FILL
XFILL_3__11276_ gnd vdd FILL
XFILL_2__14794_ gnd vdd FILL
XFILL_1__12455_ gnd vdd FILL
X_8030_ _8030_/Q _8926_/CLK _7262_/R vdd _7952_/Y gnd vdd DFFSR
XFILL_5__8377_ gnd vdd FILL
XFILL_0__15973_ gnd vdd FILL
XFILL_0__11096_ gnd vdd FILL
XFILL_6__14175_ gnd vdd FILL
XFILL_3__13015_ gnd vdd FILL
X_16079_ _16079_/A _15581_/C _15544_/A _16079_/D gnd _16079_/Y vdd OAI22X1
XFILL_5__13925_ gnd vdd FILL
XFILL_4__15354_ gnd vdd FILL
XFILL_0__7683_ gnd vdd FILL
XFILL_2__7619_ gnd vdd FILL
XSFILL89080x20050 gnd vdd FILL
XFILL_2__13745_ gnd vdd FILL
XFILL_1__11406_ gnd vdd FILL
XFILL_2__10957_ gnd vdd FILL
XFILL_1__15174_ gnd vdd FILL
XFILL_0__10047_ gnd vdd FILL
XFILL_1__12386_ gnd vdd FILL
XFILL_5__7328_ gnd vdd FILL
XFILL_2__8599_ gnd vdd FILL
XFILL_0__14924_ gnd vdd FILL
XFILL_0__9422_ gnd vdd FILL
XSFILL89320x82050 gnd vdd FILL
XSFILL53960x59050 gnd vdd FILL
XFILL_4__14305_ gnd vdd FILL
XFILL_4__11517_ gnd vdd FILL
XFILL_5__13856_ gnd vdd FILL
XFILL_4__15285_ gnd vdd FILL
XSFILL3560x23050 gnd vdd FILL
XFILL_3__9131_ gnd vdd FILL
XFILL_1__14125_ gnd vdd FILL
XFILL_4__12497_ gnd vdd FILL
XFILL_3__10158_ gnd vdd FILL
XFILL_1__11337_ gnd vdd FILL
XFILL_2__13676_ gnd vdd FILL
XFILL_0__14855_ gnd vdd FILL
XFILL_2__10888_ gnd vdd FILL
XFILL_0__9353_ gnd vdd FILL
XFILL_4__14236_ gnd vdd FILL
XSFILL28760x35050 gnd vdd FILL
XFILL_6__10269_ gnd vdd FILL
XFILL_4__11448_ gnd vdd FILL
XFILL_2__15415_ gnd vdd FILL
XFILL_2__12627_ gnd vdd FILL
XFILL_5__13787_ gnd vdd FILL
X_9981_ _9979_/B _9981_/B gnd _9982_/C vdd NAND2X1
XFILL_2__16395_ gnd vdd FILL
XSFILL54040x68050 gnd vdd FILL
XFILL_0__13806_ gnd vdd FILL
XFILL_1__14056_ gnd vdd FILL
XFILL_3__14966_ gnd vdd FILL
XFILL_1__11268_ gnd vdd FILL
XFILL_5__10999_ gnd vdd FILL
XFILL_0__11998_ gnd vdd FILL
XFILL_5__15526_ gnd vdd FILL
XFILL_0__14786_ gnd vdd FILL
XFILL_3__8013_ gnd vdd FILL
XSFILL94440x73050 gnd vdd FILL
XFILL_5__12738_ gnd vdd FILL
X_8932_ _8864_/A _8541_/CLK _7258_/R vdd _8932_/D gnd vdd DFFSR
XFILL_4__14167_ gnd vdd FILL
XFILL_0__9284_ gnd vdd FILL
XFILL_2__15346_ gnd vdd FILL
XFILL_1__13007_ gnd vdd FILL
XFILL_3__13917_ gnd vdd FILL
XFILL_4__11379_ gnd vdd FILL
XFILL_3__14897_ gnd vdd FILL
XFILL_0__10949_ gnd vdd FILL
XFILL_0__13737_ gnd vdd FILL
XFILL_1__11199_ gnd vdd FILL
XFILL_4__13118_ gnd vdd FILL
XFILL_0__8235_ gnd vdd FILL
XFILL_5__15457_ gnd vdd FILL
X_8863_ _8863_/A _8854_/B _8862_/Y gnd _8931_/D vdd OAI21X1
XFILL_2__11509_ gnd vdd FILL
XFILL_4__14098_ gnd vdd FILL
XSFILL33880x26050 gnd vdd FILL
XFILL_3__13848_ gnd vdd FILL
XFILL_2__15277_ gnd vdd FILL
XFILL_2__12489_ gnd vdd FILL
XFILL_0__13668_ gnd vdd FILL
XFILL_5__14408_ gnd vdd FILL
X_7814_ _7814_/A _6918_/B gnd _7815_/C vdd NAND2X1
XFILL_5__15388_ gnd vdd FILL
XFILL_2__14228_ gnd vdd FILL
XFILL_0__15407_ gnd vdd FILL
X_8794_ _8706_/A _9707_/CLK _8801_/R vdd _8794_/D gnd vdd DFFSR
XFILL_3__13779_ gnd vdd FILL
XSFILL48920x48050 gnd vdd FILL
XFILL_0__12619_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1081 gnd vdd FILL
XFILL_1__14958_ gnd vdd FILL
XFILL_0__7117_ gnd vdd FILL
XFILL_0__13599_ gnd vdd FILL
XFILL_0__16387_ gnd vdd FILL
XFILL_6__9673_ gnd vdd FILL
XFILL_5__14339_ gnd vdd FILL
XFILL_3__15518_ gnd vdd FILL
XFILL_0__8097_ gnd vdd FILL
X_7745_ _7791_/Q gnd _7747_/A vdd INVX1
XFILL_2__14159_ gnd vdd FILL
XFILL_1__13909_ gnd vdd FILL
XFILL_3__8915_ gnd vdd FILL
XFILL_3__9895_ gnd vdd FILL
XFILL_0__15338_ gnd vdd FILL
XFILL_6__8624_ gnd vdd FILL
XFILL_1__14889_ gnd vdd FILL
XSFILL49000x57050 gnd vdd FILL
XFILL_0__7048_ gnd vdd FILL
XFILL_1__7930_ gnd vdd FILL
XFILL_3__8846_ gnd vdd FILL
X_7676_ _7768_/Q gnd _7676_/Y vdd INVX1
XFILL_3__15449_ gnd vdd FILL
XSFILL89400x62050 gnd vdd FILL
XFILL_5__16009_ gnd vdd FILL
XFILL_0__15269_ gnd vdd FILL
X_9415_ _9457_/Q gnd _9417_/A vdd INVX1
XFILL_1__7861_ gnd vdd FILL
XFILL_4__7570_ gnd vdd FILL
XFILL_3__8777_ gnd vdd FILL
XFILL_1__9600_ gnd vdd FILL
XSFILL28840x15050 gnd vdd FILL
X_9346_ _9434_/Q gnd _9348_/A vdd INVX1
XFILL_0__8999_ gnd vdd FILL
XFILL_4_BUFX2_insert303 gnd vdd FILL
XSFILL109160x70050 gnd vdd FILL
XFILL_3__7728_ gnd vdd FILL
XFILL_4_BUFX2_insert314 gnd vdd FILL
XFILL_4_BUFX2_insert325 gnd vdd FILL
XFILL_1__9531_ gnd vdd FILL
XFILL_4_BUFX2_insert336 gnd vdd FILL
X_9277_ _9277_/A _9277_/B _9277_/C gnd _9325_/D vdd OAI21X1
XFILL_4__9240_ gnd vdd FILL
XFILL_4_BUFX2_insert347 gnd vdd FILL
XFILL_4_BUFX2_insert358 gnd vdd FILL
XFILL_4_BUFX2_insert369 gnd vdd FILL
XFILL_6__7368_ gnd vdd FILL
X_8228_ _8208_/B _8228_/B gnd _8229_/C vdd NAND2X1
XFILL_1__9462_ gnd vdd FILL
XSFILL83560x77050 gnd vdd FILL
XFILL_4__9171_ gnd vdd FILL
X_10090_ _14442_/A _8815_/CLK _8047_/R vdd _10090_/D gnd vdd DFFSR
XSFILL18760x67050 gnd vdd FILL
XSFILL8600x77050 gnd vdd FILL
XFILL_4__8122_ gnd vdd FILL
XFILL_1__9393_ gnd vdd FILL
X_8159_ _8159_/Q _8815_/CLK _8047_/R vdd _8159_/D gnd vdd DFFSR
XFILL_6__9038_ gnd vdd FILL
XSFILL39000x7050 gnd vdd FILL
XSFILL33800x70050 gnd vdd FILL
XFILL_1__8344_ gnd vdd FILL
XSFILL23880x58050 gnd vdd FILL
XFILL_1__8275_ gnd vdd FILL
X_12800_ _12800_/Q _8171_/CLK _8171_/R vdd _12724_/Y gnd vdd DFFSR
X_13780_ _9608_/A gnd _13780_/Y vdd INVX1
XFILL_1__7226_ gnd vdd FILL
X_10992_ _10991_/Y gnd _11220_/A vdd INVX2
X_12731_ _11876_/B gnd _12731_/Y vdd INVX1
XSFILL54200x28050 gnd vdd FILL
XFILL_1_BUFX2_insert226 gnd vdd FILL
XFILL_1_BUFX2_insert237 gnd vdd FILL
XFILL_1_BUFX2_insert248 gnd vdd FILL
XFILL_1_BUFX2_insert259 gnd vdd FILL
XSFILL79160x32050 gnd vdd FILL
XFILL_4__8955_ gnd vdd FILL
X_15450_ _8671_/Q gnd _15452_/C vdd INVX1
X_12662_ _12660_/Y vdd _12661_/Y gnd _12694_/D vdd OAI21X1
XFILL_2__7970_ gnd vdd FILL
XFILL_1__7088_ gnd vdd FILL
X_14401_ _14390_/Y _14401_/B gnd _14402_/B vdd NOR2X1
XFILL_0_BUFX2_insert904 gnd vdd FILL
XFILL_4__8886_ gnd vdd FILL
X_11613_ _11613_/A gnd _12494_/B vdd INVX1
X_15381_ _15381_/A _15381_/B _15381_/C gnd _15381_/Y vdd NAND3X1
XFILL_0_BUFX2_insert915 gnd vdd FILL
X_12593_ _12591_/Y vdd _12593_/C gnd _12671_/D vdd OAI21X1
XFILL_2__6921_ gnd vdd FILL
XSFILL114360x41050 gnd vdd FILL
XFILL_0_BUFX2_insert926 gnd vdd FILL
XFILL_0_BUFX2_insert937 gnd vdd FILL
XFILL_0_BUFX2_insert948 gnd vdd FILL
XFILL_4__7837_ gnd vdd FILL
XSFILL18840x47050 gnd vdd FILL
X_14332_ _14323_/Y _14324_/Y _14331_/Y gnd _14332_/Y vdd NAND3X1
XFILL_0_BUFX2_insert959 gnd vdd FILL
X_11544_ _11544_/A _11509_/B _11495_/C _11290_/A gnd _11544_/Y vdd AOI22X1
XFILL_2__9640_ gnd vdd FILL
XFILL_2__6852_ gnd vdd FILL
XFILL_5__10020_ gnd vdd FILL
X_14263_ _14263_/A _14263_/B _14260_/Y gnd _14264_/B vdd NAND3X1
X_11475_ _11454_/A _11318_/C _11475_/C gnd _11486_/C vdd OAI21X1
XSFILL28680x6050 gnd vdd FILL
XFILL_4__10750_ gnd vdd FILL
XFILL_4__9507_ gnd vdd FILL
X_16002_ _16002_/A _14551_/Y _16002_/C _16002_/D gnd _16003_/B vdd OAI22X1
XFILL_1__10570_ gnd vdd FILL
XFILL_5__9280_ gnd vdd FILL
X_13214_ _13246_/A gnd _13215_/B vdd INVX1
X_10426_ _10426_/A _10426_/B _10425_/Y gnd _10476_/D vdd OAI21X1
XFILL_4__7699_ gnd vdd FILL
XFILL_1__9729_ gnd vdd FILL
X_14194_ _14194_/A _14193_/Y _14194_/C gnd _14194_/Y vdd NAND3X1
XFILL_2__8522_ gnd vdd FILL
XFILL_6__12290_ gnd vdd FILL
XFILL_3__11130_ gnd vdd FILL
XFILL_4__10681_ gnd vdd FILL
XSFILL109720x28050 gnd vdd FILL
XFILL_5__8231_ gnd vdd FILL
XFILL_2__11860_ gnd vdd FILL
XFILL_6_CLKBUF1_insert203 gnd vdd FILL
X_13145_ _13145_/A gnd _13145_/Y vdd INVX1
XFILL_4__12420_ gnd vdd FILL
XFILL_6__11241_ gnd vdd FILL
XFILL_6_CLKBUF1_insert214 gnd vdd FILL
XFILL_4_BUFX2_insert870 gnd vdd FILL
X_10357_ _14956_/B _9205_/CLK _8433_/R vdd _10357_/D gnd vdd DFFSR
XFILL_2__10811_ gnd vdd FILL
XFILL_5__11971_ gnd vdd FILL
XFILL_1__12240_ gnd vdd FILL
XFILL_3__11061_ gnd vdd FILL
XFILL_2__8453_ gnd vdd FILL
XFILL_4_BUFX2_insert881 gnd vdd FILL
XFILL_4_BUFX2_insert892 gnd vdd FILL
XFILL_4__9369_ gnd vdd FILL
XFILL_2__11791_ gnd vdd FILL
XFILL_0__12970_ gnd vdd FILL
XFILL_5__13710_ gnd vdd FILL
XFILL_5__10922_ gnd vdd FILL
XFILL_4__12351_ gnd vdd FILL
XFILL_3__10012_ gnd vdd FILL
X_13076_ _6899_/A _7532_/CLK _8816_/R vdd _13076_/D gnd vdd DFFSR
X_10288_ _10264_/A _7856_/B gnd _10289_/C vdd NAND2X1
XFILL_5__14690_ gnd vdd FILL
XFILL_2__13530_ gnd vdd FILL
XFILL_2__8384_ gnd vdd FILL
XFILL_2__10742_ gnd vdd FILL
XFILL_1__12171_ gnd vdd FILL
XFILL_5__7113_ gnd vdd FILL
XSFILL79240x12050 gnd vdd FILL
XFILL_0__11921_ gnd vdd FILL
XSFILL3480x38050 gnd vdd FILL
X_12027_ _12031_/A _12027_/B _12031_/C gnd _12027_/Y vdd NAND3X1
XFILL_4__11302_ gnd vdd FILL
XFILL_5__8093_ gnd vdd FILL
XFILL_5__13641_ gnd vdd FILL
XFILL_4__15070_ gnd vdd FILL
XFILL_2__7335_ gnd vdd FILL
XFILL_3__14820_ gnd vdd FILL
XFILL_4__12282_ gnd vdd FILL
XFILL_1__11122_ gnd vdd FILL
XFILL_2__13461_ gnd vdd FILL
XFILL_0__14640_ gnd vdd FILL
XFILL_5__7044_ gnd vdd FILL
XFILL_2__10673_ gnd vdd FILL
XFILL_0__11852_ gnd vdd FILL
XFILL_4__14021_ gnd vdd FILL
XFILL_2__15200_ gnd vdd FILL
XFILL_5__16360_ gnd vdd FILL
XFILL_4__11233_ gnd vdd FILL
XFILL_2__12412_ gnd vdd FILL
XFILL_5__10784_ gnd vdd FILL
XFILL_3__14751_ gnd vdd FILL
XFILL_5__13572_ gnd vdd FILL
XFILL_2__16180_ gnd vdd FILL
XFILL_1__15930_ gnd vdd FILL
XFILL_3__11963_ gnd vdd FILL
XFILL_1__11053_ gnd vdd FILL
XFILL_0__10803_ gnd vdd FILL
XFILL_2__13392_ gnd vdd FILL
XFILL_0__14571_ gnd vdd FILL
XFILL_5__15311_ gnd vdd FILL
XFILL_0__11783_ gnd vdd FILL
XFILL_5__12523_ gnd vdd FILL
XFILL_2__9005_ gnd vdd FILL
XFILL_3__10914_ gnd vdd FILL
X_13978_ _15498_/D _13978_/B gnd _13978_/Y vdd NOR2X1
XFILL_5__16291_ gnd vdd FILL
XFILL_4__11164_ gnd vdd FILL
XFILL_3__13702_ gnd vdd FILL
XFILL_1__10004_ gnd vdd FILL
XFILL_2__15131_ gnd vdd FILL
XFILL_2__12343_ gnd vdd FILL
XFILL_0__16310_ gnd vdd FILL
XFILL_3__14682_ gnd vdd FILL
XFILL_3__11894_ gnd vdd FILL
XFILL_2__7197_ gnd vdd FILL
XFILL_0__13522_ gnd vdd FILL
XFILL_1__15861_ gnd vdd FILL
XSFILL69160x64050 gnd vdd FILL
XFILL_0__8020_ gnd vdd FILL
XFILL_4__10115_ gnd vdd FILL
X_15717_ _15717_/A _15197_/B gnd _15719_/C vdd NOR2X1
XFILL_5__15242_ gnd vdd FILL
X_12929_ _12929_/Q _9823_/CLK _9823_/R vdd _12855_/Y gnd vdd DFFSR
XFILL_5__8995_ gnd vdd FILL
XFILL_3__13633_ gnd vdd FILL
XFILL_5__12454_ gnd vdd FILL
XFILL_4__15972_ gnd vdd FILL
XFILL_1__14812_ gnd vdd FILL
XFILL_2__15062_ gnd vdd FILL
XFILL_4__11095_ gnd vdd FILL
XFILL_0__16241_ gnd vdd FILL
XFILL_0__13453_ gnd vdd FILL
XFILL_2__12274_ gnd vdd FILL
XFILL_1__15792_ gnd vdd FILL
XFILL_0__10665_ gnd vdd FILL
XFILL_5__7946_ gnd vdd FILL
XFILL_5__11405_ gnd vdd FILL
XFILL_6__10956_ gnd vdd FILL
XSFILL104360x73050 gnd vdd FILL
XFILL_4__10046_ gnd vdd FILL
X_15648_ _15646_/Y _15648_/B gnd _15649_/B vdd NOR2X1
XFILL_1_BUFX2_insert760 gnd vdd FILL
XFILL_5__15173_ gnd vdd FILL
XFILL_2__14013_ gnd vdd FILL
XFILL_3__16352_ gnd vdd FILL
XFILL_4__14923_ gnd vdd FILL
XFILL_5__12385_ gnd vdd FILL
XFILL_1_BUFX2_insert771 gnd vdd FILL
XFILL_3__13564_ gnd vdd FILL
XFILL_2__11225_ gnd vdd FILL
XFILL_0__12404_ gnd vdd FILL
XFILL_3__10776_ gnd vdd FILL
XFILL_3__6961_ gnd vdd FILL
XFILL_1__14743_ gnd vdd FILL
XFILL_0__16172_ gnd vdd FILL
XFILL_1__11955_ gnd vdd FILL
XFILL_0__13384_ gnd vdd FILL
XFILL_1_BUFX2_insert782 gnd vdd FILL
XSFILL89720x5050 gnd vdd FILL
XFILL_5__14124_ gnd vdd FILL
XSFILL74280x55050 gnd vdd FILL
XFILL_5__7877_ gnd vdd FILL
XFILL_1_BUFX2_insert793 gnd vdd FILL
XFILL_3__15303_ gnd vdd FILL
XFILL_3__12515_ gnd vdd FILL
XFILL_3__8700_ gnd vdd FILL
X_7530_ _7530_/Q _7530_/CLK _7523_/R vdd _7530_/D gnd vdd DFFSR
X_15579_ _15579_/A _15579_/B gnd _15579_/Y vdd NOR2X1
XFILL_5__11336_ gnd vdd FILL
XFILL_4__14854_ gnd vdd FILL
XFILL_2__9907_ gnd vdd FILL
XSFILL109400x10050 gnd vdd FILL
XFILL_3__16283_ gnd vdd FILL
XFILL_1__10906_ gnd vdd FILL
XFILL_0__12335_ gnd vdd FILL
XFILL_2__11156_ gnd vdd FILL
XFILL_0__15123_ gnd vdd FILL
XFILL_3__13495_ gnd vdd FILL
XFILL_3__9680_ gnd vdd FILL
XFILL_5__9616_ gnd vdd FILL
XFILL_3__6892_ gnd vdd FILL
XFILL_1__14674_ gnd vdd FILL
XFILL_1__11886_ gnd vdd FILL
XFILL_4_BUFX2_insert20 gnd vdd FILL
XFILL_4__13805_ gnd vdd FILL
X_7461_ _7461_/A _7460_/A _7461_/C gnd _7525_/D vdd OAI21X1
XFILL_3__15234_ gnd vdd FILL
XFILL_5__14055_ gnd vdd FILL
XFILL_4_BUFX2_insert31 gnd vdd FILL
XSFILL49080x31050 gnd vdd FILL
XFILL_5__11267_ gnd vdd FILL
XFILL_3__8631_ gnd vdd FILL
XFILL_3__12446_ gnd vdd FILL
XFILL_4_BUFX2_insert42 gnd vdd FILL
XFILL_2__10107_ gnd vdd FILL
XFILL_1__16413_ gnd vdd FILL
XSFILL3560x18050 gnd vdd FILL
XFILL_1__13625_ gnd vdd FILL
XFILL_4_BUFX2_insert53 gnd vdd FILL
XFILL_2__15964_ gnd vdd FILL
XFILL_4__14785_ gnd vdd FILL
XFILL_4__11997_ gnd vdd FILL
XFILL_0__15054_ gnd vdd FILL
XFILL_0__12266_ gnd vdd FILL
XFILL_6__8340_ gnd vdd FILL
XFILL_2__11087_ gnd vdd FILL
XFILL_1__10837_ gnd vdd FILL
XFILL_5__9547_ gnd vdd FILL
X_9200_ _9200_/Q _8289_/CLK _7649_/R vdd _9200_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert64 gnd vdd FILL
XFILL_5__13006_ gnd vdd FILL
XFILL_4_BUFX2_insert75 gnd vdd FILL
XFILL_0__8853_ gnd vdd FILL
XFILL_4_BUFX2_insert86 gnd vdd FILL
XFILL_3__15165_ gnd vdd FILL
XFILL_4__13736_ gnd vdd FILL
X_7392_ _7316_/A _9716_/CLK _8682_/R vdd _7392_/D gnd vdd DFFSR
XFILL_5__11198_ gnd vdd FILL
XFILL_4__10948_ gnd vdd FILL
XFILL_2__10038_ gnd vdd FILL
XFILL_1__16344_ gnd vdd FILL
XFILL_3__12377_ gnd vdd FILL
XFILL_0__14005_ gnd vdd FILL
XFILL_2__14915_ gnd vdd FILL
XFILL_0__11217_ gnd vdd FILL
XFILL_2__9769_ gnd vdd FILL
XFILL_4_BUFX2_insert97 gnd vdd FILL
XFILL_2__15895_ gnd vdd FILL
XFILL_1__13556_ gnd vdd FILL
XFILL_1__10768_ gnd vdd FILL
XFILL_0__12197_ gnd vdd FILL
XFILL_0__7804_ gnd vdd FILL
XFILL_5__10149_ gnd vdd FILL
XFILL_5__9478_ gnd vdd FILL
XFILL_3__14116_ gnd vdd FILL
X_9131_ _9129_/Y _9116_/B _9130_/Y gnd _9131_/Y vdd OAI21X1
XSFILL94440x68050 gnd vdd FILL
XFILL_0__8784_ gnd vdd FILL
XFILL_3__11328_ gnd vdd FILL
XFILL_2__14846_ gnd vdd FILL
XFILL_4__13667_ gnd vdd FILL
XFILL_1__12507_ gnd vdd FILL
XFILL_4__10879_ gnd vdd FILL
XSFILL49000x2050 gnd vdd FILL
XFILL_3__15096_ gnd vdd FILL
XFILL_3__8493_ gnd vdd FILL
XFILL_0__11148_ gnd vdd FILL
XFILL_1__16275_ gnd vdd FILL
XFILL_6__14227_ gnd vdd FILL
XFILL_1__13487_ gnd vdd FILL
X_9062_ _9062_/Q _7021_/CLK _9062_/R vdd _9062_/D gnd vdd DFFSR
XFILL_0__7735_ gnd vdd FILL
XFILL_4__15406_ gnd vdd FILL
XFILL_1__10699_ gnd vdd FILL
XFILL_4__12618_ gnd vdd FILL
XFILL_3__14047_ gnd vdd FILL
XFILL_5__14957_ gnd vdd FILL
XFILL_2_BUFX2_insert1003 gnd vdd FILL
XFILL_4__16386_ gnd vdd FILL
XFILL_1__15226_ gnd vdd FILL
XFILL_3__11259_ gnd vdd FILL
XFILL_3__7444_ gnd vdd FILL
XFILL_4__13598_ gnd vdd FILL
XFILL_2_BUFX2_insert1014 gnd vdd FILL
XFILL_1__12438_ gnd vdd FILL
XFILL_2__14777_ gnd vdd FILL
XSFILL68200x80050 gnd vdd FILL
XFILL_2_BUFX2_insert1025 gnd vdd FILL
XFILL_2__11989_ gnd vdd FILL
XFILL_0__15956_ gnd vdd FILL
XFILL_0__11079_ gnd vdd FILL
X_8013_ _8013_/A gnd _8015_/A vdd INVX1
XFILL_5__13908_ gnd vdd FILL
XFILL_2_BUFX2_insert1036 gnd vdd FILL
XFILL_4__15337_ gnd vdd FILL
XFILL_2_BUFX2_insert1047 gnd vdd FILL
XFILL_2__13728_ gnd vdd FILL
XFILL_5__14888_ gnd vdd FILL
XFILL_3__7375_ gnd vdd FILL
XFILL_2_BUFX2_insert1058 gnd vdd FILL
XFILL_1__15157_ gnd vdd FILL
XFILL_0__14907_ gnd vdd FILL
XFILL_1__12369_ gnd vdd FILL
XFILL_0__9405_ gnd vdd FILL
XFILL_2_BUFX2_insert1069 gnd vdd FILL
XFILL_6__7084_ gnd vdd FILL
XFILL_0__15887_ gnd vdd FILL
XFILL_5__13839_ gnd vdd FILL
XFILL_3__9114_ gnd vdd FILL
XSFILL8680x51050 gnd vdd FILL
XFILL_0__7597_ gnd vdd FILL
XFILL_1__14108_ gnd vdd FILL
XFILL_4__15268_ gnd vdd FILL
XFILL_2__13659_ gnd vdd FILL
XFILL_3__15998_ gnd vdd FILL
XFILL_0__14838_ gnd vdd FILL
XFILL_1__15088_ gnd vdd FILL
XFILL_0__9336_ gnd vdd FILL
XFILL_4__14219_ gnd vdd FILL
X_9964_ _9964_/Q _7916_/CLK _9964_/R vdd _9964_/D gnd vdd DFFSR
XFILL_3__9045_ gnd vdd FILL
XFILL_4__15199_ gnd vdd FILL
XFILL_1__14039_ gnd vdd FILL
XFILL_3__14949_ gnd vdd FILL
XFILL_2__16378_ gnd vdd FILL
XSFILL89400x57050 gnd vdd FILL
XFILL_5__15509_ gnd vdd FILL
XFILL_0__14769_ gnd vdd FILL
XFILL_0__9267_ gnd vdd FILL
XFILL_1__8060_ gnd vdd FILL
X_8915_ _8915_/A gnd _8915_/Y vdd INVX1
XFILL_2__15329_ gnd vdd FILL
X_9895_ _9920_/B _9895_/B gnd _9896_/C vdd NAND2X1
XFILL_0_BUFX2_insert1040 gnd vdd FILL
XFILL_0__8218_ gnd vdd FILL
XFILL_0_BUFX2_insert1051 gnd vdd FILL
X_8846_ _8926_/Q gnd _8846_/Y vdd INVX1
XFILL_0_BUFX2_insert1062 gnd vdd FILL
XFILL_0_BUFX2_insert1073 gnd vdd FILL
XFILL_0_BUFX2_insert1084 gnd vdd FILL
XSFILL13640x52050 gnd vdd FILL
XSFILL14120x59050 gnd vdd FILL
XFILL_0__8149_ gnd vdd FILL
XFILL_4__8740_ gnd vdd FILL
X_8777_ _8775_/Y _8788_/A _8776_/Y gnd _8817_/D vdd OAI21X1
XSFILL38680x1050 gnd vdd FILL
XFILL_6_BUFX2_insert976 gnd vdd FILL
XFILL_1__8962_ gnd vdd FILL
XFILL_6__6868_ gnd vdd FILL
X_7728_ _7729_/B _8624_/B gnd _7728_/Y vdd NAND2X1
XFILL_3__9878_ gnd vdd FILL
X_7659_ _7605_/A _7261_/CLK _8669_/R vdd _7659_/D gnd vdd DFFSR
XFILL_1__8893_ gnd vdd FILL
XSFILL104520x33050 gnd vdd FILL
XFILL_4__7622_ gnd vdd FILL
XFILL_3__8829_ gnd vdd FILL
XSFILL8760x31050 gnd vdd FILL
XFILL_1__7844_ gnd vdd FILL
XSFILL33800x65050 gnd vdd FILL
XFILL_4__7553_ gnd vdd FILL
XFILL_4_BUFX2_insert100 gnd vdd FILL
X_11260_ _11258_/Y _11259_/Y gnd _11448_/A vdd NOR2X1
X_9329_ _9329_/Q _7537_/CLK _7537_/R vdd _9289_/Y gnd vdd DFFSR
XFILL_4__7484_ gnd vdd FILL
X_10211_ _14081_/A _6999_/CLK _7011_/R vdd _10211_/D gnd vdd DFFSR
XFILL_1__9514_ gnd vdd FILL
X_11191_ _11191_/A _11191_/B gnd _11191_/Y vdd NOR2X1
XFILL_4__9223_ gnd vdd FILL
XFILL111960x75050 gnd vdd FILL
XFILL_3_BUFX2_insert800 gnd vdd FILL
XFILL_3_BUFX2_insert811 gnd vdd FILL
X_10142_ _10106_/A _7838_/B gnd _10143_/C vdd NAND2X1
XFILL_3_BUFX2_insert822 gnd vdd FILL
XSFILL38280x15050 gnd vdd FILL
XSFILL13720x32050 gnd vdd FILL
XFILL_3_BUFX2_insert833 gnd vdd FILL
XFILL_4__9154_ gnd vdd FILL
XFILL_3_BUFX2_insert844 gnd vdd FILL
X_10073_ _9983_/A _7282_/CLK _9062_/R vdd _9985_/Y gnd vdd DFFSR
X_14950_ _14946_/Y _14950_/B gnd _14950_/Y vdd NOR2X1
XFILL_3_BUFX2_insert855 gnd vdd FILL
XFILL_3_BUFX2_insert866 gnd vdd FILL
XFILL_1__9376_ gnd vdd FILL
XFILL_3_BUFX2_insert877 gnd vdd FILL
XFILL_4__8105_ gnd vdd FILL
XFILL_3_BUFX2_insert888 gnd vdd FILL
XFILL_4__9085_ gnd vdd FILL
XFILL_3_BUFX2_insert899 gnd vdd FILL
X_13901_ _7903_/Q gnd _13901_/Y vdd INVX1
X_14881_ _14881_/A _14881_/B _14597_/C gnd _13039_/B vdd AOI21X1
XFILL_1__8327_ gnd vdd FILL
XFILL_2__7120_ gnd vdd FILL
X_13832_ _7435_/A gnd _13833_/D vdd INVX1
XSFILL84280x18050 gnd vdd FILL
XFILL_2__7051_ gnd vdd FILL
XFILL_1__8258_ gnd vdd FILL
X_13763_ _13763_/A _14555_/C gnd _13769_/C vdd NOR2X1
XFILL_1__7209_ gnd vdd FILL
X_10975_ _10911_/A gnd _10977_/A vdd INVX1
XSFILL53800x3050 gnd vdd FILL
XFILL_1__8189_ gnd vdd FILL
XFILL_5__7800_ gnd vdd FILL
X_12714_ _12768_/A memoryOutData[6] gnd _12715_/C vdd NAND2X1
XFILL_5__8780_ gnd vdd FILL
X_15502_ _15756_/D gnd _16212_/A vdd INVX4
XFILL_4__9987_ gnd vdd FILL
XFILL_3__10630_ gnd vdd FILL
X_13694_ _15261_/A gnd _13694_/Y vdd INVX1
XFILL_5__7731_ gnd vdd FILL
XFILL_0__10450_ gnd vdd FILL
X_15433_ _15433_/A _15433_/B _15432_/Y gnd _15433_/Y vdd NAND3X1
X_12645_ _12645_/A gnd _12647_/A vdd INVX1
XFILL_5__12170_ gnd vdd FILL
XFILL_0_BUFX2_insert701 gnd vdd FILL
XFILL_0_BUFX2_insert712 gnd vdd FILL
XFILL_4__11920_ gnd vdd FILL
XFILL_2__11010_ gnd vdd FILL
XFILL_0_BUFX2_insert723 gnd vdd FILL
XFILL_2__7953_ gnd vdd FILL
XFILL_3__10561_ gnd vdd FILL
XFILL_1__11740_ gnd vdd FILL
XFILL_0__10381_ gnd vdd FILL
XFILL_0_CLKBUF1_insert160 gnd vdd FILL
XFILL_0_BUFX2_insert734 gnd vdd FILL
XFILL_5__11121_ gnd vdd FILL
XFILL_4__8869_ gnd vdd FILL
X_15364_ _7901_/Q gnd _15364_/Y vdd INVX1
XFILL_0_BUFX2_insert745 gnd vdd FILL
XFILL_3__12300_ gnd vdd FILL
XFILL_0_CLKBUF1_insert171 gnd vdd FILL
X_12576_ _12576_/A gnd _12578_/A vdd INVX1
XFILL_2__6904_ gnd vdd FILL
XFILL_6__10672_ gnd vdd FILL
XFILL_0_BUFX2_insert756 gnd vdd FILL
XFILL_0_CLKBUF1_insert182 gnd vdd FILL
XSFILL13800x12050 gnd vdd FILL
XFILL_3__13280_ gnd vdd FILL
XFILL_0_BUFX2_insert767 gnd vdd FILL
XFILL_0__12120_ gnd vdd FILL
XFILL_4__11851_ gnd vdd FILL
XFILL_0_CLKBUF1_insert193 gnd vdd FILL
XFILL_2__7884_ gnd vdd FILL
XFILL_5__9401_ gnd vdd FILL
XFILL_3__10492_ gnd vdd FILL
XFILL112120x64050 gnd vdd FILL
XFILL_0_BUFX2_insert778 gnd vdd FILL
X_14315_ _9320_/Q gnd _15795_/A vdd INVX1
XFILL_1__11671_ gnd vdd FILL
XFILL_0_BUFX2_insert789 gnd vdd FILL
XFILL_5__7593_ gnd vdd FILL
X_11527_ _11527_/A _11527_/B _11527_/C gnd _11527_/Y vdd OAI21X1
XFILL_5__11052_ gnd vdd FILL
XFILL_2__9623_ gnd vdd FILL
XFILL_3__12231_ gnd vdd FILL
X_15295_ _15295_/A _15276_/Y _15294_/Y gnd _15296_/B vdd NOR3X1
XFILL_4__10802_ gnd vdd FILL
XFILL_4__14570_ gnd vdd FILL
XFILL_1__13410_ gnd vdd FILL
XFILL_4__11782_ gnd vdd FILL
XFILL_2__12961_ gnd vdd FILL
XFILL_0__12051_ gnd vdd FILL
XFILL_1__10622_ gnd vdd FILL
XFILL_1__14390_ gnd vdd FILL
XFILL_5__10003_ gnd vdd FILL
X_14246_ _14555_/B _14244_/Y _13857_/C _14246_/D gnd _14250_/B vdd OAI22X1
XSFILL114440x16050 gnd vdd FILL
XFILL_2__14700_ gnd vdd FILL
X_11458_ _11194_/Y gnd _11461_/B vdd INVX1
XFILL_4__13521_ gnd vdd FILL
XFILL_5__15860_ gnd vdd FILL
XFILL_2__11912_ gnd vdd FILL
XFILL_3__12162_ gnd vdd FILL
XFILL_0__11002_ gnd vdd FILL
XFILL_2__9554_ gnd vdd FILL
XFILL_1__13341_ gnd vdd FILL
XFILL_2__15680_ gnd vdd FILL
XSFILL114440x9050 gnd vdd FILL
XFILL_2__12892_ gnd vdd FILL
XFILL_1__10553_ gnd vdd FILL
XFILL_5__9263_ gnd vdd FILL
XFILL_5__14811_ gnd vdd FILL
X_10409_ _10409_/A gnd _10409_/Y vdd INVX1
X_14177_ _8995_/A gnd _14177_/Y vdd INVX1
XFILL_4__16240_ gnd vdd FILL
XFILL_2__8505_ gnd vdd FILL
XFILL_3__11113_ gnd vdd FILL
XFILL_2__14631_ gnd vdd FILL
XFILL_4__10664_ gnd vdd FILL
XFILL_4__13452_ gnd vdd FILL
XFILL_5__15791_ gnd vdd FILL
X_11389_ _11389_/A _11389_/B gnd _11390_/C vdd NAND2X1
XFILL_2__9485_ gnd vdd FILL
XFILL_3__12093_ gnd vdd FILL
XFILL_0__15810_ gnd vdd FILL
XFILL_5__8214_ gnd vdd FILL
XFILL_1__16060_ gnd vdd FILL
XFILL_2__11843_ gnd vdd FILL
XFILL_1__13272_ gnd vdd FILL
XFILL_6__14012_ gnd vdd FILL
X_13128_ _13099_/B _12054_/Y gnd _13128_/Y vdd NAND2X1
XFILL_4__12403_ gnd vdd FILL
XFILL_5__14742_ gnd vdd FILL
XFILL_3__15921_ gnd vdd FILL
XFILL_4__16171_ gnd vdd FILL
XFILL_5__11954_ gnd vdd FILL
XFILL_4__13383_ gnd vdd FILL
XFILL_1__15011_ gnd vdd FILL
XFILL_3__11044_ gnd vdd FILL
XFILL_2__14562_ gnd vdd FILL
XFILL_1__12223_ gnd vdd FILL
XFILL_2__11774_ gnd vdd FILL
XFILL_0__15741_ gnd vdd FILL
XFILL_5__8145_ gnd vdd FILL
XSFILL84200x62050 gnd vdd FILL
XFILL_0__12953_ gnd vdd FILL
XFILL_5__10905_ gnd vdd FILL
XFILL_0__7451_ gnd vdd FILL
X_13059_ _6882_/A _8176_/CLK _8176_/R vdd _13059_/D gnd vdd DFFSR
XFILL_2__16301_ gnd vdd FILL
XFILL_4__12334_ gnd vdd FILL
XFILL_4__15122_ gnd vdd FILL
XFILL_5__14673_ gnd vdd FILL
XFILL_2__13513_ gnd vdd FILL
XSFILL104360x68050 gnd vdd FILL
XFILL_5__11885_ gnd vdd FILL
XFILL_3__7160_ gnd vdd FILL
XFILL_3__15852_ gnd vdd FILL
XFILL_2__8367_ gnd vdd FILL
XFILL_2__14493_ gnd vdd FILL
XFILL_0__11904_ gnd vdd FILL
XFILL_1__12154_ gnd vdd FILL
XFILL_0__15672_ gnd vdd FILL
XFILL_5__8076_ gnd vdd FILL
XFILL_5__16412_ gnd vdd FILL
XFILL_5__13624_ gnd vdd FILL
XFILL_0__12884_ gnd vdd FILL
XFILL_2__16232_ gnd vdd FILL
XFILL_3__14803_ gnd vdd FILL
XFILL_4__15053_ gnd vdd FILL
XFILL_4__12265_ gnd vdd FILL
XFILL_2__7318_ gnd vdd FILL
XFILL_5__10836_ gnd vdd FILL
XFILL_2__13444_ gnd vdd FILL
XFILL_1__11105_ gnd vdd FILL
XFILL_0__14623_ gnd vdd FILL
XFILL_1__12085_ gnd vdd FILL
XFILL_2__10656_ gnd vdd FILL
XFILL_3__12995_ gnd vdd FILL
XFILL_3__15783_ gnd vdd FILL
XFILL_3__7091_ gnd vdd FILL
XFILL_0__9121_ gnd vdd FILL
XFILL_0__11835_ gnd vdd FILL
XFILL_5__16343_ gnd vdd FILL
XFILL_4__14004_ gnd vdd FILL
XFILL_4__11216_ gnd vdd FILL
XFILL_6__15894_ gnd vdd FILL
XFILL_5__13555_ gnd vdd FILL
XSFILL49080x26050 gnd vdd FILL
XFILL_5__10767_ gnd vdd FILL
XSFILL74680x71050 gnd vdd FILL
XFILL_1__15913_ gnd vdd FILL
XFILL_3__11946_ gnd vdd FILL
XFILL112200x44050 gnd vdd FILL
X_6961_ _6959_/Y _6937_/B _6961_/C gnd _7017_/D vdd OAI21X1
XFILL_3__14734_ gnd vdd FILL
XFILL_4__12196_ gnd vdd FILL
XFILL_1__11036_ gnd vdd FILL
XFILL_2__7249_ gnd vdd FILL
XFILL_2__16163_ gnd vdd FILL
XFILL_2__13375_ gnd vdd FILL
XSFILL24520x43050 gnd vdd FILL
XSFILL48840x81050 gnd vdd FILL
XFILL_0__14554_ gnd vdd FILL
XFILL_5__12506_ gnd vdd FILL
X_8700_ _8700_/A gnd _8702_/A vdd INVX1
XFILL_0__11766_ gnd vdd FILL
XFILL_4__11147_ gnd vdd FILL
XFILL_2__15114_ gnd vdd FILL
XFILL_5__16274_ gnd vdd FILL
XFILL_5__13486_ gnd vdd FILL
X_9680_ _9680_/A gnd _9680_/Y vdd INVX1
XFILL_2__12326_ gnd vdd FILL
XFILL_3__11877_ gnd vdd FILL
XFILL_5__10698_ gnd vdd FILL
XFILL_2__16094_ gnd vdd FILL
X_6892_ _6892_/A gnd memoryWriteData[22] vdd BUFX2
XFILL_1__15844_ gnd vdd FILL
XFILL_3__14665_ gnd vdd FILL
XFILL_0__13505_ gnd vdd FILL
XFILL_0__8003_ gnd vdd FILL
XFILL_0__14485_ gnd vdd FILL
XFILL_5__15225_ gnd vdd FILL
XFILL_0__11697_ gnd vdd FILL
XFILL_5__12437_ gnd vdd FILL
X_8631_ _8631_/A _8589_/B _8630_/Y gnd _8631_/Y vdd OAI21X1
XFILL_3__16404_ gnd vdd FILL
XFILL_5__8978_ gnd vdd FILL
XFILL_3__13616_ gnd vdd FILL
XFILL_3__10828_ gnd vdd FILL
XFILL_2__15045_ gnd vdd FILL
XFILL_6__11988_ gnd vdd FILL
XFILL_4__15955_ gnd vdd FILL
XFILL_6_BUFX2_insert239 gnd vdd FILL
XFILL_4__11078_ gnd vdd FILL
XFILL_3__9801_ gnd vdd FILL
XFILL_3__14596_ gnd vdd FILL
XFILL_0__16224_ gnd vdd FILL
XFILL_2__12257_ gnd vdd FILL
XFILL_0__10648_ gnd vdd FILL
XFILL_3__7993_ gnd vdd FILL
XFILL_1__15775_ gnd vdd FILL
XFILL_0__13436_ gnd vdd FILL
XFILL_1__12987_ gnd vdd FILL
XFILL_5__7929_ gnd vdd FILL
XFILL_1_BUFX2_insert590 gnd vdd FILL
XFILL_4__10029_ gnd vdd FILL
XFILL_5__15156_ gnd vdd FILL
XFILL_4__14906_ gnd vdd FILL
XFILL_5__12368_ gnd vdd FILL
XFILL_3__16335_ gnd vdd FILL
X_8562_ _8522_/A _8562_/CLK _7270_/R vdd _8524_/Y gnd vdd DFFSR
XFILL_3__13547_ gnd vdd FILL
XFILL_2__11208_ gnd vdd FILL
XFILL_3__9732_ gnd vdd FILL
XFILL_3__6944_ gnd vdd FILL
XFILL_1__14726_ gnd vdd FILL
XFILL_3__10759_ gnd vdd FILL
XFILL_4__15886_ gnd vdd FILL
XFILL_5_BUFX2_insert906 gnd vdd FILL
XFILL_2__12188_ gnd vdd FILL
XFILL_1__11938_ gnd vdd FILL
XSFILL53960x9050 gnd vdd FILL
XFILL_0__16155_ gnd vdd FILL
XFILL_0__13367_ gnd vdd FILL
XFILL_5_BUFX2_insert917 gnd vdd FILL
XFILL_5__14107_ gnd vdd FILL
XFILL_0__10579_ gnd vdd FILL
X_7513_ _7513_/Q _7129_/CLK _9049_/R vdd _7425_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert928 gnd vdd FILL
XFILL_5__11319_ gnd vdd FILL
XFILL_4__14837_ gnd vdd FILL
XFILL_5_BUFX2_insert939 gnd vdd FILL
XFILL_5__15087_ gnd vdd FILL
XSFILL54040x81050 gnd vdd FILL
XFILL_3__9663_ gnd vdd FILL
XFILL_5__12299_ gnd vdd FILL
X_8493_ _8494_/B _9901_/B gnd _8493_/Y vdd NAND2X1
XFILL_2__11139_ gnd vdd FILL
XFILL_0__15106_ gnd vdd FILL
XFILL_3__13478_ gnd vdd FILL
XFILL_3__16266_ gnd vdd FILL
XFILL_3__6875_ gnd vdd FILL
XFILL_1__14657_ gnd vdd FILL
XFILL_0__12318_ gnd vdd FILL
XFILL_0__13298_ gnd vdd FILL
XFILL_6__12609_ gnd vdd FILL
XSFILL104440x48050 gnd vdd FILL
XFILL_1__11869_ gnd vdd FILL
XFILL_0__16086_ gnd vdd FILL
XFILL_5__14038_ gnd vdd FILL
XFILL_0__8905_ gnd vdd FILL
XFILL_3__12429_ gnd vdd FILL
XFILL_3__15217_ gnd vdd FILL
XFILL_0__9885_ gnd vdd FILL
X_7444_ _7520_/Q gnd _7446_/A vdd INVX1
XFILL_1__13608_ gnd vdd FILL
XFILL_3__8614_ gnd vdd FILL
XFILL_3__16197_ gnd vdd FILL
XSFILL8680x46050 gnd vdd FILL
XFILL_4__14768_ gnd vdd FILL
XFILL_0__15037_ gnd vdd FILL
XFILL_2__15947_ gnd vdd FILL
XFILL_0__12249_ gnd vdd FILL
XFILL_3__9594_ gnd vdd FILL
XFILL_1__14588_ gnd vdd FILL
XFILL_0__8836_ gnd vdd FILL
XFILL_3__15148_ gnd vdd FILL
XFILL_4__13719_ gnd vdd FILL
X_7375_ _7375_/A _7336_/B _7374_/Y gnd _7411_/D vdd OAI21X1
XFILL_1__16327_ gnd vdd FILL
XFILL_4__14699_ gnd vdd FILL
XSFILL59160x3050 gnd vdd FILL
XFILL_1__13539_ gnd vdd FILL
XFILL_2__15878_ gnd vdd FILL
X_9114_ _9186_/Q gnd _9114_/Y vdd INVX1
XFILL_0__8767_ gnd vdd FILL
XFILL_1__7560_ gnd vdd FILL
XFILL_5__15989_ gnd vdd FILL
XSFILL48920x61050 gnd vdd FILL
XFILL_3__15079_ gnd vdd FILL
XFILL_2__14829_ gnd vdd FILL
XFILL_3__8476_ gnd vdd FILL
XFILL_1__16258_ gnd vdd FILL
XFILL_3_BUFX2_insert107 gnd vdd FILL
XFILL_0__7718_ gnd vdd FILL
X_9045_ _9043_/Y _9044_/A _9045_/C gnd _9077_/D vdd OAI21X1
XFILL_3__7427_ gnd vdd FILL
XFILL_4__16369_ gnd vdd FILL
XFILL_1__15209_ gnd vdd FILL
XFILL_1__7491_ gnd vdd FILL
XFILL_0__8698_ gnd vdd FILL
XFILL_1__16189_ gnd vdd FILL
XFILL_0__15939_ gnd vdd FILL
XFILL_1__9230_ gnd vdd FILL
XSFILL13640x47050 gnd vdd FILL
XCLKBUF1_insert1074 clk gnd CLKBUF1_insert206/A vdd CLKBUF1
XFILL_3__7358_ gnd vdd FILL
XFILL_2_BUFX2_insert807 gnd vdd FILL
XFILL_2_BUFX2_insert818 gnd vdd FILL
XFILL_1__9161_ gnd vdd FILL
XFILL_2_BUFX2_insert829 gnd vdd FILL
XFILL_3__7289_ gnd vdd FILL
XFILL_0_BUFX2_insert40 gnd vdd FILL
XFILL_1__8112_ gnd vdd FILL
XFILL_0_BUFX2_insert51 gnd vdd FILL
XSFILL54120x61050 gnd vdd FILL
XFILL_1__9092_ gnd vdd FILL
XFILL_3__9028_ gnd vdd FILL
X_9947_ _9947_/Q _8663_/CLK _8664_/R vdd _9947_/D gnd vdd DFFSR
XFILL_4__9910_ gnd vdd FILL
XFILL_0_BUFX2_insert62 gnd vdd FILL
XSFILL104520x28050 gnd vdd FILL
XFILL_0_BUFX2_insert73 gnd vdd FILL
XFILL_0_BUFX2_insert84 gnd vdd FILL
XFILL_0_BUFX2_insert95 gnd vdd FILL
XSFILL8760x26050 gnd vdd FILL
X_9878_ _9876_/Y _9937_/A _9878_/C gnd _9952_/D vdd OAI21X1
X_10760_ _10844_/Q gnd _10760_/Y vdd INVX1
X_8829_ _8916_/A _8701_/B gnd _8829_/Y vdd NAND2X1
XFILL_4__9772_ gnd vdd FILL
XFILL_6_BUFX2_insert751 gnd vdd FILL
XBUFX2_insert806 _13490_/Y gnd _14185_/B vdd BUFX2
XFILL_4__6984_ gnd vdd FILL
XSFILL18760x80050 gnd vdd FILL
XBUFX2_insert817 _12384_/Y gnd _7838_/B vdd BUFX2
X_10691_ _10691_/A _10676_/B _10690_/Y gnd _10691_/Y vdd OAI21X1
XBUFX2_insert828 _13287_/Y gnd _7460_/A vdd BUFX2
XFILL_1__9994_ gnd vdd FILL
XBUFX2_insert839 _13324_/Y gnd _8655_/B vdd BUFX2
XFILL_4__8723_ gnd vdd FILL
X_12430_ _12430_/A gnd _12430_/Y vdd INVX1
XFILL_4__8654_ gnd vdd FILL
X_12361_ _12361_/A gnd _12361_/Y vdd INVX1
XFILL_1_CLKBUF1_insert200 gnd vdd FILL
XFILL_1_CLKBUF1_insert211 gnd vdd FILL
XFILL_1__8876_ gnd vdd FILL
XSFILL78920x77050 gnd vdd FILL
XFILL_4__7605_ gnd vdd FILL
XSFILL109640x61050 gnd vdd FILL
XFILL_1_CLKBUF1_insert222 gnd vdd FILL
X_14100_ _7907_/Q gnd _14101_/D vdd INVX1
XFILL_4__8585_ gnd vdd FILL
X_11312_ _11311_/Y _11111_/Y _11312_/C gnd _11312_/Y vdd OAI21X1
X_15080_ _15078_/Y _9047_/Q _9175_/Q _15079_/Y gnd _15085_/C vdd AOI22X1
X_12292_ _12216_/B _12297_/D _12300_/C gnd _12292_/Y vdd NAND3X1
XFILL_1__7827_ gnd vdd FILL
X_14031_ _14031_/A _14027_/Y gnd _14036_/C vdd NOR2X1
X_11243_ _11242_/Y gnd _11447_/B vdd INVX1
XSFILL69800x20050 gnd vdd FILL
XFILL_1__7758_ gnd vdd FILL
XFILL_4__7467_ gnd vdd FILL
X_11174_ _11195_/A _11173_/Y _11174_/C gnd _11191_/B vdd OAI21X1
XFILL_2__9270_ gnd vdd FILL
XFILL_1__7689_ gnd vdd FILL
XFILL_4__9206_ gnd vdd FILL
XFILL_3_BUFX2_insert630 gnd vdd FILL
X_10125_ _10123_/Y _10166_/A _10125_/C gnd _10125_/Y vdd OAI21X1
XFILL_3_BUFX2_insert641 gnd vdd FILL
XFILL_3_BUFX2_insert652 gnd vdd FILL
XFILL_1__9428_ gnd vdd FILL
XFILL_2__8221_ gnd vdd FILL
XFILL_4__10380_ gnd vdd FILL
X_15982_ _15982_/A _15980_/Y gnd _15983_/C vdd NOR2X1
XFILL_4__9137_ gnd vdd FILL
XFILL_3_BUFX2_insert663 gnd vdd FILL
XFILL_3_BUFX2_insert674 gnd vdd FILL
XFILL_3_BUFX2_insert685 gnd vdd FILL
XFILL_3_BUFX2_insert696 gnd vdd FILL
X_10056_ _10066_/B _7752_/B gnd _10056_/Y vdd NAND2X1
X_14933_ _8915_/A gnd _14934_/A vdd INVX1
XFILL_2__10510_ gnd vdd FILL
XFILL_1__9359_ gnd vdd FILL
XFILL_5__11670_ gnd vdd FILL
XFILL_2__11490_ gnd vdd FILL
XFILL_2__7103_ gnd vdd FILL
XFILL_6__12960_ gnd vdd FILL
XFILL_4__12050_ gnd vdd FILL
XSFILL63960x35050 gnd vdd FILL
XFILL_3__11800_ gnd vdd FILL
XFILL_5__10621_ gnd vdd FILL
X_14864_ _7539_/Q gnd _14864_/Y vdd INVX1
XFILL_3__12780_ gnd vdd FILL
XFILL_4__8019_ gnd vdd FILL
XFILL_2__10441_ gnd vdd FILL
XFILL_2__8083_ gnd vdd FILL
XFILL_0__11620_ gnd vdd FILL
XFILL_5__8901_ gnd vdd FILL
XFILL112120x59050 gnd vdd FILL
XFILL_6__11911_ gnd vdd FILL
XSFILL23160x32050 gnd vdd FILL
XFILL_4__11001_ gnd vdd FILL
XFILL_5__13340_ gnd vdd FILL
X_13815_ _13815_/A _13815_/B _13814_/Y gnd _13816_/A vdd NAND3X1
XFILL_5__9881_ gnd vdd FILL
X_14795_ _8946_/Q gnd _14795_/Y vdd INVX1
XFILL_5__10552_ gnd vdd FILL
XFILL_2__7034_ gnd vdd FILL
XFILL_3__11731_ gnd vdd FILL
XFILL_1__12910_ gnd vdd FILL
XFILL_2__13160_ gnd vdd FILL
XFILL_2__10372_ gnd vdd FILL
XSFILL64040x44050 gnd vdd FILL
XFILL_0__11551_ gnd vdd FILL
XFILL_5__8832_ gnd vdd FILL
XFILL_1__13890_ gnd vdd FILL
X_13746_ _9992_/A gnd _15299_/B vdd INVX1
XFILL_5__13271_ gnd vdd FILL
X_10958_ _10941_/Y _10957_/Y gnd _10959_/B vdd NOR2X1
XFILL_2__12111_ gnd vdd FILL
XFILL_3__14450_ gnd vdd FILL
XFILL_3__11662_ gnd vdd FILL
XFILL_0__10502_ gnd vdd FILL
XFILL112280x3050 gnd vdd FILL
XFILL_1__12841_ gnd vdd FILL
XFILL_2__13091_ gnd vdd FILL
XFILL_5__15010_ gnd vdd FILL
XFILL_0__11482_ gnd vdd FILL
XFILL_0__14270_ gnd vdd FILL
XFILL_5__8763_ gnd vdd FILL
XFILL_3__13401_ gnd vdd FILL
XFILL_5__12222_ gnd vdd FILL
X_13677_ _13675_/Y _14479_/B _14865_/C _13676_/Y gnd _13681_/B vdd OAI22X1
XFILL_4__15740_ gnd vdd FILL
XFILL_6__11773_ gnd vdd FILL
XFILL_4__12952_ gnd vdd FILL
XFILL_2__12042_ gnd vdd FILL
X_10889_ _10889_/A _10889_/B gnd _10889_/Y vdd NAND2X1
XFILL_3__14381_ gnd vdd FILL
XFILL_0__13221_ gnd vdd FILL
XSFILL3480x51050 gnd vdd FILL
XFILL_1__15560_ gnd vdd FILL
XFILL_0__10433_ gnd vdd FILL
XFILL_3__11593_ gnd vdd FILL
XFILL_1__12772_ gnd vdd FILL
XFILL_2__8985_ gnd vdd FILL
XFILL_5__7714_ gnd vdd FILL
XFILL_0_BUFX2_insert520 gnd vdd FILL
X_12628_ vdd memoryOutData[20] gnd _12629_/C vdd NAND2X1
XFILL_0_BUFX2_insert531 gnd vdd FILL
X_15416_ _15416_/A _16089_/B gnd _15416_/Y vdd NOR2X1
XFILL_3__13332_ gnd vdd FILL
XFILL_5__8694_ gnd vdd FILL
XFILL_0_BUFX2_insert542 gnd vdd FILL
XFILL_3__16120_ gnd vdd FILL
XFILL_4__11903_ gnd vdd FILL
XFILL_5__12153_ gnd vdd FILL
X_16396_ _16076_/A gnd _16396_/Y vdd INVX1
XFILL_4__15671_ gnd vdd FILL
XFILL_1__14511_ gnd vdd FILL
XFILL_3__10544_ gnd vdd FILL
XFILL_0_BUFX2_insert553 gnd vdd FILL
XFILL_2__7936_ gnd vdd FILL
XFILL_0__13152_ gnd vdd FILL
XFILL_1__11723_ gnd vdd FILL
XFILL_4__12883_ gnd vdd FILL
XFILL_0__10364_ gnd vdd FILL
XFILL_1__15491_ gnd vdd FILL
XFILL_0_BUFX2_insert564 gnd vdd FILL
X_15347_ _15347_/A _15347_/B gnd _15348_/B vdd NOR2X1
XFILL_0_BUFX2_insert575 gnd vdd FILL
XSFILL84200x57050 gnd vdd FILL
XFILL_5__11104_ gnd vdd FILL
XFILL_0__6951_ gnd vdd FILL
X_12559_ _12083_/B _12538_/CLK _12689_/R vdd _12513_/Y gnd vdd DFFSR
XFILL_4__14622_ gnd vdd FILL
XFILL_5__12084_ gnd vdd FILL
XFILL_0_BUFX2_insert586 gnd vdd FILL
XFILL_3__16051_ gnd vdd FILL
XFILL_3__13263_ gnd vdd FILL
XFILL_0__12103_ gnd vdd FILL
XFILL_2__15801_ gnd vdd FILL
XFILL_4__11834_ gnd vdd FILL
XFILL_2__7867_ gnd vdd FILL
XFILL_0_BUFX2_insert597 gnd vdd FILL
XFILL_1__14442_ gnd vdd FILL
XFILL_2__13993_ gnd vdd FILL
XFILL_0__13083_ gnd vdd FILL
XFILL_1__11654_ gnd vdd FILL
XFILL_0__10295_ gnd vdd FILL
XFILL_5__15912_ gnd vdd FILL
XFILL_3__15002_ gnd vdd FILL
XFILL_5__7576_ gnd vdd FILL
XFILL_5__11035_ gnd vdd FILL
XFILL_0__9670_ gnd vdd FILL
XSFILL59000x33050 gnd vdd FILL
XFILL_3__12214_ gnd vdd FILL
X_15278_ _15760_/A _13730_/D _15278_/C gnd _15280_/A vdd OAI21X1
XFILL_4__14553_ gnd vdd FILL
XFILL_0__6882_ gnd vdd FILL
XFILL_2__9606_ gnd vdd FILL
XFILL_2__15732_ gnd vdd FILL
XFILL_0__12034_ gnd vdd FILL
XFILL_4__11765_ gnd vdd FILL
XFILL_2__7798_ gnd vdd FILL
XFILL_1__14373_ gnd vdd FILL
X_14229_ _8038_/Q gnd _14229_/Y vdd INVX1
XFILL_0__8621_ gnd vdd FILL
XFILL_1__11585_ gnd vdd FILL
X_7160_ _7160_/A _7207_/A _7160_/C gnd _7254_/D vdd OAI21X1
XFILL_5__15843_ gnd vdd FILL
XFILL_4__13504_ gnd vdd FILL
XFILL_3__8330_ gnd vdd FILL
XFILL_1__16112_ gnd vdd FILL
XFILL_3__12145_ gnd vdd FILL
XFILL_1__13324_ gnd vdd FILL
XFILL_4__14484_ gnd vdd FILL
XFILL_2__15663_ gnd vdd FILL
XFILL_4__11696_ gnd vdd FILL
XFILL_2__9537_ gnd vdd FILL
XFILL_1__10536_ gnd vdd FILL
XFILL_2__12875_ gnd vdd FILL
XSFILL23720x7050 gnd vdd FILL
XCLKBUF1_insert210 CLKBUF1_insert206/A gnd _7268_/CLK vdd CLKBUF1
XFILL_5__9246_ gnd vdd FILL
XSFILL44040x50 gnd vdd FILL
XSFILL109800x21050 gnd vdd FILL
XFILL_4__16223_ gnd vdd FILL
XCLKBUF1_insert221 CLKBUF1_insert193/A gnd _8792_/CLK vdd CLKBUF1
XFILL_2__14614_ gnd vdd FILL
XFILL_4__13435_ gnd vdd FILL
XFILL_4__10647_ gnd vdd FILL
XFILL_5__15774_ gnd vdd FILL
X_7091_ _7124_/A _9907_/B gnd _7091_/Y vdd NAND2X1
XSFILL64120x24050 gnd vdd FILL
XFILL_1__16043_ gnd vdd FILL
XFILL_3__12076_ gnd vdd FILL
XFILL_3__8261_ gnd vdd FILL
XFILL_5__12986_ gnd vdd FILL
XFILL_2__9468_ gnd vdd FILL
XFILL_2__11826_ gnd vdd FILL
XFILL_1__13255_ gnd vdd FILL
XFILL_2__15594_ gnd vdd FILL
XFILL_0__7503_ gnd vdd FILL
XFILL_0__13985_ gnd vdd FILL
XFILL_5__14725_ gnd vdd FILL
XFILL_3__15904_ gnd vdd FILL
XFILL_0__8483_ gnd vdd FILL
XFILL_5__11937_ gnd vdd FILL
XFILL_3__7212_ gnd vdd FILL
XFILL_3__11027_ gnd vdd FILL
XFILL_4__16154_ gnd vdd FILL
XFILL_4__13366_ gnd vdd FILL
XFILL_2__14545_ gnd vdd FILL
XFILL_1__12206_ gnd vdd FILL
XFILL_4__10578_ gnd vdd FILL
XFILL_3__8192_ gnd vdd FILL
XFILL_5__8128_ gnd vdd FILL
XFILL_2__9399_ gnd vdd FILL
XFILL_0__15724_ gnd vdd FILL
XFILL_2__11757_ gnd vdd FILL
XFILL_1__10398_ gnd vdd FILL
XSFILL53960x67050 gnd vdd FILL
XFILL_0__7434_ gnd vdd FILL
XFILL_4__15105_ gnd vdd FILL
XSFILL3560x31050 gnd vdd FILL
XFILL_5__14656_ gnd vdd FILL
XFILL_4__12317_ gnd vdd FILL
XFILL_4__13297_ gnd vdd FILL
XFILL_3__15835_ gnd vdd FILL
XFILL_5__11868_ gnd vdd FILL
XFILL_2__10708_ gnd vdd FILL
XFILL_4__16085_ gnd vdd FILL
XFILL_2__14476_ gnd vdd FILL
XFILL_1__12137_ gnd vdd FILL
XFILL_0__15655_ gnd vdd FILL
XFILL_5__8059_ gnd vdd FILL
XFILL_2__11688_ gnd vdd FILL
XSFILL43400x25050 gnd vdd FILL
XFILL_5__13607_ gnd vdd FILL
XFILL_0__12867_ gnd vdd FILL
X_9801_ _9801_/A _9785_/A _9800_/Y gnd _9841_/D vdd OAI21X1
XFILL_2__16215_ gnd vdd FILL
XFILL_4__15036_ gnd vdd FILL
XFILL_4__12248_ gnd vdd FILL
XFILL_0__7365_ gnd vdd FILL
XFILL_5__10819_ gnd vdd FILL
XFILL_5__14587_ gnd vdd FILL
XFILL_2__13427_ gnd vdd FILL
XFILL_2__10639_ gnd vdd FILL
XSFILL54040x76050 gnd vdd FILL
XFILL_0__14606_ gnd vdd FILL
XFILL_3__7074_ gnd vdd FILL
X_7993_ _7970_/B _9017_/B gnd _7994_/C vdd NAND2X1
XFILL_3__15766_ gnd vdd FILL
XFILL_5__11799_ gnd vdd FILL
XFILL_0__9104_ gnd vdd FILL
XFILL_1__12068_ gnd vdd FILL
XFILL_3__12978_ gnd vdd FILL
XFILL_0__11818_ gnd vdd FILL
XFILL_5__16326_ gnd vdd FILL
XFILL_0__15586_ gnd vdd FILL
XFILL_6__8872_ gnd vdd FILL
XSFILL94440x81050 gnd vdd FILL
X_9732_ _9732_/A _9741_/B _9731_/Y gnd _9818_/D vdd OAI21X1
XFILL_5__13538_ gnd vdd FILL
XFILL_0__7296_ gnd vdd FILL
XFILL_4__12179_ gnd vdd FILL
X_6944_ _7012_/Q gnd _6946_/A vdd INVX1
XFILL_3__14717_ gnd vdd FILL
XFILL_2__16146_ gnd vdd FILL
XFILL_2__13358_ gnd vdd FILL
XFILL_3__11929_ gnd vdd FILL
XFILL_1__11019_ gnd vdd FILL
XFILL_3__15697_ gnd vdd FILL
XFILL_0__14537_ gnd vdd FILL
XFILL_0__9035_ gnd vdd FILL
XFILL_0__11749_ gnd vdd FILL
XFILL_5__16257_ gnd vdd FILL
X_9663_ _9615_/A _7231_/B gnd _9664_/C vdd NAND2X1
XFILL_5__13469_ gnd vdd FILL
XFILL_2__12309_ gnd vdd FILL
XSFILL33880x34050 gnd vdd FILL
XFILL_1__15827_ gnd vdd FILL
X_6875_ _6875_/A gnd memoryWriteData[5] vdd BUFX2
XFILL_2__16077_ gnd vdd FILL
XFILL_3__14648_ gnd vdd FILL
XFILL_2__13289_ gnd vdd FILL
XSFILL58680x79050 gnd vdd FILL
XFILL_0__14468_ gnd vdd FILL
XFILL_5__15208_ gnd vdd FILL
XFILL111800x12050 gnd vdd FILL
X_8614_ _8678_/Q gnd _8614_/Y vdd INVX1
XFILL_5__16188_ gnd vdd FILL
XFILL_2__15028_ gnd vdd FILL
XFILL_4__15938_ gnd vdd FILL
XFILL_6__14759_ gnd vdd FILL
XFILL_0__16207_ gnd vdd FILL
XSFILL48920x56050 gnd vdd FILL
X_9594_ _9628_/B _9082_/B gnd _9595_/C vdd NAND2X1
XFILL_3__14579_ gnd vdd FILL
XFILL_0__13419_ gnd vdd FILL
XFILL_1__15758_ gnd vdd FILL
XFILL_3__7976_ gnd vdd FILL
XFILL_5_BUFX2_insert703 gnd vdd FILL
XFILL_0__14399_ gnd vdd FILL
XFILL_5__15139_ gnd vdd FILL
X_8545_ _8545_/Q _9707_/CLK _8801_/R vdd _8545_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert714 gnd vdd FILL
XFILL_3__16318_ gnd vdd FILL
XFILL_1__6991_ gnd vdd FILL
XFILL_1__14709_ gnd vdd FILL
XFILL_5_BUFX2_insert725 gnd vdd FILL
XFILL_4__15869_ gnd vdd FILL
XFILL_3__6927_ gnd vdd FILL
XFILL_5_BUFX2_insert736 gnd vdd FILL
XFILL_0__16138_ gnd vdd FILL
XFILL_1__15689_ gnd vdd FILL
XFILL_5_BUFX2_insert747 gnd vdd FILL
XSFILL49000x65050 gnd vdd FILL
XFILL_1__8730_ gnd vdd FILL
XFILL_5_BUFX2_insert758 gnd vdd FILL
XFILL_0__9937_ gnd vdd FILL
XFILL_5_BUFX2_insert769 gnd vdd FILL
X_8476_ _8474_/Y _8484_/A _8476_/C gnd _8546_/D vdd OAI21X1
XFILL_3__16249_ gnd vdd FILL
XSFILL89400x70050 gnd vdd FILL
XFILL_3__6858_ gnd vdd FILL
XFILL_3__9646_ gnd vdd FILL
XFILL_0__16069_ gnd vdd FILL
XSFILL3640x11050 gnd vdd FILL
XSFILL109560x76050 gnd vdd FILL
X_7427_ _7503_/B _9859_/B gnd _7428_/C vdd NAND2X1
XFILL_1__8661_ gnd vdd FILL
XFILL_0__9868_ gnd vdd FILL
XFILL_4__8370_ gnd vdd FILL
XSFILL28840x23050 gnd vdd FILL
XFILL_1__7612_ gnd vdd FILL
XSFILL54120x56050 gnd vdd FILL
XFILL_6__9286_ gnd vdd FILL
XFILL_1__8592_ gnd vdd FILL
X_7358_ _7406_/Q gnd _7358_/Y vdd INVX1
XFILL_4__7321_ gnd vdd FILL
XFILL_0__9799_ gnd vdd FILL
XFILL_3__8528_ gnd vdd FILL
XFILL_6__8237_ gnd vdd FILL
XFILL_1__7543_ gnd vdd FILL
XFILL_3__8459_ gnd vdd FILL
X_7289_ _7383_/Q gnd _7289_/Y vdd INVX1
XFILL_4__7252_ gnd vdd FILL
XSFILL104120x25050 gnd vdd FILL
X_9028_ _9028_/A gnd _9030_/A vdd INVX1
XFILL_1__7474_ gnd vdd FILL
XFILL_4__7183_ gnd vdd FILL
XFILL_1__9213_ gnd vdd FILL
XSFILL18760x75050 gnd vdd FILL
XFILL_2_BUFX2_insert604 gnd vdd FILL
XSFILL105000x53050 gnd vdd FILL
XFILL_2_BUFX2_insert615 gnd vdd FILL
XSFILL58360x61050 gnd vdd FILL
XFILL_2_BUFX2_insert626 gnd vdd FILL
X_11930_ _11921_/A _12385_/A gnd _11930_/Y vdd NAND2X1
XFILL_2_BUFX2_insert637 gnd vdd FILL
XFILL_2_BUFX2_insert648 gnd vdd FILL
XFILL_1__9144_ gnd vdd FILL
XFILL_2_BUFX2_insert659 gnd vdd FILL
X_11861_ _12029_/A _12458_/B _12053_/A gnd _11862_/B vdd NOR3X1
XSFILL23880x66050 gnd vdd FILL
X_13600_ _7513_/Q gnd _13600_/Y vdd INVX1
X_10812_ _10831_/B _9532_/B gnd _10812_/Y vdd NAND2X1
X_14580_ _14580_/A _14580_/B _14579_/Y gnd _14596_/B vdd NAND3X1
X_11792_ _11034_/B _11778_/B _11792_/C gnd _11792_/Y vdd OAI21X1
XSFILL113880x19050 gnd vdd FILL
XFILL_5_BUFX2_insert19 gnd vdd FILL
X_13531_ _13528_/Y _13530_/Y _13531_/C gnd _13532_/B vdd NAND3X1
X_10743_ _6903_/A _10762_/B gnd _10743_/Y vdd NAND2X1
XBUFX2_insert603 BUFX2_insert570/A gnd _12692_/R vdd BUFX2
XSFILL39560x54050 gnd vdd FILL
XBUFX2_insert614 _10926_/Y gnd _11999_/A vdd BUFX2
XBUFX2_insert625 _12363_/Y gnd _9353_/B vdd BUFX2
XBUFX2_insert636 _12354_/Y gnd _9600_/B vdd BUFX2
XFILL_4__9755_ gnd vdd FILL
X_16250_ _15696_/A _10100_/Q _10192_/A _15695_/D gnd _16251_/B vdd AOI22X1
XFILL_4__6967_ gnd vdd FILL
X_13462_ _13456_/Y _13462_/B gnd _13474_/A vdd NOR2X1
XFILL_6_BUFX2_insert592 gnd vdd FILL
XBUFX2_insert647 _10915_/Y gnd _11988_/B vdd BUFX2
X_10674_ _14414_/D gnd _10676_/A vdd INVX1
XBUFX2_insert658 _11988_/Y gnd _12073_/C vdd BUFX2
XFILL_2__8770_ gnd vdd FILL
X_15201_ _15201_/A _15200_/Y gnd _15201_/Y vdd NOR2X1
XFILL_4__8706_ gnd vdd FILL
XBUFX2_insert669 _12345_/Y gnd _6903_/A vdd BUFX2
XFILL_1__9977_ gnd vdd FILL
X_12413_ _12368_/A _12413_/B gnd _12414_/C vdd NAND2X1
X_16181_ _14826_/Y _15197_/B _15197_/C _14808_/Y gnd _16184_/B vdd OAI22X1
XFILL_4__6898_ gnd vdd FILL
X_13393_ _13372_/A _13418_/A _13404_/B gnd _13393_/Y vdd NAND3X1
XFILL_2__7721_ gnd vdd FILL
XFILL_5__7430_ gnd vdd FILL
XFILL_4__8637_ gnd vdd FILL
XSFILL18840x55050 gnd vdd FILL
X_15132_ _15563_/A _15132_/B _15563_/C _15132_/D gnd _15135_/B vdd OAI22X1
X_12344_ _12663_/Q _12422_/A gnd _12345_/C vdd NAND2X1
XSFILL84280x31050 gnd vdd FILL
XFILL_3__10260_ gnd vdd FILL
XFILL_1__8859_ gnd vdd FILL
XFILL_2__10990_ gnd vdd FILL
XFILL_5__7361_ gnd vdd FILL
XFILL_4__8568_ gnd vdd FILL
X_15063_ _10358_/A gnd _15066_/B vdd INVX1
XSFILL99320x53050 gnd vdd FILL
X_12275_ _12239_/A gnd _12239_/C gnd _12278_/A vdd NAND3X1
XFILL_4__11550_ gnd vdd FILL
XFILL_3__10191_ gnd vdd FILL
XFILL_5__9100_ gnd vdd FILL
XFILL_2__7583_ gnd vdd FILL
X_14014_ _8215_/A gnd _14014_/Y vdd INVX1
XFILL_1__11370_ gnd vdd FILL
XFILL_4__10501_ gnd vdd FILL
XFILL_5__7292_ gnd vdd FILL
XFILL_4__8499_ gnd vdd FILL
X_11226_ _11220_/A _11226_/B _11223_/Y gnd _11230_/B vdd OAI21X1
XFILL_6__13090_ gnd vdd FILL
XFILL_5__12840_ gnd vdd FILL
XFILL_4__11481_ gnd vdd FILL
XFILL_2__12660_ gnd vdd FILL
XFILL_1__10321_ gnd vdd FILL
XFILL112280x13050 gnd vdd FILL
XFILL_5__9031_ gnd vdd FILL
XFILL_4__13220_ gnd vdd FILL
XFILL_4__10432_ gnd vdd FILL
X_11157_ _12298_/Y _11113_/Y gnd _11157_/Y vdd NOR2X1
XFILL_2__9253_ gnd vdd FILL
XFILL_5__12771_ gnd vdd FILL
XFILL_2__11611_ gnd vdd FILL
XFILL_1__10252_ gnd vdd FILL
XFILL_1__13040_ gnd vdd FILL
XFILL_3__13950_ gnd vdd FILL
XFILL_2__12591_ gnd vdd FILL
XFILL_3_BUFX2_insert460 gnd vdd FILL
XFILL_3_BUFX2_insert471 gnd vdd FILL
XFILL_0__13770_ gnd vdd FILL
XFILL_5__14510_ gnd vdd FILL
X_10108_ _13572_/A gnd _10108_/Y vdd INVX1
XFILL_0__10982_ gnd vdd FILL
XFILL_2__8204_ gnd vdd FILL
XFILL_4__13151_ gnd vdd FILL
XFILL_5__11722_ gnd vdd FILL
XFILL_3_BUFX2_insert482 gnd vdd FILL
X_15965_ _15965_/A _15961_/Y gnd _15965_/Y vdd NOR2X1
XFILL_3__12901_ gnd vdd FILL
XFILL_2__14330_ gnd vdd FILL
XFILL_4__10363_ gnd vdd FILL
X_11088_ _12270_/Y _11278_/B gnd _11090_/C vdd NOR2X1
XFILL_5__15490_ gnd vdd FILL
XFILL_3_BUFX2_insert493 gnd vdd FILL
XFILL_2__11542_ gnd vdd FILL
XSFILL79240x20050 gnd vdd FILL
XFILL_0__12721_ gnd vdd FILL
XFILL_3__13881_ gnd vdd FILL
XFILL_1__10183_ gnd vdd FILL
XFILL_4__12102_ gnd vdd FILL
XSFILL3480x46050 gnd vdd FILL
X_10039_ _10039_/A _9996_/A _10038_/Y gnd _10091_/D vdd OAI21X1
X_14916_ _14915_/Y _14916_/B gnd _14916_/Y vdd NOR2X1
XFILL_5__14441_ gnd vdd FILL
XFILL_3__15620_ gnd vdd FILL
XFILL_2__8135_ gnd vdd FILL
XFILL_4__13082_ gnd vdd FILL
XFILL_5__11653_ gnd vdd FILL
XFILL_4__10294_ gnd vdd FILL
X_15896_ _15893_/Y _15895_/Y _15896_/C gnd _15902_/C vdd NOR3X1
XFILL_2__14261_ gnd vdd FILL
XFILL_3__12832_ gnd vdd FILL
XFILL_0__15440_ gnd vdd FILL
XFILL_2__11473_ gnd vdd FILL
XFILL_0__12652_ gnd vdd FILL
XFILL_5__9933_ gnd vdd FILL
XFILL_1__14991_ gnd vdd FILL
XFILL_2__16000_ gnd vdd FILL
XFILL_6__15731_ gnd vdd FILL
XFILL_4__12033_ gnd vdd FILL
XFILL_2__13212_ gnd vdd FILL
X_14847_ _7885_/A _13865_/B _14847_/C _7155_/Q gnd _14858_/A vdd AOI22X1
XFILL_5__14372_ gnd vdd FILL
XFILL_3__12763_ gnd vdd FILL
XFILL_2__8066_ gnd vdd FILL
XFILL_3__15551_ gnd vdd FILL
XFILL_2__10424_ gnd vdd FILL
XFILL_5__11584_ gnd vdd FILL
XFILL_2__14192_ gnd vdd FILL
XFILL_0__11603_ gnd vdd FILL
XSFILL84360x11050 gnd vdd FILL
XFILL_1__13942_ gnd vdd FILL
XFILL_0__15371_ gnd vdd FILL
XFILL_5__16111_ gnd vdd FILL
XFILL_5__13323_ gnd vdd FILL
XFILL_0__12583_ gnd vdd FILL
XFILL_5__9864_ gnd vdd FILL
XFILL_5__10535_ gnd vdd FILL
XFILL_3__14502_ gnd vdd FILL
XFILL_3__11714_ gnd vdd FILL
XFILL_0__7081_ gnd vdd FILL
XFILL_2__13143_ gnd vdd FILL
X_14778_ _14778_/A _14778_/B _14030_/C _16151_/D gnd _14778_/Y vdd OAI22X1
XFILL_0__14322_ gnd vdd FILL
XFILL_3__15482_ gnd vdd FILL
XFILL_1__13873_ gnd vdd FILL
XSFILL99400x33050 gnd vdd FILL
XFILL_0__11534_ gnd vdd FILL
XFILL_5__16042_ gnd vdd FILL
XFILL_5__13254_ gnd vdd FILL
X_13729_ _7515_/Q gnd _13730_/D vdd INVX1
XFILL_5__9795_ gnd vdd FILL
XFILL_1__15612_ gnd vdd FILL
XFILL111720x27050 gnd vdd FILL
XFILL_3__11645_ gnd vdd FILL
XFILL_3__14433_ gnd vdd FILL
XFILL_4__13984_ gnd vdd FILL
XFILL_1__12824_ gnd vdd FILL
XFILL_3__7830_ gnd vdd FILL
XFILL_0__14253_ gnd vdd FILL
XFILL_2__10286_ gnd vdd FILL
XFILL_0__11465_ gnd vdd FILL
XFILL_6__14544_ gnd vdd FILL
XFILL_5__12205_ gnd vdd FILL
XFILL_5__8746_ gnd vdd FILL
XFILL_4__15723_ gnd vdd FILL
X_16448_ _16448_/Q _9589_/CLK _7537_/R vdd _16448_/D gnd vdd DFFSR
XSFILL104360x81050 gnd vdd FILL
XFILL_2__12025_ gnd vdd FILL
XFILL_3__14364_ gnd vdd FILL
XFILL_5__10397_ gnd vdd FILL
XSFILL64120x19050 gnd vdd FILL
XFILL_1__15543_ gnd vdd FILL
XFILL_3__11576_ gnd vdd FILL
XFILL_3__7761_ gnd vdd FILL
XFILL_1__12755_ gnd vdd FILL
XFILL_2__8968_ gnd vdd FILL
XFILL_0_BUFX2_insert350 gnd vdd FILL
XFILL_0__10416_ gnd vdd FILL
XSFILL74280x63050 gnd vdd FILL
XFILL_0__14184_ gnd vdd FILL
XFILL_0__11396_ gnd vdd FILL
XFILL_0_BUFX2_insert361 gnd vdd FILL
XFILL_5__12136_ gnd vdd FILL
X_8330_ _8328_/Y _8356_/A _8329_/Y gnd _8412_/D vdd OAI21X1
XFILL_3__16103_ gnd vdd FILL
XFILL_0_BUFX2_insert372 gnd vdd FILL
XFILL_3__13315_ gnd vdd FILL
XFILL_4__15654_ gnd vdd FILL
XFILL_3__9500_ gnd vdd FILL
X_16379_ gnd gnd gnd _16379_/Y vdd NAND2X1
XFILL_0__7983_ gnd vdd FILL
XFILL_3__10527_ gnd vdd FILL
XFILL_4__12866_ gnd vdd FILL
XFILL_1__11706_ gnd vdd FILL
XFILL_3__14295_ gnd vdd FILL
XFILL_0_BUFX2_insert383 gnd vdd FILL
XFILL_3__7692_ gnd vdd FILL
XFILL_0__13135_ gnd vdd FILL
XFILL_0_BUFX2_insert394 gnd vdd FILL
XFILL_1__15474_ gnd vdd FILL
XFILL_5__7628_ gnd vdd FILL
XFILL_2__8899_ gnd vdd FILL
XFILL_4__14605_ gnd vdd FILL
XFILL_0__6934_ gnd vdd FILL
XFILL_0__9722_ gnd vdd FILL
XFILL_3__13246_ gnd vdd FILL
XFILL_3__16034_ gnd vdd FILL
XFILL_5__12067_ gnd vdd FILL
X_8261_ _8216_/A _6981_/B gnd _8262_/C vdd NAND2X1
XFILL_4__11817_ gnd vdd FILL
XFILL_4__15585_ gnd vdd FILL
XSFILL3560x26050 gnd vdd FILL
XFILL_1__14425_ gnd vdd FILL
XFILL_2__13976_ gnd vdd FILL
XFILL_1__11637_ gnd vdd FILL
XFILL_0__10278_ gnd vdd FILL
XFILL_6__16145_ gnd vdd FILL
XFILL_6__13357_ gnd vdd FILL
XFILL_0__9653_ gnd vdd FILL
X_7212_ _7212_/A gnd _7214_/A vdd INVX1
XFILL_5__7559_ gnd vdd FILL
XFILL_5__11018_ gnd vdd FILL
XFILL_4__14536_ gnd vdd FILL
XFILL_0__6865_ gnd vdd FILL
X_8192_ _8208_/B _8576_/B gnd _8193_/C vdd NAND2X1
XFILL_2__15715_ gnd vdd FILL
XFILL_3__9362_ gnd vdd FILL
XFILL_4__11748_ gnd vdd FILL
XFILL_0__12017_ gnd vdd FILL
XFILL_1__14356_ gnd vdd FILL
XFILL_3__10389_ gnd vdd FILL
XFILL_0__8604_ gnd vdd FILL
XFILL_1__11568_ gnd vdd FILL
XSFILL33880x8050 gnd vdd FILL
XSFILL94440x76050 gnd vdd FILL
XFILL_3__12128_ gnd vdd FILL
XFILL_5__15826_ gnd vdd FILL
XFILL_3__8313_ gnd vdd FILL
X_7143_ _7081_/A _7143_/CLK _9959_/R vdd _7143_/D gnd vdd DFFSR
XFILL_1__13307_ gnd vdd FILL
XFILL_4__14467_ gnd vdd FILL
XFILL_3__9293_ gnd vdd FILL
XFILL_2__15646_ gnd vdd FILL
XFILL_1__10519_ gnd vdd FILL
XFILL_2__12858_ gnd vdd FILL
XFILL_4__11679_ gnd vdd FILL
XFILL_5__9229_ gnd vdd FILL
XFILL_1__14287_ gnd vdd FILL
XFILL_4__16206_ gnd vdd FILL
XFILL_6__12239_ gnd vdd FILL
XFILL_1__11499_ gnd vdd FILL
XFILL_4__13418_ gnd vdd FILL
X_7074_ _7074_/A _7095_/B _7073_/Y gnd _7140_/D vdd OAI21X1
XFILL_5__15757_ gnd vdd FILL
XFILL_1__16026_ gnd vdd FILL
XSFILL69240x52050 gnd vdd FILL
XFILL_3__12059_ gnd vdd FILL
XFILL_5__12969_ gnd vdd FILL
XSFILL33880x29050 gnd vdd FILL
XFILL_3__8244_ gnd vdd FILL
XFILL_2__11809_ gnd vdd FILL
XFILL_1__13238_ gnd vdd FILL
XFILL_4__14398_ gnd vdd FILL
XFILL_5_BUFX2_insert1040 gnd vdd FILL
XFILL_2__12789_ gnd vdd FILL
XFILL_5_BUFX2_insert1051 gnd vdd FILL
XFILL_2__15577_ gnd vdd FILL
XFILL_5_BUFX2_insert1062 gnd vdd FILL
XFILL_5__14708_ gnd vdd FILL
XFILL_0__13968_ gnd vdd FILL
XFILL_5_BUFX2_insert1073 gnd vdd FILL
XFILL_0__8466_ gnd vdd FILL
XFILL_4__16137_ gnd vdd FILL
XFILL_4__13349_ gnd vdd FILL
XFILL_5_BUFX2_insert1084 gnd vdd FILL
XFILL_5__15688_ gnd vdd FILL
XFILL_0__15707_ gnd vdd FILL
XFILL_2__14528_ gnd vdd FILL
XSFILL73720x77050 gnd vdd FILL
XFILL_1__13169_ gnd vdd FILL
XFILL_0__7417_ gnd vdd FILL
XFILL_5__14639_ gnd vdd FILL
XFILL_0__13899_ gnd vdd FILL
XFILL_0__8397_ gnd vdd FILL
XFILL_3__15818_ gnd vdd FILL
XFILL_1__7190_ gnd vdd FILL
XFILL_4__16068_ gnd vdd FILL
XFILL_2__14459_ gnd vdd FILL
XSFILL79240x7050 gnd vdd FILL
XFILL_0__15638_ gnd vdd FILL
XFILL_4__15019_ gnd vdd FILL
XFILL_0__7348_ gnd vdd FILL
X_7976_ _7976_/A _7948_/A _7975_/Y gnd _7976_/Y vdd OAI21X1
XFILL_3__7057_ gnd vdd FILL
XFILL_3__15749_ gnd vdd FILL
XFILL_0__15569_ gnd vdd FILL
XFILL_5__16309_ gnd vdd FILL
X_9715_ _9677_/A _8306_/CLK _7533_/R vdd _9715_/D gnd vdd DFFSR
X_6927_ _6988_/B _8719_/B gnd _6928_/C vdd NAND2X1
XFILL_2__16129_ gnd vdd FILL
XFILL_4__7870_ gnd vdd FILL
XFILL_0__9018_ gnd vdd FILL
XSFILL28840x18050 gnd vdd FILL
XFILL_1__9900_ gnd vdd FILL
X_9646_ _9644_/Y _9628_/B _9645_/Y gnd _9704_/D vdd OAI21X1
X_6858_ _6858_/A gnd memoryAddress[20] vdd BUFX2
XSFILL13640x60050 gnd vdd FILL
XSFILL79080x55050 gnd vdd FILL
XFILL_5_BUFX2_insert500 gnd vdd FILL
XSFILL28440x20050 gnd vdd FILL
XFILL_5_BUFX2_insert511 gnd vdd FILL
X_9577_ _9577_/Q _9705_/CLK _9964_/R vdd _9577_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert522 gnd vdd FILL
XFILL_4__9540_ gnd vdd FILL
XFILL_3__7959_ gnd vdd FILL
XFILL_5_BUFX2_insert533 gnd vdd FILL
XFILL_5_BUFX2_insert544 gnd vdd FILL
X_8528_ _8564_/Q gnd _8528_/Y vdd INVX1
XFILL_1__6974_ gnd vdd FILL
XFILL_1__9762_ gnd vdd FILL
XFILL_5_BUFX2_insert555 gnd vdd FILL
XFILL_5_BUFX2_insert566 gnd vdd FILL
XFILL_4__9471_ gnd vdd FILL
XFILL_5_BUFX2_insert577 gnd vdd FILL
XFILL_3_BUFX2_insert3 gnd vdd FILL
XFILL_1__8713_ gnd vdd FILL
XFILL_5_BUFX2_insert588 gnd vdd FILL
X_10390_ _10390_/A _10450_/B _10389_/Y gnd _10464_/D vdd OAI21X1
X_8459_ _8459_/A gnd _8461_/A vdd INVX1
XSFILL104520x41050 gnd vdd FILL
XFILL_5_BUFX2_insert599 gnd vdd FILL
XFILL_3__9629_ gnd vdd FILL
XFILL_6__9338_ gnd vdd FILL
XSFILL33800x73050 gnd vdd FILL
XFILL_1__8644_ gnd vdd FILL
XFILL_4__8353_ gnd vdd FILL
X_12060_ _12012_/A _12807_/Q _11996_/C gnd _12062_/B vdd NAND3X1
XFILL_1__8575_ gnd vdd FILL
XFILL_2_CLKBUF1_insert114 gnd vdd FILL
XFILL_4__7304_ gnd vdd FILL
XFILL_2_CLKBUF1_insert125 gnd vdd FILL
X_11011_ _12222_/Y _12120_/Y gnd _11011_/Y vdd OR2X2
XFILL_2_CLKBUF1_insert136 gnd vdd FILL
XFILL_2_CLKBUF1_insert147 gnd vdd FILL
XFILL_2_CLKBUF1_insert158 gnd vdd FILL
XFILL_2_CLKBUF1_insert169 gnd vdd FILL
XFILL_4__7235_ gnd vdd FILL
XFILL_1__7457_ gnd vdd FILL
XFILL_2_BUFX2_insert401 gnd vdd FILL
XSFILL13720x40050 gnd vdd FILL
XFILL_2_BUFX2_insert412 gnd vdd FILL
XFILL_4__7166_ gnd vdd FILL
XFILL_2_BUFX2_insert423 gnd vdd FILL
X_12962_ _12960_/Y vdd _12962_/C gnd _12962_/Y vdd OAI21X1
X_15750_ _15801_/A _14292_/Y _15801_/C _15749_/Y gnd _15753_/B vdd OAI22X1
XFILL_2_BUFX2_insert434 gnd vdd FILL
XFILL_2_BUFX2_insert445 gnd vdd FILL
XFILL_2_BUFX2_insert456 gnd vdd FILL
X_11913_ _11913_/A _11934_/B _11912_/Y gnd _6846_/A vdd OAI21X1
XFILL_2_BUFX2_insert467 gnd vdd FILL
XFILL_4__7097_ gnd vdd FILL
X_14701_ _14701_/A _14700_/Y gnd _14701_/Y vdd NOR2X1
XFILL_1__9127_ gnd vdd FILL
X_15681_ _14199_/Y _15681_/B _15681_/C _14198_/Y gnd _15684_/B vdd OAI22X1
X_12893_ vdd _12893_/B gnd _12894_/C vdd NAND2X1
XFILL_2_BUFX2_insert478 gnd vdd FILL
XFILL_2_BUFX2_insert489 gnd vdd FILL
XFILL_5__6930_ gnd vdd FILL
X_14632_ _10094_/Q gnd _14632_/Y vdd INVX1
XSFILL84280x26050 gnd vdd FILL
X_11844_ _11843_/Y gnd _11226_/B gnd _11844_/Y vdd OAI21X1
XFILL_2__9940_ gnd vdd FILL
X_14563_ _7917_/Q gnd _14563_/Y vdd INVX1
XFILL_5__6861_ gnd vdd FILL
XFILL_5__10320_ gnd vdd FILL
XFILL_1__8009_ gnd vdd FILL
XSFILL99320x48050 gnd vdd FILL
X_11775_ _11762_/B _11758_/B gnd _11776_/C vdd NOR2X1
XFILL_2__10140_ gnd vdd FILL
XBUFX2_insert400 _13293_/Y gnd _7577_/B vdd BUFX2
XFILL_4__9807_ gnd vdd FILL
XFILL_2__9871_ gnd vdd FILL
XFILL_5__8600_ gnd vdd FILL
XBUFX2_insert411 _13484_/Y gnd _14572_/C vdd BUFX2
XFILL_1__10870_ gnd vdd FILL
X_16302_ _16302_/A _16301_/Y gnd _16308_/A vdd NOR2X1
XFILL_6__11610_ gnd vdd FILL
XFILL_5__10251_ gnd vdd FILL
X_10726_ _15704_/B _7411_/CLK _8929_/R vdd _10726_/D gnd vdd DFFSR
XBUFX2_insert422 _14991_/Y gnd _15945_/C vdd BUFX2
X_13514_ _13843_/C _13514_/B _13514_/C _13420_/C gnd _13514_/Y vdd OAI22X1
XBUFX2_insert433 _13326_/Y gnd _8740_/A vdd BUFX2
XFILL_4__7999_ gnd vdd FILL
X_14494_ _10293_/A gnd _14496_/B vdd INVX1
XFILL_3__11430_ gnd vdd FILL
XFILL_2__8822_ gnd vdd FILL
XBUFX2_insert444 _12378_/Y gnd _8472_/B vdd BUFX2
XFILL_4__10981_ gnd vdd FILL
XBUFX2_insert455 _13442_/Y gnd _14815_/C vdd BUFX2
XFILL_0__11250_ gnd vdd FILL
XFILL_4__9738_ gnd vdd FILL
XFILL_5__8531_ gnd vdd FILL
XBUFX2_insert466 _13318_/Y gnd _8321_/B vdd BUFX2
X_16233_ _15197_/C _14864_/Y _16232_/Y gnd _16236_/A vdd OAI21X1
X_13445_ _6998_/Q gnd _13445_/Y vdd INVX1
XFILL_4__12720_ gnd vdd FILL
X_10657_ _10658_/B _7713_/B gnd _10657_/Y vdd NAND2X1
XBUFX2_insert477 _15038_/Y gnd _15920_/B vdd BUFX2
XFILL_5__10182_ gnd vdd FILL
XBUFX2_insert488 _12372_/Y gnd _7186_/B vdd BUFX2
XFILL_3__11361_ gnd vdd FILL
XBUFX2_insert499 BUFX2_insert520/A gnd _7775_/R vdd BUFX2
XFILL_2__8753_ gnd vdd FILL
XFILL_0__11181_ gnd vdd FILL
XFILL_5__8462_ gnd vdd FILL
XFILL_3__13100_ gnd vdd FILL
XFILL_4__9669_ gnd vdd FILL
X_13376_ _11881_/A _13376_/B gnd _13718_/B vdd NOR2X1
XFILL_3__10312_ gnd vdd FILL
XSFILL13800x20050 gnd vdd FILL
X_16164_ _16140_/Y _16164_/B _14791_/C gnd _16164_/Y vdd AOI21X1
XFILL_4__12651_ gnd vdd FILL
XFILL_2__13830_ gnd vdd FILL
X_10588_ _15298_/D _7534_/CLK _8156_/R vdd _10506_/Y gnd vdd DFFSR
XFILL_5__14990_ gnd vdd FILL
XFILL_2__7704_ gnd vdd FILL
XFILL_3__14080_ gnd vdd FILL
XFILL_3__11292_ gnd vdd FILL
XFILL_0__10132_ gnd vdd FILL
XFILL_1__12471_ gnd vdd FILL
X_12327_ _12327_/A gnd _12319_/C gnd _12330_/A vdd NAND3X1
X_15115_ _15760_/A _13491_/Y _15115_/C gnd _15119_/A vdd OAI21X1
XFILL_5__8393_ gnd vdd FILL
XFILL_6__14191_ gnd vdd FILL
X_16095_ _16088_/Y _16095_/B _16093_/Y gnd _16102_/B vdd NAND3X1
XFILL_3__13031_ gnd vdd FILL
XFILL_4__11602_ gnd vdd FILL
XFILL_5__13941_ gnd vdd FILL
XFILL_1__14210_ gnd vdd FILL
XFILL_4__15370_ gnd vdd FILL
XFILL_3__10243_ gnd vdd FILL
XFILL_2__7635_ gnd vdd FILL
XFILL_4__12582_ gnd vdd FILL
XFILL_2__13761_ gnd vdd FILL
XFILL_1__11422_ gnd vdd FILL
XFILL_2__10973_ gnd vdd FILL
XFILL_0__10063_ gnd vdd FILL
XFILL_1__15190_ gnd vdd FILL
XFILL_0__14940_ gnd vdd FILL
XFILL_5__7344_ gnd vdd FILL
X_15046_ _15244_/C _14981_/Y _16035_/B gnd _15046_/Y vdd NAND3X1
XSFILL114440x24050 gnd vdd FILL
XFILL_4__14321_ gnd vdd FILL
X_12258_ _12255_/Y _12258_/B _12258_/C gnd _12258_/Y vdd NAND3X1
XFILL_5__13872_ gnd vdd FILL
XFILL_2__12712_ gnd vdd FILL
XFILL_2__15500_ gnd vdd FILL
XFILL_4__11533_ gnd vdd FILL
XFILL_2__7566_ gnd vdd FILL
XFILL_3__10174_ gnd vdd FILL
XFILL_1__14141_ gnd vdd FILL
XFILL_2__13692_ gnd vdd FILL
XFILL_1__11353_ gnd vdd FILL
XFILL_0__14871_ gnd vdd FILL
XFILL_5__15611_ gnd vdd FILL
X_11209_ _12330_/Y _11208_/Y gnd _11209_/Y vdd NOR2X1
XFILL_5__12823_ gnd vdd FILL
XFILL_4__14252_ gnd vdd FILL
X_12189_ _12187_/Y _12179_/A _12189_/C gnd _12189_/Y vdd OAI21X1
XFILL_1_BUFX2_insert17 gnd vdd FILL
XSFILL89240x2050 gnd vdd FILL
XFILL_1__10304_ gnd vdd FILL
XFILL_2__12643_ gnd vdd FILL
XFILL_1_BUFX2_insert28 gnd vdd FILL
XFILL_2__15431_ gnd vdd FILL
XFILL_4__11464_ gnd vdd FILL
XFILL_0__13822_ gnd vdd FILL
XFILL_5__9014_ gnd vdd FILL
XFILL_3__14982_ gnd vdd FILL
XFILL_1__14072_ gnd vdd FILL
XFILL_2__7497_ gnd vdd FILL
XFILL_1_BUFX2_insert39 gnd vdd FILL
XFILL_0__8320_ gnd vdd FILL
XSFILL69160x67050 gnd vdd FILL
XFILL_6__12024_ gnd vdd FILL
XSFILL99400x28050 gnd vdd FILL
XFILL_1__11284_ gnd vdd FILL
XFILL_5__15542_ gnd vdd FILL
XFILL_5__12754_ gnd vdd FILL
XFILL_4__10415_ gnd vdd FILL
XFILL_2__15362_ gnd vdd FILL
XFILL_4__14183_ gnd vdd FILL
XFILL_1__13023_ gnd vdd FILL
XFILL_4__11395_ gnd vdd FILL
XFILL_3__13933_ gnd vdd FILL
XFILL_2__9236_ gnd vdd FILL
XFILL_2__12574_ gnd vdd FILL
XFILL_3_BUFX2_insert290 gnd vdd FILL
XFILL_1__10235_ gnd vdd FILL
XSFILL84200x70050 gnd vdd FILL
XFILL_0__13753_ gnd vdd FILL
XFILL_0__10965_ gnd vdd FILL
XFILL_0__8251_ gnd vdd FILL
XFILL_5__11705_ gnd vdd FILL
XFILL_4__13134_ gnd vdd FILL
X_15948_ _16106_/A _15948_/B _15947_/Y _15948_/D gnd _15948_/Y vdd OAI22X1
XFILL_2__14313_ gnd vdd FILL
XFILL_5__15473_ gnd vdd FILL
XSFILL104360x76050 gnd vdd FILL
XFILL_2__9167_ gnd vdd FILL
XFILL_2__11525_ gnd vdd FILL
XFILL_0__12704_ gnd vdd FILL
XFILL_3__13864_ gnd vdd FILL
XFILL_2__15293_ gnd vdd FILL
XFILL_1__10166_ gnd vdd FILL
XFILL_0__7202_ gnd vdd FILL
XFILL_0__13684_ gnd vdd FILL
XSFILL89720x8050 gnd vdd FILL
XSFILL23640x23050 gnd vdd FILL
XFILL_5__14424_ gnd vdd FILL
XFILL_2__8118_ gnd vdd FILL
XFILL_0__8182_ gnd vdd FILL
XFILL_6__6970_ gnd vdd FILL
XFILL_0__10896_ gnd vdd FILL
XFILL_5__11636_ gnd vdd FILL
X_7830_ _7830_/A _7892_/A _7830_/C gnd _7830_/Y vdd OAI21X1
XFILL_3__15603_ gnd vdd FILL
XFILL_4__10277_ gnd vdd FILL
XFILL_2__14244_ gnd vdd FILL
XSFILL109400x13050 gnd vdd FILL
X_15879_ _15953_/A _15878_/Y _15841_/C _15879_/D gnd _15879_/Y vdd OAI22X1
XFILL_2__9098_ gnd vdd FILL
XFILL_2__11456_ gnd vdd FILL
XFILL_0__15423_ gnd vdd FILL
XFILL_0__12635_ gnd vdd FILL
XFILL_5__9916_ gnd vdd FILL
XFILL_3__13795_ gnd vdd FILL
XFILL_2_BUFX2_insert990 gnd vdd FILL
XFILL_1__14974_ gnd vdd FILL
XFILL_3__9980_ gnd vdd FILL
XFILL_4__12016_ gnd vdd FILL
XFILL_5__14355_ gnd vdd FILL
XSFILL49080x34050 gnd vdd FILL
XFILL_2__10407_ gnd vdd FILL
XFILL112200x52050 gnd vdd FILL
XFILL_3__15534_ gnd vdd FILL
XFILL_5__11567_ gnd vdd FILL
X_7761_ _7729_/B _8273_/B gnd _7761_/Y vdd NAND2X1
XFILL_3__12746_ gnd vdd FILL
XFILL_2__14175_ gnd vdd FILL
XFILL_1__13925_ gnd vdd FILL
XFILL_0__15354_ gnd vdd FILL
XFILL_2__11387_ gnd vdd FILL
XFILL_5__13306_ gnd vdd FILL
XFILL_6__8640_ gnd vdd FILL
XFILL_5__9847_ gnd vdd FILL
X_9500_ _9500_/A _9466_/A _9500_/C gnd _9570_/D vdd OAI21X1
XFILL_0__7064_ gnd vdd FILL
XFILL_6__12857_ gnd vdd FILL
XFILL_5__10518_ gnd vdd FILL
XFILL_2__13126_ gnd vdd FILL
XFILL_5__14286_ gnd vdd FILL
X_7692_ _7759_/B _7564_/B gnd _7693_/C vdd NAND2X1
XFILL_0__14305_ gnd vdd FILL
XFILL_5__11498_ gnd vdd FILL
XFILL_3__15465_ gnd vdd FILL
XFILL_1__13856_ gnd vdd FILL
XFILL_0__11517_ gnd vdd FILL
XFILL_3__8862_ gnd vdd FILL
XFILL_5__16025_ gnd vdd FILL
XFILL_0__15285_ gnd vdd FILL
XFILL_5__13237_ gnd vdd FILL
XFILL_0__12497_ gnd vdd FILL
X_9431_ _9431_/Q _9447_/CLK _9447_/R vdd _9339_/Y gnd vdd DFFSR
XFILL_5__9778_ gnd vdd FILL
XFILL_5__10449_ gnd vdd FILL
XFILL_3__14416_ gnd vdd FILL
XFILL_3__7813_ gnd vdd FILL
XFILL_3__11628_ gnd vdd FILL
XFILL_4__13967_ gnd vdd FILL
XFILL_3__15396_ gnd vdd FILL
XFILL_0__14236_ gnd vdd FILL
XFILL_2__10269_ gnd vdd FILL
XSFILL53960x80050 gnd vdd FILL
XFILL_5__8729_ gnd vdd FILL
XFILL_1__13787_ gnd vdd FILL
XFILL_0__11448_ gnd vdd FILL
XFILL_4__15706_ gnd vdd FILL
XFILL_1__10999_ gnd vdd FILL
XFILL_5__13168_ gnd vdd FILL
XFILL_2__12008_ gnd vdd FILL
XFILL_4__12918_ gnd vdd FILL
X_9362_ _9425_/A _9362_/B gnd _9362_/Y vdd NAND2X1
XSFILL69240x47050 gnd vdd FILL
XFILL_1__15526_ gnd vdd FILL
XFILL_3__14347_ gnd vdd FILL
XFILL_3__11559_ gnd vdd FILL
XFILL_3__7744_ gnd vdd FILL
XFILL_1__12738_ gnd vdd FILL
XFILL_4__13898_ gnd vdd FILL
XFILL_0__14167_ gnd vdd FILL
X_8313_ _8407_/Q gnd _8315_/A vdd INVX1
XFILL_0__11379_ gnd vdd FILL
XFILL_5__12119_ gnd vdd FILL
XFILL_4__15637_ gnd vdd FILL
XFILL_0__7966_ gnd vdd FILL
X_9293_ _9293_/A gnd _9293_/Y vdd INVX1
XFILL_4_BUFX2_insert507 gnd vdd FILL
XFILL_4__12849_ gnd vdd FILL
XFILL_5__13099_ gnd vdd FILL
XFILL_4_BUFX2_insert518 gnd vdd FILL
XFILL_0__13118_ gnd vdd FILL
XFILL_3__7675_ gnd vdd FILL
XFILL_1__15457_ gnd vdd FILL
XFILL_3__14278_ gnd vdd FILL
XFILL_4_BUFX2_insert529 gnd vdd FILL
XSFILL104440x56050 gnd vdd FILL
XFILL_0__6917_ gnd vdd FILL
XFILL_0__14098_ gnd vdd FILL
XFILL_3__16017_ gnd vdd FILL
X_8244_ _8242_/Y _8244_/B _8244_/C gnd _8244_/Y vdd OAI21X1
XFILL_3__13229_ gnd vdd FILL
XFILL_3__9414_ gnd vdd FILL
XFILL_4__15568_ gnd vdd FILL
XSFILL73880x31050 gnd vdd FILL
XFILL_1__14408_ gnd vdd FILL
XSFILL8680x54050 gnd vdd FILL
XFILL_1__15388_ gnd vdd FILL
XFILL_2__13959_ gnd vdd FILL
XFILL_0__9636_ gnd vdd FILL
XFILL_4__14519_ gnd vdd FILL
XFILL_0__6848_ gnd vdd FILL
X_8175_ _8129_/A _7007_/CLK _9332_/R vdd _8175_/D gnd vdd DFFSR
XFILL_3__9345_ gnd vdd FILL
XFILL_4__15499_ gnd vdd FILL
XFILL_1__14339_ gnd vdd FILL
XFILL_1__8360_ gnd vdd FILL
X_7126_ _7030_/A _8562_/CLK _9430_/R vdd _7126_/D gnd vdd DFFSR
XFILL_5__15809_ gnd vdd FILL
XFILL_2__15629_ gnd vdd FILL
XFILL_3__9276_ gnd vdd FILL
XFILL_1__7311_ gnd vdd FILL
XFILL_0__8518_ gnd vdd FILL
XFILL_1__16009_ gnd vdd FILL
XFILL_0__9498_ gnd vdd FILL
X_7057_ _7135_/Q gnd _7059_/A vdd INVX1
XFILL_3__8227_ gnd vdd FILL
XSFILL13640x55050 gnd vdd FILL
XFILL_3_CLKBUF1_insert209 gnd vdd FILL
XFILL_0__8449_ gnd vdd FILL
XFILL_1__7242_ gnd vdd FILL
XFILL_3__7109_ gnd vdd FILL
XFILL_1__7173_ gnd vdd FILL
XFILL_1_BUFX2_insert408 gnd vdd FILL
XFILL_3__8089_ gnd vdd FILL
XFILL_4__8971_ gnd vdd FILL
XSFILL114280x59050 gnd vdd FILL
XFILL_1_BUFX2_insert419 gnd vdd FILL
X_7959_ _7959_/A gnd _7959_/Y vdd INVX1
XSFILL104520x36050 gnd vdd FILL
XSFILL33800x68050 gnd vdd FILL
XSFILL8760x34050 gnd vdd FILL
XFILL_4__7853_ gnd vdd FILL
X_11560_ _11116_/Y gnd _11561_/A vdd INVX1
X_9629_ _9699_/Q gnd _9629_/Y vdd INVX1
XFILL_6__8769_ gnd vdd FILL
XFILL_1_CLKBUF1_insert1076 gnd vdd FILL
X_10511_ _10511_/A _8207_/B gnd _10512_/C vdd NAND2X1
XFILL_5_BUFX2_insert330 gnd vdd FILL
X_11491_ _11511_/A _11491_/B _11181_/Y gnd _11492_/A vdd AOI21X1
XFILL_5_BUFX2_insert341 gnd vdd FILL
XBUFX2_insert20 _13443_/Y gnd _14830_/B vdd BUFX2
XBUFX2_insert31 _13320_/Y gnd _8440_/B vdd BUFX2
XFILL_4__9523_ gnd vdd FILL
XFILL_5_BUFX2_insert352 gnd vdd FILL
X_13230_ _13288_/B gnd _13230_/Y vdd INVX2
XBUFX2_insert42 _14986_/Y gnd _15524_/A vdd BUFX2
X_10442_ _10442_/A gnd _10444_/A vdd INVX1
XSFILL108760x41050 gnd vdd FILL
XFILL_5_BUFX2_insert363 gnd vdd FILL
XBUFX2_insert53 _13309_/Y gnd _8100_/A vdd BUFX2
XFILL_5_BUFX2_insert374 gnd vdd FILL
XFILL_5_BUFX2_insert385 gnd vdd FILL
XFILL_1__6957_ gnd vdd FILL
XBUFX2_insert64 _12215_/Y gnd _12301_/B vdd BUFX2
XFILL_1__9745_ gnd vdd FILL
XBUFX2_insert75 _12366_/Y gnd _7948_/B vdd BUFX2
XFILL_5_BUFX2_insert396 gnd vdd FILL
XSFILL13720x35050 gnd vdd FILL
XBUFX2_insert86 _13390_/Y gnd _14068_/C vdd BUFX2
X_13161_ _13173_/A _13161_/B gnd _13162_/C vdd NAND2X1
X_10373_ _15261_/A gnd _10373_/Y vdd INVX1
XBUFX2_insert97 _15068_/Y gnd _15958_/B vdd BUFX2
XFILL_1__9676_ gnd vdd FILL
XFILL_1__6888_ gnd vdd FILL
XFILL_4__8405_ gnd vdd FILL
X_12112_ _11988_/B _13172_/A _12096_/C gnd _12114_/B vdd NAND3X1
XFILL_4__9385_ gnd vdd FILL
X_13092_ _13099_/B _13092_/B gnd _13093_/C vdd NAND2X1
XFILL_2__7420_ gnd vdd FILL
XFILL_1__8627_ gnd vdd FILL
XFILL_4__8336_ gnd vdd FILL
X_12043_ _12031_/A _12385_/A _12031_/C gnd _12046_/A vdd NAND3X1
XFILL_2__7351_ gnd vdd FILL
XSFILL13640x1050 gnd vdd FILL
XFILL_5__7060_ gnd vdd FILL
XFILL_4__8267_ gnd vdd FILL
XFILL_1__7509_ gnd vdd FILL
XFILL_1__8489_ gnd vdd FILL
XFILL_4__7218_ gnd vdd FILL
X_15802_ _15802_/A _14341_/Y _14338_/Y _15802_/D gnd _15803_/B vdd OAI22X1
XFILL_4__8198_ gnd vdd FILL
XFILL_2__9021_ gnd vdd FILL
XFILL_4__11180_ gnd vdd FILL
XFILL_3__10930_ gnd vdd FILL
XFILL_1__10020_ gnd vdd FILL
X_13994_ _13994_/A gnd _13995_/D vdd INVX1
XFILL_2_BUFX2_insert231 gnd vdd FILL
XFILL_2_BUFX2_insert242 gnd vdd FILL
XFILL_0__10750_ gnd vdd FILL
XFILL_2_BUFX2_insert253 gnd vdd FILL
XFILL_4__10131_ gnd vdd FILL
X_15733_ _15078_/Y _9063_/Q _9191_/Q _15079_/Y gnd _15733_/Y vdd AOI22X1
XFILL_2_BUFX2_insert264 gnd vdd FILL
X_12945_ _12901_/A _7532_/CLK _8176_/R vdd _12945_/D gnd vdd DFFSR
XFILL_5__12470_ gnd vdd FILL
XFILL_2__11310_ gnd vdd FILL
XSFILL23560x38050 gnd vdd FILL
XFILL_2_BUFX2_insert275 gnd vdd FILL
XFILL_2_BUFX2_insert286 gnd vdd FILL
XFILL_2__12290_ gnd vdd FILL
XFILL_0__10681_ gnd vdd FILL
XSFILL63960x43050 gnd vdd FILL
XFILL_5__7962_ gnd vdd FILL
XFILL_2_BUFX2_insert297 gnd vdd FILL
XFILL_5__11421_ gnd vdd FILL
XFILL_3__12600_ gnd vdd FILL
XFILL_4__10062_ gnd vdd FILL
X_15664_ _8805_/Q gnd _15665_/D vdd INVX1
XFILL_1_BUFX2_insert920 gnd vdd FILL
XSFILL13800x15050 gnd vdd FILL
XFILL_3__13580_ gnd vdd FILL
X_12876_ _12874_/Y vdd _12875_/Y gnd _12876_/Y vdd OAI21X1
XFILL_2__11241_ gnd vdd FILL
XFILL_3__10792_ gnd vdd FILL
XFILL_0__12420_ gnd vdd FILL
XFILL_1_BUFX2_insert931 gnd vdd FILL
XFILL_5__6913_ gnd vdd FILL
XFILL112120x67050 gnd vdd FILL
XFILL_1__11971_ gnd vdd FILL
XFILL_1_BUFX2_insert942 gnd vdd FILL
X_14615_ _14614_/Y _14615_/B _14203_/C _14613_/Y gnd _14615_/Y vdd OAI22X1
XFILL_5__14140_ gnd vdd FILL
XFILL_1_BUFX2_insert953 gnd vdd FILL
XFILL_1_BUFX2_insert964 gnd vdd FILL
XFILL_5__7893_ gnd vdd FILL
XFILL_5__11352_ gnd vdd FILL
X_11827_ _11234_/Y _11240_/Y _11827_/C gnd _11827_/Y vdd OAI21X1
XFILL_4__14870_ gnd vdd FILL
XFILL_3__12531_ gnd vdd FILL
XFILL_2__9923_ gnd vdd FILL
XFILL_1__13710_ gnd vdd FILL
X_15595_ _15595_/A _15595_/B _15595_/C gnd _15597_/A vdd OAI21X1
XFILL_1__10922_ gnd vdd FILL
XSFILL64040x52050 gnd vdd FILL
XFILL_1_BUFX2_insert975 gnd vdd FILL
XFILL_2__11172_ gnd vdd FILL
XFILL_1_BUFX2_insert986 gnd vdd FILL
XFILL_5__9632_ gnd vdd FILL
XFILL_0__12351_ gnd vdd FILL
XFILL_1__14690_ gnd vdd FILL
XFILL_5__10303_ gnd vdd FILL
XFILL_5__6844_ gnd vdd FILL
XFILL_1_BUFX2_insert997 gnd vdd FILL
XFILL_4__13821_ gnd vdd FILL
X_14546_ _14546_/A _14545_/Y gnd _14546_/Y vdd NOR2X1
XFILL_5__14071_ gnd vdd FILL
X_11758_ _11037_/Y _11758_/B gnd _11758_/Y vdd NOR2X1
XFILL_2__10123_ gnd vdd FILL
XFILL_3__12462_ gnd vdd FILL
XFILL_3__15250_ gnd vdd FILL
XFILL_5__11283_ gnd vdd FILL
XBUFX2_insert230 _11228_/Y gnd _11682_/B vdd BUFX2
XFILL_1__13641_ gnd vdd FILL
XFILL_0__11302_ gnd vdd FILL
XFILL_2__9854_ gnd vdd FILL
XFILL_2__15980_ gnd vdd FILL
XFILL_0__15070_ gnd vdd FILL
XBUFX2_insert241 _15065_/Y gnd _15392_/B vdd BUFX2
XFILL_5__13022_ gnd vdd FILL
XBUFX2_insert252 _10922_/Y gnd _15338_/C vdd BUFX2
X_10709_ _10709_/A _10615_/B _10708_/Y gnd _10709_/Y vdd OAI21X1
XFILL_0__12282_ gnd vdd FILL
XFILL_3__14201_ gnd vdd FILL
XFILL_6__12573_ gnd vdd FILL
XFILL_5__10234_ gnd vdd FILL
XFILL_3__11413_ gnd vdd FILL
XBUFX2_insert263 _11225_/Y gnd _11226_/B vdd BUFX2
X_14477_ _9067_/Q gnd _14477_/Y vdd INVX1
XBUFX2_insert274 _13364_/Y gnd _10700_/B vdd BUFX2
XFILL_4__13752_ gnd vdd FILL
XSFILL43880x10050 gnd vdd FILL
X_11689_ _11678_/Y _11679_/Y _11689_/C gnd _11689_/Y vdd AOI21X1
XFILL_4__10964_ gnd vdd FILL
XFILL_3__15181_ gnd vdd FILL
XFILL_3__12393_ gnd vdd FILL
XFILL_0__14021_ gnd vdd FILL
XFILL_2__10054_ gnd vdd FILL
XFILL_2__14931_ gnd vdd FILL
XFILL_1__16360_ gnd vdd FILL
XBUFX2_insert285 _15003_/Y gnd _16306_/C vdd BUFX2
XFILL_2__6997_ gnd vdd FILL
XFILL_2__9785_ gnd vdd FILL
XFILL_5__8514_ gnd vdd FILL
XFILL_1__13572_ gnd vdd FILL
XFILL_0__11233_ gnd vdd FILL
XFILL_0__7820_ gnd vdd FILL
XBUFX2_insert296 _13356_/Y gnd _10304_/B vdd BUFX2
X_16216_ _12767_/A _16216_/B gnd _16216_/Y vdd NAND2X1
XFILL_5_CLKBUF1_insert120 gnd vdd FILL
XFILL_1__10784_ gnd vdd FILL
XFILL_5_CLKBUF1_insert131 gnd vdd FILL
XFILL_4__12703_ gnd vdd FILL
X_13428_ _13401_/Y _13428_/B gnd _13476_/A vdd NOR2X1
XFILL_5__9494_ gnd vdd FILL
XFILL_5_CLKBUF1_insert142 gnd vdd FILL
XFILL_5__10165_ gnd vdd FILL
XFILL_1__15311_ gnd vdd FILL
XFILL_3__14132_ gnd vdd FILL
XFILL_3__11344_ gnd vdd FILL
XFILL_4__13683_ gnd vdd FILL
XFILL_1__12523_ gnd vdd FILL
XFILL_2__8736_ gnd vdd FILL
XFILL_5_CLKBUF1_insert153 gnd vdd FILL
XFILL_2__14862_ gnd vdd FILL
XFILL_5_CLKBUF1_insert164 gnd vdd FILL
XFILL_4__10895_ gnd vdd FILL
XFILL_1__16291_ gnd vdd FILL
XFILL_0__11164_ gnd vdd FILL
XSFILL84200x65050 gnd vdd FILL
XFILL_5__8445_ gnd vdd FILL
X_13359_ _13359_/A gnd _13363_/B vdd INVX1
XFILL_5_CLKBUF1_insert175 gnd vdd FILL
XFILL_4__15422_ gnd vdd FILL
XFILL_0__7751_ gnd vdd FILL
X_16147_ _16147_/A _16147_/B gnd _16153_/A vdd NOR2X1
XFILL_4__12634_ gnd vdd FILL
XFILL_5_CLKBUF1_insert186 gnd vdd FILL
XFILL_3__14063_ gnd vdd FILL
XFILL_5__14973_ gnd vdd FILL
XFILL_2__13813_ gnd vdd FILL
XFILL_3__7460_ gnd vdd FILL
XFILL_0__10115_ gnd vdd FILL
XFILL_1__15242_ gnd vdd FILL
XFILL_3__11275_ gnd vdd FILL
XFILL_5_CLKBUF1_insert197 gnd vdd FILL
XFILL_1__12454_ gnd vdd FILL
XFILL_0__15972_ gnd vdd FILL
XFILL_2__14793_ gnd vdd FILL
XFILL_0__11095_ gnd vdd FILL
XFILL_5__8376_ gnd vdd FILL
XFILL_3__13014_ gnd vdd FILL
XSFILL59000x41050 gnd vdd FILL
XFILL_5__13924_ gnd vdd FILL
XFILL_4__15353_ gnd vdd FILL
XFILL_0__7682_ gnd vdd FILL
X_16078_ _16077_/Y _16311_/A _14999_/A _14650_/D gnd _16078_/Y vdd OAI22X1
XFILL_2__7618_ gnd vdd FILL
XFILL_1__11405_ gnd vdd FILL
XFILL_2__10956_ gnd vdd FILL
XFILL_0__10046_ gnd vdd FILL
XFILL_2__13744_ gnd vdd FILL
XFILL_1__15173_ gnd vdd FILL
XFILL_0__14923_ gnd vdd FILL
XFILL_0__9421_ gnd vdd FILL
XFILL_6__13125_ gnd vdd FILL
XFILL_1__12385_ gnd vdd FILL
XFILL_2__8598_ gnd vdd FILL
XFILL_5__7327_ gnd vdd FILL
X_15029_ _12764_/A _14984_/Y gnd _15656_/B vdd NAND2X1
XFILL_4__14304_ gnd vdd FILL
XFILL_5__13855_ gnd vdd FILL
XFILL_4__11516_ gnd vdd FILL
XFILL_1__14124_ gnd vdd FILL
XFILL112200x47050 gnd vdd FILL
XFILL_3__10157_ gnd vdd FILL
XFILL_4__15284_ gnd vdd FILL
XFILL_3__9130_ gnd vdd FILL
XFILL_2__13675_ gnd vdd FILL
XFILL_4__12496_ gnd vdd FILL
XFILL_2__7549_ gnd vdd FILL
XFILL_1__11336_ gnd vdd FILL
XFILL_0__14854_ gnd vdd FILL
XFILL_2__10887_ gnd vdd FILL
XFILL_0__9352_ gnd vdd FILL
XFILL_4__14235_ gnd vdd FILL
XSFILL64120x32050 gnd vdd FILL
XSFILL88840x4050 gnd vdd FILL
XFILL_2__15414_ gnd vdd FILL
XFILL_2__12626_ gnd vdd FILL
XFILL_5__13786_ gnd vdd FILL
X_9980_ _9980_/A gnd _9980_/Y vdd INVX1
XFILL_4__11447_ gnd vdd FILL
XFILL_0__13805_ gnd vdd FILL
XFILL_1__14055_ gnd vdd FILL
XFILL_3__14965_ gnd vdd FILL
XFILL_5__10998_ gnd vdd FILL
XFILL_1__11267_ gnd vdd FILL
XFILL_2__16394_ gnd vdd FILL
XFILL_5__15525_ gnd vdd FILL
XFILL_5__7189_ gnd vdd FILL
XFILL_0__14785_ gnd vdd FILL
XFILL_5__12737_ gnd vdd FILL
XFILL_3__8012_ gnd vdd FILL
XFILL_0__11997_ gnd vdd FILL
XFILL_0__9283_ gnd vdd FILL
X_8931_ _8931_/Q _7791_/CLK _9711_/R vdd _8931_/D gnd vdd DFFSR
XFILL_2__9219_ gnd vdd FILL
XFILL_4__14166_ gnd vdd FILL
XFILL_1__13006_ gnd vdd FILL
XFILL_3__13916_ gnd vdd FILL
XFILL_2__15345_ gnd vdd FILL
XFILL_4__11378_ gnd vdd FILL
XFILL_0__13736_ gnd vdd FILL
XFILL_3__14896_ gnd vdd FILL
XFILL_0__10948_ gnd vdd FILL
XSFILL53960x75050 gnd vdd FILL
XFILL_1__11198_ gnd vdd FILL
XFILL_0__8234_ gnd vdd FILL
XFILL_4__13117_ gnd vdd FILL
XFILL_5__15456_ gnd vdd FILL
XFILL_2__11508_ gnd vdd FILL
X_8862_ _8854_/B _9246_/B gnd _8862_/Y vdd NAND2X1
XFILL_3__13847_ gnd vdd FILL
XFILL_4__14097_ gnd vdd FILL
XFILL_2__15276_ gnd vdd FILL
XFILL_1__10149_ gnd vdd FILL
XFILL_2__12488_ gnd vdd FILL
XFILL_6__9741_ gnd vdd FILL
XFILL_0__13667_ gnd vdd FILL
XFILL_5__14407_ gnd vdd FILL
XSFILL28760x51050 gnd vdd FILL
XFILL_0__10879_ gnd vdd FILL
X_7813_ _7813_/A gnd _7815_/A vdd INVX1
XFILL_5__11619_ gnd vdd FILL
XFILL_5__15387_ gnd vdd FILL
XFILL_2__14227_ gnd vdd FILL
X_8793_ _8793_/Q _9817_/CLK _8942_/R vdd _8705_/Y gnd vdd DFFSR
XFILL_0__15406_ gnd vdd FILL
XFILL_5__12599_ gnd vdd FILL
XFILL_2__11439_ gnd vdd FILL
XFILL_0__12618_ gnd vdd FILL
XFILL_3__13778_ gnd vdd FILL
XFILL_0__7116_ gnd vdd FILL
XFILL_0__16386_ gnd vdd FILL
XFILL_1__14957_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1082 gnd vdd FILL
XFILL_0__13598_ gnd vdd FILL
XFILL_5__14338_ gnd vdd FILL
X_7744_ _7744_/A _7744_/B _7743_/Y gnd _7790_/D vdd OAI21X1
XFILL_3__15517_ gnd vdd FILL
XFILL_0__8096_ gnd vdd FILL
XFILL_3__12729_ gnd vdd FILL
XFILL_2__14158_ gnd vdd FILL
XFILL_6__13889_ gnd vdd FILL
XFILL_3__8914_ gnd vdd FILL
XFILL_0__15337_ gnd vdd FILL
XSFILL8680x49050 gnd vdd FILL
XFILL_1__13908_ gnd vdd FILL
XFILL_3__9894_ gnd vdd FILL
XFILL_1__14888_ gnd vdd FILL
XFILL_6__15628_ gnd vdd FILL
XFILL_0__7047_ gnd vdd FILL
XSFILL33880x42050 gnd vdd FILL
XFILL_2__13109_ gnd vdd FILL
XFILL_5__14269_ gnd vdd FILL
XFILL_3__15448_ gnd vdd FILL
X_7675_ _7675_/A _7723_/B _7674_/Y gnd _7675_/Y vdd OAI21X1
XSFILL105320x79050 gnd vdd FILL
XFILL_1__13839_ gnd vdd FILL
XFILL_3__8845_ gnd vdd FILL
XFILL_4__14999_ gnd vdd FILL
XFILL_2__14089_ gnd vdd FILL
XFILL_5__16008_ gnd vdd FILL
XFILL_0__15268_ gnd vdd FILL
X_9414_ _9414_/A _9398_/A _9414_/C gnd _9456_/D vdd OAI21X1
XFILL_1__7860_ gnd vdd FILL
XFILL_3__15379_ gnd vdd FILL
XFILL_0__14219_ gnd vdd FILL
XFILL_3__8776_ gnd vdd FILL
XFILL_0__15199_ gnd vdd FILL
X_9345_ _9345_/A _9359_/A _9345_/C gnd _9433_/D vdd OAI21X1
XFILL_6__8485_ gnd vdd FILL
XFILL_0__8998_ gnd vdd FILL
XFILL_4_BUFX2_insert304 gnd vdd FILL
XFILL_1__15509_ gnd vdd FILL
XFILL_3__7727_ gnd vdd FILL
XFILL_6__7436_ gnd vdd FILL
XSFILL49000x73050 gnd vdd FILL
XFILL_4_BUFX2_insert315 gnd vdd FILL
XFILL_4_BUFX2_insert326 gnd vdd FILL
XFILL_1__9530_ gnd vdd FILL
XFILL_0__7949_ gnd vdd FILL
X_9276_ _9277_/B _8764_/B gnd _9277_/C vdd NAND2X1
XFILL_4_BUFX2_insert337 gnd vdd FILL
XFILL_4_BUFX2_insert348 gnd vdd FILL
XFILL_4_BUFX2_insert359 gnd vdd FILL
X_8227_ _8293_/Q gnd _8227_/Y vdd INVX1
XSFILL28840x31050 gnd vdd FILL
XSFILL28040x12050 gnd vdd FILL
XFILL_4__9170_ gnd vdd FILL
XFILL_3__7589_ gnd vdd FILL
XSFILL54120x64050 gnd vdd FILL
XFILL_0__9619_ gnd vdd FILL
X_8158_ _8158_/Q _8025_/CLK _9566_/R vdd _8158_/D gnd vdd DFFSR
XFILL_1__9392_ gnd vdd FILL
XFILL_4__8121_ gnd vdd FILL
X_7109_ _7064_/A _8005_/B gnd _7109_/Y vdd NAND2X1
XFILL_1__8343_ gnd vdd FILL
X_8089_ _8089_/A _8118_/A _8089_/C gnd _8161_/D vdd OAI21X1
XFILL_3__9259_ gnd vdd FILL
XFILL_1__8274_ gnd vdd FILL
XSFILL18760x83050 gnd vdd FILL
XFILL_1__7225_ gnd vdd FILL
XSFILL99640x79050 gnd vdd FILL
X_10991_ _10988_/Y _10990_/Y gnd _10991_/Y vdd NOR2X1
XSFILL34040x31050 gnd vdd FILL
X_12730_ _12728_/Y _12762_/A _12730_/C gnd _12802_/D vdd OAI21X1
XFILL_1_BUFX2_insert227 gnd vdd FILL
XFILL_1_BUFX2_insert238 gnd vdd FILL
XFILL_4__8954_ gnd vdd FILL
X_12661_ vdd memoryOutData[31] gnd _12661_/Y vdd NAND2X1
XFILL_1_BUFX2_insert249 gnd vdd FILL
XFILL_1__7087_ gnd vdd FILL
X_14400_ _14400_/A _14399_/Y _14400_/C gnd _14401_/B vdd NAND3X1
X_11612_ _11612_/A _11611_/Y gnd _11613_/A vdd NOR2X1
XFILL_0_BUFX2_insert905 gnd vdd FILL
XFILL_4__8885_ gnd vdd FILL
X_12592_ vdd memoryOutData[8] gnd _12593_/C vdd NAND2X1
X_15380_ _9438_/Q _15380_/B _15380_/C _9870_/A gnd _15381_/B vdd AOI22X1
XFILL_0_BUFX2_insert916 gnd vdd FILL
XSFILL38120x77050 gnd vdd FILL
XFILL_2__6920_ gnd vdd FILL
XSFILL28920x11050 gnd vdd FILL
XFILL_0_BUFX2_insert927 gnd vdd FILL
XFILL_4__7836_ gnd vdd FILL
XFILL_0_BUFX2_insert938 gnd vdd FILL
XFILL_0_BUFX2_insert949 gnd vdd FILL
X_14331_ _14327_/Y _14331_/B gnd _14331_/Y vdd NOR2X1
X_11543_ _11571_/A _11543_/B _11543_/C gnd _11549_/A vdd NAND3X1
XFILL_2__6851_ gnd vdd FILL
X_14262_ _14262_/A _14344_/B _13865_/B _7910_/Q gnd _14263_/B vdd AOI22X1
X_11474_ _11324_/Y gnd _11475_/C vdd INVX1
XFILL_4__9506_ gnd vdd FILL
XFILL_1__7989_ gnd vdd FILL
X_13213_ _13213_/A gnd _13219_/B vdd INVX2
X_16001_ _10043_/A gnd _16002_/D vdd INVX1
X_10425_ _10426_/B _9657_/B gnd _10425_/Y vdd NAND2X1
X_14193_ _14193_/A _14193_/B gnd _14193_/Y vdd NOR2X1
XSFILL8440x11050 gnd vdd FILL
XFILL_4__7698_ gnd vdd FILL
XFILL_1__9728_ gnd vdd FILL
XFILL_2__8521_ gnd vdd FILL
XFILL_4__10680_ gnd vdd FILL
XSFILL18840x63050 gnd vdd FILL
XFILL_5__8230_ gnd vdd FILL
X_13144_ _13142_/Y _13153_/B _13144_/C gnd _13196_/D vdd OAI21X1
X_10356_ _14885_/A _7274_/CLK _9332_/R vdd _10356_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert860 gnd vdd FILL
XFILL_5__11970_ gnd vdd FILL
XFILL_2__10810_ gnd vdd FILL
XFILL_3__11060_ gnd vdd FILL
XFILL_1__9659_ gnd vdd FILL
XFILL_2__8452_ gnd vdd FILL
XFILL_4_BUFX2_insert871 gnd vdd FILL
XFILL_4_BUFX2_insert882 gnd vdd FILL
XFILL_2__11790_ gnd vdd FILL
XFILL_4_BUFX2_insert893 gnd vdd FILL
XFILL_4__9368_ gnd vdd FILL
XFILL_5__10921_ gnd vdd FILL
XSFILL99320x61050 gnd vdd FILL
XFILL_3__10011_ gnd vdd FILL
X_13075_ _6898_/A _8560_/CLK _9313_/R vdd _13075_/D gnd vdd DFFSR
XFILL_4__12350_ gnd vdd FILL
X_10287_ _14359_/D gnd _10287_/Y vdd INVX1
XFILL_2__8383_ gnd vdd FILL
XFILL_4__8319_ gnd vdd FILL
XFILL_0__11920_ gnd vdd FILL
XFILL_1__12170_ gnd vdd FILL
XFILL_5__7112_ gnd vdd FILL
XFILL_5__8092_ gnd vdd FILL
X_12026_ _12026_/A _12024_/Y _12025_/Y gnd _12026_/Y vdd NAND3X1
XFILL_5__13640_ gnd vdd FILL
XFILL_4__9299_ gnd vdd FILL
XFILL_4__11301_ gnd vdd FILL
XFILL_2__7334_ gnd vdd FILL
XSFILL38760x14050 gnd vdd FILL
XFILL_2__13460_ gnd vdd FILL
XSFILL109720x44050 gnd vdd FILL
XFILL_4__12281_ gnd vdd FILL
XFILL_1__11121_ gnd vdd FILL
XSFILL63960x7050 gnd vdd FILL
XFILL112280x21050 gnd vdd FILL
XFILL_5__7043_ gnd vdd FILL
XSFILL64040x47050 gnd vdd FILL
XFILL_2__10672_ gnd vdd FILL
XFILL_0__11851_ gnd vdd FILL
XFILL_4__14020_ gnd vdd FILL
XFILL_2__12411_ gnd vdd FILL
XFILL_5__13571_ gnd vdd FILL
XFILL_4__11232_ gnd vdd FILL
XSFILL24040x63050 gnd vdd FILL
XFILL_3__14750_ gnd vdd FILL
XFILL_5__10783_ gnd vdd FILL
XFILL_2__13391_ gnd vdd FILL
XFILL_3__11962_ gnd vdd FILL
XFILL112280x6050 gnd vdd FILL
XFILL_1__11052_ gnd vdd FILL
XFILL_0__10802_ gnd vdd FILL
XFILL_0__14570_ gnd vdd FILL
XFILL_5__15310_ gnd vdd FILL
XFILL_5__12522_ gnd vdd FILL
XFILL_0__11782_ gnd vdd FILL
XFILL_6__14861_ gnd vdd FILL
XFILL_5__16290_ gnd vdd FILL
XFILL_2__9004_ gnd vdd FILL
XFILL_4__11163_ gnd vdd FILL
XFILL_2__15130_ gnd vdd FILL
XFILL_3__13701_ gnd vdd FILL
XFILL_3__10913_ gnd vdd FILL
X_13977_ _8087_/A gnd _15498_/D vdd INVX1
XFILL_2__12342_ gnd vdd FILL
XFILL_1__10003_ gnd vdd FILL
XFILL_2__7196_ gnd vdd FILL
XFILL_3__14681_ gnd vdd FILL
XFILL_0__13521_ gnd vdd FILL
XSFILL3480x54050 gnd vdd FILL
XFILL_3__11893_ gnd vdd FILL
XFILL_1__15860_ gnd vdd FILL
XFILL_6__13812_ gnd vdd FILL
X_15716_ _7398_/Q gnd _15717_/A vdd INVX1
XFILL_4__10114_ gnd vdd FILL
XFILL_5__15241_ gnd vdd FILL
XFILL_5__8994_ gnd vdd FILL
XFILL_5__12453_ gnd vdd FILL
X_12928_ _12928_/Q _8180_/CLK _7391_/R vdd _12852_/Y gnd vdd DFFSR
XSFILL84760x17050 gnd vdd FILL
XFILL_3__13632_ gnd vdd FILL
XFILL_4__15971_ gnd vdd FILL
XFILL_2__15061_ gnd vdd FILL
XFILL_4__11094_ gnd vdd FILL
XFILL_0__16240_ gnd vdd FILL
XFILL_1__14811_ gnd vdd FILL
XFILL_2__12273_ gnd vdd FILL
XSFILL69160x1050 gnd vdd FILL
XFILL_0__13452_ gnd vdd FILL
XFILL_1__15791_ gnd vdd FILL
XFILL_5__7945_ gnd vdd FILL
XFILL_0__10664_ gnd vdd FILL
XFILL_5__11404_ gnd vdd FILL
XFILL_4__10045_ gnd vdd FILL
X_15647_ _16002_/A _14127_/Y _16002_/C _14125_/D gnd _15648_/B vdd OAI22X1
XFILL_2__14012_ gnd vdd FILL
XFILL_5__15172_ gnd vdd FILL
XFILL_4__14922_ gnd vdd FILL
XFILL_1_BUFX2_insert750 gnd vdd FILL
XFILL_5__12384_ gnd vdd FILL
X_12859_ _12859_/A gnd _12859_/Y vdd INVX1
XFILL_3__16351_ gnd vdd FILL
XFILL_2__11224_ gnd vdd FILL
XFILL_0__12403_ gnd vdd FILL
XFILL_3__10775_ gnd vdd FILL
XFILL_1_BUFX2_insert761 gnd vdd FILL
XFILL_1__14742_ gnd vdd FILL
XFILL_3__13563_ gnd vdd FILL
XSFILL44200x76050 gnd vdd FILL
XFILL_0__16171_ gnd vdd FILL
XFILL_1__11954_ gnd vdd FILL
XFILL_3__6960_ gnd vdd FILL
XFILL_1_BUFX2_insert772 gnd vdd FILL
XFILL_5__14123_ gnd vdd FILL
XFILL_0__13383_ gnd vdd FILL
XFILL_1_BUFX2_insert783 gnd vdd FILL
XFILL_3__15302_ gnd vdd FILL
XFILL_6__13674_ gnd vdd FILL
XSFILL59000x36050 gnd vdd FILL
XFILL_5__7876_ gnd vdd FILL
XFILL_5__11335_ gnd vdd FILL
XFILL_4__14853_ gnd vdd FILL
XFILL_1_BUFX2_insert794 gnd vdd FILL
XFILL_3__12514_ gnd vdd FILL
XFILL_2__9906_ gnd vdd FILL
X_15578_ _15813_/C _14111_/A _15578_/C _16155_/D gnd _15579_/A vdd OAI22X1
XFILL_1__10905_ gnd vdd FILL
XFILL_2__11155_ gnd vdd FILL
XFILL_0__15122_ gnd vdd FILL
XFILL_3__16282_ gnd vdd FILL
XFILL_5__9615_ gnd vdd FILL
XFILL_3__6891_ gnd vdd FILL
XSFILL99400x41050 gnd vdd FILL
XFILL_3__13494_ gnd vdd FILL
XFILL_0__12334_ gnd vdd FILL
XFILL_1__14673_ gnd vdd FILL
XFILL_6__15413_ gnd vdd FILL
XFILL_1__11885_ gnd vdd FILL
XFILL_4_BUFX2_insert10 gnd vdd FILL
XFILL_4__13804_ gnd vdd FILL
XFILL_4_BUFX2_insert21 gnd vdd FILL
XFILL_5__14054_ gnd vdd FILL
X_14529_ _15931_/A _14389_/B _13865_/B _7916_/Q gnd _14529_/Y vdd AOI22X1
X_7460_ _7460_/A _8356_/B gnd _7461_/C vdd NAND2X1
XFILL_3__15233_ gnd vdd FILL
XFILL_2__10106_ gnd vdd FILL
XFILL_5__11266_ gnd vdd FILL
XFILL_3__8630_ gnd vdd FILL
XFILL_1__13624_ gnd vdd FILL
XFILL_3__12445_ gnd vdd FILL
XFILL_1__16412_ gnd vdd FILL
XFILL_4_BUFX2_insert32 gnd vdd FILL
XFILL_4__14784_ gnd vdd FILL
XFILL_4_BUFX2_insert43 gnd vdd FILL
XFILL_0__15053_ gnd vdd FILL
XFILL_4__11996_ gnd vdd FILL
XFILL_2__15963_ gnd vdd FILL
XFILL_2__11086_ gnd vdd FILL
XFILL_1__10836_ gnd vdd FILL
XFILL_5__9546_ gnd vdd FILL
XFILL_0__12265_ gnd vdd FILL
XFILL_5__13005_ gnd vdd FILL
XSFILL109800x24050 gnd vdd FILL
XFILL_4_BUFX2_insert54 gnd vdd FILL
XSFILL48840x79050 gnd vdd FILL
XFILL_4_BUFX2_insert65 gnd vdd FILL
XSFILL64120x27050 gnd vdd FILL
XFILL_0__8852_ gnd vdd FILL
XFILL_4__13735_ gnd vdd FILL
XFILL_4__10947_ gnd vdd FILL
XFILL_2__10037_ gnd vdd FILL
XFILL_4_BUFX2_insert76 gnd vdd FILL
XFILL_1__16343_ gnd vdd FILL
XFILL_3__12376_ gnd vdd FILL
XFILL_0__14004_ gnd vdd FILL
XFILL_3__15164_ gnd vdd FILL
XFILL_5__11197_ gnd vdd FILL
X_7391_ _7391_/Q _8297_/CLK _7391_/R vdd _7315_/Y gnd vdd DFFSR
XFILL_2__14914_ gnd vdd FILL
XFILL_2__9768_ gnd vdd FILL
XFILL_4_BUFX2_insert87 gnd vdd FILL
XFILL_1__13555_ gnd vdd FILL
XFILL_0__11216_ gnd vdd FILL
XFILL_1__10767_ gnd vdd FILL
XFILL_2__15894_ gnd vdd FILL
XFILL_4_BUFX2_insert98 gnd vdd FILL
XFILL_6__11507_ gnd vdd FILL
XFILL_0__12196_ gnd vdd FILL
XFILL_5__9477_ gnd vdd FILL
XFILL_0__7803_ gnd vdd FILL
XFILL_6__15275_ gnd vdd FILL
X_9130_ _9116_/B _7594_/B gnd _9130_/Y vdd NAND2X1
XFILL_5__10148_ gnd vdd FILL
XFILL_0__8783_ gnd vdd FILL
XFILL_3__14115_ gnd vdd FILL
XFILL_2__8719_ gnd vdd FILL
XFILL_1__12506_ gnd vdd FILL
XFILL_4__13666_ gnd vdd FILL
XFILL_3__11327_ gnd vdd FILL
XFILL_2__14845_ gnd vdd FILL
XFILL_4__10878_ gnd vdd FILL
XFILL_3__15095_ gnd vdd FILL
XFILL_1__16274_ gnd vdd FILL
XFILL_1__13486_ gnd vdd FILL
XFILL_3__8492_ gnd vdd FILL
XFILL_0__11147_ gnd vdd FILL
XFILL_4__15405_ gnd vdd FILL
XFILL_1__10698_ gnd vdd FILL
XFILL_4__12617_ gnd vdd FILL
XFILL_0__7734_ gnd vdd FILL
X_9061_ _8995_/A _7269_/CLK _9061_/R vdd _8997_/Y gnd vdd DFFSR
XFILL_4__16385_ gnd vdd FILL
XFILL_1__15225_ gnd vdd FILL
XFILL_3__14046_ gnd vdd FILL
XSFILL3560x34050 gnd vdd FILL
XFILL_3__11258_ gnd vdd FILL
XFILL_5__14956_ gnd vdd FILL
XFILL_4__13597_ gnd vdd FILL
XFILL_1__12437_ gnd vdd FILL
XFILL_3__7443_ gnd vdd FILL
XFILL_2__11988_ gnd vdd FILL
XFILL_0__15955_ gnd vdd FILL
XFILL_2_BUFX2_insert1004 gnd vdd FILL
XFILL_0__11078_ gnd vdd FILL
XFILL_2__14776_ gnd vdd FILL
XFILL_5__8359_ gnd vdd FILL
X_8012_ _8012_/A _7997_/B _8011_/Y gnd _8012_/Y vdd OAI21X1
XFILL_2_BUFX2_insert1015 gnd vdd FILL
XFILL_4__15336_ gnd vdd FILL
XFILL_2_BUFX2_insert1026 gnd vdd FILL
XSFILL28760x46050 gnd vdd FILL
XFILL_5__13907_ gnd vdd FILL
XFILL_6__11369_ gnd vdd FILL
XSFILL53560x72050 gnd vdd FILL
XFILL_2_BUFX2_insert1037 gnd vdd FILL
XFILL_5__14887_ gnd vdd FILL
XFILL_3__7374_ gnd vdd FILL
XFILL_2_BUFX2_insert1048 gnd vdd FILL
XFILL_1__15156_ gnd vdd FILL
XFILL_3__11189_ gnd vdd FILL
XFILL_2__13727_ gnd vdd FILL
XFILL_0__14906_ gnd vdd FILL
XFILL_2__10939_ gnd vdd FILL
XFILL_1__12368_ gnd vdd FILL
XFILL_0__10029_ gnd vdd FILL
XFILL_0__9404_ gnd vdd FILL
XFILL_2_BUFX2_insert1059 gnd vdd FILL
XFILL_0__15886_ gnd vdd FILL
XFILL_6__14088_ gnd vdd FILL
XFILL_5__13838_ gnd vdd FILL
XFILL_3__9113_ gnd vdd FILL
XFILL_0__7596_ gnd vdd FILL
XFILL_1__14107_ gnd vdd FILL
XFILL_4__15267_ gnd vdd FILL
XFILL_4__12479_ gnd vdd FILL
XFILL_1__11319_ gnd vdd FILL
XFILL_0__14837_ gnd vdd FILL
XFILL_3__15997_ gnd vdd FILL
XFILL_2__13658_ gnd vdd FILL
XFILL_1__15087_ gnd vdd FILL
XFILL_1__12299_ gnd vdd FILL
XFILL_4__14218_ gnd vdd FILL
XFILL_0__9335_ gnd vdd FILL
XSFILL3560x3050 gnd vdd FILL
X_9963_ _9963_/Q _9963_/CLK _9963_/R vdd _9911_/Y gnd vdd DFFSR
XFILL_5__13769_ gnd vdd FILL
XFILL_4__15198_ gnd vdd FILL
XFILL_2__12609_ gnd vdd FILL
XFILL_1__14038_ gnd vdd FILL
XSFILL33880x37050 gnd vdd FILL
XFILL_3__14948_ gnd vdd FILL
XFILL_3__9044_ gnd vdd FILL
XFILL_2__13589_ gnd vdd FILL
XFILL_2__16377_ gnd vdd FILL
XFILL_0__14768_ gnd vdd FILL
XFILL_5__15508_ gnd vdd FILL
XFILL_0__9266_ gnd vdd FILL
X_8914_ _8912_/Y _8902_/B _8914_/C gnd _8948_/D vdd OAI21X1
XFILL_4__14149_ gnd vdd FILL
XFILL_2__15328_ gnd vdd FILL
X_9894_ _9958_/Q gnd _9896_/A vdd INVX1
XFILL_3__14879_ gnd vdd FILL
XFILL_0__13719_ gnd vdd FILL
XFILL_0__8217_ gnd vdd FILL
XFILL_0_BUFX2_insert1030 gnd vdd FILL
XFILL_0_BUFX2_insert1041 gnd vdd FILL
XFILL_0__14699_ gnd vdd FILL
X_8845_ _8845_/A _8845_/B _8844_/Y gnd _8845_/Y vdd OAI21X1
XFILL_0_BUFX2_insert1052 gnd vdd FILL
XFILL_5__15439_ gnd vdd FILL
XFILL_2__15259_ gnd vdd FILL
XFILL_0_BUFX2_insert1063 gnd vdd FILL
XSFILL89960x30050 gnd vdd FILL
XSFILL89160x11050 gnd vdd FILL
XFILL_0_BUFX2_insert1085 gnd vdd FILL
XFILL_1__15989_ gnd vdd FILL
XFILL_0__8148_ gnd vdd FILL
X_8776_ _8788_/A _8008_/B gnd _8776_/Y vdd NAND2X1
XFILL_6_BUFX2_insert955 gnd vdd FILL
XFILL_0__16369_ gnd vdd FILL
XSFILL3640x14050 gnd vdd FILL
XFILL_0__8079_ gnd vdd FILL
XSFILL109560x79050 gnd vdd FILL
XFILL_6_BUFX2_insert966 gnd vdd FILL
XSFILL110040x67050 gnd vdd FILL
X_7727_ _7727_/A gnd _7729_/A vdd INVX1
XFILL_1__8961_ gnd vdd FILL
XFILL_3__9877_ gnd vdd FILL
XSFILL28840x26050 gnd vdd FILL
XSFILL54920x78050 gnd vdd FILL
XSFILL54120x59050 gnd vdd FILL
X_7658_ _7658_/Q _7274_/CLK _7274_/R vdd _7604_/Y gnd vdd DFFSR
XFILL_1__8892_ gnd vdd FILL
XFILL_4__7621_ gnd vdd FILL
XFILL_3__8828_ gnd vdd FILL
XFILL_1__7843_ gnd vdd FILL
X_7589_ _7589_/A _7568_/B _7589_/C gnd _7589_/Y vdd OAI21X1
XSFILL95160x30050 gnd vdd FILL
XFILL_4__7552_ gnd vdd FILL
XFILL_3__8759_ gnd vdd FILL
XFILL_4_BUFX2_insert101 gnd vdd FILL
XSFILL33960x17050 gnd vdd FILL
X_9328_ _9284_/A _9328_/CLK _7152_/R vdd _9328_/D gnd vdd DFFSR
X_10210_ _10138_/A _8680_/CLK _8034_/R vdd _10210_/D gnd vdd DFFSR
XFILL_4__7483_ gnd vdd FILL
X_11190_ _11189_/Y gnd _11191_/A vdd INVX2
XFILL_1__9513_ gnd vdd FILL
X_9259_ _9259_/A _9208_/B _9258_/Y gnd _9259_/Y vdd OAI21X1
XFILL_4__9222_ gnd vdd FILL
X_10141_ _14081_/A gnd _10143_/A vdd INVX1
XSFILL33800x81050 gnd vdd FILL
XFILL_3_BUFX2_insert801 gnd vdd FILL
XFILL_3_BUFX2_insert812 gnd vdd FILL
XFILL_3_BUFX2_insert823 gnd vdd FILL
XFILL_3_BUFX2_insert834 gnd vdd FILL
XFILL_4__9153_ gnd vdd FILL
XFILL_3_BUFX2_insert845 gnd vdd FILL
X_10072_ _9980_/A _8663_/CLK _8664_/R vdd _9982_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert856 gnd vdd FILL
XFILL_4__8104_ gnd vdd FILL
XFILL_1__9375_ gnd vdd FILL
XFILL_3_BUFX2_insert867 gnd vdd FILL
XFILL_3_BUFX2_insert878 gnd vdd FILL
XSFILL109640x59050 gnd vdd FILL
XFILL_3_BUFX2_insert889 gnd vdd FILL
X_13900_ _13900_/A gnd _13902_/D vdd INVX1
XFILL_4__9084_ gnd vdd FILL
X_14880_ _14879_/Y _14880_/B gnd _14881_/B vdd NOR2X1
XFILL_1__8326_ gnd vdd FILL
X_13831_ _8459_/A gnd _13833_/B vdd INVX1
XFILL_2__7050_ gnd vdd FILL
XFILL_1__8257_ gnd vdd FILL
XFILL_1__7208_ gnd vdd FILL
X_10974_ _10972_/Y vdd _10974_/C gnd _10984_/D vdd OAI21X1
X_13762_ _7004_/Q gnd _13763_/A vdd INVX1
XFILL_1__8188_ gnd vdd FILL
X_15501_ _15978_/C _8545_/Q _8215_/A _16014_/C gnd _15504_/A vdd AOI22X1
X_12713_ _12713_/A gnd _12713_/Y vdd INVX1
XFILL_4__9986_ gnd vdd FILL
X_13693_ _13691_/Y _13879_/B _14555_/C _15279_/C gnd _13697_/A vdd OAI22X1
XSFILL33720x5050 gnd vdd FILL
XFILL_5__7730_ gnd vdd FILL
XSFILL18840x58050 gnd vdd FILL
X_15432_ _15431_/Y _15432_/B gnd _15432_/Y vdd NOR2X1
X_12644_ _12644_/A vdd _12644_/C gnd _12688_/D vdd OAI21X1
XFILL_3__10560_ gnd vdd FILL
XFILL_0_BUFX2_insert702 gnd vdd FILL
XFILL_2__7952_ gnd vdd FILL
XFILL_0_BUFX2_insert713 gnd vdd FILL
XFILL_0__10380_ gnd vdd FILL
XFILL_0_BUFX2_insert724 gnd vdd FILL
XFILL_0_CLKBUF1_insert150 gnd vdd FILL
XFILL_4__8868_ gnd vdd FILL
XFILL_5__11120_ gnd vdd FILL
XFILL_0_BUFX2_insert735 gnd vdd FILL
X_12575_ _12575_/A vdd _12574_/Y gnd _12665_/D vdd OAI21X1
X_15363_ _13820_/Y _15920_/B _15920_/C _13821_/D gnd _15367_/B vdd OAI22X1
XSFILL99320x56050 gnd vdd FILL
XFILL_0_CLKBUF1_insert161 gnd vdd FILL
XSFILL59080x10050 gnd vdd FILL
XFILL_2__6903_ gnd vdd FILL
XFILL_0_BUFX2_insert746 gnd vdd FILL
XFILL_0_CLKBUF1_insert172 gnd vdd FILL
XFILL_4__11850_ gnd vdd FILL
XFILL_5__9400_ gnd vdd FILL
XFILL_0_BUFX2_insert757 gnd vdd FILL
XFILL_0_CLKBUF1_insert183 gnd vdd FILL
XFILL_3__10491_ gnd vdd FILL
XFILL_0_CLKBUF1_insert194 gnd vdd FILL
XFILL_0_BUFX2_insert768 gnd vdd FILL
XFILL_4__7819_ gnd vdd FILL
XFILL_2__7883_ gnd vdd FILL
XFILL_1__11670_ gnd vdd FILL
XSFILL59320x72050 gnd vdd FILL
X_14314_ _7656_/Q _14185_/B _14214_/C _15797_/A gnd _14322_/B vdd AOI22X1
XFILL_0_BUFX2_insert779 gnd vdd FILL
XFILL_5__7592_ gnd vdd FILL
XFILL_3__12230_ gnd vdd FILL
XFILL_4__10801_ gnd vdd FILL
X_11526_ _11542_/B _11525_/Y _11542_/A gnd _11527_/A vdd AOI21X1
XFILL_5__11051_ gnd vdd FILL
X_15294_ _15293_/Y _15294_/B gnd _15294_/Y vdd NAND2X1
XFILL_2__9622_ gnd vdd FILL
XFILL_1__10621_ gnd vdd FILL
XFILL_4__11781_ gnd vdd FILL
XFILL_2__12960_ gnd vdd FILL
XFILL_0__12050_ gnd vdd FILL
XFILL112280x16050 gnd vdd FILL
XFILL_6__12341_ gnd vdd FILL
XFILL_5__10002_ gnd vdd FILL
X_14245_ _14245_/A gnd _14246_/D vdd INVX1
XFILL_4__13520_ gnd vdd FILL
X_11457_ _11457_/A _11420_/Y _11456_/Y gnd _12101_/A vdd NAND3X1
XFILL_3__12161_ gnd vdd FILL
XFILL_1__13340_ gnd vdd FILL
XFILL_2__11911_ gnd vdd FILL
XFILL_0__11001_ gnd vdd FILL
XFILL_2__9553_ gnd vdd FILL
XFILL_1__10552_ gnd vdd FILL
XFILL_2__12891_ gnd vdd FILL
X_10408_ _10408_/A _10423_/B _10407_/Y gnd _10408_/Y vdd OAI21X1
XFILL_6__15060_ gnd vdd FILL
XFILL_5__9262_ gnd vdd FILL
X_14176_ _14175_/Y _13868_/B gnd _14179_/A vdd NOR2X1
XFILL_5__14810_ gnd vdd FILL
XFILL_3__11112_ gnd vdd FILL
XFILL_2__8504_ gnd vdd FILL
XFILL_4__13451_ gnd vdd FILL
XFILL_5__15790_ gnd vdd FILL
X_11388_ _11387_/Y _11388_/B gnd _11389_/B vdd NOR2X1
XFILL_2__14630_ gnd vdd FILL
XFILL_4__10663_ gnd vdd FILL
XFILL_3__12092_ gnd vdd FILL
XSFILL79240x23050 gnd vdd FILL
XFILL_2__11842_ gnd vdd FILL
XFILL_2__9484_ gnd vdd FILL
XFILL_1__13271_ gnd vdd FILL
XFILL_5__8213_ gnd vdd FILL
XFILL_4__12402_ gnd vdd FILL
X_13127_ _11935_/A gnd _13129_/A vdd INVX1
XFILL_5__14741_ gnd vdd FILL
X_10339_ _14077_/C _7530_/CLK _7523_/R vdd _10271_/Y gnd vdd DFFSR
XFILL_3__15920_ gnd vdd FILL
XFILL_4__16170_ gnd vdd FILL
XFILL_5__11953_ gnd vdd FILL
XFILL_1__15010_ gnd vdd FILL
XFILL_3__11043_ gnd vdd FILL
XFILL_4_BUFX2_insert690 gnd vdd FILL
XFILL_4__13382_ gnd vdd FILL
XFILL_1__12222_ gnd vdd FILL
XFILL_2__14561_ gnd vdd FILL
XFILL_0__15740_ gnd vdd FILL
XFILL_2__11773_ gnd vdd FILL
XFILL_0__12952_ gnd vdd FILL
XFILL_5__8144_ gnd vdd FILL
XFILL_5__10904_ gnd vdd FILL
XFILL_0__7450_ gnd vdd FILL
X_13058_ _6881_/A _8176_/CLK _8176_/R vdd _13058_/D gnd vdd DFFSR
XSFILL114440x32050 gnd vdd FILL
XFILL_6__11154_ gnd vdd FILL
XFILL_4__15121_ gnd vdd FILL
XFILL_2__16300_ gnd vdd FILL
XFILL_4__12333_ gnd vdd FILL
XFILL_5__14672_ gnd vdd FILL
XFILL_5__11884_ gnd vdd FILL
XFILL_3__15851_ gnd vdd FILL
XFILL_2__13512_ gnd vdd FILL
XFILL_2__14492_ gnd vdd FILL
XFILL_0__11903_ gnd vdd FILL
XFILL_1__12153_ gnd vdd FILL
XFILL_2__8366_ gnd vdd FILL
XSFILL84360x14050 gnd vdd FILL
XFILL_0__15671_ gnd vdd FILL
X_12009_ _12009_/A _12113_/B _12113_/C gnd gnd _12010_/C vdd AOI22X1
XFILL_5__13623_ gnd vdd FILL
XFILL_5__8075_ gnd vdd FILL
XFILL_5__16411_ gnd vdd FILL
XFILL_0__12883_ gnd vdd FILL
XFILL_3__14802_ gnd vdd FILL
XFILL_4__15052_ gnd vdd FILL
XFILL_0__7381_ gnd vdd FILL
XFILL_5__10835_ gnd vdd FILL
XFILL_2__16231_ gnd vdd FILL
XFILL_2__13443_ gnd vdd FILL
XFILL_4__12264_ gnd vdd FILL
XFILL_1__11104_ gnd vdd FILL
XFILL_2__7317_ gnd vdd FILL
XFILL_0__14622_ gnd vdd FILL
XFILL_3__15782_ gnd vdd FILL
XFILL_3__7090_ gnd vdd FILL
XFILL_2__10655_ gnd vdd FILL
XFILL_1__12084_ gnd vdd FILL
XFILL_0__9120_ gnd vdd FILL
XFILL_3__12994_ gnd vdd FILL
XFILL_0__11834_ gnd vdd FILL
XSFILL69160x75050 gnd vdd FILL
XFILL_4__14003_ gnd vdd FILL
XFILL_6__10036_ gnd vdd FILL
XFILL_5__16342_ gnd vdd FILL
XFILL_5__13554_ gnd vdd FILL
XFILL_4__11215_ gnd vdd FILL
XFILL_5__10766_ gnd vdd FILL
XFILL_3__14733_ gnd vdd FILL
X_6960_ _6937_/B _6960_/B gnd _6961_/C vdd NAND2X1
XFILL_2__7248_ gnd vdd FILL
XFILL_1__15912_ gnd vdd FILL
XFILL_2__13374_ gnd vdd FILL
XFILL_3__11945_ gnd vdd FILL
XFILL_4__12195_ gnd vdd FILL
XFILL_2__16162_ gnd vdd FILL
XFILL_1__11035_ gnd vdd FILL
XFILL_0__14553_ gnd vdd FILL
XFILL_5__12505_ gnd vdd FILL
XFILL_0__11765_ gnd vdd FILL
XFILL_5__16273_ gnd vdd FILL
XFILL_4__11146_ gnd vdd FILL
XFILL_5__13485_ gnd vdd FILL
XFILL_2__15113_ gnd vdd FILL
XFILL_2__12325_ gnd vdd FILL
XFILL_2__7179_ gnd vdd FILL
X_6891_ _6891_/A gnd memoryWriteData[21] vdd BUFX2
XFILL_2__16093_ gnd vdd FILL
XFILL_3__14664_ gnd vdd FILL
XFILL_0__13504_ gnd vdd FILL
XFILL_5__10697_ gnd vdd FILL
XFILL_3__11876_ gnd vdd FILL
XFILL_1__15843_ gnd vdd FILL
XFILL_0__8002_ gnd vdd FILL
XFILL_0__14484_ gnd vdd FILL
XFILL_5__15224_ gnd vdd FILL
X_8630_ _8589_/B _8630_/B gnd _8630_/Y vdd NAND2X1
XFILL_5__12436_ gnd vdd FILL
XFILL_0__11696_ gnd vdd FILL
XFILL_3__16403_ gnd vdd FILL
XFILL_5__8977_ gnd vdd FILL
XFILL_3__13615_ gnd vdd FILL
XFILL_6_BUFX2_insert229 gnd vdd FILL
XFILL_3__9800_ gnd vdd FILL
XFILL_0__16223_ gnd vdd FILL
XFILL_3__10827_ gnd vdd FILL
XFILL_2__15044_ gnd vdd FILL
XFILL_4__15954_ gnd vdd FILL
XFILL_2__12256_ gnd vdd FILL
XFILL_4__11077_ gnd vdd FILL
XFILL_3__14595_ gnd vdd FILL
XFILL_0__13435_ gnd vdd FILL
XFILL_0__10647_ gnd vdd FILL
XFILL_3__7992_ gnd vdd FILL
XFILL_1__12986_ gnd vdd FILL
XFILL_1__15774_ gnd vdd FILL
XFILL_5__7928_ gnd vdd FILL
XSFILL49080x42050 gnd vdd FILL
XFILL_5__15155_ gnd vdd FILL
XFILL112200x60050 gnd vdd FILL
XFILL_5__12367_ gnd vdd FILL
XFILL_3__16334_ gnd vdd FILL
X_8561_ _8519_/A _7537_/CLK _7537_/R vdd _8561_/D gnd vdd DFFSR
XFILL_4__10028_ gnd vdd FILL
XFILL_2__11207_ gnd vdd FILL
XFILL_4__14905_ gnd vdd FILL
XFILL_1_BUFX2_insert580 gnd vdd FILL
XFILL_3__9731_ gnd vdd FILL
XFILL_1_BUFX2_insert591 gnd vdd FILL
XSFILL3560x29050 gnd vdd FILL
XFILL_3__13546_ gnd vdd FILL
XFILL_4__15885_ gnd vdd FILL
XFILL_2__12187_ gnd vdd FILL
XFILL_1__11937_ gnd vdd FILL
XFILL_1__14725_ gnd vdd FILL
XFILL_3__6943_ gnd vdd FILL
XFILL_3__10758_ gnd vdd FILL
XFILL_0__16154_ gnd vdd FILL
XFILL_5_BUFX2_insert907 gnd vdd FILL
XFILL_0__13366_ gnd vdd FILL
XFILL_5__14106_ gnd vdd FILL
XFILL_5__11318_ gnd vdd FILL
X_7512_ _7420_/A _8679_/CLK _7131_/R vdd _7512_/D gnd vdd DFFSR
XFILL_0__10578_ gnd vdd FILL
XFILL_5__7859_ gnd vdd FILL
XFILL_4__14836_ gnd vdd FILL
XFILL_5_BUFX2_insert918 gnd vdd FILL
XFILL_5__15086_ gnd vdd FILL
X_8492_ _8492_/A gnd _8494_/A vdd INVX1
XFILL_5_BUFX2_insert929 gnd vdd FILL
XFILL_2__11138_ gnd vdd FILL
XSFILL114520x12050 gnd vdd FILL
XFILL_0__15105_ gnd vdd FILL
XFILL_3__16265_ gnd vdd FILL
XFILL_5__12298_ gnd vdd FILL
XFILL_3__9662_ gnd vdd FILL
XFILL_3__13477_ gnd vdd FILL
XFILL_0__12317_ gnd vdd FILL
XFILL_3__6874_ gnd vdd FILL
XFILL_1__11868_ gnd vdd FILL
XFILL_1__14656_ gnd vdd FILL
XFILL_0__16085_ gnd vdd FILL
XFILL_3__10689_ gnd vdd FILL
XFILL_0__13297_ gnd vdd FILL
XFILL_5__14037_ gnd vdd FILL
XFILL_0__8904_ gnd vdd FILL
XFILL_3__15216_ gnd vdd FILL
X_7443_ _7443_/A _7472_/A _7443_/C gnd _7519_/D vdd OAI21X1
XFILL_5__11249_ gnd vdd FILL
XSFILL94440x79050 gnd vdd FILL
XFILL_3__12428_ gnd vdd FILL
XFILL_3__8613_ gnd vdd FILL
XFILL_0__9884_ gnd vdd FILL
XFILL_4__14767_ gnd vdd FILL
XFILL_1__13607_ gnd vdd FILL
XFILL_3__16196_ gnd vdd FILL
XFILL_0__15036_ gnd vdd FILL
XSFILL28360x43050 gnd vdd FILL
XFILL_2__15946_ gnd vdd FILL
XFILL_4__11979_ gnd vdd FILL
XFILL_1__10819_ gnd vdd FILL
XFILL_2__11069_ gnd vdd FILL
XFILL_1__14587_ gnd vdd FILL
XFILL_5__9529_ gnd vdd FILL
XFILL_0__12248_ gnd vdd FILL
XFILL_3__9593_ gnd vdd FILL
XFILL_1__11799_ gnd vdd FILL
XFILL_0__8835_ gnd vdd FILL
XFILL_4__13718_ gnd vdd FILL
X_7374_ _7336_/B _8526_/B gnd _7374_/Y vdd NAND2X1
XSFILL69240x55050 gnd vdd FILL
XFILL_3__15147_ gnd vdd FILL
XFILL_3__12359_ gnd vdd FILL
XFILL_4__14698_ gnd vdd FILL
XFILL_1__16326_ gnd vdd FILL
XFILL_1__13538_ gnd vdd FILL
XFILL_2__15877_ gnd vdd FILL
XFILL_0__12179_ gnd vdd FILL
X_9113_ _9111_/Y _9164_/B _9112_/Y gnd _9185_/D vdd OAI21X1
XFILL_0__8766_ gnd vdd FILL
XFILL_4__13649_ gnd vdd FILL
XFILL_5__15988_ gnd vdd FILL
XFILL_2__14828_ gnd vdd FILL
XFILL_3__15078_ gnd vdd FILL
XFILL_1__13469_ gnd vdd FILL
XFILL_3__8475_ gnd vdd FILL
XFILL_1__16257_ gnd vdd FILL
XSFILL104440x64050 gnd vdd FILL
XSFILL39080x5050 gnd vdd FILL
XFILL_0__7717_ gnd vdd FILL
XFILL_3_BUFX2_insert108 gnd vdd FILL
X_9044_ _9044_/A _9172_/B gnd _9045_/C vdd NAND2X1
XFILL_3__14029_ gnd vdd FILL
XFILL_5__14939_ gnd vdd FILL
XFILL_1__7490_ gnd vdd FILL
XFILL_4__16368_ gnd vdd FILL
XFILL_1__15208_ gnd vdd FILL
XSFILL8680x62050 gnd vdd FILL
XFILL_3__7426_ gnd vdd FILL
XFILL_0__8697_ gnd vdd FILL
XSFILL23720x11050 gnd vdd FILL
XFILL_1__16188_ gnd vdd FILL
XFILL_2__14759_ gnd vdd FILL
XFILL_0__15938_ gnd vdd FILL
XFILL_4__15319_ gnd vdd FILL
XFILL_4__16299_ gnd vdd FILL
XCLKBUF1_insert1075 clk gnd CLKBUF1_insert182/A vdd CLKBUF1
XFILL_1__15139_ gnd vdd FILL
XSFILL89400x68050 gnd vdd FILL
XFILL_3__7357_ gnd vdd FILL
XFILL_0__15869_ gnd vdd FILL
XFILL_1__9160_ gnd vdd FILL
XFILL_2_BUFX2_insert808 gnd vdd FILL
XFILL_0__7579_ gnd vdd FILL
XFILL_2_BUFX2_insert819 gnd vdd FILL
XFILL_3__7288_ gnd vdd FILL
XFILL_1__8111_ gnd vdd FILL
XFILL_0_BUFX2_insert30 gnd vdd FILL
XFILL_1__9091_ gnd vdd FILL
XFILL_0_BUFX2_insert41 gnd vdd FILL
X_9946_ _9946_/Q _9306_/CLK _9306_/R vdd _9946_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert52 gnd vdd FILL
XFILL_3__9027_ gnd vdd FILL
XFILL_0_BUFX2_insert63 gnd vdd FILL
XFILL_0_BUFX2_insert74 gnd vdd FILL
XSFILL13640x63050 gnd vdd FILL
XSFILL94520x59050 gnd vdd FILL
XFILL_0__9249_ gnd vdd FILL
XFILL_0_BUFX2_insert85 gnd vdd FILL
XSFILL79080x58050 gnd vdd FILL
XFILL_0_BUFX2_insert96 gnd vdd FILL
X_9877_ _9937_/A _8853_/B gnd _9878_/C vdd NAND2X1
XFILL_6__7968_ gnd vdd FILL
X_8828_ _8828_/A gnd _8830_/A vdd INVX1
XFILL_6_BUFX2_insert730 gnd vdd FILL
XFILL_4__9771_ gnd vdd FILL
XFILL_6_BUFX2_insert741 gnd vdd FILL
XFILL_6__6919_ gnd vdd FILL
XFILL_4__6983_ gnd vdd FILL
XBUFX2_insert807 _13490_/Y gnd _14290_/C vdd BUFX2
X_10690_ _10676_/B _9794_/B gnd _10690_/Y vdd NAND2X1
X_8759_ _8757_/Y _8759_/B _8759_/C gnd _8811_/D vdd OAI21X1
XBUFX2_insert818 _12384_/Y gnd _8606_/B vdd BUFX2
XFILL_1__9993_ gnd vdd FILL
XBUFX2_insert829 _13287_/Y gnd _7457_/A vdd BUFX2
XSFILL104520x44050 gnd vdd FILL
XFILL_4__8722_ gnd vdd FILL
XFILL_3__9929_ gnd vdd FILL
XSFILL33800x76050 gnd vdd FILL
XFILL_4__8653_ gnd vdd FILL
X_12360_ _12358_/Y _12395_/A _12360_/C gnd _12360_/Y vdd OAI21X1
XFILL_1_CLKBUF1_insert201 gnd vdd FILL
XFILL_1_CLKBUF1_insert212 gnd vdd FILL
XFILL_1__8875_ gnd vdd FILL
XFILL_4__7604_ gnd vdd FILL
X_11311_ _11115_/Y gnd _11311_/Y vdd INVX2
XFILL_1_CLKBUF1_insert223 gnd vdd FILL
XFILL_4__8584_ gnd vdd FILL
X_12291_ _12216_/A gnd _12311_/C gnd _12294_/A vdd NAND3X1
XFILL_1__7826_ gnd vdd FILL
X_14030_ _14030_/A _14029_/Y _14030_/C _14030_/D gnd _14031_/A vdd OAI22X1
X_11242_ _11236_/Y _11013_/Y _11003_/Y gnd _11242_/Y vdd OAI21X1
XFILL_1__7757_ gnd vdd FILL
XFILL_4__7466_ gnd vdd FILL
XSFILL79160x38050 gnd vdd FILL
X_11173_ _12198_/Y _12326_/Y gnd _11173_/Y vdd NOR2X1
XFILL_1__7688_ gnd vdd FILL
XFILL_3_BUFX2_insert620 gnd vdd FILL
X_10124_ _10166_/A _7180_/B gnd _10125_/C vdd NAND2X1
XSFILL94200x41050 gnd vdd FILL
XFILL_3_BUFX2_insert631 gnd vdd FILL
X_15981_ _14563_/Y _15981_/B _15410_/D _14592_/Y gnd _15982_/A vdd OAI22X1
XSFILL113880x40050 gnd vdd FILL
XFILL_2__8220_ gnd vdd FILL
XFILL_1__9427_ gnd vdd FILL
XFILL_3_BUFX2_insert642 gnd vdd FILL
XFILL_3_BUFX2_insert653 gnd vdd FILL
XFILL_4__9136_ gnd vdd FILL
XFILL_3_BUFX2_insert664 gnd vdd FILL
XFILL_3_BUFX2_insert675 gnd vdd FILL
X_14932_ _10229_/Q gnd _14932_/Y vdd INVX1
X_10055_ _14777_/A gnd _10057_/A vdd INVX1
XFILL_3_BUFX2_insert686 gnd vdd FILL
XSFILL84280x29050 gnd vdd FILL
XFILL_1__9358_ gnd vdd FILL
XFILL_3_BUFX2_insert697 gnd vdd FILL
XFILL_2__7102_ gnd vdd FILL
XSFILL98840x44050 gnd vdd FILL
XFILL_5__10620_ gnd vdd FILL
X_14863_ _8435_/Q gnd _14863_/Y vdd INVX1
XFILL_2__10440_ gnd vdd FILL
XFILL_2__8082_ gnd vdd FILL
XFILL_1__9289_ gnd vdd FILL
XFILL_5__8900_ gnd vdd FILL
XFILL_4__8018_ gnd vdd FILL
XSFILL99480x10050 gnd vdd FILL
X_13814_ _13813_/Y _13814_/B gnd _13814_/Y vdd NOR2X1
XFILL_5__9880_ gnd vdd FILL
XFILL_4__11000_ gnd vdd FILL
XFILL_5__10551_ gnd vdd FILL
XFILL_2__7033_ gnd vdd FILL
X_14794_ _9290_/A gnd _14796_/D vdd INVX1
XFILL_3__11730_ gnd vdd FILL
XFILL_2__10371_ gnd vdd FILL
XFILL_5__8831_ gnd vdd FILL
XFILL_0__11550_ gnd vdd FILL
XFILL_5__13270_ gnd vdd FILL
X_13745_ _14200_/C _13744_/Y _14636_/C _13743_/Y gnd _13749_/A vdd OAI22X1
XFILL_2__12110_ gnd vdd FILL
X_10957_ _12782_/A _10957_/B gnd _10957_/Y vdd NAND2X1
XFILL_2__13090_ gnd vdd FILL
XSFILL23560x46050 gnd vdd FILL
XFILL_0__10501_ gnd vdd FILL
XFILL_3__11661_ gnd vdd FILL
XFILL_1__12840_ gnd vdd FILL
XSFILL43880x6050 gnd vdd FILL
XFILL_5__8762_ gnd vdd FILL
XSFILL109320x36050 gnd vdd FILL
XFILL_0__11481_ gnd vdd FILL
XFILL_5__12221_ gnd vdd FILL
XFILL_3__13400_ gnd vdd FILL
XSFILL13800x23050 gnd vdd FILL
X_13676_ _7514_/Q gnd _13676_/Y vdd INVX1
XFILL_2__12041_ gnd vdd FILL
XFILL_4__12951_ gnd vdd FILL
XFILL_0__13220_ gnd vdd FILL
X_10888_ _10879_/Y _10888_/B _10878_/Y gnd _10889_/A vdd AOI21X1
XFILL_3__14380_ gnd vdd FILL
XFILL_3__11592_ gnd vdd FILL
XSFILL79240x18050 gnd vdd FILL
XFILL_0_BUFX2_insert510 gnd vdd FILL
XFILL_1__12771_ gnd vdd FILL
XFILL_0__10432_ gnd vdd FILL
XFILL_2__8984_ gnd vdd FILL
XFILL_5__7713_ gnd vdd FILL
XFILL112120x75050 gnd vdd FILL
X_15415_ _9311_/Q _15892_/B gnd _15415_/Y vdd NAND2X1
XFILL_0_BUFX2_insert521 gnd vdd FILL
X_12627_ _12683_/Q gnd _12627_/Y vdd INVX1
XFILL_4__11902_ gnd vdd FILL
XFILL_5__12152_ gnd vdd FILL
X_16395_ _16393_/Y gnd _16394_/Y gnd _16441_/D vdd OAI21X1
XFILL_0_BUFX2_insert532 gnd vdd FILL
XFILL_3__13331_ gnd vdd FILL
XFILL_4__15670_ gnd vdd FILL
XFILL_2__7935_ gnd vdd FILL
XFILL_1__14510_ gnd vdd FILL
XFILL_4__12882_ gnd vdd FILL
XFILL_3__10543_ gnd vdd FILL
XFILL_0_BUFX2_insert543 gnd vdd FILL
XFILL_1__11722_ gnd vdd FILL
XFILL_0__13151_ gnd vdd FILL
XFILL_1__15490_ gnd vdd FILL
XFILL_0_BUFX2_insert554 gnd vdd FILL
XFILL_0_BUFX2_insert565 gnd vdd FILL
XFILL_5__11103_ gnd vdd FILL
XFILL_0__10363_ gnd vdd FILL
X_15346_ _15204_/A _13823_/Y _13822_/Y _15980_/C gnd _15347_/B vdd OAI22X1
XFILL_4__14621_ gnd vdd FILL
XSFILL114440x27050 gnd vdd FILL
XFILL_0__6950_ gnd vdd FILL
XFILL_5__12083_ gnd vdd FILL
X_12558_ _12508_/A _13175_/CLK _13199_/R vdd _12510_/Y gnd vdd DFFSR
XFILL_2__15800_ gnd vdd FILL
XFILL_0_BUFX2_insert576 gnd vdd FILL
XFILL_3__16050_ gnd vdd FILL
XFILL_4__11833_ gnd vdd FILL
XFILL_3__13262_ gnd vdd FILL
XFILL_0__12102_ gnd vdd FILL
XFILL_0_BUFX2_insert587 gnd vdd FILL
XFILL_1__14441_ gnd vdd FILL
XFILL_0_BUFX2_insert598 gnd vdd FILL
XFILL_2__7866_ gnd vdd FILL
XFILL_1__11653_ gnd vdd FILL
XFILL_0__10294_ gnd vdd FILL
XFILL_2__13992_ gnd vdd FILL
XFILL_0__13082_ gnd vdd FILL
XFILL_5__15911_ gnd vdd FILL
XFILL_3__15001_ gnd vdd FILL
XFILL_5__7575_ gnd vdd FILL
X_11509_ _11181_/Y _11509_/B _11495_/C _11182_/Y gnd _11510_/C vdd AOI22X1
XFILL_5__11034_ gnd vdd FILL
XFILL_4__14552_ gnd vdd FILL
XFILL_0__6881_ gnd vdd FILL
XFILL_3__12213_ gnd vdd FILL
XFILL_2__9605_ gnd vdd FILL
X_15277_ _7301_/A _15114_/B _15114_/C gnd _15278_/C vdd NAND3X1
XFILL_2__15731_ gnd vdd FILL
X_12489_ _12489_/A vdd _12488_/Y gnd _12551_/D vdd OAI21X1
XFILL_4__11764_ gnd vdd FILL
XFILL_0__12033_ gnd vdd FILL
XFILL_1__14372_ gnd vdd FILL
XFILL_1__11584_ gnd vdd FILL
XFILL_6__15112_ gnd vdd FILL
X_14228_ _8678_/Q gnd _14228_/Y vdd INVX1
XFILL_0__8620_ gnd vdd FILL
XFILL_4__13503_ gnd vdd FILL
XFILL_5__15842_ gnd vdd FILL
XFILL_1__13323_ gnd vdd FILL
XFILL_4__14483_ gnd vdd FILL
XFILL_2__9536_ gnd vdd FILL
XFILL_1__16111_ gnd vdd FILL
XFILL_3__12144_ gnd vdd FILL
XFILL_1__10535_ gnd vdd FILL
XFILL_2__15662_ gnd vdd FILL
XFILL_4__11695_ gnd vdd FILL
XSFILL84200x73050 gnd vdd FILL
XFILL_2__12874_ gnd vdd FILL
XFILL_5__9245_ gnd vdd FILL
XFILL_4__16222_ gnd vdd FILL
XCLKBUF1_insert200 CLKBUF1_insert169/A gnd _9823_/CLK vdd CLKBUF1
X_14159_ _8036_/Q gnd _15642_/D vdd INVX1
XCLKBUF1_insert211 CLKBUF1_insert206/A gnd _8161_/CLK vdd CLKBUF1
XFILL_4__13434_ gnd vdd FILL
XFILL_1__16042_ gnd vdd FILL
XFILL_2__14613_ gnd vdd FILL
XFILL_3__12075_ gnd vdd FILL
XFILL_5__12985_ gnd vdd FILL
XCLKBUF1_insert222 CLKBUF1_insert169/A gnd _8176_/CLK vdd CLKBUF1
XFILL_5__15773_ gnd vdd FILL
X_7090_ _7090_/A gnd _7092_/A vdd INVX1
XFILL_4__10646_ gnd vdd FILL
XFILL_1__13254_ gnd vdd FILL
XFILL_3__8260_ gnd vdd FILL
XFILL_2__11825_ gnd vdd FILL
XFILL_2__9467_ gnd vdd FILL
XFILL_2__15593_ gnd vdd FILL
XFILL_0__7502_ gnd vdd FILL
XFILL_0__13984_ gnd vdd FILL
XFILL_3__15903_ gnd vdd FILL
XFILL_5__11936_ gnd vdd FILL
XFILL_0__8482_ gnd vdd FILL
XFILL_5__14724_ gnd vdd FILL
XFILL_3__11026_ gnd vdd FILL
XFILL_4__16153_ gnd vdd FILL
XFILL_4__13365_ gnd vdd FILL
XFILL_1__12205_ gnd vdd FILL
XFILL_3__7211_ gnd vdd FILL
XFILL_3__8191_ gnd vdd FILL
XFILL_2__14544_ gnd vdd FILL
XFILL_4__10577_ gnd vdd FILL
XFILL_5__8127_ gnd vdd FILL
XFILL_2__9398_ gnd vdd FILL
XFILL_0__15723_ gnd vdd FILL
XFILL_2__11756_ gnd vdd FILL
XFILL_0__7433_ gnd vdd FILL
XFILL_1__10397_ gnd vdd FILL
XFILL_4__15104_ gnd vdd FILL
XFILL_4__12316_ gnd vdd FILL
XSFILL49080x37050 gnd vdd FILL
XFILL_3__15834_ gnd vdd FILL
XFILL_5__11867_ gnd vdd FILL
XFILL_5__14655_ gnd vdd FILL
XFILL_4__16084_ gnd vdd FILL
XFILL_4__13296_ gnd vdd FILL
XFILL_1__12136_ gnd vdd FILL
XFILL112200x55050 gnd vdd FILL
XFILL_2__10707_ gnd vdd FILL
XFILL_2__8349_ gnd vdd FILL
XFILL_2__14475_ gnd vdd FILL
XFILL_0__15654_ gnd vdd FILL
XFILL_2__11687_ gnd vdd FILL
XFILL_0__12866_ gnd vdd FILL
XFILL_5__8058_ gnd vdd FILL
XFILL_5__13606_ gnd vdd FILL
XFILL_4__15035_ gnd vdd FILL
XSFILL64120x40050 gnd vdd FILL
XFILL_6__15945_ gnd vdd FILL
XFILL_0__7364_ gnd vdd FILL
XFILL_5__10818_ gnd vdd FILL
X_9800_ _9785_/A _7752_/B gnd _9800_/Y vdd NAND2X1
XFILL_2__16214_ gnd vdd FILL
XFILL_5__14586_ gnd vdd FILL
XFILL_4__12247_ gnd vdd FILL
XFILL_2__10638_ gnd vdd FILL
XFILL_0__14605_ gnd vdd FILL
XFILL_3__7073_ gnd vdd FILL
XFILL_2__13426_ gnd vdd FILL
X_7992_ _7992_/A gnd _7994_/A vdd INVX1
XFILL_3__15765_ gnd vdd FILL
XFILL_5__11798_ gnd vdd FILL
XFILL_3__12977_ gnd vdd FILL
XFILL_1__12067_ gnd vdd FILL
XFILL_0__11817_ gnd vdd FILL
XFILL_0__9103_ gnd vdd FILL
XFILL_0__15585_ gnd vdd FILL
XFILL_5__16325_ gnd vdd FILL
XFILL_5__13537_ gnd vdd FILL
XFILL_0__7295_ gnd vdd FILL
X_9731_ _9741_/B _7555_/B gnd _9731_/Y vdd NAND2X1
XFILL_3__14716_ gnd vdd FILL
X_6943_ _6943_/A _6985_/B _6943_/C gnd _7011_/D vdd OAI21X1
XFILL_5__10749_ gnd vdd FILL
XFILL_4__12178_ gnd vdd FILL
XFILL_3__11928_ gnd vdd FILL
XFILL_1__11018_ gnd vdd FILL
XFILL_2__16145_ gnd vdd FILL
XFILL_2__13357_ gnd vdd FILL
XFILL_3__15696_ gnd vdd FILL
XFILL_0__14536_ gnd vdd FILL
XFILL_2__10569_ gnd vdd FILL
XFILL_0__9034_ gnd vdd FILL
XFILL_0__11748_ gnd vdd FILL
XSFILL53960x83050 gnd vdd FILL
X_9662_ _9710_/Q gnd _9664_/A vdd INVX1
XFILL_5__13468_ gnd vdd FILL
XFILL_4__11129_ gnd vdd FILL
XFILL_5__16256_ gnd vdd FILL
XFILL_3__14647_ gnd vdd FILL
X_6874_ _6874_/A gnd memoryWriteData[4] vdd BUFX2
XFILL_2__12308_ gnd vdd FILL
XFILL_2__13288_ gnd vdd FILL
XFILL_1__15826_ gnd vdd FILL
XFILL_3__11859_ gnd vdd FILL
XFILL_2__16076_ gnd vdd FILL
XFILL_0__14467_ gnd vdd FILL
XFILL_5__15207_ gnd vdd FILL
X_8613_ _8611_/Y _8567_/B _8613_/C gnd _8677_/D vdd OAI21X1
XFILL_5__12419_ gnd vdd FILL
XFILL_0__11679_ gnd vdd FILL
XFILL_5__16187_ gnd vdd FILL
XFILL_0__16206_ gnd vdd FILL
XFILL_2__15027_ gnd vdd FILL
XFILL_5__13399_ gnd vdd FILL
XFILL_4__15937_ gnd vdd FILL
XFILL_2__12239_ gnd vdd FILL
X_9593_ _9593_/A gnd _9595_/A vdd INVX1
XFILL_3__14578_ gnd vdd FILL
XFILL_0__13418_ gnd vdd FILL
XFILL_3__7975_ gnd vdd FILL
XFILL_1__15757_ gnd vdd FILL
XSFILL104440x59050 gnd vdd FILL
XFILL_1__12969_ gnd vdd FILL
XFILL_0__14398_ gnd vdd FILL
XSFILL64200x2050 gnd vdd FILL
XFILL_5__15138_ gnd vdd FILL
XFILL_5_BUFX2_insert704 gnd vdd FILL
XFILL_6__7684_ gnd vdd FILL
XFILL_3__16317_ gnd vdd FILL
X_8544_ _8544_/Q _9716_/CLK _8682_/R vdd _8544_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert715 gnd vdd FILL
XFILL_3__13529_ gnd vdd FILL
XFILL_1__6990_ gnd vdd FILL
XFILL_5_BUFX2_insert726 gnd vdd FILL
XFILL_3__6926_ gnd vdd FILL
XFILL_1__14708_ gnd vdd FILL
XFILL_4__15868_ gnd vdd FILL
XFILL_0__16137_ gnd vdd FILL
XFILL_0__13349_ gnd vdd FILL
XFILL_1__15688_ gnd vdd FILL
XFILL_5_BUFX2_insert737 gnd vdd FILL
XFILL_5__15069_ gnd vdd FILL
XFILL_5_BUFX2_insert748 gnd vdd FILL
XFILL_0__9936_ gnd vdd FILL
XFILL_4__14819_ gnd vdd FILL
X_8475_ _8484_/A _8987_/B gnd _8476_/C vdd NAND2X1
XFILL_5_BUFX2_insert759 gnd vdd FILL
XFILL_3__16248_ gnd vdd FILL
XFILL_4__15799_ gnd vdd FILL
XFILL_3__9645_ gnd vdd FILL
XFILL_1__14639_ gnd vdd FILL
XFILL_3__6857_ gnd vdd FILL
XFILL_0__16068_ gnd vdd FILL
XSFILL49160x17050 gnd vdd FILL
X_7426_ _7514_/Q gnd _7428_/A vdd INVX1
XSFILL24600x34050 gnd vdd FILL
XSFILL48920x72050 gnd vdd FILL
XFILL_0__9867_ gnd vdd FILL
XFILL_1__8660_ gnd vdd FILL
XFILL_2__15929_ gnd vdd FILL
XFILL_3__16179_ gnd vdd FILL
XFILL_0__15019_ gnd vdd FILL
XSFILL78360x6050 gnd vdd FILL
XSFILL64200x20050 gnd vdd FILL
XFILL_1__7611_ gnd vdd FILL
X_7357_ _7357_/A _7336_/B _7356_/Y gnd _7405_/D vdd OAI21X1
XFILL_1__8591_ gnd vdd FILL
XFILL_3__8527_ gnd vdd FILL
XFILL_4__7320_ gnd vdd FILL
XFILL_0__9798_ gnd vdd FILL
XFILL_1__16309_ gnd vdd FILL
XSFILL13640x58050 gnd vdd FILL
XFILL_1__7542_ gnd vdd FILL
XFILL_0__8749_ gnd vdd FILL
X_7288_ _7286_/Y _7359_/A _7288_/C gnd _7382_/D vdd OAI21X1
XFILL_3__8458_ gnd vdd FILL
XFILL_4__7251_ gnd vdd FILL
XSFILL68840x23050 gnd vdd FILL
X_9027_ _9027_/A _9011_/A _9027_/C gnd _9027_/Y vdd OAI21X1
XSFILL39080x69050 gnd vdd FILL
XFILL_1__7473_ gnd vdd FILL
XFILL_4__7182_ gnd vdd FILL
XFILL_3__8389_ gnd vdd FILL
XFILL_1__9212_ gnd vdd FILL
XFILL_2_BUFX2_insert605 gnd vdd FILL
XFILL_2_BUFX2_insert616 gnd vdd FILL
XSFILL104520x39050 gnd vdd FILL
XFILL_2_BUFX2_insert627 gnd vdd FILL
XFILL_1__9143_ gnd vdd FILL
XFILL_2_BUFX2_insert638 gnd vdd FILL
XSFILL8760x37050 gnd vdd FILL
XFILL_2_BUFX2_insert649 gnd vdd FILL
XSFILL53880x1050 gnd vdd FILL
X_11860_ _11580_/A _11613_/A gnd _11860_/Y vdd NAND2X1
X_9929_ _9927_/Y _9941_/B _9928_/Y gnd _9969_/D vdd OAI21X1
X_10811_ _10861_/Q gnd _10813_/A vdd INVX1
X_11791_ _11026_/A _11732_/B _11764_/D _11026_/B gnd _11792_/C vdd AOI22X1
X_13530_ _13530_/A _14868_/A _14214_/C _9977_/A gnd _13530_/Y vdd AOI22X1
X_10742_ _13410_/A gnd _10742_/Y vdd INVX1
XBUFX2_insert604 BUFX2_insert556/A gnd _8801_/R vdd BUFX2
XBUFX2_insert615 _10926_/Y gnd _12047_/A vdd BUFX2
XFILL_4__9754_ gnd vdd FILL
XSFILL13720x38050 gnd vdd FILL
XFILL_4__6966_ gnd vdd FILL
XBUFX2_insert626 _12363_/Y gnd _9737_/B vdd BUFX2
XFILL_6_BUFX2_insert582 gnd vdd FILL
X_13461_ _14237_/B _13457_/Y _13461_/C _15048_/B gnd _13462_/B vdd OAI22X1
X_10673_ _10671_/Y _10658_/B _10673_/C gnd _10729_/D vdd OAI21X1
XBUFX2_insert637 _12438_/Y gnd _7380_/B vdd BUFX2
XSFILL23880x82050 gnd vdd FILL
XBUFX2_insert648 _10915_/Y gnd _12072_/A vdd BUFX2
XFILL_4__8705_ gnd vdd FILL
XFILL_1__9976_ gnd vdd FILL
XBUFX2_insert659 _11988_/Y gnd _12061_/C vdd BUFX2
X_15200_ _16026_/D _15200_/B _15899_/C _15198_/Y gnd _15200_/Y vdd OAI22X1
X_12412_ _12508_/A gnd _12412_/Y vdd INVX1
XFILL_4__9685_ gnd vdd FILL
X_16180_ _15708_/A _16180_/B _15708_/C gnd _16180_/Y vdd NOR3X1
XFILL_4__6897_ gnd vdd FILL
XFILL_2__7720_ gnd vdd FILL
X_13392_ _11881_/A _12809_/Q gnd _13418_/A vdd NOR2X1
XFILL_4__8636_ gnd vdd FILL
X_15131_ _7128_/Q gnd _15132_/B vdd INVX1
X_12343_ _12343_/A gnd _12343_/Y vdd INVX1
XFILL_1__8858_ gnd vdd FILL
XFILL_4__8567_ gnd vdd FILL
XFILL_5__7360_ gnd vdd FILL
XSFILL13640x4050 gnd vdd FILL
X_15062_ _15062_/A _15313_/B _15061_/Y gnd _15062_/Y vdd NOR3X1
X_12274_ _12271_/Y _12274_/B _12274_/C gnd _12274_/Y vdd NAND3X1
XFILL_1__7809_ gnd vdd FILL
XFILL_3__10190_ gnd vdd FILL
XFILL_2__7582_ gnd vdd FILL
XFILL_1__8789_ gnd vdd FILL
X_14013_ _8545_/Q gnd _14013_/Y vdd INVX1
X_11225_ _10889_/Y _10882_/Y _11224_/Y gnd _11225_/Y vdd NAND3X1
XFILL_4__10500_ gnd vdd FILL
XFILL_4__8498_ gnd vdd FILL
XFILL_5__7291_ gnd vdd FILL
XFILL_1__10320_ gnd vdd FILL
XFILL_4__11480_ gnd vdd FILL
XSFILL18840x71050 gnd vdd FILL
XFILL_5__9030_ gnd vdd FILL
XFILL_4__7449_ gnd vdd FILL
XSFILL19320x78050 gnd vdd FILL
X_11156_ _11156_/A _11407_/C gnd _11569_/C vdd AND2X2
XFILL_5__12770_ gnd vdd FILL
XFILL_4__10431_ gnd vdd FILL
XFILL_2__9252_ gnd vdd FILL
XFILL_2__11610_ gnd vdd FILL
XFILL_2__12590_ gnd vdd FILL
XFILL_1__10251_ gnd vdd FILL
XFILL_3_BUFX2_insert450 gnd vdd FILL
X_10107_ _10107_/A _10106_/A _10107_/C gnd _10107_/Y vdd OAI21X1
XFILL_0__10981_ gnd vdd FILL
XFILL_3_BUFX2_insert461 gnd vdd FILL
XFILL_5__11721_ gnd vdd FILL
XFILL_2__8203_ gnd vdd FILL
XFILL_4__13150_ gnd vdd FILL
X_15964_ _15070_/C _15964_/B _16199_/C _15964_/D gnd _15965_/A vdd OAI22X1
XFILL_3_BUFX2_insert472 gnd vdd FILL
X_11087_ _12156_/Y gnd _11278_/B vdd INVX2
XFILL_3__12900_ gnd vdd FILL
XSFILL13800x18050 gnd vdd FILL
XFILL_3_BUFX2_insert483 gnd vdd FILL
XFILL_2__11541_ gnd vdd FILL
XSFILL59000x3050 gnd vdd FILL
XFILL_4__10362_ gnd vdd FILL
XFILL_0__12720_ gnd vdd FILL
XFILL_3__13880_ gnd vdd FILL
XFILL_3_BUFX2_insert494 gnd vdd FILL
XFILL_4__9119_ gnd vdd FILL
XFILL_1__10182_ gnd vdd FILL
X_10038_ _9996_/A _7990_/B gnd _10038_/Y vdd NAND2X1
XFILL_4__12101_ gnd vdd FILL
X_14915_ _14700_/A _16272_/D _14711_/B _14914_/Y gnd _14915_/Y vdd OAI22X1
XFILL_5__14440_ gnd vdd FILL
XFILL_5__11652_ gnd vdd FILL
X_15895_ _15895_/A _15656_/B _15656_/C gnd _15895_/Y vdd NOR3X1
XFILL_4__13081_ gnd vdd FILL
XFILL_6__13991_ gnd vdd FILL
XFILL_2__8134_ gnd vdd FILL
XFILL_3__12831_ gnd vdd FILL
XFILL_4__10293_ gnd vdd FILL
XFILL_2__14260_ gnd vdd FILL
XFILL_2__11472_ gnd vdd FILL
XFILL_0__12651_ gnd vdd FILL
XSFILL64040x55050 gnd vdd FILL
XFILL_5__9932_ gnd vdd FILL
XFILL_1__14990_ gnd vdd FILL
X_14846_ _14846_/A _14838_/Y _14846_/C gnd _14859_/B vdd NAND3X1
XFILL_4__12032_ gnd vdd FILL
XFILL_5__14371_ gnd vdd FILL
XFILL_2__10423_ gnd vdd FILL
XFILL_2__13211_ gnd vdd FILL
XFILL_3__15550_ gnd vdd FILL
XFILL_5__11583_ gnd vdd FILL
XFILL_3__12762_ gnd vdd FILL
XFILL_2__8065_ gnd vdd FILL
XFILL_2__14191_ gnd vdd FILL
XFILL_0__11602_ gnd vdd FILL
XFILL_0__15370_ gnd vdd FILL
XFILL_1__13941_ gnd vdd FILL
XFILL_5__13322_ gnd vdd FILL
XFILL_0__12582_ gnd vdd FILL
XFILL_0_BUFX2_insert0 gnd vdd FILL
XFILL_5__16110_ gnd vdd FILL
XFILL_5__9863_ gnd vdd FILL
XFILL_5__10534_ gnd vdd FILL
XFILL_0__7080_ gnd vdd FILL
XFILL_3__14501_ gnd vdd FILL
XFILL_2__13142_ gnd vdd FILL
XFILL_3__11713_ gnd vdd FILL
X_14777_ _14777_/A gnd _16151_/D vdd INVX1
X_11989_ _12440_/A _12073_/B _12073_/C gnd gnd _11990_/C vdd AOI22X1
XFILL_0__14321_ gnd vdd FILL
XSFILL43880x13050 gnd vdd FILL
XFILL_3__15481_ gnd vdd FILL
XFILL_0__11533_ gnd vdd FILL
XFILL_1__13872_ gnd vdd FILL
XFILL_5__16041_ gnd vdd FILL
XFILL_5__13253_ gnd vdd FILL
XFILL_5__9794_ gnd vdd FILL
XFILL_6__11824_ gnd vdd FILL
X_13728_ _9221_/A gnd _13728_/Y vdd INVX1
XFILL_6__15592_ gnd vdd FILL
XFILL_3__14432_ gnd vdd FILL
XFILL_1__15611_ gnd vdd FILL
XFILL_4__13983_ gnd vdd FILL
XFILL_3__11644_ gnd vdd FILL
XFILL_0__14252_ gnd vdd FILL
XFILL_1__12823_ gnd vdd FILL
XFILL_2__10285_ gnd vdd FILL
XFILL_5__12204_ gnd vdd FILL
XFILL_5__8745_ gnd vdd FILL
XFILL_0__11464_ gnd vdd FILL
XSFILL84200x68050 gnd vdd FILL
X_16447_ _16268_/A _8815_/CLK _9056_/R vdd _16413_/Y gnd vdd DFFSR
X_13659_ _8834_/A gnd _13659_/Y vdd INVX1
XFILL_4__15722_ gnd vdd FILL
XFILL_2__12024_ gnd vdd FILL
XFILL_5__10396_ gnd vdd FILL
XFILL_3__14363_ gnd vdd FILL
XFILL_1__12754_ gnd vdd FILL
XFILL_1__15542_ gnd vdd FILL
XFILL_0__10415_ gnd vdd FILL
XFILL_2__8967_ gnd vdd FILL
XFILL_3__11575_ gnd vdd FILL
XFILL_3__7760_ gnd vdd FILL
XFILL_0__14183_ gnd vdd FILL
XFILL_0_BUFX2_insert340 gnd vdd FILL
XSFILL28840x50 gnd vdd FILL
XFILL_5__12135_ gnd vdd FILL
XFILL_3__16102_ gnd vdd FILL
XFILL_0_BUFX2_insert351 gnd vdd FILL
XFILL_0__11395_ gnd vdd FILL
XFILL_3__13314_ gnd vdd FILL
XFILL_4__15653_ gnd vdd FILL
X_16378_ _15826_/A gnd _16378_/Y vdd INVX1
XFILL_0_BUFX2_insert362 gnd vdd FILL
XFILL_6__11686_ gnd vdd FILL
XFILL_0_BUFX2_insert373 gnd vdd FILL
XFILL_4__12865_ gnd vdd FILL
XFILL_0__7982_ gnd vdd FILL
XFILL_1__11705_ gnd vdd FILL
XFILL_3__10526_ gnd vdd FILL
XFILL_0__13134_ gnd vdd FILL
XFILL_0_BUFX2_insert384 gnd vdd FILL
XFILL_3__14294_ gnd vdd FILL
XFILL_3__7691_ gnd vdd FILL
XFILL_5__7627_ gnd vdd FILL
XFILL_2__8898_ gnd vdd FILL
XFILL_1__15473_ gnd vdd FILL
XFILL_4__14604_ gnd vdd FILL
X_15329_ _15329_/A _15329_/B gnd _15336_/A vdd NOR2X1
XFILL_0__9721_ gnd vdd FILL
XFILL_0_BUFX2_insert395 gnd vdd FILL
XFILL_3__16033_ gnd vdd FILL
XFILL_5__12066_ gnd vdd FILL
X_8260_ _8304_/Q gnd _8262_/A vdd INVX1
XFILL_0__6933_ gnd vdd FILL
XFILL_4__11816_ gnd vdd FILL
XFILL_3__13245_ gnd vdd FILL
XFILL_4__15584_ gnd vdd FILL
XFILL_2__7849_ gnd vdd FILL
XFILL_1__11636_ gnd vdd FILL
XFILL_1__14424_ gnd vdd FILL
XFILL_2__13975_ gnd vdd FILL
XFILL_0__10277_ gnd vdd FILL
XFILL_5__7558_ gnd vdd FILL
XFILL_5__11017_ gnd vdd FILL
X_7211_ _7211_/A _7210_/A _7211_/C gnd _7271_/D vdd OAI21X1
XFILL_4__14535_ gnd vdd FILL
XSFILL64120x35050 gnd vdd FILL
XFILL_6__10568_ gnd vdd FILL
XFILL_0__9652_ gnd vdd FILL
X_8191_ _8191_/A gnd _8191_/Y vdd INVX1
XFILL_2__15714_ gnd vdd FILL
XFILL_0__6864_ gnd vdd FILL
XFILL_4__11747_ gnd vdd FILL
XFILL_0__12016_ gnd vdd FILL
XFILL_1__14355_ gnd vdd FILL
XFILL_3__9361_ gnd vdd FILL
XFILL_3__10388_ gnd vdd FILL
XFILL_1__11567_ gnd vdd FILL
XFILL_0__8603_ gnd vdd FILL
X_7142_ _7142_/Q _8537_/CLK _8166_/R vdd _7142_/D gnd vdd DFFSR
XFILL_5__15825_ gnd vdd FILL
XFILL_5__7489_ gnd vdd FILL
XFILL_1__13306_ gnd vdd FILL
XFILL_4__14466_ gnd vdd FILL
XFILL_3__8312_ gnd vdd FILL
XFILL_3__12127_ gnd vdd FILL
XFILL_2__9519_ gnd vdd FILL
XFILL_2__15645_ gnd vdd FILL
XFILL_4__11678_ gnd vdd FILL
XFILL_1__10518_ gnd vdd FILL
XFILL_5__9228_ gnd vdd FILL
XFILL_2__12857_ gnd vdd FILL
XFILL_3__9292_ gnd vdd FILL
XFILL_1__14286_ gnd vdd FILL
XFILL_4__16205_ gnd vdd FILL
XFILL_1__11498_ gnd vdd FILL
XFILL_4__13417_ gnd vdd FILL
X_7073_ _7095_/B _8225_/B gnd _7073_/Y vdd NAND2X1
XSFILL3560x42050 gnd vdd FILL
XFILL_4__10629_ gnd vdd FILL
XFILL_5__15756_ gnd vdd FILL
XFILL_1__13237_ gnd vdd FILL
XFILL_1__16025_ gnd vdd FILL
XFILL_3__12058_ gnd vdd FILL
XFILL_4__14397_ gnd vdd FILL
XFILL_5_BUFX2_insert1030 gnd vdd FILL
XFILL_2__11808_ gnd vdd FILL
XFILL_3__8243_ gnd vdd FILL
XFILL_5__12968_ gnd vdd FILL
XFILL_5_BUFX2_insert1041 gnd vdd FILL
XFILL_1__10449_ gnd vdd FILL
XFILL_2__15576_ gnd vdd FILL
XFILL_2__12788_ gnd vdd FILL
XFILL_5_BUFX2_insert1052 gnd vdd FILL
XFILL_5__9159_ gnd vdd FILL
XFILL_0__13967_ gnd vdd FILL
XFILL_5__14707_ gnd vdd FILL
XFILL_4__16136_ gnd vdd FILL
XFILL_4__13348_ gnd vdd FILL
XSFILL28760x54050 gnd vdd FILL
XFILL_5__11919_ gnd vdd FILL
XFILL_0__8465_ gnd vdd FILL
XFILL_5_BUFX2_insert1063 gnd vdd FILL
XFILL_3__11009_ gnd vdd FILL
XFILL_5__15687_ gnd vdd FILL
XFILL_2__14527_ gnd vdd FILL
XFILL_5__12899_ gnd vdd FILL
XFILL_5_BUFX2_insert1085 gnd vdd FILL
XFILL_1__13168_ gnd vdd FILL
XFILL_0__15706_ gnd vdd FILL
XFILL_0__12918_ gnd vdd FILL
XFILL_2__11739_ gnd vdd FILL
XFILL_0__7416_ gnd vdd FILL
XFILL_0__13898_ gnd vdd FILL
XFILL_5__14638_ gnd vdd FILL
XFILL_3__15817_ gnd vdd FILL
XFILL_4__16067_ gnd vdd FILL
XFILL_4__13279_ gnd vdd FILL
XFILL_0__8396_ gnd vdd FILL
XFILL_3__7125_ gnd vdd FILL
XFILL_1__12119_ gnd vdd FILL
XFILL_2__14458_ gnd vdd FILL
XFILL_0__12849_ gnd vdd FILL
XFILL_0__15637_ gnd vdd FILL
XFILL_1__13099_ gnd vdd FILL
XFILL_4__15018_ gnd vdd FILL
XFILL_0__7347_ gnd vdd FILL
X_7975_ _7948_/A _7975_/B gnd _7975_/Y vdd NAND2X1
XFILL_5__14569_ gnd vdd FILL
XFILL_2__13409_ gnd vdd FILL
XSFILL33880x45050 gnd vdd FILL
XFILL_3__15748_ gnd vdd FILL
XFILL_3__7056_ gnd vdd FILL
XFILL_0__15568_ gnd vdd FILL
XFILL_2__14389_ gnd vdd FILL
XSFILL59160x9050 gnd vdd FILL
XFILL_5__16308_ gnd vdd FILL
X_6926_ _6926_/A gnd _6926_/Y vdd INVX1
X_9714_ _9674_/A _8562_/CLK _9430_/R vdd _9676_/Y gnd vdd DFFSR
XFILL_6__15859_ gnd vdd FILL
XFILL_2__16128_ gnd vdd FILL
XFILL_3__15679_ gnd vdd FILL
XSFILL48920x67050 gnd vdd FILL
XFILL_0__14519_ gnd vdd FILL
XSFILL64200x15050 gnd vdd FILL
XFILL_0__15499_ gnd vdd FILL
XFILL_0__9017_ gnd vdd FILL
XFILL_5__16239_ gnd vdd FILL
X_6857_ _6857_/A gnd memoryAddress[19] vdd BUFX2
X_9645_ _9628_/B _9901_/B gnd _9645_/Y vdd NAND2X1
XFILL_1__15809_ gnd vdd FILL
XSFILL24200x31050 gnd vdd FILL
XFILL_2__16059_ gnd vdd FILL
XSFILL49000x76050 gnd vdd FILL
XFILL_5_BUFX2_insert501 gnd vdd FILL
X_9576_ _9516_/A _8680_/CLK _8034_/R vdd _9576_/D gnd vdd DFFSR
XSFILL89400x81050 gnd vdd FILL
XFILL_3__7958_ gnd vdd FILL
XFILL_5_BUFX2_insert512 gnd vdd FILL
XFILL_5_BUFX2_insert523 gnd vdd FILL
XSFILL3640x22050 gnd vdd FILL
X_8527_ _8527_/A _8503_/B _8527_/C gnd _8563_/D vdd OAI21X1
XFILL_5_BUFX2_insert534 gnd vdd FILL
XFILL_1__9761_ gnd vdd FILL
XFILL_5_BUFX2_insert545 gnd vdd FILL
XFILL_1__6973_ gnd vdd FILL
XFILL_3__6909_ gnd vdd FILL
XFILL_5_BUFX2_insert556 gnd vdd FILL
XSFILL28840x34050 gnd vdd FILL
XFILL_4__9470_ gnd vdd FILL
XFILL_5_BUFX2_insert567 gnd vdd FILL
XFILL_3_BUFX2_insert4 gnd vdd FILL
XSFILL94280x10050 gnd vdd FILL
XFILL_3__7889_ gnd vdd FILL
XFILL_5_BUFX2_insert578 gnd vdd FILL
XFILL_0__9919_ gnd vdd FILL
XFILL_1__8712_ gnd vdd FILL
XFILL112120x3050 gnd vdd FILL
XSFILL54120x67050 gnd vdd FILL
X_8458_ _8456_/Y _8484_/A _8458_/C gnd _8540_/D vdd OAI21X1
XFILL_5_BUFX2_insert589 gnd vdd FILL
XFILL_3__9628_ gnd vdd FILL
XSFILL34680x4050 gnd vdd FILL
X_7409_ _7367_/A _7537_/CLK _7537_/R vdd _7409_/D gnd vdd DFFSR
XFILL_1__8643_ gnd vdd FILL
X_8389_ _8345_/B _7877_/B gnd _8389_/Y vdd NAND2X1
XFILL_4__8352_ gnd vdd FILL
XFILL_1__8574_ gnd vdd FILL
XFILL_4__7303_ gnd vdd FILL
X_11010_ _12222_/Y _12120_/Y gnd _11010_/Y vdd NAND2X1
XFILL_2_CLKBUF1_insert115 gnd vdd FILL
XFILL_2_CLKBUF1_insert126 gnd vdd FILL
XSFILL74040x18050 gnd vdd FILL
XFILL_2_CLKBUF1_insert137 gnd vdd FILL
XFILL_2_CLKBUF1_insert148 gnd vdd FILL
XFILL_2_CLKBUF1_insert159 gnd vdd FILL
XFILL_4__7234_ gnd vdd FILL
XFILL_1__7456_ gnd vdd FILL
XFILL_2_BUFX2_insert402 gnd vdd FILL
XFILL_4__7165_ gnd vdd FILL
XFILL_2_BUFX2_insert413 gnd vdd FILL
X_12961_ vdd _12961_/B gnd _12962_/C vdd NAND2X1
XFILL_2_BUFX2_insert424 gnd vdd FILL
XSFILL23880x77050 gnd vdd FILL
XFILL_2_BUFX2_insert435 gnd vdd FILL
XFILL_2_BUFX2_insert446 gnd vdd FILL
X_14700_ _14700_/A _14700_/B _13978_/B _16098_/C gnd _14700_/Y vdd OAI22X1
XSFILL93720x24050 gnd vdd FILL
X_11912_ _11934_/B _11912_/B gnd _11912_/Y vdd NAND2X1
XFILL_4__7096_ gnd vdd FILL
XFILL_2_BUFX2_insert457 gnd vdd FILL
XFILL_2_BUFX2_insert468 gnd vdd FILL
X_15680_ _16432_/Q _15680_/B _15680_/C gnd _15689_/C vdd NAND3X1
XFILL_1__9126_ gnd vdd FILL
X_12892_ _12942_/Q gnd _12892_/Y vdd INVX1
XFILL_2_BUFX2_insert479 gnd vdd FILL
X_14631_ _10302_/A gnd _14631_/Y vdd INVX1
X_11843_ _11214_/Y _10882_/Y gnd _11843_/Y vdd OR2X2
XSFILL79160x51050 gnd vdd FILL
XFILL_5__6860_ gnd vdd FILL
X_14562_ _16390_/A gnd _14562_/Y vdd INVX1
XFILL_1__8008_ gnd vdd FILL
X_11774_ _11774_/A gnd _12461_/B vdd INVX1
XFILL_4__9806_ gnd vdd FILL
XFILL_2__9870_ gnd vdd FILL
XBUFX2_insert401 _13293_/Y gnd _7606_/A vdd BUFX2
X_16301_ _16301_/A _14946_/B _16301_/C _15948_/D gnd _16301_/Y vdd OAI22X1
XBUFX2_insert412 _13484_/Y gnd _14358_/B vdd BUFX2
X_13513_ _7383_/Q gnd _13514_/B vdd INVX1
X_10725_ _10659_/A _8025_/CLK _8025_/R vdd _10661_/Y gnd vdd DFFSR
XFILL_4__7998_ gnd vdd FILL
XFILL_5__10250_ gnd vdd FILL
XBUFX2_insert423 _14991_/Y gnd _15114_/C vdd BUFX2
X_14493_ _14491_/Y _13824_/B _14575_/C _14492_/Y gnd _14497_/B vdd OAI22X1
XSFILL8440x14050 gnd vdd FILL
XFILL_4__10980_ gnd vdd FILL
XBUFX2_insert434 _13326_/Y gnd _8765_/B vdd BUFX2
XFILL_4__9737_ gnd vdd FILL
XBUFX2_insert445 _12378_/Y gnd _6936_/B vdd BUFX2
XFILL_5__8530_ gnd vdd FILL
X_16232_ _7411_/Q _16232_/B _15202_/B gnd _16232_/Y vdd NAND3X1
XFILL_4__6949_ gnd vdd FILL
XBUFX2_insert456 _13442_/Y gnd _14575_/C vdd BUFX2
XBUFX2_insert467 _13318_/Y gnd _8356_/A vdd BUFX2
X_13444_ _13444_/A _14830_/B _14815_/C _13441_/Y gnd _13450_/B vdd OAI22X1
X_10656_ _10656_/A gnd _10656_/Y vdd INVX1
XFILL_5__10181_ gnd vdd FILL
XBUFX2_insert478 _15038_/Y gnd _15681_/B vdd BUFX2
XFILL_3__11360_ gnd vdd FILL
XFILL_2__8752_ gnd vdd FILL
XBUFX2_insert489 _13471_/Y gnd _14862_/C vdd BUFX2
XFILL_5__8461_ gnd vdd FILL
XSFILL9320x42050 gnd vdd FILL
XFILL_4__9668_ gnd vdd FILL
XFILL_0__11180_ gnd vdd FILL
XFILL_6__11471_ gnd vdd FILL
X_16163_ _16163_/A _16141_/Y _16162_/Y gnd _16164_/B vdd NOR3X1
XFILL_4__12650_ gnd vdd FILL
XSFILL99320x64050 gnd vdd FILL
X_13375_ _12809_/Q gnd _13376_/B vdd INVX1
XFILL_2__7703_ gnd vdd FILL
XFILL_3__10311_ gnd vdd FILL
X_10587_ _10501_/A _8152_/CLK _8664_/R vdd _10587_/D gnd vdd DFFSR
XFILL_3__11291_ gnd vdd FILL
XFILL_1__12470_ gnd vdd FILL
XFILL_0__10131_ gnd vdd FILL
XFILL_4__8619_ gnd vdd FILL
X_15114_ _7383_/Q _15114_/B _15114_/C gnd _15115_/C vdd NAND3X1
XFILL_4__9599_ gnd vdd FILL
XFILL_4__11601_ gnd vdd FILL
XFILL_5__8392_ gnd vdd FILL
X_12326_ _12326_/A _12326_/B _12326_/C gnd _12326_/Y vdd NAND3X1
XFILL_3__10242_ gnd vdd FILL
X_16094_ _9412_/A _15380_/B _15380_/C _9924_/A gnd _16095_/B vdd AOI22X1
XFILL_3__13030_ gnd vdd FILL
XFILL_5__13940_ gnd vdd FILL
XFILL_4__12581_ gnd vdd FILL
XFILL_1__11421_ gnd vdd FILL
XFILL_2__7634_ gnd vdd FILL
XFILL_2__13760_ gnd vdd FILL
XFILL_0__10062_ gnd vdd FILL
XFILL_2__10972_ gnd vdd FILL
XFILL_6__13141_ gnd vdd FILL
XFILL_5__7343_ gnd vdd FILL
X_15045_ _15726_/A _13399_/D _13464_/Y _15045_/D gnd _15045_/Y vdd OAI22X1
XFILL_4__14320_ gnd vdd FILL
X_12257_ _6880_/A _12249_/B _12249_/C _12719_/A gnd _12258_/C vdd AOI22X1
XFILL_4__11532_ gnd vdd FILL
XFILL_3__10173_ gnd vdd FILL
XFILL_5__13871_ gnd vdd FILL
XFILL_2__12711_ gnd vdd FILL
XFILL_1__14140_ gnd vdd FILL
XFILL_2__7565_ gnd vdd FILL
XFILL_1__11352_ gnd vdd FILL
XFILL_0__14870_ gnd vdd FILL
XFILL_2__13691_ gnd vdd FILL
XFILL_5__15610_ gnd vdd FILL
X_11208_ _12201_/Y gnd _11208_/Y vdd INVX1
XFILL_4__14251_ gnd vdd FILL
X_12188_ _12179_/A _12895_/A gnd _12189_/C vdd NAND2X1
XFILL_6__10284_ gnd vdd FILL
XFILL_1__10303_ gnd vdd FILL
XFILL_1_BUFX2_insert18 gnd vdd FILL
XSFILL79240x31050 gnd vdd FILL
XFILL_2__15430_ gnd vdd FILL
XFILL_4__11463_ gnd vdd FILL
XFILL_0__13821_ gnd vdd FILL
XFILL_5__9013_ gnd vdd FILL
XFILL_1_BUFX2_insert29 gnd vdd FILL
XFILL_2__12642_ gnd vdd FILL
XFILL_3__14981_ gnd vdd FILL
XFILL_1__14071_ gnd vdd FILL
XFILL_2__7496_ gnd vdd FILL
XFILL_1__11283_ gnd vdd FILL
XSFILL113800x74050 gnd vdd FILL
XFILL_5__12753_ gnd vdd FILL
XFILL_5__15541_ gnd vdd FILL
XFILL_4__10414_ gnd vdd FILL
X_11139_ _11149_/A _11133_/Y _11138_/Y gnd _11139_/Y vdd OAI21X1
XFILL_1__13022_ gnd vdd FILL
XFILL_4__14182_ gnd vdd FILL
XFILL_2__9235_ gnd vdd FILL
XFILL_3__13932_ gnd vdd FILL
XFILL_2__15361_ gnd vdd FILL
XFILL_1__10234_ gnd vdd FILL
XFILL_4__11394_ gnd vdd FILL
XFILL_2__12573_ gnd vdd FILL
XFILL_3_BUFX2_insert280 gnd vdd FILL
XFILL_0__13752_ gnd vdd FILL
XFILL_0__10964_ gnd vdd FILL
XFILL_3_BUFX2_insert291 gnd vdd FILL
XFILL_0__8250_ gnd vdd FILL
XFILL_4__13133_ gnd vdd FILL
X_15947_ _7020_/Q gnd _15947_/Y vdd INVX1
XFILL_5__11704_ gnd vdd FILL
XFILL_5__15472_ gnd vdd FILL
XFILL_2__14312_ gnd vdd FILL
XFILL_2__9166_ gnd vdd FILL
XFILL_0__12703_ gnd vdd FILL
XFILL_3__13863_ gnd vdd FILL
XFILL_2__11524_ gnd vdd FILL
XFILL_1__10165_ gnd vdd FILL
XFILL_2__15292_ gnd vdd FILL
XFILL_0__13683_ gnd vdd FILL
XFILL_0__7201_ gnd vdd FILL
XFILL_0__10895_ gnd vdd FILL
XFILL_5__11635_ gnd vdd FILL
XFILL_3__15602_ gnd vdd FILL
XFILL_5__14423_ gnd vdd FILL
XFILL_2__8117_ gnd vdd FILL
XSFILL59000x39050 gnd vdd FILL
X_15878_ _15878_/A gnd _15878_/Y vdd INVX1
XFILL_4__10276_ gnd vdd FILL
XFILL_2__14243_ gnd vdd FILL
XFILL_2__11455_ gnd vdd FILL
XFILL_0__15422_ gnd vdd FILL
XFILL_0__12634_ gnd vdd FILL
XFILL_3__13794_ gnd vdd FILL
XFILL_2__9097_ gnd vdd FILL
XFILL_2_BUFX2_insert980 gnd vdd FILL
XSFILL69160x83050 gnd vdd FILL
XFILL_5__9915_ gnd vdd FILL
XFILL_1__14973_ gnd vdd FILL
XFILL_2_BUFX2_insert991 gnd vdd FILL
XFILL_4__12015_ gnd vdd FILL
X_14829_ _8050_/Q gnd _14830_/D vdd INVX1
XFILL_5__14354_ gnd vdd FILL
XFILL_3__15533_ gnd vdd FILL
XFILL_5__11566_ gnd vdd FILL
X_7760_ _7796_/Q gnd _7762_/A vdd INVX1
XFILL_2__10406_ gnd vdd FILL
XFILL_3__12745_ gnd vdd FILL
XFILL111720x38050 gnd vdd FILL
XFILL_2__14174_ gnd vdd FILL
XFILL_0__15353_ gnd vdd FILL
XFILL_2__11386_ gnd vdd FILL
XFILL_1__13924_ gnd vdd FILL
XFILL_5__9846_ gnd vdd FILL
XFILL_5__13305_ gnd vdd FILL
XFILL_6__15644_ gnd vdd FILL
XFILL_0__7063_ gnd vdd FILL
XFILL_5__10517_ gnd vdd FILL
XFILL_5__14285_ gnd vdd FILL
X_7691_ _7773_/Q gnd _7691_/Y vdd INVX1
XFILL_2__13125_ gnd vdd FILL
XFILL_0__14304_ gnd vdd FILL
XFILL_3__15464_ gnd vdd FILL
XFILL_5__11497_ gnd vdd FILL
XFILL_0__11516_ gnd vdd FILL
XFILL_3__8861_ gnd vdd FILL
XFILL_1__13855_ gnd vdd FILL
XFILL_0__15284_ gnd vdd FILL
XFILL_5__13236_ gnd vdd FILL
XFILL_5__16024_ gnd vdd FILL
X_9430_ _9334_/A _9436_/CLK _9430_/R vdd _9430_/D gnd vdd DFFSR
XFILL_0__12496_ gnd vdd FILL
XFILL_5__9777_ gnd vdd FILL
XFILL_5__6989_ gnd vdd FILL
XFILL_5__10448_ gnd vdd FILL
XFILL_3__14415_ gnd vdd FILL
XFILL_3__7812_ gnd vdd FILL
XFILL_3__11627_ gnd vdd FILL
XFILL_4__13966_ gnd vdd FILL
XFILL_3__15395_ gnd vdd FILL
XFILL_0__14235_ gnd vdd FILL
XFILL_2__10268_ gnd vdd FILL
XFILL_5__8728_ gnd vdd FILL
XFILL_2__9999_ gnd vdd FILL
XFILL_0__11447_ gnd vdd FILL
XFILL_1__13786_ gnd vdd FILL
XSFILL79320x11050 gnd vdd FILL
XFILL_1__10998_ gnd vdd FILL
XFILL_4__15705_ gnd vdd FILL
XFILL_5__13167_ gnd vdd FILL
XSFILL49080x50050 gnd vdd FILL
X_9361_ _9361_/A gnd _9363_/A vdd INVX1
XFILL_5__10379_ gnd vdd FILL
XFILL_2__12007_ gnd vdd FILL
XFILL_3__14346_ gnd vdd FILL
XSFILL3560x37050 gnd vdd FILL
XFILL_4__12917_ gnd vdd FILL
XFILL_3__7743_ gnd vdd FILL
XFILL_1__15525_ gnd vdd FILL
XFILL_4__13897_ gnd vdd FILL
XFILL_3__11558_ gnd vdd FILL
XFILL_1__12737_ gnd vdd FILL
XFILL_0__14166_ gnd vdd FILL
X_8312_ _8312_/A _8356_/A _8312_/C gnd _8406_/D vdd OAI21X1
XBUFX2_insert990 _13351_/Y gnd _9993_/A vdd BUFX2
XFILL_5__12118_ gnd vdd FILL
XFILL_0__11378_ gnd vdd FILL
XFILL_5__8659_ gnd vdd FILL
XFILL_6__14457_ gnd vdd FILL
XFILL_3__10509_ gnd vdd FILL
XFILL_4__12848_ gnd vdd FILL
XFILL_4__15636_ gnd vdd FILL
XSFILL28760x49050 gnd vdd FILL
XFILL_5__13098_ gnd vdd FILL
X_9292_ _9292_/A _9301_/B _9292_/C gnd _9292_/Y vdd OAI21X1
XFILL_0__7965_ gnd vdd FILL
XFILL_0__13117_ gnd vdd FILL
XSFILL114520x20050 gnd vdd FILL
XFILL_3__14277_ gnd vdd FILL
XFILL_4_BUFX2_insert508 gnd vdd FILL
XFILL_3__11489_ gnd vdd FILL
XFILL_3__7674_ gnd vdd FILL
XFILL_1__15456_ gnd vdd FILL
XFILL_6__13408_ gnd vdd FILL
XFILL_4_BUFX2_insert519 gnd vdd FILL
XFILL_0__14097_ gnd vdd FILL
XFILL_3__16016_ gnd vdd FILL
XFILL_0__6916_ gnd vdd FILL
XFILL_5__12049_ gnd vdd FILL
X_8243_ _8244_/B _8243_/B gnd _8244_/C vdd NAND2X1
XFILL_3__13228_ gnd vdd FILL
XFILL_3__9413_ gnd vdd FILL
XFILL_4__12779_ gnd vdd FILL
XFILL_4__15567_ gnd vdd FILL
XFILL_1__14407_ gnd vdd FILL
XFILL_2__13958_ gnd vdd FILL
XFILL_1__11619_ gnd vdd FILL
XFILL_1__15387_ gnd vdd FILL
XFILL_1__12599_ gnd vdd FILL
XFILL_0__9635_ gnd vdd FILL
X_8174_ _8126_/A _8942_/CLK _8942_/R vdd _8174_/D gnd vdd DFFSR
XFILL_4__14518_ gnd vdd FILL
XFILL_0__6847_ gnd vdd FILL
XSFILL3560x6050 gnd vdd FILL
XSFILL44120x1050 gnd vdd FILL
XFILL_3__9344_ gnd vdd FILL
XSFILL69240x63050 gnd vdd FILL
XFILL_4__15498_ gnd vdd FILL
XFILL_3__13159_ gnd vdd FILL
XFILL_2__12909_ gnd vdd FILL
XFILL_1__14338_ gnd vdd FILL
XFILL_2__13889_ gnd vdd FILL
X_7125_ _7125_/A _7068_/B _7124_/Y gnd _7125_/Y vdd OAI21X1
XFILL_5__15808_ gnd vdd FILL
XFILL_6__16058_ gnd vdd FILL
XFILL_4__14449_ gnd vdd FILL
XFILL_2__15628_ gnd vdd FILL
XFILL_3__9275_ gnd vdd FILL
XFILL_6__8004_ gnd vdd FILL
XSFILL104440x72050 gnd vdd FILL
XFILL_6__15009_ gnd vdd FILL
XFILL_1__14269_ gnd vdd FILL
XFILL_1__7310_ gnd vdd FILL
XFILL_0__8517_ gnd vdd FILL
X_7056_ _7054_/Y _7055_/A _7056_/C gnd _7134_/D vdd OAI21X1
XFILL_0__14999_ gnd vdd FILL
XFILL_5__15739_ gnd vdd FILL
XFILL_1__16008_ gnd vdd FILL
XFILL_0__9497_ gnd vdd FILL
XFILL_3__8226_ gnd vdd FILL
XSFILL74360x54050 gnd vdd FILL
XFILL_2__15559_ gnd vdd FILL
XFILL_0__8448_ gnd vdd FILL
XFILL_4__16119_ gnd vdd FILL
XFILL_1__7241_ gnd vdd FILL
XSFILL89400x76050 gnd vdd FILL
XSFILL3640x17050 gnd vdd FILL
XFILL_1__7172_ gnd vdd FILL
XFILL_0__8379_ gnd vdd FILL
XFILL_3__7108_ gnd vdd FILL
XFILL_4__8970_ gnd vdd FILL
XFILL_3__8088_ gnd vdd FILL
XFILL_1_BUFX2_insert409 gnd vdd FILL
XFILL_6__9886_ gnd vdd FILL
XFILL_3__7039_ gnd vdd FILL
X_7958_ _7958_/A _7955_/B _7957_/Y gnd _8032_/D vdd OAI21X1
XSFILL13640x71050 gnd vdd FILL
XSFILL94520x67050 gnd vdd FILL
XFILL_6__8837_ gnd vdd FILL
X_6909_ _6955_/B _7037_/B gnd _6909_/Y vdd NAND2X1
X_7889_ _7878_/B _7889_/B gnd _7890_/C vdd NAND2X1
XFILL_4__7852_ gnd vdd FILL
X_9628_ _9628_/A _9628_/B _9627_/Y gnd _9628_/Y vdd OAI21X1
XFILL_1_CLKBUF1_insert1077 gnd vdd FILL
X_10510_ _10590_/Q gnd _10510_/Y vdd INVX1
XFILL_5_BUFX2_insert320 gnd vdd FILL
XFILL_1__9813_ gnd vdd FILL
X_11490_ _11490_/A _11433_/Y gnd _11491_/B vdd NAND2X1
XBUFX2_insert10 _13280_/Y gnd _7308_/A vdd BUFX2
XSFILL104520x52050 gnd vdd FILL
XFILL_4__9522_ gnd vdd FILL
XSFILL33560x22050 gnd vdd FILL
X_9559_ _9465_/A _9447_/CLK _7285_/R vdd _9559_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert331 gnd vdd FILL
XBUFX2_insert21 _13443_/Y gnd _13824_/B vdd BUFX2
XSFILL88600x28050 gnd vdd FILL
XFILL_5_BUFX2_insert342 gnd vdd FILL
XFILL_5_BUFX2_insert353 gnd vdd FILL
X_10441_ _10441_/A _10426_/B _10441_/C gnd _10481_/D vdd OAI21X1
XBUFX2_insert32 _13320_/Y gnd _8496_/A vdd BUFX2
XBUFX2_insert43 _14986_/Y gnd _16002_/C vdd BUFX2
XFILL_5_BUFX2_insert364 gnd vdd FILL
XFILL_1__9744_ gnd vdd FILL
XSFILL9240x57050 gnd vdd FILL
XBUFX2_insert54 _13309_/Y gnd _8133_/A vdd BUFX2
XSFILL98760x72050 gnd vdd FILL
XFILL_1__6956_ gnd vdd FILL
XFILL_5_BUFX2_insert375 gnd vdd FILL
XBUFX2_insert65 _12215_/Y gnd _12277_/B vdd BUFX2
XFILL_5_BUFX2_insert386 gnd vdd FILL
XFILL_5_BUFX2_insert397 gnd vdd FILL
XBUFX2_insert76 _12366_/Y gnd _7564_/B vdd BUFX2
XBUFX2_insert87 _13390_/Y gnd _14615_/B vdd BUFX2
X_10372_ _10372_/A _10372_/B _10371_/Y gnd _10372_/Y vdd OAI21X1
X_13160_ _13202_/Q gnd _13160_/Y vdd INVX1
XBUFX2_insert98 _15068_/Y gnd _15683_/B vdd BUFX2
XFILL_1__9675_ gnd vdd FILL
XFILL_4__8404_ gnd vdd FILL
XFILL_1__6887_ gnd vdd FILL
XFILL_4__9384_ gnd vdd FILL
X_12111_ _12111_/A _12436_/A _12111_/C gnd _12114_/A vdd NAND3X1
X_13091_ _12127_/A gnd _13093_/A vdd INVX1
XFILL_1__8626_ gnd vdd FILL
XFILL_4__8335_ gnd vdd FILL
X_12042_ _12042_/A _12042_/B _12042_/C gnd _13119_/B vdd NAND3X1
XFILL_2__7350_ gnd vdd FILL
XSFILL13720x51050 gnd vdd FILL
XFILL_4__8266_ gnd vdd FILL
XSFILL79160x46050 gnd vdd FILL
XFILL_1__7508_ gnd vdd FILL
XFILL_1__8488_ gnd vdd FILL
XFILL_4__7217_ gnd vdd FILL
X_15801_ _15801_/A _14325_/Y _15801_/C _14330_/D gnd _15801_/Y vdd OAI22X1
XFILL_4__8197_ gnd vdd FILL
XFILL_2__9020_ gnd vdd FILL
XSFILL109560x50 gnd vdd FILL
XFILL_1__7439_ gnd vdd FILL
X_13993_ _10465_/Q gnd _13995_/A vdd INVX1
XSFILL33720x8050 gnd vdd FILL
XFILL_2_BUFX2_insert232 gnd vdd FILL
X_15732_ _15732_/A _15732_/B _14597_/C gnd _12872_/B vdd AOI21X1
XFILL_2_BUFX2_insert243 gnd vdd FILL
XFILL_2_BUFX2_insert254 gnd vdd FILL
XSFILL84280x37050 gnd vdd FILL
XFILL_4__10130_ gnd vdd FILL
X_12944_ _12898_/A _8180_/CLK _7391_/R vdd _12900_/Y gnd vdd DFFSR
XFILL_2_BUFX2_insert265 gnd vdd FILL
XFILL_2_BUFX2_insert276 gnd vdd FILL
XFILL_4__7079_ gnd vdd FILL
XFILL_2_BUFX2_insert287 gnd vdd FILL
XSFILL98840x52050 gnd vdd FILL
XFILL_5__7961_ gnd vdd FILL
XFILL_0__10680_ gnd vdd FILL
XFILL_5__11420_ gnd vdd FILL
X_15663_ _15384_/A _15663_/B _14191_/Y _15384_/D gnd _15663_/Y vdd OAI22X1
XFILL_1__9109_ gnd vdd FILL
XFILL_2_BUFX2_insert298 gnd vdd FILL
XFILL_6__10971_ gnd vdd FILL
XFILL_4__10061_ gnd vdd FILL
XFILL_1_BUFX2_insert910 gnd vdd FILL
XSFILL99320x59050 gnd vdd FILL
X_12875_ vdd _12875_/B gnd _12875_/Y vdd NAND2X1
XSFILL59080x13050 gnd vdd FILL
XFILL_2__11240_ gnd vdd FILL
XFILL_1_BUFX2_insert921 gnd vdd FILL
XFILL_5__6912_ gnd vdd FILL
XFILL_3__10791_ gnd vdd FILL
XFILL_1__11970_ gnd vdd FILL
XFILL_1_BUFX2_insert932 gnd vdd FILL
X_14614_ _8814_/Q gnd _14614_/Y vdd INVX1
X_11826_ _11234_/Y _11240_/Y _11835_/C gnd _11827_/C vdd AOI21X1
XFILL_1_BUFX2_insert943 gnd vdd FILL
XFILL_5__11351_ gnd vdd FILL
XFILL_5__7892_ gnd vdd FILL
XFILL_1_BUFX2_insert954 gnd vdd FILL
XFILL_3__12530_ gnd vdd FILL
XFILL_2__9922_ gnd vdd FILL
X_15594_ _9373_/A _15114_/C _15764_/C gnd _15595_/C vdd NAND3X1
XFILL_1_BUFX2_insert965 gnd vdd FILL
XFILL_1__10921_ gnd vdd FILL
XFILL_2__11171_ gnd vdd FILL
XFILL_0__12350_ gnd vdd FILL
XFILL_1_BUFX2_insert976 gnd vdd FILL
XFILL_5__9631_ gnd vdd FILL
XFILL112280x19050 gnd vdd FILL
XFILL_5__10302_ gnd vdd FILL
XFILL_5__6843_ gnd vdd FILL
XFILL_1_BUFX2_insert987 gnd vdd FILL
XFILL_4__13820_ gnd vdd FILL
X_14545_ _14544_/Y _14545_/B _14489_/C _14543_/Y gnd _14545_/Y vdd OAI22X1
XFILL_5__14070_ gnd vdd FILL
XFILL_2__10122_ gnd vdd FILL
XFILL_1_BUFX2_insert998 gnd vdd FILL
XFILL_5__11282_ gnd vdd FILL
X_11757_ _11776_/B _11776_/A gnd _11758_/B vdd AND2X2
XFILL_3__12461_ gnd vdd FILL
XFILL_0__11301_ gnd vdd FILL
XFILL_2__9853_ gnd vdd FILL
XFILL_1__13640_ gnd vdd FILL
XBUFX2_insert231 _11228_/Y gnd _11349_/B vdd BUFX2
XFILL_5__13021_ gnd vdd FILL
XBUFX2_insert242 _15065_/Y gnd _15972_/B vdd BUFX2
XFILL_0__12281_ gnd vdd FILL
XFILL_3__14200_ gnd vdd FILL
X_10708_ _10681_/A _9940_/B gnd _10708_/Y vdd NAND2X1
XFILL_5__10233_ gnd vdd FILL
X_14476_ _14474_/Y _13843_/C _14200_/C _14475_/Y gnd _14480_/A vdd OAI22X1
XBUFX2_insert253 _10922_/Y gnd _14597_/C vdd BUFX2
XFILL_4__13751_ gnd vdd FILL
XFILL_3__11412_ gnd vdd FILL
XFILL_3__15180_ gnd vdd FILL
XFILL_4__10963_ gnd vdd FILL
XFILL_0__14020_ gnd vdd FILL
XBUFX2_insert264 _15024_/Y gnd _16018_/C vdd BUFX2
XFILL_2__14930_ gnd vdd FILL
XFILL_2__10053_ gnd vdd FILL
X_11688_ _11686_/Y _11688_/B _11683_/Y gnd _11689_/C vdd OAI21X1
XFILL_3__12392_ gnd vdd FILL
XFILL_2__9784_ gnd vdd FILL
XBUFX2_insert275 _13364_/Y gnd _10615_/B vdd BUFX2
XFILL_5__8513_ gnd vdd FILL
XFILL_1__13571_ gnd vdd FILL
XFILL_0__11232_ gnd vdd FILL
XSFILL79240x26050 gnd vdd FILL
XFILL112120x83050 gnd vdd FILL
X_16215_ _9933_/A gnd _16217_/A vdd INVX1
XBUFX2_insert286 _15059_/Y gnd _15386_/B vdd BUFX2
XFILL_2__6996_ gnd vdd FILL
XFILL_1__10783_ gnd vdd FILL
XFILL_4__12702_ gnd vdd FILL
X_13427_ _13426_/Y _13427_/B gnd _13428_/B vdd NAND2X1
XFILL_5_CLKBUF1_insert121 gnd vdd FILL
XFILL_6__11523_ gnd vdd FILL
XFILL_5__9493_ gnd vdd FILL
XBUFX2_insert297 _13356_/Y gnd _10271_/B vdd BUFX2
X_10639_ _10661_/B _9487_/B gnd _10640_/C vdd NAND2X1
XFILL_3__14131_ gnd vdd FILL
XFILL_5_CLKBUF1_insert132 gnd vdd FILL
XFILL_5__10164_ gnd vdd FILL
XFILL_6__15291_ gnd vdd FILL
XFILL_1__15310_ gnd vdd FILL
XFILL_4__13682_ gnd vdd FILL
XFILL_1__12522_ gnd vdd FILL
XFILL_2__8735_ gnd vdd FILL
XFILL_3__11343_ gnd vdd FILL
XFILL_2__14861_ gnd vdd FILL
XFILL_5_CLKBUF1_insert143 gnd vdd FILL
XFILL_4__10894_ gnd vdd FILL
XFILL_1__16290_ gnd vdd FILL
XFILL_0__11163_ gnd vdd FILL
XFILL_5_CLKBUF1_insert154 gnd vdd FILL
XFILL_5__8444_ gnd vdd FILL
XFILL_6__14242_ gnd vdd FILL
XSFILL114440x35050 gnd vdd FILL
XFILL_5_CLKBUF1_insert165 gnd vdd FILL
X_16146_ _16144_/Y _15792_/B _15948_/D _16145_/Y gnd _16147_/B vdd OAI22X1
XFILL_4__12633_ gnd vdd FILL
X_13358_ _13274_/A _13365_/B gnd _13361_/A vdd NAND2X1
XFILL_5_CLKBUF1_insert176 gnd vdd FILL
XFILL_4__15421_ gnd vdd FILL
XFILL_0__7750_ gnd vdd FILL
XFILL_5_CLKBUF1_insert187 gnd vdd FILL
XFILL_2__13812_ gnd vdd FILL
XFILL_3__14062_ gnd vdd FILL
XFILL_5__14972_ gnd vdd FILL
XFILL_0__10114_ gnd vdd FILL
XFILL_1__15241_ gnd vdd FILL
XFILL_1__12453_ gnd vdd FILL
XFILL_3__11274_ gnd vdd FILL
XSFILL83880x10050 gnd vdd FILL
XFILL_2__14792_ gnd vdd FILL
XFILL_5_CLKBUF1_insert198 gnd vdd FILL
XFILL_5__8375_ gnd vdd FILL
XFILL_0__15971_ gnd vdd FILL
X_12309_ _6893_/A _12277_/B _12309_/C _11885_/B gnd _12310_/C vdd AOI22X1
XFILL_0__11094_ gnd vdd FILL
XFILL_4__15352_ gnd vdd FILL
XFILL_5__13923_ gnd vdd FILL
X_16077_ _7279_/Q gnd _16077_/Y vdd INVX1
XFILL_3__13013_ gnd vdd FILL
XFILL_0__7681_ gnd vdd FILL
X_13289_ _13342_/B _13289_/B gnd _13289_/Y vdd OR2X2
XFILL_2__7617_ gnd vdd FILL
XFILL_1__11404_ gnd vdd FILL
XFILL_2__13743_ gnd vdd FILL
XSFILL44360x33050 gnd vdd FILL
XFILL_1__15172_ gnd vdd FILL
XFILL_2__10955_ gnd vdd FILL
XFILL_0__10045_ gnd vdd FILL
XFILL_1__12384_ gnd vdd FILL
XFILL_2__8597_ gnd vdd FILL
XFILL_5__7326_ gnd vdd FILL
XFILL_0__14922_ gnd vdd FILL
XFILL_0__9420_ gnd vdd FILL
X_15028_ _15028_/A _15028_/B gnd _15077_/A vdd NOR2X1
XSFILL99400x39050 gnd vdd FILL
XFILL_4__14303_ gnd vdd FILL
XFILL_4__11515_ gnd vdd FILL
XFILL_5__13854_ gnd vdd FILL
XFILL_4__15283_ gnd vdd FILL
XFILL_1__14123_ gnd vdd FILL
XFILL_4__12495_ gnd vdd FILL
XFILL_3__10156_ gnd vdd FILL
XFILL_2__7548_ gnd vdd FILL
XFILL_1__11335_ gnd vdd FILL
XFILL_2__13674_ gnd vdd FILL
XSFILL84200x81050 gnd vdd FILL
XFILL_0__14853_ gnd vdd FILL
XFILL_2__10886_ gnd vdd FILL
XFILL_4__14234_ gnd vdd FILL
XFILL_0__9351_ gnd vdd FILL
XFILL_2__15413_ gnd vdd FILL
XFILL_4__11446_ gnd vdd FILL
XFILL_2__12625_ gnd vdd FILL
XFILL_5__13785_ gnd vdd FILL
XFILL_1__14054_ gnd vdd FILL
XFILL_3__14964_ gnd vdd FILL
XFILL_5__10997_ gnd vdd FILL
XFILL_2__7479_ gnd vdd FILL
XFILL_0__13804_ gnd vdd FILL
XFILL_2__16393_ gnd vdd FILL
XFILL_1__11266_ gnd vdd FILL
XFILL_0__14784_ gnd vdd FILL
XSFILL74280x69050 gnd vdd FILL
XFILL_0__11996_ gnd vdd FILL
XFILL_5__15524_ gnd vdd FILL
XFILL_5__7188_ gnd vdd FILL
XFILL_5__12736_ gnd vdd FILL
XFILL_2__9218_ gnd vdd FILL
XFILL_3__8011_ gnd vdd FILL
XFILL_4__14165_ gnd vdd FILL
X_8930_ _8930_/Q _8680_/CLK _8424_/R vdd _8860_/Y gnd vdd DFFSR
XFILL_1__13005_ gnd vdd FILL
XFILL_0__9282_ gnd vdd FILL
XFILL_3__13915_ gnd vdd FILL
XFILL_2__15344_ gnd vdd FILL
XSFILL68760x6050 gnd vdd FILL
XFILL_4__11377_ gnd vdd FILL
XFILL_3__14895_ gnd vdd FILL
XFILL_0__10947_ gnd vdd FILL
XFILL_0__13735_ gnd vdd FILL
XFILL_1__11197_ gnd vdd FILL
XFILL_4__13116_ gnd vdd FILL
XFILL_0__8233_ gnd vdd FILL
XFILL_5__15455_ gnd vdd FILL
XFILL_2__9149_ gnd vdd FILL
XFILL_3__13846_ gnd vdd FILL
XFILL112200x63050 gnd vdd FILL
X_8861_ _8931_/Q gnd _8863_/A vdd INVX1
XFILL_2__11507_ gnd vdd FILL
XFILL_4__14096_ gnd vdd FILL
XFILL_1__10148_ gnd vdd FILL
XFILL_2__15275_ gnd vdd FILL
XFILL_0__13666_ gnd vdd FILL
XFILL_2__12487_ gnd vdd FILL
XFILL_0__10878_ gnd vdd FILL
XFILL_5__14406_ gnd vdd FILL
X_7812_ _7812_/A _7887_/B _7811_/Y gnd _7898_/D vdd OAI21X1
XFILL_5__11618_ gnd vdd FILL
XFILL_5__15386_ gnd vdd FILL
XFILL_2__14226_ gnd vdd FILL
XFILL_5__12598_ gnd vdd FILL
XFILL_4__10259_ gnd vdd FILL
X_8792_ _8700_/A _8792_/CLK _7896_/R vdd _8792_/D gnd vdd DFFSR
XFILL_0__12617_ gnd vdd FILL
XFILL_0__15405_ gnd vdd FILL
XFILL_3__13777_ gnd vdd FILL
XFILL_2__11438_ gnd vdd FILL
XFILL_3__10989_ gnd vdd FILL
XFILL_1__14956_ gnd vdd FILL
XFILL_0__13597_ gnd vdd FILL
XFILL_0__7115_ gnd vdd FILL
XFILL_0__16385_ gnd vdd FILL
XFILL_6__12908_ gnd vdd FILL
X_7743_ _7744_/B _7743_/B gnd _7743_/Y vdd NAND2X1
XFILL_0_CLKBUF1_insert1083 gnd vdd FILL
XFILL_3__15516_ gnd vdd FILL
XFILL_5__14337_ gnd vdd FILL
XFILL_5__11549_ gnd vdd FILL
XFILL_6__6883_ gnd vdd FILL
XFILL_0__8095_ gnd vdd FILL
XFILL_3__12728_ gnd vdd FILL
XSFILL43800x47050 gnd vdd FILL
XFILL_3__8913_ gnd vdd FILL
XFILL_2__14157_ gnd vdd FILL
XFILL_1__13907_ gnd vdd FILL
XFILL_3__9893_ gnd vdd FILL
XFILL_0__15336_ gnd vdd FILL
XFILL_2__11369_ gnd vdd FILL
XFILL_0__7046_ gnd vdd FILL
XFILL_1__14887_ gnd vdd FILL
XSFILL4040x62050 gnd vdd FILL
XFILL_2__13108_ gnd vdd FILL
X_7674_ _7723_/B _9978_/B gnd _7674_/Y vdd NAND2X1
XFILL_3__15447_ gnd vdd FILL
XSFILL18600x23050 gnd vdd FILL
XFILL_5__14268_ gnd vdd FILL
XFILL_3__12659_ gnd vdd FILL
XFILL_3__8844_ gnd vdd FILL
XSFILL69240x58050 gnd vdd FILL
XFILL_1__13838_ gnd vdd FILL
XFILL_4__14998_ gnd vdd FILL
XFILL_2__14088_ gnd vdd FILL
XFILL_0__15267_ gnd vdd FILL
XFILL_5__16007_ gnd vdd FILL
XFILL_0__12479_ gnd vdd FILL
XFILL_5__13219_ gnd vdd FILL
X_9413_ _9398_/A _9413_/B gnd _9414_/C vdd NAND2X1
XFILL_5__14199_ gnd vdd FILL
XFILL_0__14218_ gnd vdd FILL
XFILL_3__15378_ gnd vdd FILL
XFILL_2__13039_ gnd vdd FILL
XFILL_4__13949_ gnd vdd FILL
XSFILL103960x60050 gnd vdd FILL
XFILL_3__8775_ gnd vdd FILL
XSFILL104440x67050 gnd vdd FILL
XFILL_0__15198_ gnd vdd FILL
XFILL_1__13769_ gnd vdd FILL
X_9344_ _9359_/A _9344_/B gnd _9345_/C vdd NAND2X1
XFILL_3__14329_ gnd vdd FILL
XFILL_0__8997_ gnd vdd FILL
XFILL_1__15508_ gnd vdd FILL
XFILL_3__7726_ gnd vdd FILL
XFILL_0__14149_ gnd vdd FILL
XSFILL23720x14050 gnd vdd FILL
XFILL_4_BUFX2_insert305 gnd vdd FILL
XFILL_4_BUFX2_insert316 gnd vdd FILL
XFILL_0__7948_ gnd vdd FILL
X_9275_ _9325_/Q gnd _9277_/A vdd INVX1
XFILL_4__15619_ gnd vdd FILL
XFILL_4_BUFX2_insert327 gnd vdd FILL
XFILL_4_BUFX2_insert338 gnd vdd FILL
XFILL_1__15439_ gnd vdd FILL
XFILL_4_BUFX2_insert349 gnd vdd FILL
X_8226_ _8224_/Y _8246_/A _8226_/C gnd _8292_/D vdd OAI21X1
XFILL_0__7879_ gnd vdd FILL
XFILL_6__9105_ gnd vdd FILL
XFILL_3__7588_ gnd vdd FILL
XFILL_0__9618_ gnd vdd FILL
X_8157_ _8157_/Q _8171_/CLK _8171_/R vdd _8157_/D gnd vdd DFFSR
XFILL_4__8120_ gnd vdd FILL
XFILL_1__9391_ gnd vdd FILL
XSFILL13640x66050 gnd vdd FILL
X_7108_ _7108_/A gnd _7110_/A vdd INVX1
XFILL_0__9549_ gnd vdd FILL
XFILL_1__8342_ gnd vdd FILL
X_8088_ _8118_/A _8088_/B gnd _8089_/C vdd NAND2X1
XFILL_3__9258_ gnd vdd FILL
X_7039_ _7039_/A gnd _7041_/A vdd INVX1
XFILL_3__8209_ gnd vdd FILL
XFILL_1__8273_ gnd vdd FILL
XSFILL54120x80050 gnd vdd FILL
XFILL_1__7224_ gnd vdd FILL
X_10990_ _10989_/Y gnd _10990_/Y vdd INVX1
XSFILL104520x47050 gnd vdd FILL
XFILL_1_BUFX2_insert228 gnd vdd FILL
XFILL_4__8953_ gnd vdd FILL
XFILL_1_BUFX2_insert239 gnd vdd FILL
X_12660_ _12694_/Q gnd _12660_/Y vdd INVX1
XFILL_1__7086_ gnd vdd FILL
XSFILL74040x31050 gnd vdd FILL
X_11611_ _11610_/Y _11835_/C _11608_/Y gnd _11611_/Y vdd OAI21X1
XFILL_4__8884_ gnd vdd FILL
XFILL_0_BUFX2_insert906 gnd vdd FILL
X_12591_ _12591_/A gnd _12591_/Y vdd INVX1
XFILL_0_BUFX2_insert917 gnd vdd FILL
XFILL_4__7835_ gnd vdd FILL
XFILL_0_BUFX2_insert928 gnd vdd FILL
X_14330_ _14330_/A _14946_/A _13876_/C _14330_/D gnd _14331_/B vdd OAI22X1
XFILL_0_BUFX2_insert939 gnd vdd FILL
X_11542_ _11542_/A _11542_/B _11525_/Y gnd _11543_/B vdd NAND3X1
XFILL_2__6850_ gnd vdd FILL
XSFILL13720x46050 gnd vdd FILL
X_14261_ _13865_/C _7782_/Q _7142_/Q _13592_/D gnd _14263_/A vdd AOI22X1
X_11473_ _11167_/Y _11320_/Y _11473_/C gnd _11478_/B vdd NAND3X1
XFILL_4__9505_ gnd vdd FILL
X_16000_ _16000_/A _16000_/B _14591_/Y _15169_/A gnd _16003_/A vdd OAI22X1
XFILL_1__7988_ gnd vdd FILL
X_13212_ _13209_/Y _13302_/C gnd _13213_/A vdd AND2X2
X_10424_ _15931_/A gnd _10426_/A vdd INVX1
XFILL_4__7697_ gnd vdd FILL
XFILL_1__9727_ gnd vdd FILL
X_14192_ _14190_/Y _13860_/B _13857_/B _14191_/Y gnd _14193_/A vdd OAI22X1
XFILL_2__8520_ gnd vdd FILL
XSFILL80040x50050 gnd vdd FILL
XFILL_1__6939_ gnd vdd FILL
XSFILL54200x60050 gnd vdd FILL
X_13143_ _13153_/B _13143_/B gnd _13144_/C vdd NAND2X1
X_10355_ _10355_/Q _8429_/CLK _9203_/R vdd _10319_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert850 gnd vdd FILL
XFILL_2__8451_ gnd vdd FILL
XFILL_1__9658_ gnd vdd FILL
XFILL_4_BUFX2_insert861 gnd vdd FILL
XFILL_4__9367_ gnd vdd FILL
XFILL_4_BUFX2_insert872 gnd vdd FILL
XFILL_4_BUFX2_insert883 gnd vdd FILL
XFILL_6__11170_ gnd vdd FILL
XFILL_4_BUFX2_insert894 gnd vdd FILL
XFILL_5__10920_ gnd vdd FILL
XFILL_1__8609_ gnd vdd FILL
XFILL_3__10010_ gnd vdd FILL
X_10286_ _10284_/Y _10285_/A _10286_/C gnd _10344_/D vdd OAI21X1
X_13074_ _6897_/A _8169_/CLK _8937_/R vdd _13074_/D gnd vdd DFFSR
XFILL_2__8382_ gnd vdd FILL
XFILL_5__7111_ gnd vdd FILL
XFILL_4__8318_ gnd vdd FILL
XSFILL83560x8050 gnd vdd FILL
XFILL_5__8091_ gnd vdd FILL
X_12025_ _12467_/B _12025_/B _12025_/C gnd gnd _12025_/Y vdd AOI22X1
XFILL_4__9298_ gnd vdd FILL
XSFILL79320x50 gnd vdd FILL
XFILL_4__11300_ gnd vdd FILL
XSFILL99480x13050 gnd vdd FILL
XSFILL74120x11050 gnd vdd FILL
XFILL_2__7333_ gnd vdd FILL
XFILL_4__12280_ gnd vdd FILL
XFILL_1__11120_ gnd vdd FILL
XFILL_2__10671_ gnd vdd FILL
XFILL_4__8249_ gnd vdd FILL
XFILL_5__7042_ gnd vdd FILL
XFILL_0__11850_ gnd vdd FILL
XFILL_4__11231_ gnd vdd FILL
XFILL_2__12410_ gnd vdd FILL
XFILL_5__10782_ gnd vdd FILL
XFILL_5__13570_ gnd vdd FILL
XFILL_3__11961_ gnd vdd FILL
XFILL_0__10801_ gnd vdd FILL
XFILL_1__11051_ gnd vdd FILL
XFILL_2__13390_ gnd vdd FILL
XFILL_0__11781_ gnd vdd FILL
XFILL_5__12521_ gnd vdd FILL
XFILL_3__13700_ gnd vdd FILL
XFILL_2__9003_ gnd vdd FILL
XFILL_3__10912_ gnd vdd FILL
X_13976_ _7319_/A _13818_/A _14847_/C _7137_/Q gnd _13987_/A vdd AOI22X1
XFILL_1__10002_ gnd vdd FILL
XFILL_4__11162_ gnd vdd FILL
XSFILL13800x26050 gnd vdd FILL
XFILL_2__12341_ gnd vdd FILL
XFILL_3__14680_ gnd vdd FILL
XFILL_0__13520_ gnd vdd FILL
XFILL_2__7195_ gnd vdd FILL
XFILL_3__11892_ gnd vdd FILL
XFILL112120x78050 gnd vdd FILL
XSFILL23960x70050 gnd vdd FILL
X_15715_ _14232_/Y _12770_/A _15715_/C gnd _15719_/B vdd NOR3X1
XFILL_4__10113_ gnd vdd FILL
XFILL_5__8993_ gnd vdd FILL
XFILL_5__15240_ gnd vdd FILL
X_12927_ _12847_/A _9060_/CLK _9060_/R vdd _12927_/D gnd vdd DFFSR
XFILL_5__12452_ gnd vdd FILL
XFILL_3__13631_ gnd vdd FILL
XFILL_4__15970_ gnd vdd FILL
XFILL_1__14810_ gnd vdd FILL
XFILL_2__15060_ gnd vdd FILL
XFILL_4__11093_ gnd vdd FILL
XFILL_0__13451_ gnd vdd FILL
XFILL_2__12272_ gnd vdd FILL
XFILL_5__7944_ gnd vdd FILL
XFILL_0__10663_ gnd vdd FILL
XFILL_1__15790_ gnd vdd FILL
XFILL_5__11403_ gnd vdd FILL
X_15646_ _15920_/C _14151_/Y _15646_/C _15646_/D gnd _15646_/Y vdd OAI22X1
XFILL_4__10044_ gnd vdd FILL
XFILL_5__15171_ gnd vdd FILL
XFILL_5__12383_ gnd vdd FILL
XFILL_2__14011_ gnd vdd FILL
X_12858_ _12856_/Y vdd _12858_/C gnd _12930_/D vdd OAI21X1
XFILL_4__14921_ gnd vdd FILL
XFILL_1_BUFX2_insert740 gnd vdd FILL
XFILL_3__16350_ gnd vdd FILL
XFILL_1_BUFX2_insert751 gnd vdd FILL
XFILL_0__12402_ gnd vdd FILL
XFILL_3__13562_ gnd vdd FILL
XFILL_2__11223_ gnd vdd FILL
XFILL_0__16170_ gnd vdd FILL
XFILL_1_BUFX2_insert762 gnd vdd FILL
XFILL_1__14741_ gnd vdd FILL
XFILL_3__10774_ gnd vdd FILL
XFILL_1__11953_ gnd vdd FILL
XFILL_0__13382_ gnd vdd FILL
XSFILL49080x3050 gnd vdd FILL
XFILL_1_BUFX2_insert773 gnd vdd FILL
XFILL_3__15301_ gnd vdd FILL
XFILL_5__7875_ gnd vdd FILL
XFILL_5__14122_ gnd vdd FILL
X_11809_ _11012_/Y _11008_/Y _11809_/C gnd _11810_/C vdd OAI21X1
XFILL_5__11334_ gnd vdd FILL
XFILL_3__12513_ gnd vdd FILL
X_15577_ _9955_/Q gnd _15578_/C vdd INVX1
XFILL_1_BUFX2_insert784 gnd vdd FILL
X_12789_ _12789_/A memoryOutData[31] gnd _12790_/C vdd NAND2X1
XFILL_4__14852_ gnd vdd FILL
XFILL_1_BUFX2_insert795 gnd vdd FILL
XFILL_2__9905_ gnd vdd FILL
XFILL_2__11154_ gnd vdd FILL
XFILL_0__15121_ gnd vdd FILL
XFILL_3__16281_ gnd vdd FILL
XSFILL43880x21050 gnd vdd FILL
XFILL_1__10904_ gnd vdd FILL
XFILL_0__12333_ gnd vdd FILL
XFILL_3__13493_ gnd vdd FILL
XFILL_5__9614_ gnd vdd FILL
XFILL_1__14672_ gnd vdd FILL
XFILL_3__6890_ gnd vdd FILL
XFILL_1__11884_ gnd vdd FILL
XFILL_6__12624_ gnd vdd FILL
XFILL_5__14053_ gnd vdd FILL
X_14528_ _10348_/Q _13621_/B _14214_/C _15962_/A gnd _14528_/Y vdd AOI22X1
XFILL_4_BUFX2_insert11 gnd vdd FILL
XFILL_4__13803_ gnd vdd FILL
XFILL_3__15232_ gnd vdd FILL
XFILL_2__10105_ gnd vdd FILL
XFILL_5__11265_ gnd vdd FILL
XFILL_3__12444_ gnd vdd FILL
XFILL_1__16411_ gnd vdd FILL
XFILL_4_BUFX2_insert22 gnd vdd FILL
XFILL_1__13623_ gnd vdd FILL
XFILL_4__11995_ gnd vdd FILL
XFILL_2__15962_ gnd vdd FILL
XFILL_0__15052_ gnd vdd FILL
XFILL_2__11085_ gnd vdd FILL
XFILL_4_BUFX2_insert33 gnd vdd FILL
XFILL_4__14783_ gnd vdd FILL
XFILL_4_BUFX2_insert44 gnd vdd FILL
XFILL_0__12264_ gnd vdd FILL
XFILL_5__9545_ gnd vdd FILL
XFILL_1__10835_ gnd vdd FILL
XFILL_5__13004_ gnd vdd FILL
XSFILL84200x76050 gnd vdd FILL
X_14459_ _14868_/A _10677_/A _7787_/Q _13865_/C gnd _14460_/B vdd AOI22X1
XFILL_4_BUFX2_insert55 gnd vdd FILL
XFILL_0__8851_ gnd vdd FILL
X_7390_ _7390_/Q _7790_/CLK _9566_/R vdd _7390_/D gnd vdd DFFSR
XFILL_4__10946_ gnd vdd FILL
XFILL_0__14003_ gnd vdd FILL
XFILL_4_BUFX2_insert66 gnd vdd FILL
XFILL_2__10036_ gnd vdd FILL
XFILL_3__15163_ gnd vdd FILL
XFILL_4__13734_ gnd vdd FILL
XFILL_5__11196_ gnd vdd FILL
XFILL_2__14913_ gnd vdd FILL
XFILL_2__9767_ gnd vdd FILL
XFILL_1__16342_ gnd vdd FILL
XSFILL19400x66050 gnd vdd FILL
XFILL_4_BUFX2_insert77 gnd vdd FILL
XFILL_3__12375_ gnd vdd FILL
XFILL_0__11215_ gnd vdd FILL
XFILL_1__10766_ gnd vdd FILL
XFILL_2__15893_ gnd vdd FILL
XFILL_4_BUFX2_insert88 gnd vdd FILL
XFILL_2__6979_ gnd vdd FILL
XFILL_1__13554_ gnd vdd FILL
XFILL_5__9476_ gnd vdd FILL
XFILL_0__12195_ gnd vdd FILL
XFILL_0__7802_ gnd vdd FILL
XFILL_5__10147_ gnd vdd FILL
XFILL_4_BUFX2_insert99 gnd vdd FILL
XSFILL23640x29050 gnd vdd FILL
XFILL_3__14114_ gnd vdd FILL
XFILL_2__8718_ gnd vdd FILL
XFILL_0__8782_ gnd vdd FILL
XFILL_4__13665_ gnd vdd FILL
XFILL_3__11326_ gnd vdd FILL
XFILL_2__14844_ gnd vdd FILL
XFILL_1__12505_ gnd vdd FILL
XFILL_4__10877_ gnd vdd FILL
XFILL_3__15094_ gnd vdd FILL
XSFILL109400x19050 gnd vdd FILL
XFILL_3__8491_ gnd vdd FILL
XFILL_0__11146_ gnd vdd FILL
XFILL_1__16273_ gnd vdd FILL
X_16129_ _16293_/A _7153_/Q _9671_/A _15652_/D gnd _16131_/A vdd AOI22X1
XFILL_1__13485_ gnd vdd FILL
XFILL_1__10697_ gnd vdd FILL
XFILL_4__12616_ gnd vdd FILL
XFILL_0__7733_ gnd vdd FILL
XFILL_4__15404_ gnd vdd FILL
X_9060_ _8992_/A _9060_/CLK _9060_/R vdd _9060_/D gnd vdd DFFSR
XFILL_3__14045_ gnd vdd FILL
XFILL_5__14955_ gnd vdd FILL
XFILL_4__16384_ gnd vdd FILL
XFILL_4__13596_ gnd vdd FILL
XFILL112200x58050 gnd vdd FILL
XFILL_1__15224_ gnd vdd FILL
XFILL_3__11257_ gnd vdd FILL
XFILL_3__7442_ gnd vdd FILL
XFILL_2__8649_ gnd vdd FILL
XFILL_1__12436_ gnd vdd FILL
XFILL_2__14775_ gnd vdd FILL
XFILL_5__8358_ gnd vdd FILL
X_8011_ _7997_/B _8011_/B gnd _8011_/Y vdd NAND2X1
XFILL_2__11987_ gnd vdd FILL
XFILL_0__15954_ gnd vdd FILL
XFILL_2_BUFX2_insert1005 gnd vdd FILL
XFILL_0__11077_ gnd vdd FILL
XFILL_2_BUFX2_insert1016 gnd vdd FILL
XFILL_5__13906_ gnd vdd FILL
XFILL_4__15335_ gnd vdd FILL
XSFILL64120x43050 gnd vdd FILL
XFILL_2__13726_ gnd vdd FILL
XFILL_2_BUFX2_insert1027 gnd vdd FILL
XFILL_5__14886_ gnd vdd FILL
XFILL_2__10938_ gnd vdd FILL
XFILL_2_BUFX2_insert1038 gnd vdd FILL
XFILL_5__7309_ gnd vdd FILL
XFILL_3__7373_ gnd vdd FILL
XFILL_1__12367_ gnd vdd FILL
XFILL_0__10028_ gnd vdd FILL
XFILL_1__15155_ gnd vdd FILL
XFILL_3__11188_ gnd vdd FILL
XFILL_0__14905_ gnd vdd FILL
XFILL_0__9403_ gnd vdd FILL
XFILL_2_BUFX2_insert1049 gnd vdd FILL
XFILL_0__15885_ gnd vdd FILL
XFILL_5__13837_ gnd vdd FILL
XFILL_3__9112_ gnd vdd FILL
XFILL_4__15266_ gnd vdd FILL
XFILL_4__12478_ gnd vdd FILL
XFILL_0__7595_ gnd vdd FILL
XFILL_1__11318_ gnd vdd FILL
XFILL_3__10139_ gnd vdd FILL
XFILL_1__14106_ gnd vdd FILL
XFILL_2__13657_ gnd vdd FILL
XFILL_0__14836_ gnd vdd FILL
XFILL_3__15996_ gnd vdd FILL
XFILL_1__15086_ gnd vdd FILL
XFILL_1__12298_ gnd vdd FILL
XFILL_4__14217_ gnd vdd FILL
XFILL_0__9334_ gnd vdd FILL
XFILL_4__11429_ gnd vdd FILL
XFILL_4__15197_ gnd vdd FILL
XFILL_2__12608_ gnd vdd FILL
XFILL_5__13768_ gnd vdd FILL
X_9962_ _9906_/A _7020_/CLK _8053_/R vdd _9908_/Y gnd vdd DFFSR
XFILL_3__9043_ gnd vdd FILL
XFILL_1__14037_ gnd vdd FILL
XFILL_3__14947_ gnd vdd FILL
XFILL_2__16376_ gnd vdd FILL
XFILL_1__11249_ gnd vdd FILL
XFILL_2__13588_ gnd vdd FILL
XFILL_5__15507_ gnd vdd FILL
XFILL_0__11979_ gnd vdd FILL
XFILL_0__14767_ gnd vdd FILL
XFILL_5__12719_ gnd vdd FILL
XFILL_4__14148_ gnd vdd FILL
XFILL_0__9265_ gnd vdd FILL
X_8913_ _8902_/B _9041_/B gnd _8914_/C vdd NAND2X1
XFILL_2__15327_ gnd vdd FILL
X_9893_ _9891_/Y _9920_/B _9893_/C gnd _9893_/Y vdd OAI21X1
XFILL_3__14878_ gnd vdd FILL
XFILL_5__13699_ gnd vdd FILL
XSFILL44040x10050 gnd vdd FILL
XFILL_0_BUFX2_insert1020 gnd vdd FILL
XFILL_0__13718_ gnd vdd FILL
XFILL_0__8216_ gnd vdd FILL
XFILL_0_BUFX2_insert1031 gnd vdd FILL
XFILL_0__14698_ gnd vdd FILL
XFILL_5__15438_ gnd vdd FILL
XFILL_0_BUFX2_insert1042 gnd vdd FILL
XFILL_3__13829_ gnd vdd FILL
X_8844_ _8845_/B _6924_/B gnd _8844_/Y vdd NAND2X1
XFILL_6__14989_ gnd vdd FILL
XFILL_4__14079_ gnd vdd FILL
XFILL_0_BUFX2_insert1053 gnd vdd FILL
XFILL_2__15258_ gnd vdd FILL
XSFILL94280x50 gnd vdd FILL
XFILL_0_BUFX2_insert1064 gnd vdd FILL
XFILL_1__15988_ gnd vdd FILL
XFILL_0__13649_ gnd vdd FILL
XFILL_0__8147_ gnd vdd FILL
XFILL_0_BUFX2_insert1086 gnd vdd FILL
XFILL_5__15369_ gnd vdd FILL
XFILL_2__14209_ gnd vdd FILL
XSFILL33880x53050 gnd vdd FILL
X_8775_ _8817_/Q gnd _8775_/Y vdd INVX1
XFILL_2__15189_ gnd vdd FILL
XFILL_1__14939_ gnd vdd FILL
XFILL_6_BUFX2_insert945 gnd vdd FILL
XFILL_0__16368_ gnd vdd FILL
XFILL_1__8960_ gnd vdd FILL
XFILL_0__8078_ gnd vdd FILL
X_7726_ _7724_/Y _7672_/B _7726_/C gnd _7784_/D vdd OAI21X1
XSFILL48920x75050 gnd vdd FILL
XFILL_0__15319_ gnd vdd FILL
XFILL_3__9876_ gnd vdd FILL
XSFILL64200x23050 gnd vdd FILL
XFILL_0__16299_ gnd vdd FILL
XFILL_1__8891_ gnd vdd FILL
XFILL_4__7620_ gnd vdd FILL
X_7657_ _7599_/A _7664_/CLK _7920_/R vdd _7601_/Y gnd vdd DFFSR
XFILL_3__8827_ gnd vdd FILL
XFILL_1__7842_ gnd vdd FILL
X_7588_ _7568_/B _9380_/B gnd _7589_/C vdd NAND2X1
XFILL_4__7551_ gnd vdd FILL
XFILL_3__8758_ gnd vdd FILL
XSFILL3640x30050 gnd vdd FILL
XFILL_4_BUFX2_insert102 gnd vdd FILL
X_9327_ _9281_/A _7274_/CLK _7274_/R vdd _9283_/Y gnd vdd DFFSR
XFILL_3__7709_ gnd vdd FILL
XFILL_4__7482_ gnd vdd FILL
XFILL_1__9512_ gnd vdd FILL
XSFILL54120x75050 gnd vdd FILL
X_9258_ _9208_/B _9258_/B gnd _9258_/Y vdd NAND2X1
XFILL_4__9221_ gnd vdd FILL
X_10140_ _10140_/A _10140_/B _10139_/Y gnd _10210_/D vdd OAI21X1
XFILL_3_BUFX2_insert802 gnd vdd FILL
X_8209_ _8209_/A gnd _8209_/Y vdd INVX1
X_9189_ _9123_/A _8537_/CLK _9054_/R vdd _9189_/D gnd vdd DFFSR
XSFILL53880x4050 gnd vdd FILL
XFILL_3_BUFX2_insert813 gnd vdd FILL
XFILL_4__9152_ gnd vdd FILL
XFILL_3_BUFX2_insert824 gnd vdd FILL
XFILL_3_BUFX2_insert835 gnd vdd FILL
XSFILL33960x33050 gnd vdd FILL
XSFILL33160x14050 gnd vdd FILL
X_10071_ _9977_/A _8679_/CLK _7131_/R vdd _9979_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert846 gnd vdd FILL
XFILL_4__8103_ gnd vdd FILL
XFILL_1__9374_ gnd vdd FILL
XFILL_3_BUFX2_insert857 gnd vdd FILL
XFILL_3_BUFX2_insert868 gnd vdd FILL
XFILL_4__9083_ gnd vdd FILL
XFILL_3_BUFX2_insert879 gnd vdd FILL
XFILL_1__8325_ gnd vdd FILL
XSFILL88600x41050 gnd vdd FILL
X_13830_ _9995_/A _14214_/C _13830_/C gnd _13838_/B vdd AOI21X1
XFILL_1__8256_ gnd vdd FILL
X_13761_ _13761_/A _13761_/B gnd _13789_/A vdd NOR2X1
XFILL_1__7207_ gnd vdd FILL
X_10973_ _10973_/A vdd gnd _10974_/C vdd NAND2X1
XSFILL3720x10050 gnd vdd FILL
XFILL_1__8187_ gnd vdd FILL
X_15500_ _15500_/A _15500_/B gnd _15504_/C vdd NOR2X1
X_12712_ _12710_/Y _12718_/B _12711_/Y gnd _12796_/D vdd OAI21X1
XFILL_4__9985_ gnd vdd FILL
XSFILL94200x39050 gnd vdd FILL
XSFILL113880x38050 gnd vdd FILL
X_13692_ _6917_/A gnd _15279_/C vdd INVX1
XSFILL28920x22050 gnd vdd FILL
XSFILL49000x50 gnd vdd FILL
X_15431_ _13905_/A _16099_/B _16099_/C _15431_/D gnd _15431_/Y vdd OAI22X1
X_12643_ vdd memoryOutData[25] gnd _12644_/C vdd NAND2X1
XFILL_2__7951_ gnd vdd FILL
XFILL_0_BUFX2_insert703 gnd vdd FILL
XFILL_1__7069_ gnd vdd FILL
XFILL_0_CLKBUF1_insert140 gnd vdd FILL
XFILL_0_BUFX2_insert714 gnd vdd FILL
XFILL_4__8867_ gnd vdd FILL
X_15362_ _16342_/A _15680_/B _15680_/C gnd _15371_/C vdd NAND3X1
XFILL_0_BUFX2_insert725 gnd vdd FILL
XFILL_0_CLKBUF1_insert151 gnd vdd FILL
X_12574_ vdd memoryOutData[2] gnd _12574_/Y vdd NAND2X1
XFILL_0_CLKBUF1_insert162 gnd vdd FILL
XFILL_2__6902_ gnd vdd FILL
XFILL_0_BUFX2_insert736 gnd vdd FILL
XFILL_0_CLKBUF1_insert173 gnd vdd FILL
XFILL_0_BUFX2_insert747 gnd vdd FILL
XFILL_2__7882_ gnd vdd FILL
XFILL_4__7818_ gnd vdd FILL
XFILL_0_BUFX2_insert758 gnd vdd FILL
XFILL_3__10490_ gnd vdd FILL
XFILL_0_CLKBUF1_insert184 gnd vdd FILL
X_14313_ _8620_/A _13864_/B _13771_/D _8492_/A gnd _14322_/A vdd AOI22X1
XFILL_0_CLKBUF1_insert195 gnd vdd FILL
XFILL_5__7591_ gnd vdd FILL
XFILL_0_BUFX2_insert769 gnd vdd FILL
XFILL_4__10800_ gnd vdd FILL
X_11525_ _11562_/A _11562_/B _11118_/Y gnd _11525_/Y vdd OAI21X1
XFILL_5__11050_ gnd vdd FILL
X_15293_ _15293_/A _15292_/Y gnd _15293_/Y vdd NOR2X1
XFILL_2__9621_ gnd vdd FILL
XFILL_1__10620_ gnd vdd FILL
XFILL_4__11780_ gnd vdd FILL
XSFILL18840x74050 gnd vdd FILL
XFILL_5__10001_ gnd vdd FILL
XFILL_4__7749_ gnd vdd FILL
X_14244_ _15704_/B gnd _14244_/Y vdd INVX1
X_11456_ _11553_/C _11441_/Y _11455_/Y gnd _11456_/Y vdd NAND3X1
XFILL_2__11910_ gnd vdd FILL
XFILL_3__12160_ gnd vdd FILL
XFILL_0__11000_ gnd vdd FILL
XFILL_2__9552_ gnd vdd FILL
XFILL_1__10551_ gnd vdd FILL
XSFILL9320x50050 gnd vdd FILL
XFILL_2__12890_ gnd vdd FILL
XFILL_5__9261_ gnd vdd FILL
X_10407_ _10423_/B _7975_/B gnd _10407_/Y vdd NAND2X1
X_14175_ _8293_/Q gnd _14175_/Y vdd INVX1
XFILL_2__8503_ gnd vdd FILL
XSFILL63960x49050 gnd vdd FILL
XFILL_4__13450_ gnd vdd FILL
XFILL_3__11111_ gnd vdd FILL
XFILL_4__10662_ gnd vdd FILL
X_11387_ _11732_/A _11267_/Y _11386_/Y gnd _11387_/Y vdd OAI21X1
XFILL_2__9483_ gnd vdd FILL
XFILL_1__13270_ gnd vdd FILL
XFILL_4__9419_ gnd vdd FILL
XFILL_3__12091_ gnd vdd FILL
XFILL_5__8212_ gnd vdd FILL
XFILL_2__11841_ gnd vdd FILL
X_13126_ _13126_/A _13168_/B _13125_/Y gnd _13190_/D vdd OAI21X1
XFILL_4__12401_ gnd vdd FILL
XFILL_4_BUFX2_insert680 gnd vdd FILL
XFILL_5__14740_ gnd vdd FILL
X_10338_ _15537_/B _8680_/CLK _8034_/R vdd _10338_/D gnd vdd DFFSR
XFILL_5__11952_ gnd vdd FILL
XFILL_4__13381_ gnd vdd FILL
XFILL_3__11042_ gnd vdd FILL
XFILL_4_BUFX2_insert691 gnd vdd FILL
XFILL_1__12221_ gnd vdd FILL
XFILL_2__14560_ gnd vdd FILL
XFILL112280x32050 gnd vdd FILL
XFILL_5__8143_ gnd vdd FILL
XSFILL64040x58050 gnd vdd FILL
XFILL_2__11772_ gnd vdd FILL
XFILL_0__12951_ gnd vdd FILL
XSFILL113960x18050 gnd vdd FILL
XFILL_4__15120_ gnd vdd FILL
XFILL_5__10903_ gnd vdd FILL
XFILL_4__12332_ gnd vdd FILL
X_13057_ _6880_/A _9823_/CLK _9056_/R vdd _13057_/D gnd vdd DFFSR
X_10269_ _14077_/C gnd _10269_/Y vdd INVX1
XFILL_5__14671_ gnd vdd FILL
XFILL_2__13511_ gnd vdd FILL
XFILL_5__11883_ gnd vdd FILL
XFILL_1__12152_ gnd vdd FILL
XFILL_3__15850_ gnd vdd FILL
XFILL_2__8365_ gnd vdd FILL
XFILL_2__14491_ gnd vdd FILL
XFILL_6__10104_ gnd vdd FILL
XFILL_0__11902_ gnd vdd FILL
XFILL_5__16410_ gnd vdd FILL
XFILL_0__15670_ gnd vdd FILL
XFILL_5__8074_ gnd vdd FILL
X_12008_ _11988_/B _12704_/A _12096_/C gnd _12010_/B vdd NAND3X1
XFILL_0__12882_ gnd vdd FILL
XFILL_5__13622_ gnd vdd FILL
XFILL_4__15051_ gnd vdd FILL
XFILL_6__15961_ gnd vdd FILL
XFILL_2__16230_ gnd vdd FILL
XFILL_3__14801_ gnd vdd FILL
XFILL_0__7380_ gnd vdd FILL
XFILL_4__12263_ gnd vdd FILL
XFILL_1__11103_ gnd vdd FILL
XFILL_2__7316_ gnd vdd FILL
XFILL_5__10834_ gnd vdd FILL
XFILL_2__13442_ gnd vdd FILL
XSFILL114840x46050 gnd vdd FILL
XFILL_3__15781_ gnd vdd FILL
XSFILL43880x16050 gnd vdd FILL
XFILL_0__14621_ gnd vdd FILL
XFILL_1__12083_ gnd vdd FILL
XFILL_3__12993_ gnd vdd FILL
XFILL_2__10654_ gnd vdd FILL
XFILL_0__11833_ gnd vdd FILL
XFILL_4__14002_ gnd vdd FILL
XFILL_6__14912_ gnd vdd FILL
XFILL_5__16341_ gnd vdd FILL
XFILL_4__11214_ gnd vdd FILL
XFILL_5__10765_ gnd vdd FILL
XFILL_3__14732_ gnd vdd FILL
XFILL_5__13553_ gnd vdd FILL
XFILL_2__7247_ gnd vdd FILL
XFILL_1__15911_ gnd vdd FILL
XFILL_3__11944_ gnd vdd FILL
XFILL_4__12194_ gnd vdd FILL
XFILL_2__16161_ gnd vdd FILL
XFILL_1__11034_ gnd vdd FILL
XFILL_2__13373_ gnd vdd FILL
XFILL_0__14552_ gnd vdd FILL
XFILL_0__11764_ gnd vdd FILL
XFILL_5__12504_ gnd vdd FILL
XFILL_4__11145_ gnd vdd FILL
X_13959_ _13959_/A _14697_/B _14752_/C _13959_/D gnd _13959_/Y vdd OAI22X1
XFILL_2__15112_ gnd vdd FILL
XFILL_5__16272_ gnd vdd FILL
XFILL_5__13484_ gnd vdd FILL
XFILL_2__12324_ gnd vdd FILL
XFILL_3__14663_ gnd vdd FILL
XFILL_5__10696_ gnd vdd FILL
X_6890_ _6890_/A gnd memoryWriteData[20] vdd BUFX2
XFILL_2__7178_ gnd vdd FILL
XFILL_3__11875_ gnd vdd FILL
XFILL_2__16092_ gnd vdd FILL
XSFILL84360x30050 gnd vdd FILL
XFILL_1__15842_ gnd vdd FILL
XFILL_0__13503_ gnd vdd FILL
XFILL_0__14483_ gnd vdd FILL
XFILL_0__8001_ gnd vdd FILL
XFILL_5__15223_ gnd vdd FILL
XFILL_0__11695_ gnd vdd FILL
XFILL_5__8976_ gnd vdd FILL
XFILL_3__13614_ gnd vdd FILL
XSFILL59000x47050 gnd vdd FILL
XFILL_5__12435_ gnd vdd FILL
XFILL_3__16402_ gnd vdd FILL
XFILL_6__14774_ gnd vdd FILL
XFILL_3__10826_ gnd vdd FILL
XFILL_2__15043_ gnd vdd FILL
XFILL_4__15953_ gnd vdd FILL
XFILL_4__11076_ gnd vdd FILL
XFILL_3__14594_ gnd vdd FILL
XFILL_0__16222_ gnd vdd FILL
XFILL_0__13434_ gnd vdd FILL
XFILL_2__12255_ gnd vdd FILL
XFILL_3__7991_ gnd vdd FILL
XFILL_1__15773_ gnd vdd FILL
XFILL_0__10646_ gnd vdd FILL
XFILL_1__12985_ gnd vdd FILL
XFILL_5__7927_ gnd vdd FILL
XFILL_6__13725_ gnd vdd FILL
XFILL_1_BUFX2_insert570 gnd vdd FILL
XFILL_5__12366_ gnd vdd FILL
XFILL_3__16333_ gnd vdd FILL
X_15629_ _15629_/A _15629_/B gnd _15651_/A vdd NOR2X1
XFILL_5__15154_ gnd vdd FILL
XFILL_4__14904_ gnd vdd FILL
XFILL_4__10027_ gnd vdd FILL
XFILL_1_BUFX2_insert581 gnd vdd FILL
XFILL_3__9730_ gnd vdd FILL
X_8560_ _8560_/Q _8560_/CLK _8676_/R vdd _8560_/D gnd vdd DFFSR
XFILL_3__13545_ gnd vdd FILL
XFILL_2__11206_ gnd vdd FILL
XFILL_1__14724_ gnd vdd FILL
XFILL_3__6942_ gnd vdd FILL
XFILL_3__10757_ gnd vdd FILL
XSFILL23240x26050 gnd vdd FILL
XFILL_4__15884_ gnd vdd FILL
XFILL_0__13365_ gnd vdd FILL
XFILL_1_BUFX2_insert592 gnd vdd FILL
XFILL_2__12186_ gnd vdd FILL
XFILL_1__11936_ gnd vdd FILL
XFILL_0__16153_ gnd vdd FILL
XFILL_5__14105_ gnd vdd FILL
XFILL_0__10577_ gnd vdd FILL
XFILL_5__7858_ gnd vdd FILL
XFILL_5_BUFX2_insert908 gnd vdd FILL
XFILL_5__11317_ gnd vdd FILL
XFILL112360x12050 gnd vdd FILL
X_7511_ _7511_/Q _8679_/CLK _7131_/R vdd _7511_/D gnd vdd DFFSR
XFILL_4__14835_ gnd vdd FILL
XSFILL64120x38050 gnd vdd FILL
XFILL_5_BUFX2_insert919 gnd vdd FILL
X_8491_ _8489_/Y _8494_/B _8491_/C gnd _8551_/D vdd OAI21X1
XFILL_5__15085_ gnd vdd FILL
XFILL_3__16264_ gnd vdd FILL
XFILL_5__12297_ gnd vdd FILL
XFILL_3__9661_ gnd vdd FILL
XFILL_3__13476_ gnd vdd FILL
XFILL_0__12316_ gnd vdd FILL
XFILL_2__11137_ gnd vdd FILL
XFILL_0__15104_ gnd vdd FILL
XFILL_3__6873_ gnd vdd FILL
XFILL_3__10688_ gnd vdd FILL
XFILL_1__14655_ gnd vdd FILL
XFILL_0__16084_ gnd vdd FILL
XFILL_0__13296_ gnd vdd FILL
XFILL_1__11867_ gnd vdd FILL
XFILL_0__8903_ gnd vdd FILL
XFILL_3__15215_ gnd vdd FILL
XFILL_5__14036_ gnd vdd FILL
XFILL_6__16375_ gnd vdd FILL
XFILL_5__11248_ gnd vdd FILL
X_7442_ _7472_/A _7314_/B gnd _7443_/C vdd NAND2X1
XFILL_6__13587_ gnd vdd FILL
XFILL_3__12427_ gnd vdd FILL
XFILL_3__8612_ gnd vdd FILL
XFILL_0__9883_ gnd vdd FILL
XFILL_1__13606_ gnd vdd FILL
XFILL_3__16195_ gnd vdd FILL
XFILL_0__15035_ gnd vdd FILL
XFILL_2__15945_ gnd vdd FILL
XFILL_4__11978_ gnd vdd FILL
XFILL_4__14766_ gnd vdd FILL
XFILL_2__11068_ gnd vdd FILL
XFILL_3__9592_ gnd vdd FILL
XFILL_0__12247_ gnd vdd FILL
XFILL_1__10818_ gnd vdd FILL
XFILL_1__14586_ gnd vdd FILL
XFILL_6__15326_ gnd vdd FILL
XFILL_5__9528_ gnd vdd FILL
XFILL_0__8834_ gnd vdd FILL
XFILL_1__11798_ gnd vdd FILL
X_7373_ _7411_/Q gnd _7375_/A vdd INVX1
XSFILL3560x45050 gnd vdd FILL
XFILL_4__13717_ gnd vdd FILL
XFILL_5__11179_ gnd vdd FILL
XFILL_3__15146_ gnd vdd FILL
XFILL_2__10019_ gnd vdd FILL
XFILL_4__10929_ gnd vdd FILL
XFILL_3__12358_ gnd vdd FILL
XFILL_1__16325_ gnd vdd FILL
XFILL_4__14697_ gnd vdd FILL
XFILL_1__13537_ gnd vdd FILL
XFILL_2__15876_ gnd vdd FILL
XFILL_6__8252_ gnd vdd FILL
XFILL_0__12178_ gnd vdd FILL
XFILL_1__10749_ gnd vdd FILL
X_9112_ _9112_/A _6936_/B gnd _9112_/Y vdd NAND2X1
XFILL_0__8765_ gnd vdd FILL
XSFILL28760x57050 gnd vdd FILL
XFILL_6__12469_ gnd vdd FILL
XFILL_3__11309_ gnd vdd FILL
XFILL_5__15987_ gnd vdd FILL
XFILL_4__13648_ gnd vdd FILL
XFILL_2__14827_ gnd vdd FILL
XFILL_3__15077_ gnd vdd FILL
XFILL_6__7203_ gnd vdd FILL
XFILL_3__8474_ gnd vdd FILL
XFILL_3__12289_ gnd vdd FILL
XFILL_0__11129_ gnd vdd FILL
XFILL_1__16256_ gnd vdd FILL
XFILL_1__13468_ gnd vdd FILL
XFILL_0__7716_ gnd vdd FILL
X_9043_ _9043_/A gnd _9043_/Y vdd INVX1
XFILL_6__15188_ gnd vdd FILL
XFILL_3__14028_ gnd vdd FILL
XFILL_5__14938_ gnd vdd FILL
XFILL_3__7425_ gnd vdd FILL
XFILL_4__16367_ gnd vdd FILL
XFILL_1__15207_ gnd vdd FILL
XFILL_0__8696_ gnd vdd FILL
XFILL_3_BUFX2_insert109 gnd vdd FILL
XFILL_4__13579_ gnd vdd FILL
XFILL_1__12419_ gnd vdd FILL
XFILL_2__14758_ gnd vdd FILL
XFILL_1__16187_ gnd vdd FILL
XFILL_0__15937_ gnd vdd FILL
XFILL_1__13399_ gnd vdd FILL
XFILL_4__15318_ gnd vdd FILL
XSFILL69240x71050 gnd vdd FILL
XFILL_5__14869_ gnd vdd FILL
XSFILL33880x48050 gnd vdd FILL
XFILL_2__13709_ gnd vdd FILL
XFILL_3__7356_ gnd vdd FILL
XFILL_4__16298_ gnd vdd FILL
XFILL_1__15138_ gnd vdd FILL
XFILL_2__14689_ gnd vdd FILL
XCLKBUF1_insert1076 clk gnd CLKBUF1_insert169/A vdd CLKBUF1
XFILL_0__15868_ gnd vdd FILL
XFILL_2_BUFX2_insert809 gnd vdd FILL
XFILL_4__15249_ gnd vdd FILL
XFILL_0__7578_ gnd vdd FILL
XFILL_3__15979_ gnd vdd FILL
XFILL_3__7287_ gnd vdd FILL
XFILL_0__14819_ gnd vdd FILL
XFILL_1__15069_ gnd vdd FILL
XFILL_0_BUFX2_insert20 gnd vdd FILL
XFILL_1__8110_ gnd vdd FILL
XSFILL64200x18050 gnd vdd FILL
XFILL_0_BUFX2_insert31 gnd vdd FILL
XFILL_0__15799_ gnd vdd FILL
XFILL_1__9090_ gnd vdd FILL
X_9945_ _9945_/Q _8306_/CLK _7533_/R vdd _9945_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert42 gnd vdd FILL
XFILL_3__9026_ gnd vdd FILL
XFILL_2__16359_ gnd vdd FILL
XSFILL74360x62050 gnd vdd FILL
XFILL_0_BUFX2_insert53 gnd vdd FILL
XFILL_0_BUFX2_insert64 gnd vdd FILL
XSFILL49000x79050 gnd vdd FILL
XFILL_0_BUFX2_insert75 gnd vdd FILL
XFILL_0__9248_ gnd vdd FILL
XFILL_0_BUFX2_insert86 gnd vdd FILL
XSFILL23640x2050 gnd vdd FILL
X_9876_ _9952_/Q gnd _9876_/Y vdd INVX1
XFILL_0_BUFX2_insert97 gnd vdd FILL
XSFILL3640x25050 gnd vdd FILL
X_8827_ _8827_/A _8916_/A _8827_/C gnd _8919_/D vdd OAI21X1
XFILL_4__9770_ gnd vdd FILL
XFILL_6_BUFX2_insert720 gnd vdd FILL
XSFILL28840x37050 gnd vdd FILL
XFILL_4__6982_ gnd vdd FILL
XSFILL94280x13050 gnd vdd FILL
XBUFX2_insert808 _13490_/Y gnd _13848_/C vdd BUFX2
XFILL112120x6050 gnd vdd FILL
X_8758_ _8759_/B _7094_/B gnd _8759_/C vdd NAND2X1
XFILL_1__9992_ gnd vdd FILL
XFILL_4__8721_ gnd vdd FILL
XBUFX2_insert819 _12384_/Y gnd _9246_/B vdd BUFX2
XFILL_3__9928_ gnd vdd FILL
XFILL_6__9637_ gnd vdd FILL
X_7709_ _7709_/A gnd _7711_/A vdd INVX1
XFILL_6_BUFX2_insert797 gnd vdd FILL
XFILL_4__8652_ gnd vdd FILL
X_8689_ _8647_/A _8433_/CLK _7921_/R vdd _8689_/D gnd vdd DFFSR
XFILL_3__9859_ gnd vdd FILL
XFILL_1__8874_ gnd vdd FILL
XFILL_4__7603_ gnd vdd FILL
XFILL_1_CLKBUF1_insert202 gnd vdd FILL
XFILL_1_CLKBUF1_insert213 gnd vdd FILL
X_11310_ _11110_/Y gnd _11312_/C vdd INVX1
XFILL_4__8583_ gnd vdd FILL
XFILL_1_CLKBUF1_insert224 gnd vdd FILL
X_12290_ _12287_/Y _12290_/B _12289_/Y gnd _12290_/Y vdd NAND3X1
XFILL_1__7825_ gnd vdd FILL
X_11241_ _11240_/Y _11234_/Y _11241_/C gnd _11241_/Y vdd NAND3X1
XFILL_1__7756_ gnd vdd FILL
XFILL_4__7465_ gnd vdd FILL
X_11172_ _11171_/Y gnd _11195_/A vdd INVX2
XFILL_1__7687_ gnd vdd FILL
XFILL_3_BUFX2_insert610 gnd vdd FILL
X_10123_ _10205_/Q gnd _10123_/Y vdd INVX1
XSFILL110120x58050 gnd vdd FILL
XFILL_3_BUFX2_insert621 gnd vdd FILL
XFILL_3_BUFX2_insert632 gnd vdd FILL
X_15980_ _15899_/A _15979_/Y _15980_/C _14573_/Y gnd _15980_/Y vdd OAI22X1
XFILL_1__9426_ gnd vdd FILL
XFILL_3_BUFX2_insert643 gnd vdd FILL
XFILL_4__9135_ gnd vdd FILL
XFILL_3_BUFX2_insert654 gnd vdd FILL
X_10054_ _10054_/A _10054_/B _10053_/Y gnd _10054_/Y vdd OAI21X1
X_14931_ _8437_/Q _14037_/B _14868_/D _9205_/Q gnd _14931_/Y vdd AOI22X1
XFILL_3_BUFX2_insert665 gnd vdd FILL
XSFILL109240x72050 gnd vdd FILL
XSFILL38280x42050 gnd vdd FILL
XFILL_3_BUFX2_insert676 gnd vdd FILL
XFILL_1__9357_ gnd vdd FILL
XFILL_3_BUFX2_insert687 gnd vdd FILL
XFILL_3_BUFX2_insert698 gnd vdd FILL
XSFILL79160x54050 gnd vdd FILL
XFILL_2__7101_ gnd vdd FILL
X_14862_ _14862_/A _13614_/C _14862_/C _14860_/Y gnd _14866_/A vdd OAI22X1
XFILL_1__9288_ gnd vdd FILL
XFILL_2__8081_ gnd vdd FILL
XFILL_4__8017_ gnd vdd FILL
XSFILL104200x19050 gnd vdd FILL
X_13813_ _13811_/Y _13813_/B _14567_/D _13813_/D gnd _13813_/Y vdd OAI22X1
XFILL_5__10550_ gnd vdd FILL
XSFILL83640x79050 gnd vdd FILL
X_14793_ _13864_/B _8690_/Q _14793_/C _14572_/C gnd _14801_/B vdd AOI22X1
XFILL_2__7032_ gnd vdd FILL
XFILL_1__8239_ gnd vdd FILL
XFILL_2__10370_ gnd vdd FILL
XFILL_5__8830_ gnd vdd FILL
X_13744_ _7048_/A gnd _13744_/Y vdd INVX1
XSFILL84280x45050 gnd vdd FILL
XSFILL104600x40050 gnd vdd FILL
XFILL_6__11840_ gnd vdd FILL
X_10956_ _10946_/Y _10955_/Y _10956_/C gnd _10976_/B vdd NAND3X1
XFILL_0__10500_ gnd vdd FILL
XFILL_3__11660_ gnd vdd FILL
XFILL_5__8761_ gnd vdd FILL
XFILL_5__12220_ gnd vdd FILL
XFILL_0__11480_ gnd vdd FILL
X_13675_ _7810_/A gnd _13675_/Y vdd INVX1
XSFILL99320x67050 gnd vdd FILL
XSFILL59080x21050 gnd vdd FILL
XFILL_2__12040_ gnd vdd FILL
X_10887_ _10887_/A _10888_/B _10887_/C gnd _10889_/B vdd OAI21X1
XFILL_0__10431_ gnd vdd FILL
XFILL_2__8983_ gnd vdd FILL
XFILL_5__7712_ gnd vdd FILL
XFILL_3__11591_ gnd vdd FILL
X_15414_ _15414_/A _15414_/B _14265_/C gnd _12848_/B vdd AOI21X1
XFILL_1__12770_ gnd vdd FILL
XFILL_0_BUFX2_insert500 gnd vdd FILL
XFILL_6__13510_ gnd vdd FILL
XFILL_0_BUFX2_insert511 gnd vdd FILL
X_12626_ _12626_/A vdd _12626_/C gnd _12682_/D vdd OAI21X1
XFILL_5__12151_ gnd vdd FILL
XFILL_3__13330_ gnd vdd FILL
XFILL_0_BUFX2_insert522 gnd vdd FILL
XFILL_4__11901_ gnd vdd FILL
X_16394_ gnd gnd gnd _16394_/Y vdd NAND2X1
XFILL_4__9899_ gnd vdd FILL
XFILL_0_BUFX2_insert533 gnd vdd FILL
XFILL_3__10542_ gnd vdd FILL
XFILL_4__12881_ gnd vdd FILL
XFILL_2__7934_ gnd vdd FILL
XFILL_0__13150_ gnd vdd FILL
XFILL112280x27050 gnd vdd FILL
XFILL_1__11721_ gnd vdd FILL
XFILL_0_BUFX2_insert544 gnd vdd FILL
XFILL_5__11102_ gnd vdd FILL
XFILL_0__10362_ gnd vdd FILL
X_15345_ _15899_/A _15345_/B _15899_/C _13793_/Y gnd _15347_/A vdd OAI22X1
XFILL_0_BUFX2_insert555 gnd vdd FILL
XFILL_4__14620_ gnd vdd FILL
XFILL_0_BUFX2_insert566 gnd vdd FILL
XFILL_5__12082_ gnd vdd FILL
X_12557_ _12409_/A _13175_/CLK _13199_/R vdd _12557_/D gnd vdd DFFSR
XFILL_4__11832_ gnd vdd FILL
XFILL_3__13261_ gnd vdd FILL
XFILL_0__12101_ gnd vdd FILL
XFILL_0_BUFX2_insert577 gnd vdd FILL
XFILL_2__7865_ gnd vdd FILL
XFILL_1__14440_ gnd vdd FILL
XFILL_0__13081_ gnd vdd FILL
XFILL_2__13991_ gnd vdd FILL
XFILL_0_BUFX2_insert588 gnd vdd FILL
XFILL_1__11652_ gnd vdd FILL
XFILL_0__10293_ gnd vdd FILL
XFILL_5__15910_ gnd vdd FILL
XFILL_3__15000_ gnd vdd FILL
XFILL_0_BUFX2_insert599 gnd vdd FILL
X_11508_ _11621_/C gnd _11846_/C vdd INVX8
XFILL_5__7574_ gnd vdd FILL
XFILL_6__16160_ gnd vdd FILL
XFILL_5__11033_ gnd vdd FILL
XFILL_2__9604_ gnd vdd FILL
XFILL_6__13372_ gnd vdd FILL
XFILL_3__12212_ gnd vdd FILL
X_15276_ _16141_/A _15276_/B _16141_/C gnd _15276_/Y vdd NOR3X1
XFILL_4__14551_ gnd vdd FILL
XFILL_2__15730_ gnd vdd FILL
X_12488_ vdd _12053_/A gnd _12488_/Y vdd NAND2X1
XFILL_0__6880_ gnd vdd FILL
XSFILL113560x15050 gnd vdd FILL
XFILL_4__11763_ gnd vdd FILL
XFILL_0__12032_ gnd vdd FILL
XSFILL79240x34050 gnd vdd FILL
XFILL_1__14371_ gnd vdd FILL
XFILL_1__11583_ gnd vdd FILL
X_14227_ _14227_/A _14227_/B _14224_/Y gnd _14243_/A vdd NAND3X1
XSFILL113800x77050 gnd vdd FILL
XFILL_5__15841_ gnd vdd FILL
X_11439_ _11490_/A _11433_/Y _11331_/B gnd _11439_/Y vdd AOI21X1
XFILL_4__13502_ gnd vdd FILL
XFILL_4__14482_ gnd vdd FILL
XFILL_2__9535_ gnd vdd FILL
XFILL_1__16110_ gnd vdd FILL
XFILL_3__12143_ gnd vdd FILL
XFILL_1__10534_ gnd vdd FILL
XFILL_1__13322_ gnd vdd FILL
XFILL_2__15661_ gnd vdd FILL
XFILL_4__11694_ gnd vdd FILL
XSFILL69160x7050 gnd vdd FILL
XFILL_5__9244_ gnd vdd FILL
XFILL_2__12873_ gnd vdd FILL
XFILL_4__16221_ gnd vdd FILL
XCLKBUF1_insert201 CLKBUF1_insert218/A gnd _7411_/CLK vdd CLKBUF1
X_14158_ _16363_/A gnd _14160_/A vdd INVX1
XFILL_4__13433_ gnd vdd FILL
XFILL_6__12254_ gnd vdd FILL
XCLKBUF1_insert212 CLKBUF1_insert206/A gnd _8171_/CLK vdd CLKBUF1
XFILL_2__14612_ gnd vdd FILL
XFILL_5__15772_ gnd vdd FILL
XFILL_4__10645_ gnd vdd FILL
XFILL_1__16041_ gnd vdd FILL
XFILL_3__12074_ gnd vdd FILL
XFILL_5__12984_ gnd vdd FILL
XFILL_2__11824_ gnd vdd FILL
XFILL_2__9466_ gnd vdd FILL
XCLKBUF1_insert223 CLKBUF1_insert192/A gnd _8921_/CLK vdd CLKBUF1
XFILL_1__13253_ gnd vdd FILL
XFILL_2__15592_ gnd vdd FILL
XSFILL84360x25050 gnd vdd FILL
XFILL_0__7501_ gnd vdd FILL
X_13109_ _13185_/Q gnd _13111_/A vdd INVX1
XFILL_6__11205_ gnd vdd FILL
XFILL_0__13983_ gnd vdd FILL
XFILL_5__14723_ gnd vdd FILL
XFILL_4__13364_ gnd vdd FILL
XFILL_3__15902_ gnd vdd FILL
XFILL_0__8481_ gnd vdd FILL
XFILL_5__11935_ gnd vdd FILL
X_14089_ _10595_/Q gnd _14089_/Y vdd INVX1
XFILL_3__11025_ gnd vdd FILL
XFILL_4__16152_ gnd vdd FILL
XFILL_3__7210_ gnd vdd FILL
XFILL_1__12204_ gnd vdd FILL
XFILL_2__14543_ gnd vdd FILL
XFILL_4__10576_ gnd vdd FILL
XFILL_5__8126_ gnd vdd FILL
XFILL_2__9397_ gnd vdd FILL
XFILL_0__15722_ gnd vdd FILL
XFILL_3__8190_ gnd vdd FILL
XFILL_2__11755_ gnd vdd FILL
XFILL_1__10396_ gnd vdd FILL
XFILL_0__7432_ gnd vdd FILL
XFILL_4__12315_ gnd vdd FILL
XFILL_4__15103_ gnd vdd FILL
XFILL_5__14654_ gnd vdd FILL
XFILL_4__16083_ gnd vdd FILL
XFILL_4__13295_ gnd vdd FILL
XFILL_2__8348_ gnd vdd FILL
XFILL_3__15833_ gnd vdd FILL
XFILL_5__11866_ gnd vdd FILL
XFILL_2__10706_ gnd vdd FILL
XFILL_2__14474_ gnd vdd FILL
XFILL_1__12135_ gnd vdd FILL
XFILL_0__15653_ gnd vdd FILL
XFILL_5__8057_ gnd vdd FILL
XSFILL18920x9050 gnd vdd FILL
XFILL_2__11686_ gnd vdd FILL
XFILL_5__13605_ gnd vdd FILL
XFILL_0__12865_ gnd vdd FILL
XFILL_2__16213_ gnd vdd FILL
XFILL_4__15034_ gnd vdd FILL
XFILL_4__12246_ gnd vdd FILL
XFILL_5__10817_ gnd vdd FILL
XFILL_6__11067_ gnd vdd FILL
XFILL_0__7363_ gnd vdd FILL
XFILL_5__14585_ gnd vdd FILL
XFILL_2__13425_ gnd vdd FILL
X_7991_ _7989_/Y _7948_/A _7991_/C gnd _8043_/D vdd OAI21X1
XFILL_2__10637_ gnd vdd FILL
XFILL_3__12976_ gnd vdd FILL
XFILL_0__14604_ gnd vdd FILL
XFILL_3__7072_ gnd vdd FILL
XFILL_1__12066_ gnd vdd FILL
XFILL_3__15764_ gnd vdd FILL
XFILL_5__11797_ gnd vdd FILL
XFILL_0__9102_ gnd vdd FILL
XFILL_0__11816_ gnd vdd FILL
XFILL_5__16324_ gnd vdd FILL
XFILL_0__15584_ gnd vdd FILL
X_9730_ _9818_/Q gnd _9732_/A vdd INVX1
XFILL_5__13536_ gnd vdd FILL
XFILL_3__14715_ gnd vdd FILL
XFILL_3__11927_ gnd vdd FILL
XSFILL109400x32050 gnd vdd FILL
X_6942_ _6985_/B _9374_/B gnd _6943_/C vdd NAND2X1
XFILL_5__10748_ gnd vdd FILL
XFILL_0__7294_ gnd vdd FILL
XFILL_4__12177_ gnd vdd FILL
XFILL_1__11017_ gnd vdd FILL
XFILL_2__16144_ gnd vdd FILL
XFILL_2__13356_ gnd vdd FILL
XFILL_3__15695_ gnd vdd FILL
XFILL_0__14535_ gnd vdd FILL
XFILL_2__10568_ gnd vdd FILL
XFILL_0__11747_ gnd vdd FILL
XFILL_0__9033_ gnd vdd FILL
XFILL_3_CLKBUF1_insert190 gnd vdd FILL
XSFILL49080x53050 gnd vdd FILL
XFILL_4__11128_ gnd vdd FILL
XSFILL79320x14050 gnd vdd FILL
XFILL_5__16255_ gnd vdd FILL
X_9661_ _9659_/Y _9639_/A _9660_/Y gnd _9709_/D vdd OAI21X1
XFILL112200x71050 gnd vdd FILL
XFILL_5__13467_ gnd vdd FILL
XFILL_2__12307_ gnd vdd FILL
X_6873_ _6873_/A gnd memoryWriteData[3] vdd BUFX2
XFILL_5__10679_ gnd vdd FILL
XFILL_3__14646_ gnd vdd FILL
XFILL_1__15825_ gnd vdd FILL
XFILL_2__16075_ gnd vdd FILL
XFILL_3__11858_ gnd vdd FILL
XFILL_2__13287_ gnd vdd FILL
XFILL_0__14466_ gnd vdd FILL
XFILL_5__15206_ gnd vdd FILL
XFILL_2__10499_ gnd vdd FILL
XFILL_0__11678_ gnd vdd FILL
XFILL_5__8959_ gnd vdd FILL
X_8612_ _8567_/B _7972_/B gnd _8613_/C vdd NAND2X1
XFILL_5__12418_ gnd vdd FILL
XFILL_5__16186_ gnd vdd FILL
XFILL_2__15026_ gnd vdd FILL
XFILL_4__15936_ gnd vdd FILL
XFILL_3__10809_ gnd vdd FILL
XFILL_4__11059_ gnd vdd FILL
XFILL_3__14577_ gnd vdd FILL
XFILL_0__16205_ gnd vdd FILL
XFILL_5__13398_ gnd vdd FILL
X_9592_ _9590_/Y _9675_/A _9591_/Y gnd _9686_/D vdd OAI21X1
XFILL_2__12238_ gnd vdd FILL
XSFILL114520x23050 gnd vdd FILL
XFILL_3__7974_ gnd vdd FILL
XFILL_0__13417_ gnd vdd FILL
XFILL_0__10629_ gnd vdd FILL
XFILL_3__11789_ gnd vdd FILL
XFILL_1__15756_ gnd vdd FILL
XFILL_0__14397_ gnd vdd FILL
XFILL_1__12968_ gnd vdd FILL
XFILL_5__15137_ gnd vdd FILL
XFILL_5__12349_ gnd vdd FILL
XFILL_3__16316_ gnd vdd FILL
X_8543_ _8465_/A _9716_/CLK _8682_/R vdd _8543_/D gnd vdd DFFSR
XFILL_3__13528_ gnd vdd FILL
XFILL_3__6925_ gnd vdd FILL
XFILL_5_BUFX2_insert705 gnd vdd FILL
XFILL_1__14707_ gnd vdd FILL
XFILL_4__15867_ gnd vdd FILL
XFILL_5_BUFX2_insert716 gnd vdd FILL
XFILL_1__11919_ gnd vdd FILL
XFILL_2__12169_ gnd vdd FILL
XFILL_0__16136_ gnd vdd FILL
XFILL_0__13348_ gnd vdd FILL
XFILL_5_BUFX2_insert727 gnd vdd FILL
XFILL_1__15687_ gnd vdd FILL
XFILL_0__9935_ gnd vdd FILL
XFILL_5_BUFX2_insert738 gnd vdd FILL
XFILL_1__12899_ gnd vdd FILL
XFILL_5_BUFX2_insert749 gnd vdd FILL
XFILL_4__14818_ gnd vdd FILL
XFILL_5__15068_ gnd vdd FILL
XSFILL3560x9050 gnd vdd FILL
XSFILL69240x66050 gnd vdd FILL
XFILL_3__13459_ gnd vdd FILL
X_8474_ _8474_/A gnd _8474_/Y vdd INVX1
XFILL_3__9644_ gnd vdd FILL
XFILL_3__16247_ gnd vdd FILL
XFILL_1__14638_ gnd vdd FILL
XFILL_3__6856_ gnd vdd FILL
XFILL_4__15798_ gnd vdd FILL
XFILL_0__13279_ gnd vdd FILL
XFILL_6__9353_ gnd vdd FILL
XFILL_0__16067_ gnd vdd FILL
XFILL_5__14019_ gnd vdd FILL
X_7425_ _7425_/A _7425_/B _7424_/Y gnd _7425_/Y vdd OAI21X1
XFILL_0__9866_ gnd vdd FILL
XFILL_3__16178_ gnd vdd FILL
XFILL_4__14749_ gnd vdd FILL
XFILL_2__15928_ gnd vdd FILL
XFILL_0__15018_ gnd vdd FILL
XFILL_1__14569_ gnd vdd FILL
XSFILL104440x75050 gnd vdd FILL
XFILL_1__7610_ gnd vdd FILL
XFILL_3__15129_ gnd vdd FILL
XFILL_1__8590_ gnd vdd FILL
XFILL_3__8526_ gnd vdd FILL
X_7356_ _7336_/B _8764_/B gnd _7356_/Y vdd NAND2X1
XFILL_1__16308_ gnd vdd FILL
XFILL_0__9797_ gnd vdd FILL
XSFILL8680x73050 gnd vdd FILL
XSFILL23720x22050 gnd vdd FILL
XFILL_2__15859_ gnd vdd FILL
XFILL_0__8748_ gnd vdd FILL
X_7287_ _8567_/A _7359_/A gnd _7288_/C vdd NAND2X1
XFILL_1__16239_ gnd vdd FILL
XFILL_3__8457_ gnd vdd FILL
XFILL_4__7250_ gnd vdd FILL
XSFILL49160x33050 gnd vdd FILL
X_9026_ _9011_/A _9794_/B gnd _9027_/C vdd NAND2X1
XFILL_1__7472_ gnd vdd FILL
XFILL_4__7181_ gnd vdd FILL
XFILL_3__8388_ gnd vdd FILL
XFILL_1__9211_ gnd vdd FILL
XFILL_6__8097_ gnd vdd FILL
XFILL_3__7339_ gnd vdd FILL
XFILL_2_BUFX2_insert606 gnd vdd FILL
XSFILL13640x74050 gnd vdd FILL
XFILL_6__7048_ gnd vdd FILL
XFILL_2_BUFX2_insert617 gnd vdd FILL
XFILL_1__9142_ gnd vdd FILL
XFILL_2_BUFX2_insert628 gnd vdd FILL
XFILL_2_BUFX2_insert639 gnd vdd FILL
XFILL_3__9009_ gnd vdd FILL
X_9928_ _9941_/B _7240_/B gnd _9928_/Y vdd NAND2X1
XSFILL29320x62050 gnd vdd FILL
X_10810_ _10810_/A _10809_/A _10810_/C gnd _10860_/D vdd OAI21X1
X_11790_ _11762_/B _11790_/B _11790_/C gnd _11799_/B vdd NOR3X1
X_9859_ _9868_/A _9859_/B gnd _9859_/Y vdd NAND2X1
XSFILL104520x55050 gnd vdd FILL
XSFILL8760x53050 gnd vdd FILL
X_10741_ _10741_/Q _7537_/CLK _7537_/R vdd _10709_/Y gnd vdd DFFSR
XBUFX2_insert605 BUFX2_insert518/A gnd _7915_/R vdd BUFX2
XFILL_4__6965_ gnd vdd FILL
XFILL_4__9753_ gnd vdd FILL
XBUFX2_insert616 _10926_/Y gnd _11987_/A vdd BUFX2
XFILL_6_BUFX2_insert561 gnd vdd FILL
X_13460_ _13381_/A _13418_/A _13423_/B gnd _13460_/Y vdd NAND3X1
XBUFX2_insert627 _13465_/Y gnd _14640_/C vdd BUFX2
XFILL_6_BUFX2_insert572 gnd vdd FILL
X_10672_ _10681_/A _8496_/B gnd _10673_/C vdd NAND2X1
XFILL_1__9975_ gnd vdd FILL
XBUFX2_insert638 _12438_/Y gnd _7508_/B vdd BUFX2
XFILL_4__8704_ gnd vdd FILL
XBUFX2_insert649 _10915_/Y gnd _12012_/A vdd BUFX2
X_12411_ _12409_/Y _12371_/A _12411_/C gnd _12411_/Y vdd OAI21X1
XFILL_4__9684_ gnd vdd FILL
XFILL_4__6896_ gnd vdd FILL
X_13391_ _12808_/Q _12807_/Q gnd _13404_/B vdd AND2X2
XSFILL79160x2050 gnd vdd FILL
XFILL_4__8635_ gnd vdd FILL
XSFILL110280x12050 gnd vdd FILL
XSFILL53720x38050 gnd vdd FILL
X_15130_ _15916_/B _15130_/B _7548_/A _15087_/B gnd _15130_/Y vdd AOI22X1
X_12342_ _12342_/A _12342_/B _12342_/C gnd _10988_/B vdd NAND3X1
XFILL_1__8857_ gnd vdd FILL
XSFILL13720x54050 gnd vdd FILL
XFILL_4__8566_ gnd vdd FILL
X_15061_ _12767_/A _16216_/B _15061_/C gnd _15061_/Y vdd NAND3X1
XFILL_1__7808_ gnd vdd FILL
X_12273_ _6884_/A _12249_/B _12249_/C _11876_/B gnd _12274_/C vdd AOI22X1
XFILL_2__7581_ gnd vdd FILL
XSFILL39480x3050 gnd vdd FILL
XFILL_1__8788_ gnd vdd FILL
X_14012_ _14012_/A _14012_/B _14012_/C gnd _14023_/A vdd NAND3X1
XFILL_4__8497_ gnd vdd FILL
XFILL_5__7290_ gnd vdd FILL
X_11224_ gnd _10896_/Y gnd _11224_/Y vdd NOR2X1
XSFILL79640x8050 gnd vdd FILL
XFILL_1__7739_ gnd vdd FILL
XSFILL28920x4050 gnd vdd FILL
XFILL_4__7448_ gnd vdd FILL
XFILL_4__10430_ gnd vdd FILL
X_11155_ _11153_/Y _11129_/Y _11154_/Y gnd _11407_/C vdd AOI21X1
XFILL_2__9251_ gnd vdd FILL
XFILL_1__10250_ gnd vdd FILL
XFILL_3_BUFX2_insert440 gnd vdd FILL
XFILL_3_BUFX2_insert451 gnd vdd FILL
XFILL_0__10980_ gnd vdd FILL
XFILL_4__7379_ gnd vdd FILL
X_10106_ _10106_/A _9978_/B gnd _10107_/C vdd NAND2X1
XFILL_2__8202_ gnd vdd FILL
XFILL_3_BUFX2_insert462 gnd vdd FILL
XFILL_5__11720_ gnd vdd FILL
XFILL_1__9409_ gnd vdd FILL
X_15963_ _9144_/A gnd _15964_/B vdd INVX1
XFILL_4__10361_ gnd vdd FILL
X_11086_ _11086_/A _11388_/B _11085_/Y gnd _11086_/Y vdd OAI21X1
XSFILL59080x16050 gnd vdd FILL
XFILL_3_BUFX2_insert473 gnd vdd FILL
XFILL_4__9118_ gnd vdd FILL
XFILL_2__11540_ gnd vdd FILL
XFILL_1__10181_ gnd vdd FILL
XFILL_3_BUFX2_insert484 gnd vdd FILL
XFILL_4__12100_ gnd vdd FILL
XFILL_3_BUFX2_insert495 gnd vdd FILL
XSFILL99480x21050 gnd vdd FILL
X_10037_ _10091_/Q gnd _10039_/A vdd INVX1
X_14914_ _7504_/A gnd _14914_/Y vdd INVX1
X_15894_ _14477_/Y _15169_/A gnd _15896_/C vdd NOR2X1
XFILL_4__13080_ gnd vdd FILL
XFILL_2__8133_ gnd vdd FILL
XFILL_5__11651_ gnd vdd FILL
XFILL_3__12830_ gnd vdd FILL
XFILL_4__10292_ gnd vdd FILL
XFILL_0__12650_ gnd vdd FILL
XFILL_2__11471_ gnd vdd FILL
XFILL_5__9931_ gnd vdd FILL
XFILL_4__12031_ gnd vdd FILL
XFILL_2__13210_ gnd vdd FILL
X_14845_ _14844_/Y _14841_/Y gnd _14846_/C vdd NOR2X1
XFILL_5__14370_ gnd vdd FILL
XFILL_5__11582_ gnd vdd FILL
XFILL_2__10422_ gnd vdd FILL
XFILL_3__12761_ gnd vdd FILL
XFILL_2__8064_ gnd vdd FILL
XFILL_2__14190_ gnd vdd FILL
XFILL_0__11601_ gnd vdd FILL
XFILL_1__13940_ gnd vdd FILL
XFILL_0__12581_ gnd vdd FILL
XFILL_5__13321_ gnd vdd FILL
XFILL_5__9862_ gnd vdd FILL
XFILL_5__10533_ gnd vdd FILL
XFILL_3__14500_ gnd vdd FILL
XFILL_6__12872_ gnd vdd FILL
XFILL_0_BUFX2_insert1 gnd vdd FILL
XSFILL13800x34050 gnd vdd FILL
XFILL_3__11712_ gnd vdd FILL
X_14776_ _14776_/A gnd _14778_/A vdd INVX1
XFILL_2__13141_ gnd vdd FILL
X_11988_ _12007_/A _11988_/B gnd _11988_/Y vdd AND2X2
XFILL_3__15480_ gnd vdd FILL
XFILL_0__14320_ gnd vdd FILL
XSFILL79240x29050 gnd vdd FILL
XFILL_0__11532_ gnd vdd FILL
XFILL_1__13871_ gnd vdd FILL
XFILL_5__16040_ gnd vdd FILL
X_13727_ _13717_/Y _13719_/Y _13726_/Y gnd _13727_/Y vdd NAND3X1
XFILL_5__13252_ gnd vdd FILL
X_10939_ _12785_/A gnd _10939_/Y vdd INVX1
XFILL_5__9793_ gnd vdd FILL
XFILL_3__14431_ gnd vdd FILL
XFILL_3__11643_ gnd vdd FILL
XFILL_1__15610_ gnd vdd FILL
XSFILL64040x71050 gnd vdd FILL
XFILL_0__14251_ gnd vdd FILL
XFILL_4__13982_ gnd vdd FILL
XFILL_2__10284_ gnd vdd FILL
XFILL_0__11463_ gnd vdd FILL
XFILL_5__8744_ gnd vdd FILL
XFILL_5__12203_ gnd vdd FILL
X_16446_ _16408_/A _8306_/CLK _9054_/R vdd _16410_/Y gnd vdd DFFSR
XFILL_4__15721_ gnd vdd FILL
X_13658_ _13657_/Y _14567_/A _14862_/C _15211_/A gnd _13662_/B vdd OAI22X1
XSFILL3080x57050 gnd vdd FILL
XFILL_2__12023_ gnd vdd FILL
XFILL_5__10395_ gnd vdd FILL
XFILL_3__14362_ gnd vdd FILL
XFILL_1__15541_ gnd vdd FILL
XFILL_0__10414_ gnd vdd FILL
XFILL_2__8966_ gnd vdd FILL
XFILL_3__11574_ gnd vdd FILL
XFILL_0__14182_ gnd vdd FILL
XFILL_1__12753_ gnd vdd FILL
XFILL_0_BUFX2_insert330 gnd vdd FILL
X_12609_ _12609_/A gnd _12611_/A vdd INVX1
XFILL_0_BUFX2_insert341 gnd vdd FILL
XFILL_0__11394_ gnd vdd FILL
XFILL_3__13313_ gnd vdd FILL
XFILL_5__12134_ gnd vdd FILL
XFILL_3__16101_ gnd vdd FILL
X_16377_ _16375_/Y gnd _16377_/C gnd _16435_/D vdd OAI21X1
XFILL_0_BUFX2_insert352 gnd vdd FILL
XFILL_4__15652_ gnd vdd FILL
X_13589_ _9689_/Q gnd _13590_/C vdd INVX1
XFILL_0__7981_ gnd vdd FILL
XFILL_3__10525_ gnd vdd FILL
XFILL_0__13133_ gnd vdd FILL
XFILL_1__11704_ gnd vdd FILL
XFILL_0_BUFX2_insert363 gnd vdd FILL
XFILL_4__12864_ gnd vdd FILL
XFILL_3__14293_ gnd vdd FILL
XFILL_3__7690_ gnd vdd FILL
XFILL_6__16212_ gnd vdd FILL
XFILL_2__8897_ gnd vdd FILL
XFILL_1__15472_ gnd vdd FILL
XFILL_0_BUFX2_insert374 gnd vdd FILL
XFILL_0_BUFX2_insert385 gnd vdd FILL
X_15328_ _13764_/Y _15328_/B _15683_/C _15328_/D gnd _15329_/A vdd OAI22X1
XFILL_0__9720_ gnd vdd FILL
XFILL_5__7626_ gnd vdd FILL
XFILL_6__10636_ gnd vdd FILL
XFILL_4__14603_ gnd vdd FILL
XFILL_3__16032_ gnd vdd FILL
XFILL_0_BUFX2_insert396 gnd vdd FILL
XFILL_5__12065_ gnd vdd FILL
XFILL_0__6932_ gnd vdd FILL
XFILL_3__13244_ gnd vdd FILL
XFILL_4__11815_ gnd vdd FILL
XFILL_2__7848_ gnd vdd FILL
XFILL_4__15583_ gnd vdd FILL
XFILL_1__14423_ gnd vdd FILL
XFILL_1__11635_ gnd vdd FILL
XFILL_2__13974_ gnd vdd FILL
XFILL_0__10276_ gnd vdd FILL
XFILL_5__7557_ gnd vdd FILL
XFILL_5__11016_ gnd vdd FILL
X_15259_ _15258_/Y _15259_/B _14597_/C gnd _12836_/B vdd AOI21X1
XFILL_0__9651_ gnd vdd FILL
X_7210_ _7210_/A _9258_/B gnd _7211_/C vdd NAND2X1
XFILL_0__6863_ gnd vdd FILL
XFILL_4__14534_ gnd vdd FILL
X_8190_ _8190_/A _8187_/B _8189_/Y gnd _8280_/D vdd OAI21X1
XFILL_3__9360_ gnd vdd FILL
XFILL_2__15713_ gnd vdd FILL
XFILL_0__12015_ gnd vdd FILL
XFILL_4__11746_ gnd vdd FILL
XFILL_1__14354_ gnd vdd FILL
XFILL_3__10387_ gnd vdd FILL
XFILL_0__8602_ gnd vdd FILL
XFILL_1__11566_ gnd vdd FILL
X_7141_ _7141_/Q _8926_/CLK _7262_/R vdd _7077_/Y gnd vdd DFFSR
XFILL_5__7488_ gnd vdd FILL
XSFILL59000x60050 gnd vdd FILL
XFILL_5__15824_ gnd vdd FILL
XFILL_3__12126_ gnd vdd FILL
XFILL_3__8311_ gnd vdd FILL
XFILL_1__13305_ gnd vdd FILL
XFILL_4__14465_ gnd vdd FILL
XFILL_2__15644_ gnd vdd FILL
XFILL_2__9518_ gnd vdd FILL
XSFILL109400x27050 gnd vdd FILL
XFILL_4__11677_ gnd vdd FILL
XFILL_3__9291_ gnd vdd FILL
XFILL_2__12856_ gnd vdd FILL
XFILL_1__10517_ gnd vdd FILL
XFILL_5__9227_ gnd vdd FILL
XFILL_6__15025_ gnd vdd FILL
XFILL_1__14285_ gnd vdd FILL
XFILL_4__16204_ gnd vdd FILL
XFILL_0__8533_ gnd vdd FILL
XFILL_1__11497_ gnd vdd FILL
X_7072_ _7072_/A gnd _7074_/A vdd INVX1
XFILL_4__13416_ gnd vdd FILL
XSFILL49080x48050 gnd vdd FILL
XFILL_4__10628_ gnd vdd FILL
XFILL_5__15755_ gnd vdd FILL
XFILL112200x66050 gnd vdd FILL
XFILL_1__16024_ gnd vdd FILL
XFILL_5_BUFX2_insert1020 gnd vdd FILL
XFILL_3__12057_ gnd vdd FILL
XFILL_2__11807_ gnd vdd FILL
XFILL_3__8242_ gnd vdd FILL
XFILL_5__12967_ gnd vdd FILL
XFILL_1__13236_ gnd vdd FILL
XFILL_4__14396_ gnd vdd FILL
XFILL_2__15575_ gnd vdd FILL
XFILL_2__12787_ gnd vdd FILL
XFILL_5__9158_ gnd vdd FILL
XFILL_5_BUFX2_insert1031 gnd vdd FILL
XFILL_1__10448_ gnd vdd FILL
XFILL_5_BUFX2_insert1042 gnd vdd FILL
XFILL_5__14706_ gnd vdd FILL
XFILL_0__13966_ gnd vdd FILL
XFILL_0__8464_ gnd vdd FILL
XFILL_5_BUFX2_insert1053 gnd vdd FILL
XSFILL64120x51050 gnd vdd FILL
XFILL_5__11918_ gnd vdd FILL
XFILL_4__16135_ gnd vdd FILL
XFILL_3__11008_ gnd vdd FILL
XFILL_4__13347_ gnd vdd FILL
XFILL_4__10559_ gnd vdd FILL
XFILL_5__15686_ gnd vdd FILL
XFILL_5_BUFX2_insert1064 gnd vdd FILL
XFILL_2__14526_ gnd vdd FILL
XFILL_0__15705_ gnd vdd FILL
XFILL_5__8109_ gnd vdd FILL
XFILL_2__11738_ gnd vdd FILL
XFILL_5__12898_ gnd vdd FILL
XFILL_1__10379_ gnd vdd FILL
XFILL_1__13167_ gnd vdd FILL
XFILL_0__12917_ gnd vdd FILL
XFILL_5__9089_ gnd vdd FILL
XFILL_5_BUFX2_insert1086 gnd vdd FILL
XFILL_0__7415_ gnd vdd FILL
XFILL_5__14637_ gnd vdd FILL
XFILL_0__13897_ gnd vdd FILL
XFILL_4__13278_ gnd vdd FILL
XFILL_0__8395_ gnd vdd FILL
XFILL_3__7124_ gnd vdd FILL
XFILL_3__15816_ gnd vdd FILL
XFILL_4__16066_ gnd vdd FILL
XFILL_5__11849_ gnd vdd FILL
XFILL_2__14457_ gnd vdd FILL
XFILL_1__12118_ gnd vdd FILL
XFILL_0__15636_ gnd vdd FILL
XFILL_2__11669_ gnd vdd FILL
XFILL_0__12848_ gnd vdd FILL
XFILL_1__13098_ gnd vdd FILL
XFILL_4__15017_ gnd vdd FILL
XFILL_4__12229_ gnd vdd FILL
XFILL_0__7346_ gnd vdd FILL
XFILL_5__14568_ gnd vdd FILL
XFILL_2__13408_ gnd vdd FILL
X_7974_ _8038_/Q gnd _7976_/A vdd INVX1
XFILL_3__7055_ gnd vdd FILL
XFILL_3__15747_ gnd vdd FILL
XFILL_1__12049_ gnd vdd FILL
XFILL_2__14388_ gnd vdd FILL
XFILL_3__12959_ gnd vdd FILL
XFILL_0__15567_ gnd vdd FILL
XFILL_5__16307_ gnd vdd FILL
XFILL_0__12779_ gnd vdd FILL
XSFILL28760x70050 gnd vdd FILL
X_9713_ _9671_/A _7537_/CLK _7537_/R vdd _9713_/D gnd vdd DFFSR
XFILL_5__13519_ gnd vdd FILL
X_6925_ _6923_/Y _6967_/B _6925_/C gnd _6925_/Y vdd OAI21X1
XFILL_2__16127_ gnd vdd FILL
XFILL_2__13339_ gnd vdd FILL
XFILL_5__14499_ gnd vdd FILL
XFILL_3__15678_ gnd vdd FILL
XFILL_0__14518_ gnd vdd FILL
XFILL_0__9016_ gnd vdd FILL
XFILL_5__16238_ gnd vdd FILL
XFILL_0__15498_ gnd vdd FILL
X_9644_ _9644_/A gnd _9644_/Y vdd INVX1
XFILL_6__8784_ gnd vdd FILL
XFILL_3__14629_ gnd vdd FILL
X_6856_ _6856_/A gnd memoryAddress[18] vdd BUFX2
XFILL_1__15808_ gnd vdd FILL
XFILL_3_BUFX2_insert1090 gnd vdd FILL
XFILL_2__16058_ gnd vdd FILL
XSFILL8680x68050 gnd vdd FILL
XSFILL23720x17050 gnd vdd FILL
XFILL_0__14449_ gnd vdd FILL
XFILL_6__7735_ gnd vdd FILL
XFILL_4__15919_ gnd vdd FILL
XSFILL33880x61050 gnd vdd FILL
XFILL_5__16169_ gnd vdd FILL
XFILL_2__15009_ gnd vdd FILL
X_9575_ _9575_/Q _8551_/CLK _7015_/R vdd _9515_/Y gnd vdd DFFSR
XFILL_1__15739_ gnd vdd FILL
XFILL_5_BUFX2_insert502 gnd vdd FILL
XFILL_3__7957_ gnd vdd FILL
XFILL_5_BUFX2_insert513 gnd vdd FILL
X_8526_ _8503_/B _8526_/B gnd _8527_/C vdd NAND2X1
XFILL_1__9760_ gnd vdd FILL
XFILL_5_BUFX2_insert524 gnd vdd FILL
XSFILL48920x83050 gnd vdd FILL
XFILL_5_BUFX2_insert535 gnd vdd FILL
XFILL_1__6972_ gnd vdd FILL
XSFILL89560x33050 gnd vdd FILL
XSFILL54280x5050 gnd vdd FILL
XFILL_5_BUFX2_insert546 gnd vdd FILL
XFILL_0__16119_ gnd vdd FILL
XFILL_3__6908_ gnd vdd FILL
XFILL_6__9405_ gnd vdd FILL
XFILL_5_BUFX2_insert557 gnd vdd FILL
XSFILL64200x31050 gnd vdd FILL
XFILL_3__7888_ gnd vdd FILL
XFILL_5_BUFX2_insert568 gnd vdd FILL
XFILL_1__8711_ gnd vdd FILL
XFILL_0__9918_ gnd vdd FILL
XFILL_3_BUFX2_insert5 gnd vdd FILL
X_8457_ _8484_/A _9993_/B gnd _8458_/C vdd NAND2X1
XFILL_5_BUFX2_insert579 gnd vdd FILL
XFILL_3__9627_ gnd vdd FILL
XFILL_3__6839_ gnd vdd FILL
XSFILL13640x69050 gnd vdd FILL
X_7408_ _7364_/A _9328_/CLK _7408_/R vdd _7366_/Y gnd vdd DFFSR
XFILL_1__8642_ gnd vdd FILL
XSFILL28440x29050 gnd vdd FILL
XFILL_0__9849_ gnd vdd FILL
X_8388_ _8432_/Q gnd _8390_/A vdd INVX1
XFILL_4__8351_ gnd vdd FILL
XFILL_3_BUFX2_insert90 gnd vdd FILL
X_7339_ _7337_/Y _7323_/A _7339_/C gnd _7399_/D vdd OAI21X1
XFILL_1__8573_ gnd vdd FILL
XFILL_4__7302_ gnd vdd FILL
XFILL_3__8509_ gnd vdd FILL
XFILL_2_CLKBUF1_insert116 gnd vdd FILL
XFILL_3__9489_ gnd vdd FILL
XSFILL54120x83050 gnd vdd FILL
XFILL_2_CLKBUF1_insert127 gnd vdd FILL
XFILL_2_CLKBUF1_insert138 gnd vdd FILL
XFILL_2_CLKBUF1_insert149 gnd vdd FILL
XFILL_4__7233_ gnd vdd FILL
X_9009_ _9009_/A _9017_/A _9008_/Y gnd _9009_/Y vdd OAI21X1
XSFILL8760x48050 gnd vdd FILL
XFILL_1__7455_ gnd vdd FILL
XFILL_4__7164_ gnd vdd FILL
XFILL_2_BUFX2_insert403 gnd vdd FILL
XSFILL33960x41050 gnd vdd FILL
X_12960_ _6873_/A gnd _12960_/Y vdd INVX1
XFILL_2_BUFX2_insert414 gnd vdd FILL
XFILL_2_BUFX2_insert425 gnd vdd FILL
XFILL_2_BUFX2_insert436 gnd vdd FILL
XFILL_4__7095_ gnd vdd FILL
X_11911_ _13103_/A gnd _11913_/A vdd INVX1
XFILL_2_BUFX2_insert447 gnd vdd FILL
XFILL_1__9125_ gnd vdd FILL
XFILL_2_BUFX2_insert458 gnd vdd FILL
X_12891_ _12889_/Y vdd _12891_/C gnd _12941_/D vdd OAI21X1
XFILL_2_BUFX2_insert469 gnd vdd FILL
X_14630_ _14630_/A _14630_/B _14625_/Y gnd _14646_/B vdd NAND3X1
X_11842_ _12218_/Y _11009_/Y gnd _11845_/B vdd NOR2X1
XSFILL13720x49050 gnd vdd FILL
X_14561_ _9837_/Q _14213_/A _14214_/C _10043_/A gnd _14561_/Y vdd AOI22X1
XFILL_1__8007_ gnd vdd FILL
X_11773_ _11772_/Y _11763_/Y gnd _11774_/A vdd NOR2X1
XFILL_4__9805_ gnd vdd FILL
X_16300_ _7029_/Q gnd _16301_/C vdd INVX1
X_13512_ _7895_/Q gnd _13514_/C vdd INVX1
XBUFX2_insert402 _10920_/Y gnd _12407_/A vdd BUFX2
X_10724_ _10656_/A _9818_/CLK _9441_/R vdd _10724_/D gnd vdd DFFSR
X_14492_ _9579_/Q gnd _14492_/Y vdd INVX1
XFILL_4__7997_ gnd vdd FILL
XBUFX2_insert413 _13484_/Y gnd _14877_/D vdd BUFX2
XBUFX2_insert424 _14991_/Y gnd _15202_/B vdd BUFX2
XSFILL28920x30050 gnd vdd FILL
XBUFX2_insert435 _13326_/Y gnd _8753_/B vdd BUFX2
X_16231_ _16231_/A _16231_/B gnd _16231_/Y vdd NAND2X1
XFILL_4__9736_ gnd vdd FILL
XBUFX2_insert446 _12378_/Y gnd _9624_/B vdd BUFX2
XFILL_4__6948_ gnd vdd FILL
X_13443_ _13443_/A _13423_/B _13718_/B gnd _13443_/Y vdd NAND3X1
XFILL_5__10180_ gnd vdd FILL
XBUFX2_insert457 _13442_/Y gnd _14342_/B vdd BUFX2
X_10655_ _10655_/A _10619_/B _10655_/C gnd _10723_/D vdd OAI21X1
XBUFX2_insert468 _13318_/Y gnd _8360_/B vdd BUFX2
XFILL_2__8751_ gnd vdd FILL
XBUFX2_insert479 _15038_/Y gnd _16311_/A vdd BUFX2
XFILL_5__8460_ gnd vdd FILL
XFILL_4__9667_ gnd vdd FILL
XFILL_4__6879_ gnd vdd FILL
X_16162_ _16161_/Y _16162_/B gnd _16162_/Y vdd NAND2X1
X_13374_ _15002_/C _14868_/A _14180_/C _10486_/A gnd _13374_/Y vdd AOI22X1
XFILL_3__10310_ gnd vdd FILL
XFILL_2__7702_ gnd vdd FILL
XFILL_1__8909_ gnd vdd FILL
X_10586_ _13682_/B _9818_/CLK _9441_/R vdd _10500_/Y gnd vdd DFFSR
XFILL_3__11290_ gnd vdd FILL
XFILL_0__10130_ gnd vdd FILL
XFILL_1__9889_ gnd vdd FILL
XSFILL34520x28050 gnd vdd FILL
X_15113_ _15113_/A _15113_/B gnd _15126_/C vdd NAND2X1
XFILL_4__8618_ gnd vdd FILL
XSFILL99480x16050 gnd vdd FILL
XFILL_5__8391_ gnd vdd FILL
X_12325_ _6897_/A _12289_/B _12289_/C _12297_/D gnd _12326_/C vdd AOI22X1
X_16093_ _16093_/A _16093_/B _16093_/C gnd _16093_/Y vdd NOR3X1
XFILL_4__9598_ gnd vdd FILL
XFILL_4__11600_ gnd vdd FILL
XFILL_3__10241_ gnd vdd FILL
XFILL_4__12580_ gnd vdd FILL
XSFILL74120x14050 gnd vdd FILL
XFILL_2__7633_ gnd vdd FILL
XFILL_1__11420_ gnd vdd FILL
XSFILL18840x82050 gnd vdd FILL
XFILL_2__10971_ gnd vdd FILL
XFILL_0__10061_ gnd vdd FILL
XFILL_5__7342_ gnd vdd FILL
X_15044_ _15244_/C _14981_/Y _15044_/C gnd _15044_/Y vdd NAND3X1
X_12256_ _12272_/A _12801_/Q _12248_/C gnd _12258_/B vdd NAND3X1
XFILL_4__11531_ gnd vdd FILL
XFILL_5__13870_ gnd vdd FILL
XFILL_2__12710_ gnd vdd FILL
XFILL_3__10172_ gnd vdd FILL
XFILL_2__7564_ gnd vdd FILL
XFILL_2__13690_ gnd vdd FILL
XFILL_1__11351_ gnd vdd FILL
X_11207_ _11419_/A _11207_/B _11206_/Y gnd _11212_/A vdd AOI21X1
XFILL_4__14250_ gnd vdd FILL
X_12187_ _11959_/A gnd _12187_/Y vdd INVX1
XFILL_4__11462_ gnd vdd FILL
XFILL_1__10302_ gnd vdd FILL
XFILL_2__12641_ gnd vdd FILL
XFILL_5__9012_ gnd vdd FILL
XFILL_0__13820_ gnd vdd FILL
XFILL_3__14980_ gnd vdd FILL
XFILL_1__14070_ gnd vdd FILL
XFILL_2__7495_ gnd vdd FILL
XFILL_1_BUFX2_insert19 gnd vdd FILL
XFILL_1__11282_ gnd vdd FILL
XSFILL23160x54050 gnd vdd FILL
XFILL_5__15540_ gnd vdd FILL
XFILL_4__10413_ gnd vdd FILL
X_11138_ _11634_/A _11137_/Y gnd _11138_/Y vdd NAND2X1
XFILL_5__12752_ gnd vdd FILL
XFILL_4__14181_ gnd vdd FILL
XFILL_6_BUFX2_insert9 gnd vdd FILL
XFILL_2__9234_ gnd vdd FILL
XFILL_1__13021_ gnd vdd FILL
XFILL_2__15360_ gnd vdd FILL
XFILL_4__11393_ gnd vdd FILL
XFILL_1__10233_ gnd vdd FILL
XFILL_3__13931_ gnd vdd FILL
XFILL_3_BUFX2_insert270 gnd vdd FILL
XFILL_2__12572_ gnd vdd FILL
XSFILL64040x66050 gnd vdd FILL
XFILL_3_BUFX2_insert281 gnd vdd FILL
XFILL_0__13751_ gnd vdd FILL
XFILL_0__10963_ gnd vdd FILL
XFILL_4__13132_ gnd vdd FILL
XFILL_5__11703_ gnd vdd FILL
XFILL_3_BUFX2_insert292 gnd vdd FILL
X_15946_ _15632_/A _14518_/D _15946_/C gnd _15946_/Y vdd OAI21X1
XFILL_2__14311_ gnd vdd FILL
X_11069_ _12262_/Y _12150_/Y gnd _11074_/C vdd XNOR2X1
XFILL_5__15471_ gnd vdd FILL
XFILL_2__9165_ gnd vdd FILL
XFILL_2__11523_ gnd vdd FILL
XFILL_0__12702_ gnd vdd FILL
XFILL_3__13862_ gnd vdd FILL
XFILL_1__10164_ gnd vdd FILL
XFILL_2__15291_ gnd vdd FILL
XFILL_0__7200_ gnd vdd FILL
XFILL_0__13682_ gnd vdd FILL
XFILL_0__10894_ gnd vdd FILL
XFILL_5__14422_ gnd vdd FILL
XFILL_2__8116_ gnd vdd FILL
XFILL_5__11634_ gnd vdd FILL
XFILL_3__15601_ gnd vdd FILL
XFILL_4__10275_ gnd vdd FILL
XFILL_2__14242_ gnd vdd FILL
XSFILL43880x24050 gnd vdd FILL
X_15877_ _15877_/A _15877_/B gnd _15890_/A vdd NAND2X1
XFILL_3__13793_ gnd vdd FILL
XFILL_2__9096_ gnd vdd FILL
XFILL_2__11454_ gnd vdd FILL
XFILL_0__15421_ gnd vdd FILL
XFILL_0__12633_ gnd vdd FILL
XFILL_2_BUFX2_insert970 gnd vdd FILL
XFILL_5__9914_ gnd vdd FILL
XFILL_1__14972_ gnd vdd FILL
XFILL_4__12014_ gnd vdd FILL
XFILL_2_BUFX2_insert981 gnd vdd FILL
XFILL_2_BUFX2_insert992 gnd vdd FILL
X_14828_ _9674_/A gnd _14830_/A vdd INVX1
XFILL_5__14353_ gnd vdd FILL
XFILL_3__12744_ gnd vdd FILL
XFILL_2__10405_ gnd vdd FILL
XFILL_3__15532_ gnd vdd FILL
XFILL_5__11565_ gnd vdd FILL
XFILL_2__14173_ gnd vdd FILL
XFILL_1__13923_ gnd vdd FILL
XFILL_0__15352_ gnd vdd FILL
XFILL_2__11385_ gnd vdd FILL
XFILL_5__13304_ gnd vdd FILL
XFILL_5__10516_ gnd vdd FILL
XFILL_0__7062_ gnd vdd FILL
XFILL_2__13124_ gnd vdd FILL
X_14759_ _9159_/A gnd _14760_/A vdd INVX1
XFILL_5__14284_ gnd vdd FILL
X_7690_ _7688_/Y _7690_/B _7690_/C gnd _7772_/D vdd OAI21X1
XFILL_3__8860_ gnd vdd FILL
XFILL_0__14303_ gnd vdd FILL
XFILL_3__15463_ gnd vdd FILL
XFILL_5__11496_ gnd vdd FILL
XFILL_1__13854_ gnd vdd FILL
XFILL_0__11515_ gnd vdd FILL
XFILL_5__16023_ gnd vdd FILL
XFILL_0__12495_ gnd vdd FILL
XFILL_0__15283_ gnd vdd FILL
XFILL_5__13235_ gnd vdd FILL
XSFILL59000x55050 gnd vdd FILL
XFILL_5__9776_ gnd vdd FILL
XFILL_5__10447_ gnd vdd FILL
XFILL_5__6988_ gnd vdd FILL
XFILL_3__11626_ gnd vdd FILL
XFILL_3__14414_ gnd vdd FILL
XFILL_3__7811_ gnd vdd FILL
XFILL_3__15394_ gnd vdd FILL
XFILL_4__13965_ gnd vdd FILL
XSFILL99400x60050 gnd vdd FILL
XFILL_0__14234_ gnd vdd FILL
XFILL_2__10267_ gnd vdd FILL
XFILL_0__11446_ gnd vdd FILL
XFILL_1__13785_ gnd vdd FILL
XFILL_5__8727_ gnd vdd FILL
XFILL_2__9998_ gnd vdd FILL
XFILL_4__15704_ gnd vdd FILL
X_16429_ _14043_/A _8680_/CLK _8034_/R vdd _16429_/D gnd vdd DFFSR
XFILL_6__11737_ gnd vdd FILL
XFILL_1__10997_ gnd vdd FILL
X_9360_ _9358_/Y _9359_/A _9360_/C gnd _9360_/Y vdd OAI21X1
XFILL_5__13166_ gnd vdd FILL
XFILL_5__10378_ gnd vdd FILL
XFILL_2__12006_ gnd vdd FILL
XFILL_3__14345_ gnd vdd FILL
XFILL_4__12916_ gnd vdd FILL
XFILL_3__7742_ gnd vdd FILL
XFILL_1__15524_ gnd vdd FILL
XFILL_3__11557_ gnd vdd FILL
XFILL_1__12736_ gnd vdd FILL
XFILL_4__13896_ gnd vdd FILL
XFILL_0__14165_ gnd vdd FILL
XSFILL89480x48050 gnd vdd FILL
XFILL_6__7451_ gnd vdd FILL
XBUFX2_insert980 _13455_/Y gnd _13456_/A vdd BUFX2
XFILL_0__11377_ gnd vdd FILL
XBUFX2_insert991 _12408_/Y gnd _7094_/B vdd BUFX2
X_8311_ _8951_/A _8356_/A gnd _8312_/C vdd NAND2X1
XFILL_5__12117_ gnd vdd FILL
XFILL_5__8658_ gnd vdd FILL
XFILL112360x20050 gnd vdd FILL
XFILL_3__10508_ gnd vdd FILL
XFILL_4__15635_ gnd vdd FILL
XSFILL64120x46050 gnd vdd FILL
XFILL_0__7964_ gnd vdd FILL
XFILL_4__12847_ gnd vdd FILL
XFILL_5__13097_ gnd vdd FILL
X_9291_ _9301_/B _8011_/B gnd _9292_/C vdd NAND2X1
XFILL_3__14276_ gnd vdd FILL
XFILL_0__13116_ gnd vdd FILL
XFILL_1__15455_ gnd vdd FILL
XFILL_3__7673_ gnd vdd FILL
XFILL_3__11488_ gnd vdd FILL
XFILL_5__7609_ gnd vdd FILL
XFILL_0__14096_ gnd vdd FILL
XFILL_4_BUFX2_insert509 gnd vdd FILL
XFILL_0__6915_ gnd vdd FILL
XFILL_3__13227_ gnd vdd FILL
XFILL_5__8589_ gnd vdd FILL
XFILL_3__16015_ gnd vdd FILL
XFILL_5__12048_ gnd vdd FILL
X_8242_ _8242_/A gnd _8242_/Y vdd INVX1
XFILL_3__9412_ gnd vdd FILL
XFILL_4__15566_ gnd vdd FILL
XFILL_3__10439_ gnd vdd FILL
XFILL_6__11599_ gnd vdd FILL
XFILL_1__14406_ gnd vdd FILL
XFILL_4__12778_ gnd vdd FILL
XFILL_2__13957_ gnd vdd FILL
XFILL_1__11618_ gnd vdd FILL
XFILL_1__15386_ gnd vdd FILL
XFILL_6__9121_ gnd vdd FILL
XFILL_0__10259_ gnd vdd FILL
XFILL_0__9634_ gnd vdd FILL
XFILL_1__12598_ gnd vdd FILL
XFILL_0__6846_ gnd vdd FILL
XFILL_4__14517_ gnd vdd FILL
X_8173_ _8173_/Q _7021_/CLK _9062_/R vdd _8173_/D gnd vdd DFFSR
XFILL_3__9343_ gnd vdd FILL
XSFILL3560x53050 gnd vdd FILL
XFILL_2__12908_ gnd vdd FILL
XFILL_3__13158_ gnd vdd FILL
XFILL_4__11729_ gnd vdd FILL
XFILL_1__14337_ gnd vdd FILL
XFILL_4__15497_ gnd vdd FILL
XFILL_1__11549_ gnd vdd FILL
XFILL_2__13888_ gnd vdd FILL
XFILL_5__15807_ gnd vdd FILL
XFILL_3__12109_ gnd vdd FILL
X_7124_ _7124_/A _7508_/B gnd _7124_/Y vdd NAND2X1
XFILL_4__14448_ gnd vdd FILL
XFILL_3__13089_ gnd vdd FILL
XFILL_2__15627_ gnd vdd FILL
XFILL_5__13999_ gnd vdd FILL
XFILL_3__9274_ gnd vdd FILL
XFILL_2__12839_ gnd vdd FILL
XSFILL44040x13050 gnd vdd FILL
XFILL_1__14268_ gnd vdd FILL
XFILL_0__8516_ gnd vdd FILL
X_7055_ _7055_/A _9615_/B gnd _7056_/C vdd NAND2X1
XFILL_0__14998_ gnd vdd FILL
XFILL_5__15738_ gnd vdd FILL
XFILL_1__16007_ gnd vdd FILL
XFILL_0__9496_ gnd vdd FILL
XFILL_3__8225_ gnd vdd FILL
XFILL_1__13219_ gnd vdd FILL
XFILL_2__15558_ gnd vdd FILL
XFILL_4__14379_ gnd vdd FILL
XFILL_1__14199_ gnd vdd FILL
XFILL_0__13949_ gnd vdd FILL
XFILL_0__8447_ gnd vdd FILL
XFILL_4__16118_ gnd vdd FILL
XFILL_1__7240_ gnd vdd FILL
XFILL_5__15669_ gnd vdd FILL
XSFILL33880x56050 gnd vdd FILL
XFILL_2__14509_ gnd vdd FILL
XFILL_2__15489_ gnd vdd FILL
XFILL_0__8378_ gnd vdd FILL
XFILL_1__7171_ gnd vdd FILL
XFILL_3__7107_ gnd vdd FILL
XFILL_4__16049_ gnd vdd FILL
XSFILL48920x78050 gnd vdd FILL
XFILL_0__15619_ gnd vdd FILL
XFILL_3__8087_ gnd vdd FILL
XSFILL64200x26050 gnd vdd FILL
XFILL_0__7329_ gnd vdd FILL
XSFILL74360x70050 gnd vdd FILL
X_7957_ _7955_/B _7445_/B gnd _7957_/Y vdd NAND2X1
XFILL_3__7038_ gnd vdd FILL
XSFILL48520x80050 gnd vdd FILL
X_6908_ _6908_/A gnd _6910_/A vdd INVX1
X_7888_ _7888_/A gnd _7890_/A vdd INVX1
XSFILL3640x33050 gnd vdd FILL
XFILL_4__7851_ gnd vdd FILL
X_9627_ _9628_/B _8091_/B gnd _9627_/Y vdd NAND2X1
X_6839_ _6839_/A gnd memoryAddress[1] vdd BUFX2
XFILL_1_CLKBUF1_insert1078 gnd vdd FILL
XFILL_3__8989_ gnd vdd FILL
XFILL_1__9812_ gnd vdd FILL
XFILL_5_BUFX2_insert310 gnd vdd FILL
X_9558_ _9558_/Q _8022_/CLK _8674_/R vdd _9558_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert321 gnd vdd FILL
XBUFX2_insert11 _13280_/Y gnd _7297_/B vdd BUFX2
XFILL_4__9521_ gnd vdd FILL
XFILL_5_BUFX2_insert332 gnd vdd FILL
XSFILL94520x83050 gnd vdd FILL
XFILL_5_BUFX2_insert343 gnd vdd FILL
XBUFX2_insert22 _11344_/Y gnd _11743_/A vdd BUFX2
X_10440_ _10426_/B _8136_/B gnd _10441_/C vdd NAND2X1
XBUFX2_insert33 _13320_/Y gnd _8494_/B vdd BUFX2
XFILL_5_BUFX2_insert354 gnd vdd FILL
X_8509_ _8507_/Y _8508_/A _8509_/C gnd _8557_/D vdd OAI21X1
XFILL_1__9743_ gnd vdd FILL
XFILL_5_BUFX2_insert365 gnd vdd FILL
XBUFX2_insert44 _14986_/Y gnd _16199_/C vdd BUFX2
XFILL_1__6955_ gnd vdd FILL
XBUFX2_insert55 _13309_/Y gnd _8118_/A vdd BUFX2
XFILL_5_BUFX2_insert376 gnd vdd FILL
X_9489_ _9567_/Q gnd _9489_/Y vdd INVX1
XFILL_5_BUFX2_insert387 gnd vdd FILL
XBUFX2_insert66 _12215_/Y gnd _12289_/B vdd BUFX2
XBUFX2_insert77 _15015_/Y gnd _15644_/D vdd BUFX2
XSFILL33960x36050 gnd vdd FILL
X_10371_ _10372_/B _7555_/B gnd _10371_/Y vdd NAND2X1
XFILL_5_BUFX2_insert398 gnd vdd FILL
XBUFX2_insert88 _13390_/Y gnd _14567_/A vdd BUFX2
XFILL_1__9674_ gnd vdd FILL
XBUFX2_insert99 _15009_/Y gnd _15544_/A vdd BUFX2
XFILL_1__6886_ gnd vdd FILL
XFILL_4__8403_ gnd vdd FILL
XFILL_4__9383_ gnd vdd FILL
X_12110_ _12110_/A _12110_/B _12110_/C gnd _12110_/Y vdd NAND3X1
X_13090_ _13090_/A _13168_/B _13089_/Y gnd _13090_/Y vdd OAI21X1
XFILL_1__8625_ gnd vdd FILL
XFILL_4__8334_ gnd vdd FILL
X_12041_ _12041_/A _12025_/B _12025_/C gnd gnd _12042_/C vdd AOI22X1
XFILL_4__8265_ gnd vdd FILL
XFILL_1__7507_ gnd vdd FILL
XFILL_1__8487_ gnd vdd FILL
XFILL_4__7216_ gnd vdd FILL
XSFILL3720x13050 gnd vdd FILL
XFILL_4__8196_ gnd vdd FILL
X_15800_ _15793_/Y _15799_/Y gnd _15811_/A vdd NAND2X1
XFILL_1__7438_ gnd vdd FILL
X_13992_ _13991_/Y _13813_/B _13824_/B _13990_/Y gnd _13996_/B vdd OAI22X1
XFILL_2_BUFX2_insert233 gnd vdd FILL
X_12943_ _12895_/A _9050_/CLK _8171_/R vdd _12943_/D gnd vdd DFFSR
X_15731_ _15708_/Y _15731_/B _15731_/C gnd _15732_/B vdd NOR3X1
XFILL_2_BUFX2_insert244 gnd vdd FILL
XFILL_2_BUFX2_insert255 gnd vdd FILL
XFILL_1__7369_ gnd vdd FILL
XFILL_2_BUFX2_insert266 gnd vdd FILL
XSFILL79160x62050 gnd vdd FILL
XFILL_4__7078_ gnd vdd FILL
XFILL_2_BUFX2_insert277 gnd vdd FILL
XSFILL114760x69050 gnd vdd FILL
XFILL_5__7960_ gnd vdd FILL
XFILL_1__9108_ gnd vdd FILL
X_15662_ _15662_/A _7653_/Q _7459_/A _15383_/D gnd _15662_/Y vdd AOI22X1
XFILL_4__10060_ gnd vdd FILL
XFILL_1_BUFX2_insert900 gnd vdd FILL
XFILL_2_BUFX2_insert288 gnd vdd FILL
X_12874_ _12936_/Q gnd _12874_/Y vdd INVX1
XFILL_2_BUFX2_insert299 gnd vdd FILL
XFILL_3__10790_ gnd vdd FILL
XSFILL104200x27050 gnd vdd FILL
XFILL_1_BUFX2_insert911 gnd vdd FILL
XFILL_5__6911_ gnd vdd FILL
XFILL_1_BUFX2_insert922 gnd vdd FILL
X_14613_ _9534_/A gnd _14613_/Y vdd INVX1
X_11825_ _11376_/A _11848_/A _11846_/C _11015_/A gnd _11828_/B vdd AOI22X1
XFILL_1_BUFX2_insert933 gnd vdd FILL
XFILL_1__9039_ gnd vdd FILL
XFILL_5__7891_ gnd vdd FILL
X_15593_ _15593_/A _15593_/B gnd _15598_/A vdd NOR2X1
XFILL_1_BUFX2_insert944 gnd vdd FILL
XFILL_5__11350_ gnd vdd FILL
XFILL_1_BUFX2_insert955 gnd vdd FILL
XSFILL114360x71050 gnd vdd FILL
XFILL_2__9921_ gnd vdd FILL
XFILL_1__10920_ gnd vdd FILL
XFILL_2__11170_ gnd vdd FILL
XFILL_1_BUFX2_insert966 gnd vdd FILL
XSFILL18840x77050 gnd vdd FILL
XFILL_5__9630_ gnd vdd FILL
XFILL_5__10301_ gnd vdd FILL
XSFILL84280x53050 gnd vdd FILL
XFILL_1_BUFX2_insert977 gnd vdd FILL
X_14544_ _7992_/A gnd _14544_/Y vdd INVX1
XFILL_5__6842_ gnd vdd FILL
XFILL_1_BUFX2_insert988 gnd vdd FILL
XFILL_5__11281_ gnd vdd FILL
X_11756_ _11801_/B _11027_/B _11041_/A gnd _11776_/B vdd OAI21X1
XFILL_2__10121_ gnd vdd FILL
XFILL_3__12460_ gnd vdd FILL
XFILL_1_BUFX2_insert999 gnd vdd FILL
XFILL_0__11300_ gnd vdd FILL
XFILL_2__9852_ gnd vdd FILL
XFILL_0__12280_ gnd vdd FILL
XFILL_5__13020_ gnd vdd FILL
XFILL_5__10232_ gnd vdd FILL
X_10707_ _10741_/Q gnd _10709_/A vdd INVX1
XBUFX2_insert232 _11228_/Y gnd _11621_/C vdd BUFX2
XSFILL99320x75050 gnd vdd FILL
X_14475_ _7093_/A gnd _14475_/Y vdd INVX1
XBUFX2_insert243 _13460_/Y gnd _14897_/D vdd BUFX2
XFILL_3__11411_ gnd vdd FILL
XBUFX2_insert254 _10922_/Y gnd _13274_/A vdd BUFX2
XFILL_4__13750_ gnd vdd FILL
X_11687_ _11687_/A _11743_/A _11687_/C gnd _11688_/B vdd NAND3X1
XFILL_4__10962_ gnd vdd FILL
XFILL_3__12391_ gnd vdd FILL
XBUFX2_insert265 _15024_/Y gnd _15369_/D vdd BUFX2
XFILL_2__10052_ gnd vdd FILL
XSFILL59000x9050 gnd vdd FILL
XFILL_0__11231_ gnd vdd FILL
XFILL_2__9783_ gnd vdd FILL
XFILL_5__8512_ gnd vdd FILL
XFILL_4__9719_ gnd vdd FILL
XFILL_2__6995_ gnd vdd FILL
XFILL_1__13570_ gnd vdd FILL
X_16214_ _15177_/B _7245_/A gnd _16218_/C vdd AND2X2
X_13426_ _13420_/Y _13426_/B gnd _13426_/Y vdd NOR2X1
XFILL_1__10782_ gnd vdd FILL
XBUFX2_insert276 _13364_/Y gnd _10619_/B vdd BUFX2
X_10638_ _10638_/A gnd _10638_/Y vdd INVX1
XFILL_4__12701_ gnd vdd FILL
XFILL_3__14130_ gnd vdd FILL
XBUFX2_insert287 _15059_/Y gnd _16213_/B vdd BUFX2
XFILL_5__10163_ gnd vdd FILL
XFILL_5__9492_ gnd vdd FILL
XFILL_5_CLKBUF1_insert111 gnd vdd FILL
XFILL_5_CLKBUF1_insert122 gnd vdd FILL
XFILL_3__11342_ gnd vdd FILL
XBUFX2_insert298 _13356_/Y gnd _10285_/A vdd BUFX2
XFILL_2__14860_ gnd vdd FILL
XFILL_5_CLKBUF1_insert133 gnd vdd FILL
XFILL_4__13681_ gnd vdd FILL
XFILL_1__12521_ gnd vdd FILL
XFILL_4__10893_ gnd vdd FILL
XFILL_2__8734_ gnd vdd FILL
XFILL_5_CLKBUF1_insert144 gnd vdd FILL
XFILL112280x35050 gnd vdd FILL
XFILL_0__11162_ gnd vdd FILL
XFILL_5_CLKBUF1_insert155 gnd vdd FILL
XFILL_5__8443_ gnd vdd FILL
X_16145_ _7025_/Q gnd _16145_/Y vdd INVX1
X_13357_ _13289_/B _13242_/B gnd _13365_/B vdd NAND2X1
XFILL_4__15420_ gnd vdd FILL
XFILL_4__12632_ gnd vdd FILL
XFILL_2__13811_ gnd vdd FILL
XFILL_5_CLKBUF1_insert166 gnd vdd FILL
XFILL_3__14061_ gnd vdd FILL
XFILL_5__14971_ gnd vdd FILL
X_10569_ _10569_/A _10581_/B _10569_/C gnd _10609_/D vdd OAI21X1
XFILL_0__10113_ gnd vdd FILL
XFILL_1__15240_ gnd vdd FILL
XFILL_5_CLKBUF1_insert177 gnd vdd FILL
XFILL_3__11273_ gnd vdd FILL
XFILL_5_CLKBUF1_insert188 gnd vdd FILL
XFILL_1__12452_ gnd vdd FILL
XFILL_2__14791_ gnd vdd FILL
XFILL_5__8374_ gnd vdd FILL
XFILL_0__15970_ gnd vdd FILL
XFILL_5_CLKBUF1_insert199 gnd vdd FILL
X_12308_ _12224_/A _12308_/B _12224_/C gnd _12310_/B vdd NAND3X1
XSFILL74200x3050 gnd vdd FILL
XFILL_0__11093_ gnd vdd FILL
XFILL_5__13922_ gnd vdd FILL
X_16076_ _16076_/A _15680_/B _15680_/C gnd _16085_/C vdd NAND3X1
XFILL_3__13012_ gnd vdd FILL
XFILL_0__7680_ gnd vdd FILL
X_13288_ _13266_/A _13288_/B gnd _13342_/B vdd NAND2X1
XFILL_4__15351_ gnd vdd FILL
XFILL_2__7616_ gnd vdd FILL
XFILL_6__11384_ gnd vdd FILL
XFILL_2__13742_ gnd vdd FILL
XSFILL79240x42050 gnd vdd FILL
XFILL_1__11403_ gnd vdd FILL
XSFILL43880x19050 gnd vdd FILL
XFILL_2__10954_ gnd vdd FILL
XFILL_0__10044_ gnd vdd FILL
XFILL_1__15171_ gnd vdd FILL
XFILL_0__14921_ gnd vdd FILL
XFILL_2__8596_ gnd vdd FILL
XFILL_5__7325_ gnd vdd FILL
XFILL_1__12383_ gnd vdd FILL
X_15027_ _15011_/Y _15027_/B _15027_/C gnd _15028_/A vdd NAND3X1
X_12239_ _12239_/A gnd _12239_/C gnd _12239_/Y vdd NAND3X1
XFILL_4__14302_ gnd vdd FILL
XFILL_5__13853_ gnd vdd FILL
XFILL_4__11514_ gnd vdd FILL
XFILL_4__12494_ gnd vdd FILL
XFILL_3__10155_ gnd vdd FILL
XFILL_2__7547_ gnd vdd FILL
XFILL_1__14122_ gnd vdd FILL
XFILL_4__15282_ gnd vdd FILL
XFILL_2__13673_ gnd vdd FILL
XFILL_1__11334_ gnd vdd FILL
XFILL_0__14852_ gnd vdd FILL
XSFILL114440x51050 gnd vdd FILL
XFILL_2__10885_ gnd vdd FILL
XFILL_0__9350_ gnd vdd FILL
XFILL_2__15412_ gnd vdd FILL
XFILL_4__14233_ gnd vdd FILL
XSFILL34520x4050 gnd vdd FILL
XFILL_4__11445_ gnd vdd FILL
XFILL_2__12624_ gnd vdd FILL
XFILL_5__13784_ gnd vdd FILL
XFILL_2__7478_ gnd vdd FILL
XFILL_0__13803_ gnd vdd FILL
XFILL_1__14053_ gnd vdd FILL
XFILL_3__14963_ gnd vdd FILL
XFILL_5__10996_ gnd vdd FILL
XFILL_2__16392_ gnd vdd FILL
XFILL_1__11265_ gnd vdd FILL
XFILL_5__15523_ gnd vdd FILL
XFILL_5__7187_ gnd vdd FILL
XFILL_0__14783_ gnd vdd FILL
XFILL_2__9217_ gnd vdd FILL
XFILL_5__12735_ gnd vdd FILL
XFILL_3__8010_ gnd vdd FILL
XFILL_0__11995_ gnd vdd FILL
XFILL_0__9281_ gnd vdd FILL
XFILL_2__15343_ gnd vdd FILL
XFILL_4__14164_ gnd vdd FILL
XFILL_3__13914_ gnd vdd FILL
XFILL_4__11376_ gnd vdd FILL
XFILL_1__13004_ gnd vdd FILL
XSFILL99400x55050 gnd vdd FILL
XFILL_0__13734_ gnd vdd FILL
XFILL_1__11196_ gnd vdd FILL
XFILL_3__14894_ gnd vdd FILL
XFILL_0__10946_ gnd vdd FILL
XFILL_0__8232_ gnd vdd FILL
X_15929_ _15929_/A _15929_/B _13274_/A gnd _12887_/B vdd AOI21X1
XFILL_4__13115_ gnd vdd FILL
XFILL_5__15454_ gnd vdd FILL
XFILL_2__9148_ gnd vdd FILL
XFILL111720x49050 gnd vdd FILL
X_8860_ _8860_/A _8859_/A _8860_/C gnd _8860_/Y vdd OAI21X1
XFILL_2__11506_ gnd vdd FILL
XFILL_4__14095_ gnd vdd FILL
XFILL_3__13845_ gnd vdd FILL
XFILL_1__10147_ gnd vdd FILL
XFILL_2__15274_ gnd vdd FILL
XFILL_2__12486_ gnd vdd FILL
XFILL_0__13665_ gnd vdd FILL
XFILL_5__14405_ gnd vdd FILL
X_7811_ _7887_/B _9475_/B gnd _7811_/Y vdd NAND2X1
XFILL_0__10877_ gnd vdd FILL
XSFILL63640x34050 gnd vdd FILL
XFILL_5__11617_ gnd vdd FILL
XFILL112360x15050 gnd vdd FILL
XFILL_5__15385_ gnd vdd FILL
XFILL_2__14225_ gnd vdd FILL
XFILL_4__13046_ gnd vdd FILL
XFILL_4__10258_ gnd vdd FILL
XFILL_0__15404_ gnd vdd FILL
XFILL_5__12597_ gnd vdd FILL
XFILL_2__9079_ gnd vdd FILL
XFILL_2__11437_ gnd vdd FILL
X_8791_ _8791_/Q _7515_/CLK _7665_/R vdd _8699_/Y gnd vdd DFFSR
XFILL_0__12616_ gnd vdd FILL
XFILL_3__13776_ gnd vdd FILL
XFILL_3__10988_ gnd vdd FILL
XFILL_1__14955_ gnd vdd FILL
XFILL_0__7114_ gnd vdd FILL
XFILL_0__16384_ gnd vdd FILL
XFILL_0__13596_ gnd vdd FILL
XFILL_5__14336_ gnd vdd FILL
X_7742_ _7790_/Q gnd _7744_/A vdd INVX1
XFILL_3__15515_ gnd vdd FILL
XSFILL109400x40050 gnd vdd FILL
XFILL_5__11548_ gnd vdd FILL
XFILL_0__8094_ gnd vdd FILL
XFILL_4__10189_ gnd vdd FILL
XFILL_3__12727_ gnd vdd FILL
XFILL_2__14156_ gnd vdd FILL
XFILL_1__13906_ gnd vdd FILL
XFILL_3__8912_ gnd vdd FILL
XFILL_0__15335_ gnd vdd FILL
XFILL_2__11368_ gnd vdd FILL
XFILL_3__9892_ gnd vdd FILL
XFILL_1__14886_ gnd vdd FILL
XSFILL49080x61050 gnd vdd FILL
XFILL_0__7045_ gnd vdd FILL
XSFILL79320x22050 gnd vdd FILL
XFILL_2__13107_ gnd vdd FILL
XFILL_5__14267_ gnd vdd FILL
XFILL_2__10319_ gnd vdd FILL
X_7673_ _7673_/A gnd _7675_/A vdd INVX1
XFILL_3__15446_ gnd vdd FILL
XFILL_5__11479_ gnd vdd FILL
XFILL_3__12658_ gnd vdd FILL
XFILL_3__8843_ gnd vdd FILL
XFILL_1__13837_ gnd vdd FILL
XFILL_4__14997_ gnd vdd FILL
XFILL_2__14087_ gnd vdd FILL
XFILL_5__16006_ gnd vdd FILL
XFILL_2__11299_ gnd vdd FILL
XFILL_0__15266_ gnd vdd FILL
XFILL_5__13218_ gnd vdd FILL
X_9412_ _9412_/A gnd _9414_/A vdd INVX1
XFILL_0__12478_ gnd vdd FILL
XFILL_5__9759_ gnd vdd FILL
XFILL_6__15557_ gnd vdd FILL
XFILL_5__14198_ gnd vdd FILL
XFILL_2__13038_ gnd vdd FILL
XSFILL114520x31050 gnd vdd FILL
XFILL_3__11609_ gnd vdd FILL
XFILL_4__13948_ gnd vdd FILL
XFILL_3__12589_ gnd vdd FILL
XFILL_3__15377_ gnd vdd FILL
XFILL_0__14217_ gnd vdd FILL
XFILL_1__13768_ gnd vdd FILL
XFILL_3__8774_ gnd vdd FILL
XFILL_0__11429_ gnd vdd FILL
XFILL_0__15197_ gnd vdd FILL
XFILL_6__14508_ gnd vdd FILL
X_9343_ _9343_/A gnd _9345_/A vdd INVX1
XFILL_5__13149_ gnd vdd FILL
XFILL_0__8996_ gnd vdd FILL
XFILL_1__15507_ gnd vdd FILL
XFILL_3__14328_ gnd vdd FILL
XFILL_1__12719_ gnd vdd FILL
XFILL_4__13879_ gnd vdd FILL
XFILL_3__7725_ gnd vdd FILL
XFILL_0__14148_ gnd vdd FILL
XFILL_1__13699_ gnd vdd FILL
XFILL_0__7947_ gnd vdd FILL
XFILL_4__15618_ gnd vdd FILL
XFILL_4_BUFX2_insert306 gnd vdd FILL
XFILL_4_BUFX2_insert317 gnd vdd FILL
X_9274_ _9272_/Y _9301_/B _9274_/C gnd _9324_/D vdd OAI21X1
XFILL_3__14259_ gnd vdd FILL
XFILL_4_BUFX2_insert328 gnd vdd FILL
XFILL_1__15438_ gnd vdd FILL
XFILL_4_BUFX2_insert339 gnd vdd FILL
XFILL_2__14989_ gnd vdd FILL
XFILL_0__14079_ gnd vdd FILL
X_8225_ _8246_/A _8225_/B gnd _8226_/C vdd NAND2X1
XFILL_4__15549_ gnd vdd FILL
XFILL_0__7878_ gnd vdd FILL
XFILL_3__7587_ gnd vdd FILL
XFILL_1__15369_ gnd vdd FILL
XFILL_6__16109_ gnd vdd FILL
XFILL_6__7296_ gnd vdd FILL
XFILL_0__9617_ gnd vdd FILL
X_8156_ _8156_/Q _7534_/CLK _8156_/R vdd _8156_/D gnd vdd DFFSR
XFILL_1__9390_ gnd vdd FILL
XSFILL8680x81050 gnd vdd FILL
XSFILL23720x30050 gnd vdd FILL
XFILL_0__9548_ gnd vdd FILL
X_7107_ _7105_/Y _7061_/A _7107_/C gnd _7151_/D vdd OAI21X1
XFILL_1__8341_ gnd vdd FILL
X_8087_ _8087_/A gnd _8089_/A vdd INVX1
XFILL_3__9257_ gnd vdd FILL
XSFILL23640x5050 gnd vdd FILL
XFILL_0__9479_ gnd vdd FILL
X_7038_ _7038_/A _7067_/A _7037_/Y gnd _7038_/Y vdd OAI21X1
XFILL_1__8272_ gnd vdd FILL
XFILL_3__8208_ gnd vdd FILL
XFILL_1__7223_ gnd vdd FILL
XFILL_3__8139_ gnd vdd FILL
XSFILL13640x82050 gnd vdd FILL
XFILL_6__9937_ gnd vdd FILL
X_8989_ _9059_/Q gnd _8991_/A vdd INVX1
XFILL_1_BUFX2_insert229 gnd vdd FILL
XFILL_4__8952_ gnd vdd FILL
XFILL_1__7085_ gnd vdd FILL
X_11610_ _11609_/Y _11595_/C gnd _11610_/Y vdd NAND2X1
XFILL_4__8883_ gnd vdd FILL
X_12590_ _12590_/A vdd _12590_/C gnd _12670_/D vdd OAI21X1
XFILL_0_BUFX2_insert907 gnd vdd FILL
XSFILL104520x63050 gnd vdd FILL
XFILL_0_BUFX2_insert918 gnd vdd FILL
XFILL_4__7834_ gnd vdd FILL
X_11541_ _11541_/A _11531_/Y _11540_/Y gnd _12081_/A vdd NAND3X1
XFILL_0_BUFX2_insert929 gnd vdd FILL
XSFILL8760x61050 gnd vdd FILL
XSFILL23800x10050 gnd vdd FILL
X_14260_ _14256_/Y _14260_/B gnd _14260_/Y vdd NOR2X1
XFILL_4__7765_ gnd vdd FILL
X_11472_ _11471_/Y _11472_/B _11480_/A gnd _11473_/C vdd OAI21X1
XFILL_4__9504_ gnd vdd FILL
XFILL_1__7987_ gnd vdd FILL
X_13211_ _13239_/B gnd _13302_/C vdd INVX2
X_10423_ _10423_/A _10423_/B _10422_/Y gnd _10475_/D vdd OAI21X1
XFILL_4__7696_ gnd vdd FILL
X_14191_ _8165_/Q gnd _14191_/Y vdd INVX1
XFILL_1__6938_ gnd vdd FILL
XFILL_1__9726_ gnd vdd FILL
X_13142_ _13196_/Q gnd _13142_/Y vdd INVX1
X_10354_ _10354_/Q _7129_/CLK _8542_/R vdd _10316_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert840 gnd vdd FILL
XFILL_2__8450_ gnd vdd FILL
XSFILL13720x62050 gnd vdd FILL
XFILL_1__6869_ gnd vdd FILL
XFILL_4_BUFX2_insert851 gnd vdd FILL
XFILL_1__9657_ gnd vdd FILL
XFILL_4_BUFX2_insert862 gnd vdd FILL
XSFILL79160x57050 gnd vdd FILL
XFILL_4_BUFX2_insert873 gnd vdd FILL
XFILL_4__9366_ gnd vdd FILL
XFILL_4_BUFX2_insert884 gnd vdd FILL
X_13073_ _6896_/A _13184_/CLK _8176_/R vdd _13073_/D gnd vdd DFFSR
XFILL_1__8608_ gnd vdd FILL
X_10285_ _10285_/A _9517_/B gnd _10286_/C vdd NAND2X1
XFILL_2__8381_ gnd vdd FILL
XFILL_4_BUFX2_insert895 gnd vdd FILL
XFILL_5__7110_ gnd vdd FILL
XFILL_4__8317_ gnd vdd FILL
XFILL_5__8090_ gnd vdd FILL
X_12024_ _12028_/A _12716_/A _12024_/C gnd _12024_/Y vdd NAND3X1
XFILL_4__9297_ gnd vdd FILL
XFILL_2__7332_ gnd vdd FILL
XFILL_5__7041_ gnd vdd FILL
XFILL_2__10670_ gnd vdd FILL
XFILL_4__8248_ gnd vdd FILL
XFILL_6__10051_ gnd vdd FILL
XFILL_4__11230_ gnd vdd FILL
XSFILL84280x48050 gnd vdd FILL
XFILL_3__11960_ gnd vdd FILL
XFILL_5__10781_ gnd vdd FILL
XFILL_1__11050_ gnd vdd FILL
XFILL_0__10800_ gnd vdd FILL
XFILL_5__12520_ gnd vdd FILL
XFILL_0__11780_ gnd vdd FILL
XFILL_2__9002_ gnd vdd FILL
XFILL_3__10911_ gnd vdd FILL
XFILL_4__11161_ gnd vdd FILL
XFILL_1__10001_ gnd vdd FILL
XSFILL59080x24050 gnd vdd FILL
XFILL_2__12340_ gnd vdd FILL
X_13975_ _13975_/A _13975_/B _14791_/C gnd _12982_/B vdd AOI21X1
XFILL_2__7194_ gnd vdd FILL
XFILL_3__11891_ gnd vdd FILL
XFILL_4__10112_ gnd vdd FILL
X_15714_ _15714_/A _15713_/Y gnd _15720_/B vdd NOR2X1
X_12926_ _12844_/A _9050_/CLK _8171_/R vdd _12926_/D gnd vdd DFFSR
XFILL_5__8992_ gnd vdd FILL
XFILL_5__12451_ gnd vdd FILL
XFILL_3__13630_ gnd vdd FILL
XFILL_4__11092_ gnd vdd FILL
XFILL_2__12271_ gnd vdd FILL
XFILL_0__10662_ gnd vdd FILL
XFILL_0__13450_ gnd vdd FILL
XFILL_6__13741_ gnd vdd FILL
XFILL_5__7943_ gnd vdd FILL
XFILL_5__11402_ gnd vdd FILL
XFILL_4__10043_ gnd vdd FILL
XFILL_5__15170_ gnd vdd FILL
XFILL_2__14010_ gnd vdd FILL
X_15645_ _15645_/A _15642_/Y gnd _15645_/Y vdd NOR2X1
XFILL_1_BUFX2_insert730 gnd vdd FILL
XFILL_4__14920_ gnd vdd FILL
X_12857_ vdd _12857_/B gnd _12858_/C vdd NAND2X1
XFILL_5__12382_ gnd vdd FILL
XFILL_3__13561_ gnd vdd FILL
XFILL_2__11222_ gnd vdd FILL
XFILL_0__12401_ gnd vdd FILL
XFILL_1_BUFX2_insert741 gnd vdd FILL
XFILL_1__14740_ gnd vdd FILL
XFILL_3__10773_ gnd vdd FILL
XFILL_1_BUFX2_insert752 gnd vdd FILL
XFILL_1__11952_ gnd vdd FILL
XFILL_0__13381_ gnd vdd FILL
XFILL_1_BUFX2_insert763 gnd vdd FILL
XFILL_5__14121_ gnd vdd FILL
XFILL_1_BUFX2_insert774 gnd vdd FILL
XFILL_3__15300_ gnd vdd FILL
XFILL_5__7874_ gnd vdd FILL
X_11808_ _11808_/A _11808_/B _11808_/C gnd _12005_/A vdd NAND3X1
XFILL_5__11333_ gnd vdd FILL
X_12788_ _12788_/A gnd _12788_/Y vdd INVX1
XFILL_4__14851_ gnd vdd FILL
XFILL_3__12512_ gnd vdd FILL
XFILL_2__9904_ gnd vdd FILL
XFILL_6__10884_ gnd vdd FILL
X_15576_ _16261_/A _14115_/D _14115_/A _16261_/D gnd _15579_/B vdd OAI22X1
XFILL_1__10903_ gnd vdd FILL
XFILL_1_BUFX2_insert785 gnd vdd FILL
XSFILL79240x37050 gnd vdd FILL
XFILL_2__11153_ gnd vdd FILL
XFILL_3__13492_ gnd vdd FILL
XFILL_3__16280_ gnd vdd FILL
XFILL_0__15120_ gnd vdd FILL
XFILL_5__9613_ gnd vdd FILL
XFILL_0__12332_ gnd vdd FILL
XFILL_1__14671_ gnd vdd FILL
XFILL_1_BUFX2_insert796 gnd vdd FILL
XFILL_1__11883_ gnd vdd FILL
XFILL_4__13802_ gnd vdd FILL
XFILL_5__14052_ gnd vdd FILL
X_14527_ _14512_/Y _14527_/B gnd _14527_/Y vdd NOR2X1
XFILL_6__16391_ gnd vdd FILL
X_11739_ _11739_/A _11739_/B gnd _11739_/Y vdd NOR2X1
XFILL_1__16410_ gnd vdd FILL
XFILL_3__15231_ gnd vdd FILL
XFILL_2__10104_ gnd vdd FILL
XFILL_4_BUFX2_insert12 gnd vdd FILL
XFILL_3__12443_ gnd vdd FILL
XFILL_5__11264_ gnd vdd FILL
XFILL_1__13622_ gnd vdd FILL
XFILL_4__14782_ gnd vdd FILL
XFILL_0__15051_ gnd vdd FILL
XFILL_2__15961_ gnd vdd FILL
XFILL_4__11994_ gnd vdd FILL
XFILL_0__12263_ gnd vdd FILL
XFILL_2__11084_ gnd vdd FILL
XFILL_4_BUFX2_insert23 gnd vdd FILL
XFILL_1__10834_ gnd vdd FILL
XFILL_4_BUFX2_insert34 gnd vdd FILL
XFILL_6__15342_ gnd vdd FILL
XFILL_5__9544_ gnd vdd FILL
XFILL_5__13003_ gnd vdd FILL
XFILL_4_BUFX2_insert45 gnd vdd FILL
XFILL_0__8850_ gnd vdd FILL
X_14458_ _16438_/Q _14344_/B _14458_/C _7275_/Q gnd _14458_/Y vdd AOI22X1
XFILL_4_BUFX2_insert56 gnd vdd FILL
XFILL_3__15162_ gnd vdd FILL
XFILL_4__13733_ gnd vdd FILL
XFILL_4__10945_ gnd vdd FILL
XFILL_1__16341_ gnd vdd FILL
XFILL_0__14002_ gnd vdd FILL
XFILL_3__12374_ gnd vdd FILL
XFILL_2__10035_ gnd vdd FILL
XFILL_5__11195_ gnd vdd FILL
XFILL_2__14912_ gnd vdd FILL
XFILL_2__9766_ gnd vdd FILL
XSFILL84360x28050 gnd vdd FILL
XFILL_4_BUFX2_insert67 gnd vdd FILL
XFILL_2__6978_ gnd vdd FILL
XFILL_1__13553_ gnd vdd FILL
XFILL_0__11214_ gnd vdd FILL
XFILL_1__10765_ gnd vdd FILL
XFILL_2__15892_ gnd vdd FILL
XFILL_4_BUFX2_insert78 gnd vdd FILL
XFILL_0__12194_ gnd vdd FILL
XFILL_0__7801_ gnd vdd FILL
XFILL_5__9475_ gnd vdd FILL
XFILL_4_BUFX2_insert89 gnd vdd FILL
X_13409_ _13403_/Y _13879_/B _13876_/C _13402_/Y gnd _13415_/B vdd OAI22X1
XFILL_0__8781_ gnd vdd FILL
XFILL_5__10146_ gnd vdd FILL
X_14389_ _15822_/B _14389_/B _14712_/B _9833_/Q gnd _14390_/B vdd AOI22X1
XFILL_3__14113_ gnd vdd FILL
XFILL_3__11325_ gnd vdd FILL
XFILL_2__8717_ gnd vdd FILL
XFILL_1__12504_ gnd vdd FILL
XFILL_4__13664_ gnd vdd FILL
XFILL_3__15093_ gnd vdd FILL
XFILL_2__14843_ gnd vdd FILL
XFILL_4__10876_ gnd vdd FILL
XFILL_3__8490_ gnd vdd FILL
XFILL_0__11145_ gnd vdd FILL
XFILL_1__16272_ gnd vdd FILL
XFILL_1__13484_ gnd vdd FILL
XFILL_4__15403_ gnd vdd FILL
XFILL_0__7732_ gnd vdd FILL
X_16128_ _16128_/A _16127_/Y gnd _16128_/Y vdd NOR2X1
XSFILL84360x4050 gnd vdd FILL
XFILL_6__11436_ gnd vdd FILL
XFILL_1__10696_ gnd vdd FILL
XFILL_4__12615_ gnd vdd FILL
XFILL_3__14044_ gnd vdd FILL
XFILL_5__14954_ gnd vdd FILL
XFILL_4__16383_ gnd vdd FILL
XFILL_1__15223_ gnd vdd FILL
XFILL_3__7441_ gnd vdd FILL
XFILL_3__11256_ gnd vdd FILL
XFILL_4__13595_ gnd vdd FILL
XFILL_1__12435_ gnd vdd FILL
XFILL_2__8648_ gnd vdd FILL
XFILL_2__14774_ gnd vdd FILL
XFILL_2__11986_ gnd vdd FILL
XFILL_0__15953_ gnd vdd FILL
XFILL_0__11076_ gnd vdd FILL
XFILL_5__8357_ gnd vdd FILL
X_8010_ _8050_/Q gnd _8012_/A vdd INVX1
XFILL_6__14155_ gnd vdd FILL
XFILL_5__13905_ gnd vdd FILL
XFILL_4__15334_ gnd vdd FILL
XFILL_2_BUFX2_insert1006 gnd vdd FILL
X_16059_ _16047_/Y _16058_/Y _16059_/C gnd _16059_/Y vdd NAND3X1
XFILL_2_BUFX2_insert1017 gnd vdd FILL
XFILL_5__14885_ gnd vdd FILL
XFILL_2__10937_ gnd vdd FILL
XFILL_3__7372_ gnd vdd FILL
XFILL_2__8579_ gnd vdd FILL
XFILL_2_BUFX2_insert1028 gnd vdd FILL
XFILL_1__15154_ gnd vdd FILL
XFILL_3__11187_ gnd vdd FILL
XFILL_2__13725_ gnd vdd FILL
XFILL_0__14904_ gnd vdd FILL
XFILL_0__10027_ gnd vdd FILL
XFILL_1__12366_ gnd vdd FILL
XFILL_5__7308_ gnd vdd FILL
XFILL_2_BUFX2_insert1039 gnd vdd FILL
XFILL_0__9402_ gnd vdd FILL
XFILL_0__15884_ gnd vdd FILL
XFILL_5__13836_ gnd vdd FILL
XFILL_3__9111_ gnd vdd FILL
XFILL_3__10138_ gnd vdd FILL
XFILL_0__7594_ gnd vdd FILL
XFILL_6__11298_ gnd vdd FILL
XFILL_4__15265_ gnd vdd FILL
XFILL_1__14105_ gnd vdd FILL
XFILL_2__13656_ gnd vdd FILL
XFILL_4__12477_ gnd vdd FILL
XFILL_1__11317_ gnd vdd FILL
XFILL_0__14835_ gnd vdd FILL
XFILL_3__15995_ gnd vdd FILL
XFILL_1__15085_ gnd vdd FILL
XFILL_6__13037_ gnd vdd FILL
XFILL_5__7239_ gnd vdd FILL
XFILL_1__12297_ gnd vdd FILL
XFILL_4__14216_ gnd vdd FILL
XFILL_5__13767_ gnd vdd FILL
XFILL_2__12607_ gnd vdd FILL
XSFILL49080x56050 gnd vdd FILL
X_9961_ _9961_/Q _9953_/CLK _7276_/R vdd _9961_/D gnd vdd DFFSR
XFILL_3__9042_ gnd vdd FILL
XFILL_4__11428_ gnd vdd FILL
XFILL_5__10979_ gnd vdd FILL
XFILL_4__15196_ gnd vdd FILL
XFILL_1__14036_ gnd vdd FILL
XFILL_3__10069_ gnd vdd FILL
XFILL_3__14946_ gnd vdd FILL
XFILL_2__13587_ gnd vdd FILL
XFILL_2__16375_ gnd vdd FILL
XFILL_1__11248_ gnd vdd FILL
XFILL_5__15506_ gnd vdd FILL
XFILL_2__10799_ gnd vdd FILL
XFILL_0__14766_ gnd vdd FILL
XFILL_5__12718_ gnd vdd FILL
XFILL_0__9264_ gnd vdd FILL
XFILL_0__11978_ gnd vdd FILL
X_8912_ _8912_/A gnd _8912_/Y vdd INVX1
XFILL_4__14147_ gnd vdd FILL
X_9892_ _9920_/B _9380_/B gnd _9893_/C vdd NAND2X1
XFILL_2__15326_ gnd vdd FILL
XFILL_5__13698_ gnd vdd FILL
XFILL_4__11359_ gnd vdd FILL
XFILL_3__14877_ gnd vdd FILL
XSFILL114520x26050 gnd vdd FILL
XFILL_0__13717_ gnd vdd FILL
XFILL_0__10929_ gnd vdd FILL
XFILL_0_BUFX2_insert1010 gnd vdd FILL
XFILL_0__8215_ gnd vdd FILL
XFILL_1__11179_ gnd vdd FILL
XFILL_0__14697_ gnd vdd FILL
XFILL_5__15437_ gnd vdd FILL
XFILL_0_BUFX2_insert1021 gnd vdd FILL
XFILL_5__12649_ gnd vdd FILL
X_8843_ _8925_/Q gnd _8845_/A vdd INVX1
XFILL_0_BUFX2_insert1032 gnd vdd FILL
XFILL_6__7983_ gnd vdd FILL
XFILL_3__13828_ gnd vdd FILL
XFILL_0_BUFX2_insert1043 gnd vdd FILL
XFILL_2__15257_ gnd vdd FILL
XFILL_4__14078_ gnd vdd FILL
XFILL_2__12469_ gnd vdd FILL
XFILL_0_BUFX2_insert1054 gnd vdd FILL
XFILL_0__13648_ gnd vdd FILL
XFILL_1__15987_ gnd vdd FILL
XFILL_6__6934_ gnd vdd FILL
XFILL_0_BUFX2_insert1065 gnd vdd FILL
XFILL_0__8146_ gnd vdd FILL
XFILL_5__15368_ gnd vdd FILL
XFILL_2__14208_ gnd vdd FILL
XFILL_4__13029_ gnd vdd FILL
XFILL_0_BUFX2_insert1087 gnd vdd FILL
X_8774_ _8772_/Y _8759_/B _8774_/C gnd _8816_/D vdd OAI21X1
XSFILL44120x7050 gnd vdd FILL
XFILL_2__15188_ gnd vdd FILL
XFILL_3__13759_ gnd vdd FILL
XSFILL84040x10050 gnd vdd FILL
XFILL_0__16367_ gnd vdd FILL
XFILL_6_BUFX2_insert935 gnd vdd FILL
XFILL_1__14938_ gnd vdd FILL
XFILL_6__9653_ gnd vdd FILL
XFILL_5__14319_ gnd vdd FILL
XFILL_0__13579_ gnd vdd FILL
XFILL_0__8077_ gnd vdd FILL
X_7725_ _7672_/B _6957_/B gnd _7726_/C vdd NAND2X1
XFILL_5__15299_ gnd vdd FILL
XFILL_2__14139_ gnd vdd FILL
XFILL_0__15318_ gnd vdd FILL
XFILL_1__14869_ gnd vdd FILL
XFILL_6__8604_ gnd vdd FILL
XFILL_3__9875_ gnd vdd FILL
XSFILL104440x78050 gnd vdd FILL
XFILL_0__16298_ gnd vdd FILL
XFILL_1__8890_ gnd vdd FILL
X_7656_ _7656_/Q _7016_/CLK _8424_/R vdd _7598_/Y gnd vdd DFFSR
XFILL_3__15429_ gnd vdd FILL
XSFILL8680x76050 gnd vdd FILL
XFILL_3__8826_ gnd vdd FILL
XSFILL23720x25050 gnd vdd FILL
XFILL_0__15249_ gnd vdd FILL
XFILL_1__7841_ gnd vdd FILL
XSFILL33080x50050 gnd vdd FILL
XSFILL88920x75050 gnd vdd FILL
X_7587_ _7653_/Q gnd _7589_/A vdd INVX1
XFILL_4__7550_ gnd vdd FILL
XFILL_3__8757_ gnd vdd FILL
X_9326_ _9326_/Q _8942_/CLK _9561_/R vdd _9326_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert103 gnd vdd FILL
XSFILL3720x50 gnd vdd FILL
XFILL_3__7708_ gnd vdd FILL
XFILL_0__8979_ gnd vdd FILL
XSFILL39400x13050 gnd vdd FILL
XFILL_4__7481_ gnd vdd FILL
XFILL_1__9511_ gnd vdd FILL
XFILL_6__8397_ gnd vdd FILL
X_9257_ _9257_/A gnd _9259_/A vdd INVX1
XFILL_4__9220_ gnd vdd FILL
X_8208_ _8208_/A _8208_/B _8208_/C gnd _8286_/D vdd OAI21X1
XSFILL13640x77050 gnd vdd FILL
XFILL_6__7348_ gnd vdd FILL
XFILL_4__9151_ gnd vdd FILL
X_9188_ _9188_/Q _9188_/CLK _8801_/R vdd _9188_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert803 gnd vdd FILL
XFILL_3_BUFX2_insert814 gnd vdd FILL
XFILL_3_BUFX2_insert825 gnd vdd FILL
X_10070_ _9974_/A _8165_/CLK _8165_/R vdd _9976_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert836 gnd vdd FILL
XSFILL69320x49050 gnd vdd FILL
X_8139_ _8098_/B _8011_/B gnd _8139_/Y vdd NAND2X1
XFILL_1__9373_ gnd vdd FILL
XFILL_4__8102_ gnd vdd FILL
XFILL_3_BUFX2_insert847 gnd vdd FILL
XFILL_4__9082_ gnd vdd FILL
XFILL_3_BUFX2_insert858 gnd vdd FILL
XFILL_3_BUFX2_insert869 gnd vdd FILL
XFILL_1__8324_ gnd vdd FILL
XSFILL104520x58050 gnd vdd FILL
XFILL_1__8255_ gnd vdd FILL
XSFILL8760x56050 gnd vdd FILL
XSFILL73400x76050 gnd vdd FILL
X_13760_ _13751_/Y _13760_/B _13759_/Y gnd _13761_/B vdd NAND3X1
XFILL_1__7206_ gnd vdd FILL
X_10972_ _10984_/Q gnd _10972_/Y vdd INVX1
XFILL_1__8186_ gnd vdd FILL
XSFILL74040x42050 gnd vdd FILL
XFILL_4__9984_ gnd vdd FILL
X_12711_ _12718_/B memoryOutData[5] gnd _12711_/Y vdd NAND2X1
X_13691_ _9733_/A gnd _13691_/Y vdd INVX1
XSFILL79160x5050 gnd vdd FILL
X_12642_ _12642_/A gnd _12644_/A vdd INVX1
X_15430_ _8799_/Q gnd _15431_/D vdd INVX1
XSFILL108760x63050 gnd vdd FILL
XFILL_1__7068_ gnd vdd FILL
XFILL_2__7950_ gnd vdd FILL
XSFILL13720x57050 gnd vdd FILL
XFILL_0_BUFX2_insert704 gnd vdd FILL
XFILL_0_CLKBUF1_insert130 gnd vdd FILL
X_15361_ _15361_/A _15357_/Y _15361_/C gnd _15372_/A vdd NAND3X1
XFILL_0_CLKBUF1_insert141 gnd vdd FILL
XFILL_4__8866_ gnd vdd FILL
XFILL_0_BUFX2_insert715 gnd vdd FILL
XFILL_0_BUFX2_insert726 gnd vdd FILL
X_12573_ _12573_/A gnd _12575_/A vdd INVX1
XFILL_2__6901_ gnd vdd FILL
XFILL_0_CLKBUF1_insert152 gnd vdd FILL
XFILL_0_BUFX2_insert737 gnd vdd FILL
XFILL_0_CLKBUF1_insert163 gnd vdd FILL
XFILL_2__7881_ gnd vdd FILL
XFILL_4__7817_ gnd vdd FILL
XFILL_0_BUFX2_insert748 gnd vdd FILL
XFILL_0_CLKBUF1_insert174 gnd vdd FILL
XFILL_5__7590_ gnd vdd FILL
XFILL_0_CLKBUF1_insert185 gnd vdd FILL
XFILL_0_BUFX2_insert759 gnd vdd FILL
X_11524_ _11142_/A _11057_/Y _11569_/B gnd _11562_/A vdd AOI21X1
X_14312_ _14312_/A _14288_/Y _15812_/C gnd _13003_/B vdd AOI21X1
XFILL_0_CLKBUF1_insert196 gnd vdd FILL
X_15292_ _16314_/D _13733_/D _16309_/A _13696_/D gnd _15292_/Y vdd OAI22X1
XFILL_2__9620_ gnd vdd FILL
XSFILL28920x7050 gnd vdd FILL
X_14243_ _14243_/A _14243_/B gnd _14265_/A vdd NOR2X1
XFILL_5__10000_ gnd vdd FILL
XFILL_4__7748_ gnd vdd FILL
X_11455_ _11334_/A _11440_/A _11454_/Y gnd _11455_/Y vdd NAND3X1
XFILL_2__9551_ gnd vdd FILL
XFILL_1__10550_ gnd vdd FILL
X_10406_ _10406_/A gnd _10408_/A vdd INVX1
XFILL_5__9260_ gnd vdd FILL
XFILL_4__7679_ gnd vdd FILL
X_14174_ _14583_/B _15674_/A _14174_/C _14174_/D gnd _14179_/B vdd OAI22X1
XSFILL17960x62050 gnd vdd FILL
XFILL_6__12270_ gnd vdd FILL
XFILL_3__11110_ gnd vdd FILL
XFILL_2__8502_ gnd vdd FILL
X_11386_ _12250_/Y _12141_/Y gnd _11386_/Y vdd XNOR2X1
XFILL_4__10661_ gnd vdd FILL
XFILL_2__9482_ gnd vdd FILL
XFILL_3__12090_ gnd vdd FILL
XSFILL59880x38050 gnd vdd FILL
XSFILL59080x19050 gnd vdd FILL
XFILL_2__11840_ gnd vdd FILL
XFILL_4__9418_ gnd vdd FILL
XFILL_5__8211_ gnd vdd FILL
X_13125_ _13168_/B _12050_/Y gnd _13125_/Y vdd NAND2X1
XFILL_6__11221_ gnd vdd FILL
XSFILL99480x24050 gnd vdd FILL
XFILL_4__12400_ gnd vdd FILL
X_10337_ _15509_/D _9953_/CLK _7649_/R vdd _10265_/Y gnd vdd DFFSR
XFILL_5__11951_ gnd vdd FILL
XFILL_4_BUFX2_insert670 gnd vdd FILL
XFILL_3__11041_ gnd vdd FILL
XSFILL74120x22050 gnd vdd FILL
XFILL_4__13380_ gnd vdd FILL
XFILL_1__12220_ gnd vdd FILL
XFILL_4_BUFX2_insert681 gnd vdd FILL
XFILL_4_BUFX2_insert692 gnd vdd FILL
XFILL_2__11771_ gnd vdd FILL
XFILL_5__8142_ gnd vdd FILL
XFILL_4__9349_ gnd vdd FILL
XFILL_5__10902_ gnd vdd FILL
X_13056_ _6879_/A _9823_/CLK _9056_/R vdd _13056_/D gnd vdd DFFSR
XFILL_4__12331_ gnd vdd FILL
X_10268_ _10268_/A _10285_/A _10267_/Y gnd _10338_/D vdd OAI21X1
XFILL_5__14670_ gnd vdd FILL
XFILL_2__13510_ gnd vdd FILL
XFILL_5__11882_ gnd vdd FILL
XFILL_2__8364_ gnd vdd FILL
XFILL_2__14490_ gnd vdd FILL
XFILL_0__11901_ gnd vdd FILL
XFILL_1__12151_ gnd vdd FILL
XFILL_5__8073_ gnd vdd FILL
X_12007_ _12007_/A _12454_/A _12111_/C gnd _12010_/A vdd NAND3X1
XFILL_5__13621_ gnd vdd FILL
XFILL_0__12881_ gnd vdd FILL
XFILL_3__14800_ gnd vdd FILL
XFILL_4__15050_ gnd vdd FILL
XSFILL13800x37050 gnd vdd FILL
XFILL_6__11083_ gnd vdd FILL
XFILL_2__7315_ gnd vdd FILL
XFILL_5__10833_ gnd vdd FILL
XFILL_2__13441_ gnd vdd FILL
XFILL_4__12262_ gnd vdd FILL
XFILL_1__11102_ gnd vdd FILL
X_10199_ _13523_/A _8152_/CLK _9944_/R vdd _10107_/Y gnd vdd DFFSR
XFILL_0__14620_ gnd vdd FILL
XFILL_3__15780_ gnd vdd FILL
XFILL_2__10653_ gnd vdd FILL
XFILL_1__12082_ gnd vdd FILL
XFILL_3__12992_ gnd vdd FILL
XFILL_0__11832_ gnd vdd FILL
XFILL_5__16340_ gnd vdd FILL
XFILL_4__14001_ gnd vdd FILL
XFILL_5__13552_ gnd vdd FILL
XFILL_4__11213_ gnd vdd FILL
XFILL_2__7246_ gnd vdd FILL
XFILL_5__10764_ gnd vdd FILL
XFILL_3__14731_ gnd vdd FILL
XFILL_4__12193_ gnd vdd FILL
XFILL_2__16160_ gnd vdd FILL
XSFILL64040x74050 gnd vdd FILL
XFILL_1__15910_ gnd vdd FILL
XFILL_2__13372_ gnd vdd FILL
XFILL_3__11943_ gnd vdd FILL
XFILL_1__11033_ gnd vdd FILL
XFILL_0__14551_ gnd vdd FILL
XFILL_5__12503_ gnd vdd FILL
XFILL_0__11763_ gnd vdd FILL
XFILL_4__11144_ gnd vdd FILL
XFILL_2__15111_ gnd vdd FILL
XFILL_5__16271_ gnd vdd FILL
XFILL_2__12323_ gnd vdd FILL
X_13958_ _8160_/Q gnd _13959_/D vdd INVX1
XFILL_5__13483_ gnd vdd FILL
XFILL_2__7177_ gnd vdd FILL
XFILL_2__16091_ gnd vdd FILL
XFILL_3__14662_ gnd vdd FILL
XFILL_0__13502_ gnd vdd FILL
XFILL_5__10695_ gnd vdd FILL
XFILL_3__11874_ gnd vdd FILL
XFILL_0__8000_ gnd vdd FILL
XFILL_1__15841_ gnd vdd FILL
XFILL_0__14482_ gnd vdd FILL
XFILL_5__15222_ gnd vdd FILL
XFILL_5__12434_ gnd vdd FILL
XFILL_5__8975_ gnd vdd FILL
XFILL_3__16401_ gnd vdd FILL
X_12909_ _12907_/Y vdd _12909_/C gnd _12947_/D vdd OAI21X1
XFILL_0__11694_ gnd vdd FILL
XFILL_3__13613_ gnd vdd FILL
XFILL_2__15042_ gnd vdd FILL
XFILL_4__15952_ gnd vdd FILL
XFILL_4__11075_ gnd vdd FILL
XFILL_0__16221_ gnd vdd FILL
XFILL_2__12254_ gnd vdd FILL
X_13889_ _9055_/Q gnd _15416_/A vdd INVX1
XFILL_3__10825_ gnd vdd FILL
XFILL_3__14593_ gnd vdd FILL
XFILL_0__13433_ gnd vdd FILL
XFILL_1__15772_ gnd vdd FILL
XFILL_3__7990_ gnd vdd FILL
XSFILL68680x77050 gnd vdd FILL
XFILL_5__7926_ gnd vdd FILL
XFILL_1__12984_ gnd vdd FILL
XFILL_0__10645_ gnd vdd FILL
X_15628_ _15619_/Y _15628_/B _15628_/C gnd _15629_/B vdd NAND3X1
XFILL_5__15153_ gnd vdd FILL
XFILL_4__14903_ gnd vdd FILL
XFILL_4__10026_ gnd vdd FILL
XFILL_5__12365_ gnd vdd FILL
XFILL_3__16332_ gnd vdd FILL
XFILL_2__11205_ gnd vdd FILL
XFILL_1_BUFX2_insert560 gnd vdd FILL
XFILL_3__10756_ gnd vdd FILL
XFILL_1__14723_ gnd vdd FILL
XFILL_1_BUFX2_insert571 gnd vdd FILL
XFILL_3__13544_ gnd vdd FILL
XFILL_4__15883_ gnd vdd FILL
XFILL_1_BUFX2_insert582 gnd vdd FILL
XFILL_2__12185_ gnd vdd FILL
XFILL_1__11935_ gnd vdd FILL
XFILL_3__6941_ gnd vdd FILL
XFILL_0__16152_ gnd vdd FILL
XFILL_0__13364_ gnd vdd FILL
XFILL_1_BUFX2_insert593 gnd vdd FILL
XFILL_5__14104_ gnd vdd FILL
X_7510_ _7510_/Q _8022_/CLK _9046_/R vdd _7416_/Y gnd vdd DFFSR
XFILL_5__7857_ gnd vdd FILL
XFILL_5__11316_ gnd vdd FILL
XFILL_0__10576_ gnd vdd FILL
XSFILL18920x70050 gnd vdd FILL
XFILL_4__14834_ gnd vdd FILL
X_15559_ _15559_/A _15558_/Y gnd _15559_/Y vdd NOR2X1
XFILL_5__15084_ gnd vdd FILL
XFILL_5_BUFX2_insert909 gnd vdd FILL
XFILL_3__16263_ gnd vdd FILL
X_8490_ _8494_/B _8874_/B gnd _8491_/C vdd NAND2X1
XFILL_5__12296_ gnd vdd FILL
XFILL_2__11136_ gnd vdd FILL
XFILL_0__15103_ gnd vdd FILL
XFILL_3__10687_ gnd vdd FILL
XFILL_3__9660_ gnd vdd FILL
XFILL_3__13475_ gnd vdd FILL
XFILL_0__12315_ gnd vdd FILL
XFILL_1__14654_ gnd vdd FILL
XFILL_3__6872_ gnd vdd FILL
XFILL_1__11866_ gnd vdd FILL
XFILL_0__16083_ gnd vdd FILL
XFILL_0__13295_ gnd vdd FILL
XSFILL59000x63050 gnd vdd FILL
XFILL_5__14035_ gnd vdd FILL
XFILL_0__8902_ gnd vdd FILL
XFILL_3__15214_ gnd vdd FILL
X_7441_ _7441_/A gnd _7443_/A vdd INVX1
XFILL_5__11247_ gnd vdd FILL
XFILL_1__13605_ gnd vdd FILL
XFILL_0__9882_ gnd vdd FILL
XFILL_3__12426_ gnd vdd FILL
XFILL_3__8611_ gnd vdd FILL
XFILL_4__14765_ gnd vdd FILL
XFILL_3__16194_ gnd vdd FILL
XFILL_2__15944_ gnd vdd FILL
XFILL_0__15034_ gnd vdd FILL
XFILL_4__11977_ gnd vdd FILL
XFILL_2__11067_ gnd vdd FILL
XFILL_1__10817_ gnd vdd FILL
XFILL_5__9527_ gnd vdd FILL
XFILL_6__8320_ gnd vdd FILL
XFILL_1__14585_ gnd vdd FILL
XFILL_3__9591_ gnd vdd FILL
XFILL_0__12246_ gnd vdd FILL
XFILL_1__11797_ gnd vdd FILL
XFILL_0__8833_ gnd vdd FILL
XFILL111720x62050 gnd vdd FILL
XFILL_4__13716_ gnd vdd FILL
X_7372_ _7372_/A _7297_/B _7372_/C gnd _7372_/Y vdd OAI21X1
XFILL_4__10928_ gnd vdd FILL
XFILL_2__10018_ gnd vdd FILL
XFILL_3__12357_ gnd vdd FILL
XFILL_1__16324_ gnd vdd FILL
XFILL_5__11178_ gnd vdd FILL
XFILL_3__15145_ gnd vdd FILL
XFILL112200x69050 gnd vdd FILL
XFILL_4__14696_ gnd vdd FILL
XFILL_2__9749_ gnd vdd FILL
XFILL_1__13536_ gnd vdd FILL
XFILL_1__10748_ gnd vdd FILL
XSFILL38840x21050 gnd vdd FILL
XFILL_2__15875_ gnd vdd FILL
X_9111_ _9185_/Q gnd _9111_/Y vdd INVX1
XFILL_0__12177_ gnd vdd FILL
XFILL_0__8764_ gnd vdd FILL
XSFILL64120x54050 gnd vdd FILL
XFILL_3__11308_ gnd vdd FILL
XFILL_5__10129_ gnd vdd FILL
XFILL_4__13647_ gnd vdd FILL
XFILL_2__14826_ gnd vdd FILL
XFILL_5__15986_ gnd vdd FILL
XFILL_3__8473_ gnd vdd FILL
XFILL_3__15076_ gnd vdd FILL
XFILL_3__12288_ gnd vdd FILL
XFILL_1__16255_ gnd vdd FILL
XFILL_1__13467_ gnd vdd FILL
XFILL_0__11128_ gnd vdd FILL
XFILL_1__10679_ gnd vdd FILL
XFILL_0__7715_ gnd vdd FILL
X_9042_ _9042_/A _9017_/A _9041_/Y gnd _9076_/D vdd OAI21X1
XFILL_5__9389_ gnd vdd FILL
XFILL_1__15206_ gnd vdd FILL
XFILL_0__8695_ gnd vdd FILL
XFILL_3__14027_ gnd vdd FILL
XFILL_5__14937_ gnd vdd FILL
XFILL_3__11239_ gnd vdd FILL
XFILL_4__16366_ gnd vdd FILL
XFILL_3__7424_ gnd vdd FILL
XFILL_1__12418_ gnd vdd FILL
XFILL_4__13578_ gnd vdd FILL
XFILL_1__16186_ gnd vdd FILL
XFILL_0__15936_ gnd vdd FILL
XFILL_2__11969_ gnd vdd FILL
XFILL_0__11059_ gnd vdd FILL
XFILL_2__14757_ gnd vdd FILL
XFILL_1__13398_ gnd vdd FILL
XSFILL43960x12050 gnd vdd FILL
XFILL_4__15317_ gnd vdd FILL
XFILL_5__14868_ gnd vdd FILL
XSFILL3560x61050 gnd vdd FILL
XFILL_4__12529_ gnd vdd FILL
XFILL_3__7355_ gnd vdd FILL
XFILL_4__16297_ gnd vdd FILL
XFILL_2__13708_ gnd vdd FILL
XFILL_1__15137_ gnd vdd FILL
XFILL_1__12349_ gnd vdd FILL
XCLKBUF1_insert1077 clk gnd CLKBUF1_insert192/A vdd CLKBUF1
XFILL_6__7064_ gnd vdd FILL
XFILL_0__15867_ gnd vdd FILL
XFILL_2__14688_ gnd vdd FILL
XFILL_5__13819_ gnd vdd FILL
XFILL_4__15248_ gnd vdd FILL
XFILL_0__7577_ gnd vdd FILL
XFILL_5__14799_ gnd vdd FILL
XFILL_3__15978_ gnd vdd FILL
XFILL_2__13639_ gnd vdd FILL
XFILL_0__14818_ gnd vdd FILL
XFILL_3__7286_ gnd vdd FILL
XFILL_1__15068_ gnd vdd FILL
XFILL_0_BUFX2_insert10 gnd vdd FILL
XFILL_0__15798_ gnd vdd FILL
XFILL_0_BUFX2_insert21 gnd vdd FILL
X_9944_ _9852_/A _8663_/CLK _9944_/R vdd _9944_/D gnd vdd DFFSR
XFILL_4__15179_ gnd vdd FILL
XFILL_1__14019_ gnd vdd FILL
XFILL_3__9025_ gnd vdd FILL
XFILL_0_BUFX2_insert32 gnd vdd FILL
XFILL_3__14929_ gnd vdd FILL
XFILL_0_BUFX2_insert43 gnd vdd FILL
XFILL_2__16358_ gnd vdd FILL
XFILL_0__14749_ gnd vdd FILL
XFILL_0_BUFX2_insert54 gnd vdd FILL
XFILL_0_BUFX2_insert65 gnd vdd FILL
XFILL_0__9247_ gnd vdd FILL
XFILL_0_BUFX2_insert76 gnd vdd FILL
XSFILL33880x64050 gnd vdd FILL
XFILL_2__15309_ gnd vdd FILL
X_9875_ _9875_/A _9937_/A _9874_/Y gnd _9951_/D vdd OAI21X1
XFILL_0_BUFX2_insert87 gnd vdd FILL
XFILL_0_BUFX2_insert98 gnd vdd FILL
XFILL_2__16289_ gnd vdd FILL
X_8826_ _8916_/A _8314_/B gnd _8827_/C vdd NAND2X1
XFILL_6_BUFX2_insert710 gnd vdd FILL
XFILL_4__6981_ gnd vdd FILL
XFILL_0__8129_ gnd vdd FILL
XSFILL38920x2050 gnd vdd FILL
X_8757_ _8811_/Q gnd _8757_/Y vdd INVX1
XFILL_4__8720_ gnd vdd FILL
XBUFX2_insert809 _13329_/Y gnd _8969_/A vdd BUFX2
XFILL_1__9991_ gnd vdd FILL
XFILL_3__9927_ gnd vdd FILL
XFILL_6_BUFX2_insert776 gnd vdd FILL
X_7708_ _7708_/A _7672_/B _7708_/C gnd _7778_/D vdd OAI21X1
XFILL_6_BUFX2_insert787 gnd vdd FILL
X_8688_ _8688_/Q _7268_/CLK _8688_/R vdd _8646_/Y gnd vdd DFFSR
XFILL_4__8651_ gnd vdd FILL
XFILL_3__9858_ gnd vdd FILL
XSFILL3640x41050 gnd vdd FILL
X_7639_ _7639_/Q _7515_/CLK _7515_/R vdd _7639_/D gnd vdd DFFSR
XFILL_1__8873_ gnd vdd FILL
XFILL_4__7602_ gnd vdd FILL
XFILL_1_CLKBUF1_insert203 gnd vdd FILL
XSFILL28840x53050 gnd vdd FILL
XFILL_3__9789_ gnd vdd FILL
XFILL_4__8582_ gnd vdd FILL
XFILL_1_CLKBUF1_insert214 gnd vdd FILL
XFILL_1__7824_ gnd vdd FILL
XFILL_6__9498_ gnd vdd FILL
X_11240_ _11238_/Y _11239_/Y _11010_/Y gnd _11240_/Y vdd OAI21X1
XFILL_6__8449_ gnd vdd FILL
X_9309_ _9309_/Q _7147_/CLK _7531_/R vdd _9309_/D gnd vdd DFFSR
XFILL_1__7755_ gnd vdd FILL
XFILL_4__7464_ gnd vdd FILL
X_11171_ _12198_/Y _12326_/Y gnd _11171_/Y vdd NAND2X1
XFILL_1__7686_ gnd vdd FILL
XFILL_3_BUFX2_insert600 gnd vdd FILL
X_10122_ _10122_/A _10127_/A _10122_/C gnd _10204_/D vdd OAI21X1
XFILL_3_BUFX2_insert611 gnd vdd FILL
XFILL_3_BUFX2_insert622 gnd vdd FILL
XFILL_1__9425_ gnd vdd FILL
XFILL_3_BUFX2_insert633 gnd vdd FILL
XSFILL34040x53050 gnd vdd FILL
XFILL_3_BUFX2_insert644 gnd vdd FILL
XFILL_4__9134_ gnd vdd FILL
XFILL_3_BUFX2_insert655 gnd vdd FILL
X_14930_ _9461_/Q _13883_/B _13771_/D _8531_/A gnd _14939_/A vdd AOI22X1
X_10053_ _10054_/B _6981_/B gnd _10053_/Y vdd NAND2X1
XFILL_3_BUFX2_insert666 gnd vdd FILL
XFILL_1__9356_ gnd vdd FILL
XFILL_3_BUFX2_insert677 gnd vdd FILL
XFILL_3_BUFX2_insert688 gnd vdd FILL
XFILL_3_BUFX2_insert699 gnd vdd FILL
XFILL_2__7100_ gnd vdd FILL
X_14861_ _8653_/A gnd _14862_/A vdd INVX1
XFILL_2__8080_ gnd vdd FILL
XFILL_1__9287_ gnd vdd FILL
XSFILL3720x21050 gnd vdd FILL
XFILL_4__8016_ gnd vdd FILL
X_13812_ _8157_/Q gnd _13813_/D vdd INVX1
XFILL_2__7031_ gnd vdd FILL
XFILL_1__8238_ gnd vdd FILL
X_14792_ _8394_/A _13848_/B _13592_/D _7114_/A gnd _14801_/A vdd AOI22X1
XSFILL28920x33050 gnd vdd FILL
X_10955_ _10955_/A _10943_/C _10955_/C gnd _10955_/Y vdd NAND3X1
X_13743_ _10120_/A gnd _13743_/Y vdd INVX1
XSFILL79160x70050 gnd vdd FILL
XFILL_5__8760_ gnd vdd FILL
X_13674_ _13665_/Y _13666_/Y _13674_/C gnd _13674_/Y vdd NAND3X1
X_10886_ _10892_/C _10871_/Y gnd _10888_/B vdd NOR2X1
XFILL_3__11590_ gnd vdd FILL
XFILL_0__10430_ gnd vdd FILL
XFILL_2__8982_ gnd vdd FILL
XFILL_5__7711_ gnd vdd FILL
XFILL_0_BUFX2_insert501 gnd vdd FILL
X_15413_ _15413_/A _15413_/B gnd _15414_/A vdd NOR2X1
X_12625_ vdd memoryOutData[19] gnd _12626_/C vdd NAND2X1
XFILL_4__11900_ gnd vdd FILL
XFILL_5__12150_ gnd vdd FILL
XSFILL99480x19050 gnd vdd FILL
XFILL_4__9898_ gnd vdd FILL
X_16393_ _16393_/A gnd _16393_/Y vdd INVX1
XFILL_3__10541_ gnd vdd FILL
XFILL_0_BUFX2_insert512 gnd vdd FILL
XSFILL74120x17050 gnd vdd FILL
XFILL_0_BUFX2_insert523 gnd vdd FILL
XSFILL74920x36050 gnd vdd FILL
XFILL_4__12880_ gnd vdd FILL
XFILL_1__11720_ gnd vdd FILL
XFILL_2__7933_ gnd vdd FILL
XFILL_0_BUFX2_insert534 gnd vdd FILL
XFILL_0__10361_ gnd vdd FILL
XFILL_0_BUFX2_insert545 gnd vdd FILL
XFILL_4__8849_ gnd vdd FILL
XFILL_5__11101_ gnd vdd FILL
X_15344_ _9821_/Q gnd _15345_/B vdd INVX1
X_12556_ _12406_/A _12538_/CLK _12689_/R vdd _12504_/Y gnd vdd DFFSR
XFILL_3__13260_ gnd vdd FILL
XFILL_0_BUFX2_insert556 gnd vdd FILL
XFILL_5__12081_ gnd vdd FILL
XFILL_4__11831_ gnd vdd FILL
XFILL_0_BUFX2_insert567 gnd vdd FILL
XFILL_0__12100_ gnd vdd FILL
XFILL_0_BUFX2_insert578 gnd vdd FILL
XFILL_2__7864_ gnd vdd FILL
XFILL_1__11651_ gnd vdd FILL
XFILL_0__13080_ gnd vdd FILL
XFILL_2__13990_ gnd vdd FILL
XFILL_0_BUFX2_insert589 gnd vdd FILL
X_11507_ _11505_/Y _11498_/A _11507_/C gnd _11507_/Y vdd AOI21X1
XFILL_0__10292_ gnd vdd FILL
XSFILL99320x83050 gnd vdd FILL
XFILL_3__12211_ gnd vdd FILL
XFILL_5__7573_ gnd vdd FILL
XFILL_5__11032_ gnd vdd FILL
XFILL_4__14550_ gnd vdd FILL
XFILL_2__9603_ gnd vdd FILL
X_12487_ _11936_/B gnd _12489_/A vdd INVX1
X_15275_ _15275_/A gnd _15276_/B vdd INVX1
XFILL_4__11762_ gnd vdd FILL
XFILL_0__12031_ gnd vdd FILL
XFILL_1__14370_ gnd vdd FILL
XFILL_1__11582_ gnd vdd FILL
X_14226_ _7206_/A _13619_/B _13592_/A _8230_/A gnd _14227_/B vdd AOI22X1
X_11438_ _11435_/Y _11550_/C _11437_/Y gnd _11490_/A vdd AOI21X1
XFILL_4__13501_ gnd vdd FILL
XFILL_3__12142_ gnd vdd FILL
XSFILL38760x36050 gnd vdd FILL
XFILL_5__15840_ gnd vdd FILL
XFILL_1__13321_ gnd vdd FILL
XFILL_4__14481_ gnd vdd FILL
XFILL_2__9534_ gnd vdd FILL
XFILL_1__10533_ gnd vdd FILL
XFILL_2__15660_ gnd vdd FILL
XFILL_2__12872_ gnd vdd FILL
XFILL112280x43050 gnd vdd FILL
XFILL_4__11693_ gnd vdd FILL
XSFILL64040x69050 gnd vdd FILL
XFILL_5__9243_ gnd vdd FILL
XFILL_4__16220_ gnd vdd FILL
X_14157_ _14555_/B _15633_/B _14157_/C _13630_/B gnd _14157_/Y vdd OAI22X1
XFILL_4__13432_ gnd vdd FILL
XFILL_5__15771_ gnd vdd FILL
X_11369_ _11209_/Y gnd _11369_/Y vdd INVX1
XFILL_1__16040_ gnd vdd FILL
XFILL_2__14611_ gnd vdd FILL
XFILL_3__12073_ gnd vdd FILL
XCLKBUF1_insert202 CLKBUF1_insert169/A gnd _13184_/CLK vdd CLKBUF1
XFILL_5__12983_ gnd vdd FILL
XFILL_4__10644_ gnd vdd FILL
XFILL_2__11823_ gnd vdd FILL
XFILL_1__13252_ gnd vdd FILL
XCLKBUF1_insert213 CLKBUF1_insert206/A gnd _9188_/CLK vdd CLKBUF1
XFILL_2__9465_ gnd vdd FILL
XCLKBUF1_insert224 CLKBUF1_insert192/A gnd _7129_/CLK vdd CLKBUF1
XFILL_0__7500_ gnd vdd FILL
XFILL_2__15591_ gnd vdd FILL
XFILL_0__13982_ gnd vdd FILL
X_13108_ _13108_/A _13108_/B _13107_/Y gnd _13184_/D vdd OAI21X1
XFILL_5__14722_ gnd vdd FILL
XFILL_3__15901_ gnd vdd FILL
XFILL_5__11934_ gnd vdd FILL
XFILL_0__8480_ gnd vdd FILL
X_14088_ _14088_/A _14045_/A _13879_/B _14088_/D gnd _14092_/A vdd OAI22X1
XFILL_3__11024_ gnd vdd FILL
XFILL_4__16151_ gnd vdd FILL
XFILL_4__13363_ gnd vdd FILL
XFILL_1__12203_ gnd vdd FILL
XFILL_4__10575_ gnd vdd FILL
XFILL_0__15721_ gnd vdd FILL
XFILL_2__14542_ gnd vdd FILL
XFILL_2__11754_ gnd vdd FILL
XSFILL114040x38050 gnd vdd FILL
XSFILL43880x27050 gnd vdd FILL
XFILL_5__8125_ gnd vdd FILL
XFILL_2__9396_ gnd vdd FILL
X_13039_ vdd _13039_/B gnd _13040_/C vdd NAND2X1
XFILL_1__10395_ gnd vdd FILL
XFILL_0__7431_ gnd vdd FILL
XFILL_4__15102_ gnd vdd FILL
XFILL_4__12314_ gnd vdd FILL
XFILL_5__14653_ gnd vdd FILL
XFILL_3__15832_ gnd vdd FILL
XFILL_5__11865_ gnd vdd FILL
XFILL_4__16082_ gnd vdd FILL
XFILL_2__10705_ gnd vdd FILL
XFILL_4__13294_ gnd vdd FILL
XFILL_2__14473_ gnd vdd FILL
XSFILL58920x49050 gnd vdd FILL
XFILL_1__12134_ gnd vdd FILL
XFILL_2__8347_ gnd vdd FILL
XFILL_0__15652_ gnd vdd FILL
XFILL_2__11685_ gnd vdd FILL
XFILL_5__13604_ gnd vdd FILL
XFILL_5__8056_ gnd vdd FILL
XFILL_0__12864_ gnd vdd FILL
XFILL_5__10816_ gnd vdd FILL
XFILL_4__15033_ gnd vdd FILL
XFILL_0__7362_ gnd vdd FILL
XFILL_2__16212_ gnd vdd FILL
XFILL_5__14584_ gnd vdd FILL
XFILL_2__13424_ gnd vdd FILL
XFILL_4__12245_ gnd vdd FILL
X_7990_ _7948_/A _7990_/B gnd _7991_/C vdd NAND2X1
XFILL_2__10636_ gnd vdd FILL
XFILL_0__14603_ gnd vdd FILL
XSFILL84360x41050 gnd vdd FILL
XFILL_3__15763_ gnd vdd FILL
XFILL_3__7071_ gnd vdd FILL
XFILL_5__11796_ gnd vdd FILL
XFILL_0__9101_ gnd vdd FILL
XFILL_3__12975_ gnd vdd FILL
XFILL_1__12065_ gnd vdd FILL
XSFILL34200x13050 gnd vdd FILL
XFILL_0__11815_ gnd vdd FILL
XFILL_5__16323_ gnd vdd FILL
XFILL_0__15583_ gnd vdd FILL
XFILL_5__13535_ gnd vdd FILL
XFILL_2__7229_ gnd vdd FILL
XFILL_3__14714_ gnd vdd FILL
X_6941_ _7011_/Q gnd _6943_/A vdd INVX1
XFILL_5__10747_ gnd vdd FILL
XFILL_0__7293_ gnd vdd FILL
XFILL_6__15874_ gnd vdd FILL
XFILL_2__13355_ gnd vdd FILL
XFILL_3__11926_ gnd vdd FILL
XFILL_2__16143_ gnd vdd FILL
XFILL_4__12176_ gnd vdd FILL
XFILL_1__11016_ gnd vdd FILL
XSFILL99400x63050 gnd vdd FILL
XFILL_3__15694_ gnd vdd FILL
XFILL_0__14534_ gnd vdd FILL
XFILL_2__10567_ gnd vdd FILL
XFILL_0__11746_ gnd vdd FILL
XFILL_0__9032_ gnd vdd FILL
XFILL_3_CLKBUF1_insert180 gnd vdd FILL
XFILL_6__14825_ gnd vdd FILL
XFILL_5__16254_ gnd vdd FILL
X_9660_ _9639_/A _8636_/B gnd _9660_/Y vdd NAND2X1
XFILL_5__13466_ gnd vdd FILL
XFILL_2__12306_ gnd vdd FILL
XFILL_4__11127_ gnd vdd FILL
XFILL_5__10678_ gnd vdd FILL
XFILL_3_CLKBUF1_insert191 gnd vdd FILL
XFILL_3__14645_ gnd vdd FILL
XFILL_2__16074_ gnd vdd FILL
X_6872_ _6872_/A gnd memoryWriteData[2] vdd BUFX2
XFILL_2__13286_ gnd vdd FILL
XFILL_1__15824_ gnd vdd FILL
XFILL_3__11857_ gnd vdd FILL
XFILL_0__14465_ gnd vdd FILL
XFILL_5__15205_ gnd vdd FILL
XFILL_2__10498_ gnd vdd FILL
XSFILL38840x16050 gnd vdd FILL
XFILL_5__12417_ gnd vdd FILL
X_8611_ _8611_/A gnd _8611_/Y vdd INVX1
XFILL_5__8958_ gnd vdd FILL
XFILL_0__11677_ gnd vdd FILL
XFILL_6__7751_ gnd vdd FILL
XFILL_5__16185_ gnd vdd FILL
XFILL_2__15025_ gnd vdd FILL
XFILL_4__15935_ gnd vdd FILL
XFILL_6__11968_ gnd vdd FILL
XFILL_4__11058_ gnd vdd FILL
XFILL112360x23050 gnd vdd FILL
XFILL_0__16204_ gnd vdd FILL
XFILL_5__13397_ gnd vdd FILL
XSFILL64120x49050 gnd vdd FILL
X_9591_ _8183_/A _9675_/A gnd _9591_/Y vdd NAND2X1
XFILL_3__10808_ gnd vdd FILL
XFILL_2__12237_ gnd vdd FILL
XFILL_3__14576_ gnd vdd FILL
XFILL_0__13416_ gnd vdd FILL
XFILL_3__7973_ gnd vdd FILL
XFILL_0__10628_ gnd vdd FILL
XFILL_3__11788_ gnd vdd FILL
XFILL_1__12967_ gnd vdd FILL
XFILL_1__15755_ gnd vdd FILL
XFILL_0__14396_ gnd vdd FILL
XFILL_5__15136_ gnd vdd FILL
X_8542_ _8542_/Q _9817_/CLK _8542_/R vdd _8542_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert390 gnd vdd FILL
XFILL_5__8889_ gnd vdd FILL
XFILL_4__10009_ gnd vdd FILL
XFILL_5__12348_ gnd vdd FILL
XFILL_3__16315_ gnd vdd FILL
XFILL_3__13527_ gnd vdd FILL
XFILL_6__14687_ gnd vdd FILL
XFILL_4__15866_ gnd vdd FILL
XFILL_3__6924_ gnd vdd FILL
XFILL_5_BUFX2_insert706 gnd vdd FILL
XFILL_1__14706_ gnd vdd FILL
XFILL_1__11918_ gnd vdd FILL
XFILL_2__12168_ gnd vdd FILL
XFILL_0__16135_ gnd vdd FILL
XFILL_0__13347_ gnd vdd FILL
XFILL_1__15686_ gnd vdd FILL
XFILL_5_BUFX2_insert717 gnd vdd FILL
XFILL_0__10559_ gnd vdd FILL
XSFILL79320x30050 gnd vdd FILL
XFILL_1__12898_ gnd vdd FILL
XFILL_0__9934_ gnd vdd FILL
XFILL_6__13638_ gnd vdd FILL
XFILL_4__14817_ gnd vdd FILL
XFILL_5__15067_ gnd vdd FILL
XFILL_5_BUFX2_insert728 gnd vdd FILL
X_8473_ _8471_/Y _8503_/B _8473_/C gnd _8545_/D vdd OAI21X1
XSFILL3560x56050 gnd vdd FILL
XFILL_5_BUFX2_insert739 gnd vdd FILL
XFILL_5__12279_ gnd vdd FILL
XFILL_2__11119_ gnd vdd FILL
XFILL_3__16246_ gnd vdd FILL
XFILL_1__14637_ gnd vdd FILL
XFILL_3__13458_ gnd vdd FILL
XFILL_4__15797_ gnd vdd FILL
XFILL_3__9643_ gnd vdd FILL
XSFILL93560x78050 gnd vdd FILL
XFILL_2__12099_ gnd vdd FILL
XFILL_3__6855_ gnd vdd FILL
XFILL_0__16066_ gnd vdd FILL
XFILL_1__11849_ gnd vdd FILL
XFILL_0__13278_ gnd vdd FILL
XFILL_5__14018_ gnd vdd FILL
X_7424_ _7425_/B _7424_/B gnd _7424_/Y vdd NAND2X1
XSFILL28760x68050 gnd vdd FILL
XFILL_3__12409_ gnd vdd FILL
XFILL_0__9865_ gnd vdd FILL
XFILL_4__14748_ gnd vdd FILL
XFILL_2__15927_ gnd vdd FILL
XFILL_3__16177_ gnd vdd FILL
XFILL_0__15017_ gnd vdd FILL
XSFILL44040x16050 gnd vdd FILL
XFILL_1__14568_ gnd vdd FILL
XFILL_3__13389_ gnd vdd FILL
XSFILL115000x46050 gnd vdd FILL
XFILL_0__12229_ gnd vdd FILL
X_7355_ _7355_/A gnd _7357_/A vdd INVX1
XFILL_6__16288_ gnd vdd FILL
XFILL_3__15128_ gnd vdd FILL
XFILL_3__8525_ gnd vdd FILL
XFILL_0__9796_ gnd vdd FILL
XFILL_1__16307_ gnd vdd FILL
XFILL_4__14679_ gnd vdd FILL
XFILL_1__13519_ gnd vdd FILL
XFILL_2__15858_ gnd vdd FILL
XFILL_1__14499_ gnd vdd FILL
XFILL_6__15239_ gnd vdd FILL
XFILL_0__8747_ gnd vdd FILL
XFILL_5__15969_ gnd vdd FILL
XFILL_2__14809_ gnd vdd FILL
XSFILL33880x59050 gnd vdd FILL
X_7286_ _7286_/A gnd _7286_/Y vdd INVX1
XFILL_3__15059_ gnd vdd FILL
XFILL_1__16238_ gnd vdd FILL
XFILL_3__8456_ gnd vdd FILL
XFILL_2__15789_ gnd vdd FILL
X_9025_ _9025_/A gnd _9027_/A vdd INVX1
XFILL_1__7471_ gnd vdd FILL
XFILL_4__16349_ gnd vdd FILL
XFILL_4__7180_ gnd vdd FILL
XFILL_1__16169_ gnd vdd FILL
XFILL_0__15919_ gnd vdd FILL
XFILL_3__8387_ gnd vdd FILL
XFILL_1__9210_ gnd vdd FILL
XFILL_0__7629_ gnd vdd FILL
XFILL_3__7338_ gnd vdd FILL
XFILL_2_BUFX2_insert607 gnd vdd FILL
XFILL_1__9141_ gnd vdd FILL
XSFILL89960x52050 gnd vdd FILL
XFILL_2_BUFX2_insert618 gnd vdd FILL
XFILL_2_BUFX2_insert629 gnd vdd FILL
XSFILL3640x36050 gnd vdd FILL
XFILL_3__9008_ gnd vdd FILL
X_9927_ _9969_/Q gnd _9927_/Y vdd INVX1
XSFILL28840x48050 gnd vdd FILL
X_9858_ _9946_/Q gnd _9858_/Y vdd INVX1
X_10740_ _14882_/A _8180_/CLK _7391_/R vdd _10740_/D gnd vdd DFFSR
XSFILL28440x50050 gnd vdd FILL
X_8809_ _8809_/Q _7664_/CLK _7920_/R vdd _8753_/Y gnd vdd DFFSR
X_9789_ _9787_/Y _9789_/B _9788_/Y gnd _9789_/Y vdd OAI21X1
XFILL_4__9752_ gnd vdd FILL
XBUFX2_insert606 BUFX2_insert570/A gnd _8285_/R vdd BUFX2
XFILL_6_BUFX2_insert551 gnd vdd FILL
XFILL_4__6964_ gnd vdd FILL
XBUFX2_insert617 _10926_/Y gnd _12007_/A vdd BUFX2
XSFILL33960x39050 gnd vdd FILL
X_10671_ _10671_/A gnd _10671_/Y vdd INVX1
XBUFX2_insert628 _13465_/Y gnd _14865_/C vdd BUFX2
XFILL_4__8703_ gnd vdd FILL
XFILL_1__9974_ gnd vdd FILL
XBUFX2_insert639 _12438_/Y gnd _9556_/B vdd BUFX2
X_12410_ _12368_/A _12633_/A gnd _12411_/C vdd NAND2X1
XFILL_4__9683_ gnd vdd FILL
X_13390_ _13423_/A _13390_/B gnd _13390_/Y vdd NAND2X1
XFILL_4__6895_ gnd vdd FILL
XSFILL104520x71050 gnd vdd FILL
XFILL_4__8634_ gnd vdd FILL
X_12341_ _6901_/A _12301_/B _12301_/C _12313_/D gnd _12342_/C vdd AOI22X1
XFILL_1__8856_ gnd vdd FILL
XSFILL89240x13050 gnd vdd FILL
XSFILL59080x4050 gnd vdd FILL
X_15060_ _13421_/Y _15386_/B gnd _15067_/B vdd NOR2X1
X_12272_ _12272_/A _11882_/B _12272_/C gnd _12274_/B vdd NAND3X1
XFILL_1__7807_ gnd vdd FILL
XFILL_2__7580_ gnd vdd FILL
X_14011_ _14011_/A _14010_/Y gnd _14012_/C vdd NOR2X1
XSFILL3720x16050 gnd vdd FILL
XFILL_1__8787_ gnd vdd FILL
X_11223_ _10988_/Y _11223_/B gnd _11223_/Y vdd NAND2X1
XFILL_4__8496_ gnd vdd FILL
XFILL_1__7738_ gnd vdd FILL
XSFILL28920x28050 gnd vdd FILL
XFILL_4__7447_ gnd vdd FILL
X_11154_ _12294_/Y _11125_/A gnd _11154_/Y vdd NOR2X1
XSFILL13720x70050 gnd vdd FILL
XFILL_2__9250_ gnd vdd FILL
XFILL_3_BUFX2_insert430 gnd vdd FILL
X_10105_ _13523_/A gnd _10107_/A vdd INVX1
XSFILL79160x65050 gnd vdd FILL
XFILL_3_BUFX2_insert441 gnd vdd FILL
XFILL_4__7378_ gnd vdd FILL
XFILL_1__9408_ gnd vdd FILL
XFILL_2__8201_ gnd vdd FILL
XFILL_4__10360_ gnd vdd FILL
X_15962_ _15962_/A gnd _15964_/D vdd INVX1
X_11085_ _11393_/A _11074_/C _11085_/C gnd _11085_/Y vdd AOI21X1
XFILL_3_BUFX2_insert452 gnd vdd FILL
XFILL_3_BUFX2_insert463 gnd vdd FILL
XFILL_4__9117_ gnd vdd FILL
XFILL_3_BUFX2_insert474 gnd vdd FILL
XFILL_1__10180_ gnd vdd FILL
X_10036_ _10034_/Y _10054_/B _10036_/C gnd _10090_/D vdd OAI21X1
XFILL_3_BUFX2_insert485 gnd vdd FILL
X_14913_ _7796_/Q gnd _16272_/D vdd INVX1
XFILL_3_BUFX2_insert496 gnd vdd FILL
XFILL_2__8132_ gnd vdd FILL
XFILL_5__11650_ gnd vdd FILL
X_15893_ _14495_/Y _16002_/A gnd _15893_/Y vdd NOR2X1
XSFILL8440x28050 gnd vdd FILL
XFILL_1__9339_ gnd vdd FILL
XFILL_4__10291_ gnd vdd FILL
XFILL_2__11470_ gnd vdd FILL
XFILL_5__9930_ gnd vdd FILL
X_14844_ _14842_/Y _14583_/B _14555_/C _14843_/Y gnd _14844_/Y vdd OAI22X1
XSFILL84280x56050 gnd vdd FILL
XFILL_4__12030_ gnd vdd FILL
XFILL_2__10421_ gnd vdd FILL
XFILL_2__8063_ gnd vdd FILL
XFILL_5__11581_ gnd vdd FILL
XFILL_3__12760_ gnd vdd FILL
XFILL_0__11600_ gnd vdd FILL
XFILL_5__13320_ gnd vdd FILL
XFILL_0__12580_ gnd vdd FILL
XFILL_5__9861_ gnd vdd FILL
XFILL_5__10532_ gnd vdd FILL
XSFILL99320x78050 gnd vdd FILL
XFILL_2__13140_ gnd vdd FILL
XSFILL59080x32050 gnd vdd FILL
XFILL_3__11711_ gnd vdd FILL
X_14775_ _14775_/A _14774_/Y _14772_/Y gnd _14790_/B vdd NAND3X1
X_11987_ _11987_/A _12072_/A gnd _11987_/Y vdd NOR2X1
XFILL_0_BUFX2_insert2 gnd vdd FILL
XFILL_1__13870_ gnd vdd FILL
XFILL_0__11531_ gnd vdd FILL
XFILL_6__14610_ gnd vdd FILL
XFILL_5__13251_ gnd vdd FILL
XFILL_5__9792_ gnd vdd FILL
X_13726_ _13722_/Y _13726_/B gnd _13726_/Y vdd NOR2X1
X_10938_ _10938_/A _10938_/B gnd _10943_/C vdd NOR2X1
XFILL_3__14430_ gnd vdd FILL
XFILL_4_CLKBUF1_insert220 gnd vdd FILL
XFILL_4__13981_ gnd vdd FILL
XFILL_3__11642_ gnd vdd FILL
XFILL_0__14250_ gnd vdd FILL
XFILL112280x38050 gnd vdd FILL
XFILL_2__10283_ gnd vdd FILL
XFILL_5__8743_ gnd vdd FILL
XFILL_5__12202_ gnd vdd FILL
XFILL_0__11462_ gnd vdd FILL
XFILL_4__15720_ gnd vdd FILL
X_16445_ _14816_/A _8562_/CLK _7270_/R vdd _16407_/Y gnd vdd DFFSR
XFILL_6__11753_ gnd vdd FILL
X_13657_ _8706_/A gnd _13657_/Y vdd INVX1
XFILL_2__12022_ gnd vdd FILL
X_10869_ _10869_/Q _9447_/CLK _9447_/R vdd _10869_/D gnd vdd DFFSR
XFILL_1__15540_ gnd vdd FILL
XFILL_5__10394_ gnd vdd FILL
XFILL_3__14361_ gnd vdd FILL
XFILL_3__11573_ gnd vdd FILL
XFILL_1__12752_ gnd vdd FILL
XFILL_0_BUFX2_insert320 gnd vdd FILL
XFILL_0__10413_ gnd vdd FILL
XFILL_2__8965_ gnd vdd FILL
XFILL_0__14181_ gnd vdd FILL
XFILL_6__14472_ gnd vdd FILL
X_12608_ _12606_/Y vdd _12608_/C gnd _12608_/Y vdd OAI21X1
XSFILL13800x50050 gnd vdd FILL
XFILL_5__12133_ gnd vdd FILL
XFILL_3__16100_ gnd vdd FILL
XSFILL74200x6050 gnd vdd FILL
XFILL_0__11393_ gnd vdd FILL
XFILL_0_BUFX2_insert331 gnd vdd FILL
XFILL_3__13312_ gnd vdd FILL
XFILL_4__15651_ gnd vdd FILL
XFILL_3__10524_ gnd vdd FILL
XFILL_0__7980_ gnd vdd FILL
X_16376_ gnd gnd gnd _16377_/C vdd NAND2X1
XFILL_0_BUFX2_insert342 gnd vdd FILL
XFILL_0_BUFX2_insert353 gnd vdd FILL
X_13588_ _10201_/Q gnd _13588_/Y vdd INVX1
XFILL_1__11703_ gnd vdd FILL
XFILL_4__12863_ gnd vdd FILL
XSFILL79240x45050 gnd vdd FILL
XFILL_0__13132_ gnd vdd FILL
XFILL_0_BUFX2_insert364 gnd vdd FILL
XFILL_1__15471_ gnd vdd FILL
XFILL_3__14292_ gnd vdd FILL
XFILL_2__8896_ gnd vdd FILL
XFILL_0_BUFX2_insert375 gnd vdd FILL
XFILL_5__7625_ gnd vdd FILL
XFILL_4__14602_ gnd vdd FILL
X_15327_ _7688_/A gnd _15328_/D vdd INVX1
XFILL_6__13423_ gnd vdd FILL
XFILL_3__16031_ gnd vdd FILL
XFILL_0_BUFX2_insert386 gnd vdd FILL
XFILL_5__12064_ gnd vdd FILL
X_12539_ _12355_/A _12537_/CLK _12536_/R vdd _12539_/D gnd vdd DFFSR
XFILL_0__6931_ gnd vdd FILL
XFILL_4__11814_ gnd vdd FILL
XFILL_3__13243_ gnd vdd FILL
XFILL_0_BUFX2_insert397 gnd vdd FILL
XFILL_4__15582_ gnd vdd FILL
XFILL_1__14422_ gnd vdd FILL
XFILL_2__7847_ gnd vdd FILL
XFILL_1__11634_ gnd vdd FILL
XFILL_0__10275_ gnd vdd FILL
XFILL_2__13973_ gnd vdd FILL
XFILL_5__7556_ gnd vdd FILL
XSFILL114440x54050 gnd vdd FILL
XFILL_5__11015_ gnd vdd FILL
XFILL_0__6862_ gnd vdd FILL
XFILL_4__14533_ gnd vdd FILL
X_15258_ _15241_/Y _15258_/B gnd _15258_/Y vdd NOR2X1
XFILL_0__9650_ gnd vdd FILL
XFILL_2__15712_ gnd vdd FILL
XFILL_3__13174_ gnd vdd FILL
XFILL_4__11745_ gnd vdd FILL
XFILL_0__12014_ gnd vdd FILL
XFILL_1__14353_ gnd vdd FILL
XFILL_3__10386_ gnd vdd FILL
XFILL_6__12305_ gnd vdd FILL
XFILL_1__11565_ gnd vdd FILL
X_14209_ _7971_/A gnd _15663_/B vdd INVX1
XFILL_0__8601_ gnd vdd FILL
XFILL_6__16073_ gnd vdd FILL
XFILL_6__13285_ gnd vdd FILL
XFILL_5__7487_ gnd vdd FILL
X_7140_ _7072_/A _8541_/CLK _7140_/R vdd _7140_/D gnd vdd DFFSR
XFILL_5__15823_ gnd vdd FILL
XFILL_1__13304_ gnd vdd FILL
XFILL_6__10497_ gnd vdd FILL
XFILL_4__14464_ gnd vdd FILL
X_15189_ _10623_/A gnd _15191_/C vdd INVX1
XFILL_3__12125_ gnd vdd FILL
XFILL_3__8310_ gnd vdd FILL
XFILL_2__9517_ gnd vdd FILL
XFILL_2__15643_ gnd vdd FILL
XFILL_4__11676_ gnd vdd FILL
XFILL_1__10516_ gnd vdd FILL
XFILL_5__9226_ gnd vdd FILL
XFILL_3__9290_ gnd vdd FILL
XSFILL59160x12050 gnd vdd FILL
XFILL_2__12855_ gnd vdd FILL
XFILL_1__14284_ gnd vdd FILL
XSFILL99400x58050 gnd vdd FILL
XFILL_4__16203_ gnd vdd FILL
XFILL_1__11496_ gnd vdd FILL
XFILL_4__13415_ gnd vdd FILL
XFILL_0__8532_ gnd vdd FILL
XFILL_1__16023_ gnd vdd FILL
XFILL_4__10627_ gnd vdd FILL
XFILL_3__12056_ gnd vdd FILL
X_7071_ _7069_/Y _7061_/A _7071_/C gnd _7139_/D vdd OAI21X1
XFILL_5__15754_ gnd vdd FILL
XFILL_5__12966_ gnd vdd FILL
XFILL_1__13235_ gnd vdd FILL
XFILL_5_BUFX2_insert1010 gnd vdd FILL
XFILL_4__14395_ gnd vdd FILL
XFILL_2__11806_ gnd vdd FILL
XFILL_3__8241_ gnd vdd FILL
XFILL_2__12786_ gnd vdd FILL
XFILL_1__10447_ gnd vdd FILL
XFILL_2__15574_ gnd vdd FILL
XFILL_5_BUFX2_insert1021 gnd vdd FILL
XFILL_5_BUFX2_insert1032 gnd vdd FILL
XFILL_5__9157_ gnd vdd FILL
XFILL_0__13965_ gnd vdd FILL
XFILL_5_BUFX2_insert1043 gnd vdd FILL
XFILL_0__8463_ gnd vdd FILL
XFILL_5__14705_ gnd vdd FILL
XFILL_5__11917_ gnd vdd FILL
XFILL_6__12167_ gnd vdd FILL
XFILL111880x11050 gnd vdd FILL
XFILL_3__11007_ gnd vdd FILL
XFILL_4__16134_ gnd vdd FILL
XFILL_4__13346_ gnd vdd FILL
XFILL_5__15685_ gnd vdd FILL
XFILL112360x18050 gnd vdd FILL
XFILL_4__10558_ gnd vdd FILL
XFILL_5_BUFX2_insert1054 gnd vdd FILL
XFILL_5__12897_ gnd vdd FILL
XFILL_2__14525_ gnd vdd FILL
XFILL_2__9379_ gnd vdd FILL
XFILL_1__13166_ gnd vdd FILL
XFILL_0__15704_ gnd vdd FILL
XFILL_0__12916_ gnd vdd FILL
XFILL_5__8108_ gnd vdd FILL
XFILL_2__11737_ gnd vdd FILL
XFILL_5_BUFX2_insert1065 gnd vdd FILL
XFILL_1__10378_ gnd vdd FILL
XFILL_0__7414_ gnd vdd FILL
XFILL_6__11118_ gnd vdd FILL
XFILL_5_BUFX2_insert1087 gnd vdd FILL
XFILL_5__9088_ gnd vdd FILL
XFILL_0__13896_ gnd vdd FILL
XFILL_5__14636_ gnd vdd FILL
XFILL_0__8394_ gnd vdd FILL
XFILL_3__7123_ gnd vdd FILL
XFILL_3__15815_ gnd vdd FILL
XFILL_4__16065_ gnd vdd FILL
XFILL_5__11848_ gnd vdd FILL
XFILL_4__13277_ gnd vdd FILL
XSFILL109400x43050 gnd vdd FILL
XFILL_1__12117_ gnd vdd FILL
XFILL_2__14456_ gnd vdd FILL
XFILL_0__15635_ gnd vdd FILL
XFILL_4__10489_ gnd vdd FILL
XFILL_2__11668_ gnd vdd FILL
XFILL_0__12847_ gnd vdd FILL
XFILL_1__13097_ gnd vdd FILL
XFILL_0__7345_ gnd vdd FILL
XFILL_4__15016_ gnd vdd FILL
XSFILL79320x25050 gnd vdd FILL
XFILL_5__14567_ gnd vdd FILL
XFILL_4__12228_ gnd vdd FILL
XFILL_3__7054_ gnd vdd FILL
X_7973_ _7973_/A _7972_/A _7973_/C gnd _8037_/D vdd OAI21X1
XFILL_2__13407_ gnd vdd FILL
XFILL_3__15746_ gnd vdd FILL
XFILL_2__10619_ gnd vdd FILL
XFILL_5__11779_ gnd vdd FILL
XFILL_1__12048_ gnd vdd FILL
XFILL_3__12958_ gnd vdd FILL
XFILL_0__15566_ gnd vdd FILL
XFILL_2__14387_ gnd vdd FILL
XFILL_2__11599_ gnd vdd FILL
XFILL_0__12778_ gnd vdd FILL
X_9712_ _9712_/Q _9953_/CLK _7276_/R vdd _9712_/D gnd vdd DFFSR
XFILL_5__16306_ gnd vdd FILL
XFILL_6__8852_ gnd vdd FILL
XFILL_5__13518_ gnd vdd FILL
X_6924_ _6967_/B _6924_/B gnd _6925_/C vdd NAND2X1
XFILL_5__14498_ gnd vdd FILL
XFILL_3__11909_ gnd vdd FILL
XFILL_4__12159_ gnd vdd FILL
XFILL_2__16126_ gnd vdd FILL
XFILL_2__13338_ gnd vdd FILL
XFILL_3__15677_ gnd vdd FILL
XFILL_0__14517_ gnd vdd FILL
XFILL_0__9015_ gnd vdd FILL
XFILL_3__12889_ gnd vdd FILL
XFILL_6__7803_ gnd vdd FILL
XFILL_0__11729_ gnd vdd FILL
XFILL_0__15497_ gnd vdd FILL
XFILL_5__16237_ gnd vdd FILL
XFILL_5__13449_ gnd vdd FILL
X_9643_ _9641_/Y _9628_/B _9642_/Y gnd _9703_/D vdd OAI21X1
XFILL_3__14628_ gnd vdd FILL
X_6855_ _6855_/A gnd memoryAddress[17] vdd BUFX2
XFILL_2__13269_ gnd vdd FILL
XFILL_1__15807_ gnd vdd FILL
XFILL_2__16057_ gnd vdd FILL
XFILL_3_BUFX2_insert1091 gnd vdd FILL
XFILL_0__14448_ gnd vdd FILL
XFILL_1__13999_ gnd vdd FILL
XFILL_5__16168_ gnd vdd FILL
XFILL_4__15918_ gnd vdd FILL
X_9574_ _9574_/Q _7411_/CLK _7411_/R vdd _9512_/Y gnd vdd DFFSR
XFILL_2__15008_ gnd vdd FILL
XFILL_3__14559_ gnd vdd FILL
XFILL_1__15738_ gnd vdd FILL
XFILL_3__7956_ gnd vdd FILL
XFILL_5_BUFX2_insert503 gnd vdd FILL
XFILL_0__14379_ gnd vdd FILL
XFILL_5__15119_ gnd vdd FILL
X_8525_ _8525_/A gnd _8527_/A vdd INVX1
XFILL_5_BUFX2_insert514 gnd vdd FILL
XFILL_5__16099_ gnd vdd FILL
XFILL_5_BUFX2_insert525 gnd vdd FILL
XFILL_1__6971_ gnd vdd FILL
XFILL_5_BUFX2_insert536 gnd vdd FILL
XFILL_0__16118_ gnd vdd FILL
XFILL_4__15849_ gnd vdd FILL
XFILL_3__6907_ gnd vdd FILL
XFILL_3__7887_ gnd vdd FILL
XFILL_5_BUFX2_insert547 gnd vdd FILL
XFILL_1__15669_ gnd vdd FILL
XFILL_0__9917_ gnd vdd FILL
XFILL_5_BUFX2_insert558 gnd vdd FILL
XFILL_1__8710_ gnd vdd FILL
XFILL_3__16229_ gnd vdd FILL
X_8456_ _8540_/Q gnd _8456_/Y vdd INVX1
XFILL_5_BUFX2_insert569 gnd vdd FILL
XFILL_6__7596_ gnd vdd FILL
XFILL_3_BUFX2_insert6 gnd vdd FILL
XFILL_3__9626_ gnd vdd FILL
XFILL_3__6838_ gnd vdd FILL
XFILL_0__16049_ gnd vdd FILL
X_7407_ _7361_/A _7535_/CLK _8682_/R vdd _7407_/D gnd vdd DFFSR
XFILL_0__9848_ gnd vdd FILL
XFILL_1__8641_ gnd vdd FILL
X_8387_ _8385_/Y _8372_/B _8387_/C gnd _8387_/Y vdd OAI21X1
XSFILL18840x1050 gnd vdd FILL
XFILL_3__9557_ gnd vdd FILL
XFILL_4__8350_ gnd vdd FILL
X_7338_ _7323_/A _8874_/B gnd _7339_/C vdd NAND2X1
XFILL_3_BUFX2_insert80 gnd vdd FILL
XFILL_3__8508_ gnd vdd FILL
XFILL_1__8572_ gnd vdd FILL
XFILL_4__7301_ gnd vdd FILL
XFILL_0__9779_ gnd vdd FILL
XFILL_3_BUFX2_insert91 gnd vdd FILL
XFILL_3__9488_ gnd vdd FILL
XFILL_2_CLKBUF1_insert117 gnd vdd FILL
XFILL_2_CLKBUF1_insert128 gnd vdd FILL
XSFILL94280x19050 gnd vdd FILL
X_7269_ _7269_/Q _7269_/CLK _7262_/R vdd _7269_/D gnd vdd DFFSR
XFILL_2_CLKBUF1_insert139 gnd vdd FILL
XFILL_4__7232_ gnd vdd FILL
XFILL_3__8439_ gnd vdd FILL
XFILL_6__8148_ gnd vdd FILL
X_9008_ _9017_/A _9008_/B gnd _9008_/Y vdd NAND2X1
XFILL_1__7454_ gnd vdd FILL
XFILL_4__7163_ gnd vdd FILL
XFILL_2_BUFX2_insert404 gnd vdd FILL
XFILL_2_BUFX2_insert415 gnd vdd FILL
XFILL_2_BUFX2_insert426 gnd vdd FILL
XFILL_4__7094_ gnd vdd FILL
X_11910_ _11910_/A _11909_/A _11910_/C gnd _6845_/A vdd OAI21X1
XFILL_2_BUFX2_insert437 gnd vdd FILL
XFILL_1__9124_ gnd vdd FILL
XFILL_2_BUFX2_insert448 gnd vdd FILL
X_12890_ vdd _12890_/B gnd _12891_/C vdd NAND2X1
XFILL_2_BUFX2_insert459 gnd vdd FILL
XSFILL104520x66050 gnd vdd FILL
XSFILL73960x41050 gnd vdd FILL
XSFILL8760x64050 gnd vdd FILL
XSFILL23800x13050 gnd vdd FILL
X_11841_ _11840_/Y _11841_/B gnd _11993_/A vdd OR2X2
XSFILL84200x1050 gnd vdd FILL
X_14560_ _9453_/Q _13883_/B _13621_/B _10349_/Q gnd _14560_/Y vdd AOI22X1
XFILL_1__8006_ gnd vdd FILL
X_11772_ _11772_/A _11765_/Y _11772_/C gnd _11772_/Y vdd NAND3X1
XFILL_4__9804_ gnd vdd FILL
X_10723_ _15590_/A _9077_/CLK _7665_/R vdd _10723_/D gnd vdd DFFSR
X_13511_ _13511_/A _13510_/Y gnd _13519_/B vdd NOR2X1
XFILL_4__7996_ gnd vdd FILL
XBUFX2_insert403 _10920_/Y gnd _12359_/A vdd BUFX2
X_14491_ _9653_/A gnd _14491_/Y vdd INVX1
XBUFX2_insert414 _13484_/Y gnd _14956_/D vdd BUFX2
XBUFX2_insert425 _15047_/Y gnd _15384_/D vdd BUFX2
XFILL_4__9735_ gnd vdd FILL
X_16230_ _16230_/A _16230_/B gnd _16231_/B vdd NOR2X1
XFILL_4__6947_ gnd vdd FILL
XBUFX2_insert436 _13326_/Y gnd _8695_/B vdd BUFX2
X_13442_ _13443_/A _13718_/B _13465_/C gnd _13442_/Y vdd NAND3X1
X_10654_ _10619_/B _9374_/B gnd _10655_/C vdd NAND2X1
XBUFX2_insert447 _13276_/Y gnd _7210_/A vdd BUFX2
XBUFX2_insert458 _13442_/Y gnd _14203_/C vdd BUFX2
XFILL_2__8750_ gnd vdd FILL
XBUFX2_insert469 _13318_/Y gnd _8365_/A vdd BUFX2
XFILL_4__9666_ gnd vdd FILL
X_13373_ _14506_/A gnd _14868_/A vdd INVX8
X_16161_ _16161_/A _16160_/Y gnd _16161_/Y vdd NOR2X1
XFILL_4__6878_ gnd vdd FILL
X_10585_ _10495_/A _8942_/CLK _9561_/R vdd _10585_/D gnd vdd DFFSR
XFILL_1__8908_ gnd vdd FILL
XFILL_2__7701_ gnd vdd FILL
XFILL_4__8617_ gnd vdd FILL
XFILL_1__9888_ gnd vdd FILL
X_15112_ _15111_/Y _15110_/Y gnd _15113_/B vdd NOR2X1
XFILL_5__8390_ gnd vdd FILL
X_12324_ _12312_/A _12340_/B _12300_/C gnd _12326_/B vdd NAND3X1
XFILL_4__9597_ gnd vdd FILL
XFILL_3__10240_ gnd vdd FILL
X_16092_ _16091_/Y _15070_/C gnd _16093_/C vdd NOR2X1
XFILL_1__8839_ gnd vdd FILL
XFILL_2__7632_ gnd vdd FILL
XFILL_2__10970_ gnd vdd FILL
XFILL_0__10060_ gnd vdd FILL
XFILL_5__7341_ gnd vdd FILL
X_15043_ _14989_/A _15636_/B _15024_/C gnd _15726_/A vdd NAND3X1
X_12255_ _12255_/A gnd _12255_/C gnd _12255_/Y vdd NAND3X1
XFILL_4__11530_ gnd vdd FILL
XFILL_3__10171_ gnd vdd FILL
XFILL_2__7563_ gnd vdd FILL
XFILL_1__11350_ gnd vdd FILL
X_11206_ _11200_/Y _11201_/Y _11334_/A gnd _11206_/Y vdd OAI21X1
XFILL_4__8479_ gnd vdd FILL
X_12186_ _12184_/Y _12179_/A _12186_/C gnd _12186_/Y vdd OAI21X1
XFILL_2__12640_ gnd vdd FILL
XFILL_1__10301_ gnd vdd FILL
XSFILL59080x27050 gnd vdd FILL
XFILL_4__11461_ gnd vdd FILL
XFILL_2__7494_ gnd vdd FILL
XFILL_5__9011_ gnd vdd FILL
XFILL_1__11281_ gnd vdd FILL
XSFILL99480x32050 gnd vdd FILL
X_11137_ _11617_/A _11617_/B gnd _11137_/Y vdd NAND2X1
XFILL_5__12751_ gnd vdd FILL
XFILL_4__10412_ gnd vdd FILL
XSFILL74120x30050 gnd vdd FILL
XFILL_1__13020_ gnd vdd FILL
XFILL_4__14180_ gnd vdd FILL
XFILL_2__9233_ gnd vdd FILL
XFILL_3__13930_ gnd vdd FILL
XFILL_2__12571_ gnd vdd FILL
XFILL_1__10232_ gnd vdd FILL
XFILL_4__11392_ gnd vdd FILL
XFILL_0__13750_ gnd vdd FILL
XFILL_3_BUFX2_insert260 gnd vdd FILL
XFILL_0__10962_ gnd vdd FILL
XFILL_3_BUFX2_insert271 gnd vdd FILL
XFILL_5__11702_ gnd vdd FILL
XFILL_3_BUFX2_insert282 gnd vdd FILL
X_15945_ _7404_/Q _15631_/B _15945_/C gnd _15946_/C vdd NAND3X1
XFILL_4__13131_ gnd vdd FILL
X_11068_ _11096_/B _11067_/Y gnd _11389_/A vdd NOR2X1
XFILL_5__15470_ gnd vdd FILL
XFILL_2__14310_ gnd vdd FILL
XFILL_2__11522_ gnd vdd FILL
XFILL_3_BUFX2_insert293 gnd vdd FILL
XFILL_0__12701_ gnd vdd FILL
XFILL_3__13861_ gnd vdd FILL
XFILL_2__9164_ gnd vdd FILL
XFILL_2__15290_ gnd vdd FILL
XFILL_1__10163_ gnd vdd FILL
X_10019_ _10019_/A gnd _10019_/Y vdd INVX1
XFILL_0__13681_ gnd vdd FILL
XFILL_5__14421_ gnd vdd FILL
XSFILL63960x73050 gnd vdd FILL
XFILL_0__10893_ gnd vdd FILL
XFILL_5__11633_ gnd vdd FILL
XFILL_3__15600_ gnd vdd FILL
XSFILL13800x45050 gnd vdd FILL
XFILL_2__8115_ gnd vdd FILL
X_15876_ _15876_/A _15875_/Y gnd _15877_/B vdd NOR2X1
XFILL_2__14241_ gnd vdd FILL
XFILL_4__10274_ gnd vdd FILL
XFILL_2__9095_ gnd vdd FILL
XFILL_2__11453_ gnd vdd FILL
XFILL_0__15420_ gnd vdd FILL
XFILL_0__12632_ gnd vdd FILL
XFILL_3__13792_ gnd vdd FILL
XFILL_5__9913_ gnd vdd FILL
XFILL_2_BUFX2_insert960 gnd vdd FILL
XFILL_2_BUFX2_insert971 gnd vdd FILL
XFILL_1__14971_ gnd vdd FILL
X_14827_ _13843_/C _14826_/Y _14825_/Y _13617_/D gnd _14831_/A vdd OAI22X1
XFILL_4__12013_ gnd vdd FILL
XFILL_5__14352_ gnd vdd FILL
XFILL_2__10404_ gnd vdd FILL
XFILL_3__15531_ gnd vdd FILL
XFILL_2_BUFX2_insert982 gnd vdd FILL
XFILL_5__11564_ gnd vdd FILL
XFILL_2_BUFX2_insert993 gnd vdd FILL
XFILL_3__12743_ gnd vdd FILL
XFILL_2__14172_ gnd vdd FILL
XFILL_0__15351_ gnd vdd FILL
XFILL_1__13922_ gnd vdd FILL
XFILL_2__11384_ gnd vdd FILL
XFILL_5__13303_ gnd vdd FILL
XFILL_5__10515_ gnd vdd FILL
XFILL_0__7061_ gnd vdd FILL
XFILL_2__13123_ gnd vdd FILL
X_14758_ _9969_/Q gnd _16155_/C vdd INVX1
XFILL_5__14283_ gnd vdd FILL
XFILL_5__11495_ gnd vdd FILL
XFILL_3__15462_ gnd vdd FILL
XFILL_0__14302_ gnd vdd FILL
XFILL_1__13853_ gnd vdd FILL
XFILL_0__11514_ gnd vdd FILL
XFILL_5__16022_ gnd vdd FILL
XFILL_0__15282_ gnd vdd FILL
XFILL_5__13234_ gnd vdd FILL
XFILL_0__12494_ gnd vdd FILL
XFILL_5__9775_ gnd vdd FILL
X_13709_ _9051_/Q gnd _13711_/D vdd INVX1
XFILL_5__10446_ gnd vdd FILL
XFILL_5__6987_ gnd vdd FILL
XFILL_3__14413_ gnd vdd FILL
XFILL_3__7810_ gnd vdd FILL
XSFILL43880x40050 gnd vdd FILL
XFILL_3__11625_ gnd vdd FILL
X_14689_ _14868_/A _14689_/B _9199_/Q _14868_/D gnd _14690_/B vdd AOI22X1
XFILL_4__13964_ gnd vdd FILL
XFILL_3__15393_ gnd vdd FILL
XFILL_0__14233_ gnd vdd FILL
XFILL_2__10266_ gnd vdd FILL
XFILL_2__9997_ gnd vdd FILL
XFILL_1__13784_ gnd vdd FILL
XFILL_5__8726_ gnd vdd FILL
XFILL_0__11445_ gnd vdd FILL
X_16428_ _13980_/A _8161_/CLK _8033_/R vdd _16428_/D gnd vdd DFFSR
XFILL_1__10996_ gnd vdd FILL
XFILL_4__15703_ gnd vdd FILL
XFILL_5__13165_ gnd vdd FILL
XFILL_2__12005_ gnd vdd FILL
XFILL_4__12915_ gnd vdd FILL
XSFILL58920x62050 gnd vdd FILL
XFILL_5__10377_ gnd vdd FILL
XFILL_3__14344_ gnd vdd FILL
XFILL_3__7741_ gnd vdd FILL
XFILL_1__12735_ gnd vdd FILL
XFILL_1__15523_ gnd vdd FILL
XFILL_4__13895_ gnd vdd FILL
XFILL_3__11556_ gnd vdd FILL
XFILL_0__14164_ gnd vdd FILL
XFILL_2__10197_ gnd vdd FILL
XSFILL74200x10050 gnd vdd FILL
XBUFX2_insert970 _12417_/Y gnd _8511_/B vdd BUFX2
X_8310_ _8310_/A gnd _8312_/A vdd INVX1
XFILL_5__12116_ gnd vdd FILL
XFILL_5__8657_ gnd vdd FILL
XFILL_0__11376_ gnd vdd FILL
X_16359_ _16357_/Y gnd _16358_/Y gnd _16429_/D vdd OAI21X1
XFILL_4__15634_ gnd vdd FILL
XBUFX2_insert981 _13455_/Y gnd _14887_/B vdd BUFX2
XFILL_3__10507_ gnd vdd FILL
XBUFX2_insert992 _12408_/Y gnd _7222_/B vdd BUFX2
XFILL_4__12846_ gnd vdd FILL
X_9290_ _9290_/A gnd _9292_/A vdd INVX1
XFILL_5__13096_ gnd vdd FILL
XFILL_0__7963_ gnd vdd FILL
XFILL_0__13115_ gnd vdd FILL
XFILL_3__14275_ gnd vdd FILL
XFILL_5__7608_ gnd vdd FILL
XFILL_3__7672_ gnd vdd FILL
XFILL_3__11487_ gnd vdd FILL
XFILL_1__15454_ gnd vdd FILL
XFILL_2__8879_ gnd vdd FILL
XSFILL59000x71050 gnd vdd FILL
XFILL_0__14095_ gnd vdd FILL
XFILL_5__8588_ gnd vdd FILL
XFILL_3__16014_ gnd vdd FILL
XFILL_0__6914_ gnd vdd FILL
XFILL_5__12047_ gnd vdd FILL
X_8241_ _8241_/A _8216_/A _8241_/C gnd _8297_/D vdd OAI21X1
XFILL_3__13226_ gnd vdd FILL
XFILL_4__15565_ gnd vdd FILL
XFILL_3__9411_ gnd vdd FILL
XFILL_4__12777_ gnd vdd FILL
XFILL_3__10438_ gnd vdd FILL
XFILL_1__14405_ gnd vdd FILL
XFILL_1__11617_ gnd vdd FILL
XFILL_1__15385_ gnd vdd FILL
XFILL_0__13046_ gnd vdd FILL
XFILL_2__13956_ gnd vdd FILL
XFILL_1__12597_ gnd vdd FILL
XFILL_6__16125_ gnd vdd FILL
XFILL_0__10258_ gnd vdd FILL
XFILL_0__9633_ gnd vdd FILL
XFILL_4__14516_ gnd vdd FILL
XFILL_0__6845_ gnd vdd FILL
X_8172_ _8120_/A _9453_/CLK _9453_/R vdd _8172_/D gnd vdd DFFSR
XSFILL23240x50050 gnd vdd FILL
XFILL_4__11728_ gnd vdd FILL
XFILL_3__10369_ gnd vdd FILL
XFILL_3__13157_ gnd vdd FILL
XFILL_2__12907_ gnd vdd FILL
XFILL_1__14336_ gnd vdd FILL
XFILL_3__9342_ gnd vdd FILL
XFILL_4__15496_ gnd vdd FILL
XFILL_1__11548_ gnd vdd FILL
XFILL_2__13887_ gnd vdd FILL
XFILL_0__10189_ gnd vdd FILL
X_7123_ _7157_/Q gnd _7125_/A vdd INVX1
XFILL_5__15806_ gnd vdd FILL
XFILL_3__12108_ gnd vdd FILL
XFILL_4__14447_ gnd vdd FILL
XFILL_2__15626_ gnd vdd FILL
XFILL_4__11659_ gnd vdd FILL
XFILL_3__13088_ gnd vdd FILL
XFILL_3__9273_ gnd vdd FILL
XFILL_5__13998_ gnd vdd FILL
XFILL_2__12838_ gnd vdd FILL
XFILL_5__9209_ gnd vdd FILL
XFILL_1__14267_ gnd vdd FILL
XFILL_1__11479_ gnd vdd FILL
XFILL_0__14997_ gnd vdd FILL
XFILL_0__8515_ gnd vdd FILL
X_7054_ _7054_/A gnd _7054_/Y vdd INVX1
XFILL_5__15737_ gnd vdd FILL
XFILL_1__13218_ gnd vdd FILL
XFILL_1__16006_ gnd vdd FILL
XFILL_0__9495_ gnd vdd FILL
XFILL_3__8224_ gnd vdd FILL
XFILL_3__12039_ gnd vdd FILL
XFILL_4__14378_ gnd vdd FILL
XFILL_2__15557_ gnd vdd FILL
XFILL_1__14198_ gnd vdd FILL
XFILL_2__12769_ gnd vdd FILL
XFILL_0__13948_ gnd vdd FILL
XSFILL43960x20050 gnd vdd FILL
XFILL_4__16117_ gnd vdd FILL
XFILL_4__13329_ gnd vdd FILL
XSFILL39320x3050 gnd vdd FILL
XFILL_0__8446_ gnd vdd FILL
XFILL_5__15668_ gnd vdd FILL
XFILL_2__14508_ gnd vdd FILL
XFILL_1__13149_ gnd vdd FILL
XFILL_2__15488_ gnd vdd FILL
XFILL_0__13879_ gnd vdd FILL
XFILL_0__8377_ gnd vdd FILL
XFILL_5__14619_ gnd vdd FILL
XFILL_1__7170_ gnd vdd FILL
XFILL_4__16048_ gnd vdd FILL
XFILL_3__7106_ gnd vdd FILL
XFILL_5__15599_ gnd vdd FILL
XFILL_2__14439_ gnd vdd FILL
XFILL_0__15618_ gnd vdd FILL
XFILL_3__8086_ gnd vdd FILL
XFILL_0__7328_ gnd vdd FILL
XFILL_3__15729_ gnd vdd FILL
X_7956_ _7956_/A gnd _7958_/A vdd INVX1
XSFILL8680x79050 gnd vdd FILL
XFILL_3__7037_ gnd vdd FILL
XFILL_0__15549_ gnd vdd FILL
XSFILL23720x28050 gnd vdd FILL
X_6907_ _6905_/Y _6955_/B _6907_/C gnd _6999_/D vdd OAI21X1
XSFILL33880x72050 gnd vdd FILL
XFILL_2__16109_ gnd vdd FILL
X_7887_ _7887_/A _7887_/B _7887_/C gnd _7923_/D vdd OAI21X1
XFILL_4__7850_ gnd vdd FILL
X_6838_ _6838_/A gnd memoryAddress[0] vdd BUFX2
X_9626_ _9698_/Q gnd _9628_/A vdd INVX1
XSFILL64200x42050 gnd vdd FILL
XFILL_3__8988_ gnd vdd FILL
XFILL_5_BUFX2_insert300 gnd vdd FILL
XFILL_1__9811_ gnd vdd FILL
XFILL_1_CLKBUF1_insert1079 gnd vdd FILL
X_9557_ _9555_/Y _9466_/A _9557_/C gnd _9589_/D vdd OAI21X1
XFILL_6__8697_ gnd vdd FILL
XFILL_5_BUFX2_insert311 gnd vdd FILL
XFILL_4__9520_ gnd vdd FILL
XFILL_5_BUFX2_insert322 gnd vdd FILL
XFILL_3__7939_ gnd vdd FILL
XBUFX2_insert12 _13280_/Y gnd _7323_/A vdd BUFX2
XFILL_5_BUFX2_insert333 gnd vdd FILL
X_8508_ _8508_/A _8636_/B gnd _8509_/C vdd NAND2X1
XFILL_5_BUFX2_insert344 gnd vdd FILL
XBUFX2_insert23 _11344_/Y gnd _11415_/C vdd BUFX2
XFILL_1__9742_ gnd vdd FILL
XBUFX2_insert34 _13265_/Y gnd _6967_/B vdd BUFX2
XFILL_5_BUFX2_insert355 gnd vdd FILL
X_9488_ _9488_/A _9548_/B _9488_/C gnd _9566_/D vdd OAI21X1
XBUFX2_insert45 _14986_/Y gnd _16309_/A vdd BUFX2
XFILL_1__6954_ gnd vdd FILL
XBUFX2_insert56 _13309_/Y gnd _8098_/B vdd BUFX2
XFILL_5_BUFX2_insert366 gnd vdd FILL
XFILL_5_BUFX2_insert377 gnd vdd FILL
XFILL_5_BUFX2_insert388 gnd vdd FILL
X_10370_ _15234_/A gnd _10372_/A vdd INVX1
XBUFX2_insert67 _12215_/Y gnd _12237_/B vdd BUFX2
XBUFX2_insert78 _15015_/Y gnd _16000_/A vdd BUFX2
X_8439_ _8183_/A _8440_/B gnd _8439_/Y vdd NAND2X1
XFILL_5_BUFX2_insert399 gnd vdd FILL
XFILL_3__9609_ gnd vdd FILL
XBUFX2_insert89 _12357_/Y gnd _7555_/B vdd BUFX2
XFILL_1__9673_ gnd vdd FILL
XFILL_4__8402_ gnd vdd FILL
XFILL_1__6885_ gnd vdd FILL
XFILL_4__9382_ gnd vdd FILL
XFILL_1__8624_ gnd vdd FILL
XFILL_4__8333_ gnd vdd FILL
XSFILL65000x4050 gnd vdd FILL
X_12040_ _12028_/A _12802_/Q _12024_/C gnd _12042_/B vdd NAND3X1
XSFILL8760x59050 gnd vdd FILL
XFILL_4__8264_ gnd vdd FILL
XSFILL33960x52050 gnd vdd FILL
XFILL_1__7506_ gnd vdd FILL
XFILL_1__8486_ gnd vdd FILL
XFILL_4__7215_ gnd vdd FILL
XSFILL49240x19050 gnd vdd FILL
XFILL_4__8195_ gnd vdd FILL
XFILL_1__7437_ gnd vdd FILL
X_13991_ _8855_/A gnd _13991_/Y vdd INVX1
X_15730_ _15725_/Y _15730_/B gnd _15731_/C vdd NAND2X1
XSFILL108760x66050 gnd vdd FILL
X_12942_ _12942_/Q _12669_/CLK _9050_/R vdd _12894_/Y gnd vdd DFFSR
XFILL_2_BUFX2_insert234 gnd vdd FILL
XFILL_2_BUFX2_insert245 gnd vdd FILL
XFILL_1__7368_ gnd vdd FILL
XFILL_2_BUFX2_insert256 gnd vdd FILL
XFILL_4__7077_ gnd vdd FILL
XFILL_2_BUFX2_insert267 gnd vdd FILL
X_15661_ _6947_/A _15382_/B _16096_/C _7397_/Q gnd _15667_/A vdd AOI22X1
XFILL_2_BUFX2_insert278 gnd vdd FILL
XFILL_1__9107_ gnd vdd FILL
X_12873_ _12871_/Y vdd _12873_/C gnd _12935_/D vdd OAI21X1
XFILL_2_BUFX2_insert289 gnd vdd FILL
XFILL_1__7299_ gnd vdd FILL
XFILL_1_BUFX2_insert901 gnd vdd FILL
XSFILL110120x82050 gnd vdd FILL
XFILL_1_BUFX2_insert912 gnd vdd FILL
XFILL_5__6910_ gnd vdd FILL
X_14612_ _14583_/B _14611_/Y _14174_/C _14610_/Y gnd _14616_/A vdd OAI22X1
XFILL_1_BUFX2_insert923 gnd vdd FILL
XSFILL94360x2050 gnd vdd FILL
XFILL_5__7890_ gnd vdd FILL
X_11824_ _11764_/A _11234_/Y _11376_/B _11764_/D gnd _11828_/A vdd AOI22X1
XFILL_1__9038_ gnd vdd FILL
XFILL_2__9920_ gnd vdd FILL
X_15592_ _16301_/A _15590_/Y _15591_/Y _15761_/D gnd _15593_/B vdd OAI22X1
XFILL_1_BUFX2_insert934 gnd vdd FILL
XFILL_1_BUFX2_insert945 gnd vdd FILL
XFILL_1_BUFX2_insert956 gnd vdd FILL
XFILL_5__10300_ gnd vdd FILL
XFILL_1_BUFX2_insert967 gnd vdd FILL
XFILL_5__6841_ gnd vdd FILL
XFILL_1_BUFX2_insert978 gnd vdd FILL
X_14543_ _9400_/A gnd _14543_/Y vdd INVX1
XFILL_2__10120_ gnd vdd FILL
XFILL_5__11280_ gnd vdd FILL
X_11755_ _11379_/B _11377_/Y gnd _11801_/B vdd NOR2X1
XFILL_1_BUFX2_insert989 gnd vdd FILL
XFILL_2__9851_ gnd vdd FILL
XFILL_5__10231_ gnd vdd FILL
XBUFX2_insert233 _11228_/Y gnd _11423_/B vdd BUFX2
X_10706_ _10706_/A _10676_/B _10705_/Y gnd _10740_/D vdd OAI21X1
XFILL_4__7979_ gnd vdd FILL
X_14474_ _7403_/Q gnd _14474_/Y vdd INVX1
XFILL_3__11410_ gnd vdd FILL
XFILL_4__10961_ gnd vdd FILL
XFILL_3__12390_ gnd vdd FILL
XBUFX2_insert244 _13460_/Y gnd _14237_/B vdd BUFX2
XFILL_2__10051_ gnd vdd FILL
X_11686_ _11686_/A _11684_/Y gnd _11686_/Y vdd NOR2X1
XFILL_2__9782_ gnd vdd FILL
XFILL_5__8511_ gnd vdd FILL
XFILL_4__9718_ gnd vdd FILL
XBUFX2_insert255 _12423_/Y gnd _9413_/B vdd BUFX2
XFILL_0__11230_ gnd vdd FILL
X_16213_ _14852_/Y _16213_/B _15924_/B _14863_/Y gnd _16218_/A vdd OAI22X1
XFILL_1__10781_ gnd vdd FILL
XBUFX2_insert266 _15024_/Y gnd _16137_/C vdd BUFX2
XFILL_2__6994_ gnd vdd FILL
XFILL_4__12700_ gnd vdd FILL
X_13425_ _13421_/Y _13775_/B _13857_/B _13422_/Y gnd _13426_/B vdd OAI22X1
XBUFX2_insert277 _13419_/Y gnd _13420_/C vdd BUFX2
XSFILL99480x27050 gnd vdd FILL
XFILL_5__9491_ gnd vdd FILL
X_10637_ _10635_/Y _10678_/A _10637_/C gnd _10717_/D vdd OAI21X1
XFILL_5_CLKBUF1_insert112 gnd vdd FILL
XBUFX2_insert288 _15059_/Y gnd _15565_/B vdd BUFX2
XFILL_5__10162_ gnd vdd FILL
XFILL_4__13680_ gnd vdd FILL
XFILL_1__12520_ gnd vdd FILL
XFILL_5_CLKBUF1_insert123 gnd vdd FILL
XFILL_2__8733_ gnd vdd FILL
XFILL_3__11341_ gnd vdd FILL
XBUFX2_insert299 _12414_/Y gnd _8764_/B vdd BUFX2
XFILL_4__10892_ gnd vdd FILL
XFILL_4__9649_ gnd vdd FILL
XFILL_0__11161_ gnd vdd FILL
XFILL_5__8442_ gnd vdd FILL
XFILL_5_CLKBUF1_insert134 gnd vdd FILL
XFILL_5_CLKBUF1_insert145 gnd vdd FILL
X_16144_ _10481_/Q gnd _16144_/Y vdd INVX1
XFILL_4__12631_ gnd vdd FILL
XFILL_5_CLKBUF1_insert156 gnd vdd FILL
X_13356_ _13355_/Y _13356_/B gnd _13356_/Y vdd NOR2X1
X_10568_ _10581_/B _7752_/B gnd _10569_/C vdd NAND2X1
XFILL_2__13810_ gnd vdd FILL
XFILL_3__14060_ gnd vdd FILL
XFILL_5__14970_ gnd vdd FILL
XFILL_5_CLKBUF1_insert167 gnd vdd FILL
XFILL_3__11272_ gnd vdd FILL
XFILL_0__10112_ gnd vdd FILL
XFILL_5_CLKBUF1_insert178 gnd vdd FILL
XFILL_1__12451_ gnd vdd FILL
XFILL_6__10403_ gnd vdd FILL
XFILL_2__14790_ gnd vdd FILL
XFILL_5__8373_ gnd vdd FILL
X_12307_ _12227_/A gnd _12307_/C gnd _12307_/Y vdd NAND3X1
XFILL_5_CLKBUF1_insert189 gnd vdd FILL
XFILL_0__11092_ gnd vdd FILL
XFILL_4__15350_ gnd vdd FILL
X_16075_ _16075_/A _16075_/B _16070_/Y gnd _16086_/A vdd NAND3X1
XFILL_5__13921_ gnd vdd FILL
XFILL_3__13011_ gnd vdd FILL
X_13287_ _13297_/C _13287_/B gnd _13287_/Y vdd NOR2X1
XFILL_2__7615_ gnd vdd FILL
X_10499_ _10500_/B _7555_/B gnd _10499_/Y vdd NAND2X1
XSFILL99240x50 gnd vdd FILL
XFILL_1__11402_ gnd vdd FILL
XFILL_1__15170_ gnd vdd FILL
XFILL_2__13741_ gnd vdd FILL
XFILL_2__10953_ gnd vdd FILL
XFILL_0__10043_ gnd vdd FILL
XFILL_5__7324_ gnd vdd FILL
XFILL_1__12382_ gnd vdd FILL
XFILL_2__8595_ gnd vdd FILL
XFILL_0__14920_ gnd vdd FILL
X_15026_ _15025_/Y _15026_/B gnd _15027_/C vdd NOR2X1
XFILL_4__14301_ gnd vdd FILL
XSFILL8760x3050 gnd vdd FILL
X_12238_ _12238_/A _12238_/B _12237_/Y gnd _12238_/Y vdd NAND3X1
XSFILL54120x5050 gnd vdd FILL
XFILL_4__11513_ gnd vdd FILL
XFILL_5__13852_ gnd vdd FILL
XFILL_3__10154_ gnd vdd FILL
XFILL_1__14121_ gnd vdd FILL
XFILL_4__15281_ gnd vdd FILL
XFILL112280x51050 gnd vdd FILL
XFILL_4__12493_ gnd vdd FILL
XFILL_2__7546_ gnd vdd FILL
XFILL_1__11333_ gnd vdd FILL
XSFILL64040x77050 gnd vdd FILL
XFILL_0__14851_ gnd vdd FILL
XFILL_2__13672_ gnd vdd FILL
XFILL_2__10884_ gnd vdd FILL
XFILL_4__14232_ gnd vdd FILL
X_12169_ _13133_/A gnd _12171_/A vdd INVX1
XFILL_2__15411_ gnd vdd FILL
XFILL_5__13783_ gnd vdd FILL
XFILL_4__11444_ gnd vdd FILL
XFILL_2__12623_ gnd vdd FILL
XFILL_0__13802_ gnd vdd FILL
XFILL_1__14052_ gnd vdd FILL
XFILL_3__14962_ gnd vdd FILL
XFILL_5__10995_ gnd vdd FILL
XFILL_2__7477_ gnd vdd FILL
XFILL_6__12004_ gnd vdd FILL
XFILL_2__16391_ gnd vdd FILL
XFILL_1__11264_ gnd vdd FILL
XFILL_0__14782_ gnd vdd FILL
XFILL_0__9280_ gnd vdd FILL
XFILL_5__12734_ gnd vdd FILL
XFILL_5__15522_ gnd vdd FILL
XFILL_0__11994_ gnd vdd FILL
XFILL_5__7186_ gnd vdd FILL
XFILL_2__9216_ gnd vdd FILL
XFILL_4__14163_ gnd vdd FILL
XFILL_6__10196_ gnd vdd FILL
XFILL_1__13003_ gnd vdd FILL
XFILL_3__13913_ gnd vdd FILL
XFILL_2__15342_ gnd vdd FILL
XSFILL43880x35050 gnd vdd FILL
XFILL_4__11375_ gnd vdd FILL
XFILL_0__13733_ gnd vdd FILL
XFILL_3__14893_ gnd vdd FILL
XFILL_0__10945_ gnd vdd FILL
XFILL_0__8231_ gnd vdd FILL
XFILL_1__11195_ gnd vdd FILL
X_15928_ _15928_/A _15928_/B gnd _15929_/A vdd NOR2X1
XFILL_4__13114_ gnd vdd FILL
XFILL_5__15453_ gnd vdd FILL
XFILL_3__13844_ gnd vdd FILL
XFILL_2__9147_ gnd vdd FILL
XFILL_2__11505_ gnd vdd FILL
XFILL_4__14094_ gnd vdd FILL
XFILL_2__12485_ gnd vdd FILL
XFILL_1__10146_ gnd vdd FILL
XSFILL18680x11050 gnd vdd FILL
XFILL_2__15273_ gnd vdd FILL
XFILL_0__13664_ gnd vdd FILL
XFILL_6__6950_ gnd vdd FILL
X_7810_ _7810_/A gnd _7812_/A vdd INVX1
XFILL_0__10876_ gnd vdd FILL
XFILL_5__11616_ gnd vdd FILL
XFILL_5__14404_ gnd vdd FILL
XFILL_5__15384_ gnd vdd FILL
XFILL_4__13045_ gnd vdd FILL
XFILL_6__13955_ gnd vdd FILL
X_15859_ _8626_/A _16212_/A gnd _15860_/B vdd NAND2X1
XFILL_0__15403_ gnd vdd FILL
XFILL_5__12596_ gnd vdd FILL
XFILL_2__14224_ gnd vdd FILL
X_8790_ _8790_/Q _6998_/CLK _7644_/R vdd _8696_/Y gnd vdd DFFSR
XFILL_4__10257_ gnd vdd FILL
XFILL_2__11436_ gnd vdd FILL
XFILL_0__12615_ gnd vdd FILL
XFILL_3__13775_ gnd vdd FILL
XFILL_2__9078_ gnd vdd FILL
XFILL_2_BUFX2_insert790 gnd vdd FILL
XFILL_0__16383_ gnd vdd FILL
XFILL_0__7113_ gnd vdd FILL
XFILL_1__14954_ gnd vdd FILL
XFILL_0__13595_ gnd vdd FILL
XFILL_5__14335_ gnd vdd FILL
X_7741_ _7741_/A _7759_/B _7741_/C gnd _7789_/D vdd OAI21X1
XSFILL59000x66050 gnd vdd FILL
XFILL_3__15514_ gnd vdd FILL
XFILL_5__11547_ gnd vdd FILL
XFILL_0__8093_ gnd vdd FILL
XFILL_3__8911_ gnd vdd FILL
XFILL_3__12726_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1074 gnd vdd FILL
XSFILL99400x71050 gnd vdd FILL
XFILL_4__10188_ gnd vdd FILL
XFILL_0__15334_ gnd vdd FILL
XFILL_2__14155_ gnd vdd FILL
XFILL_1__13905_ gnd vdd FILL
XFILL_2__11367_ gnd vdd FILL
XFILL_3__9891_ gnd vdd FILL
XFILL_0__7044_ gnd vdd FILL
XFILL_1__14885_ gnd vdd FILL
XFILL_5__14266_ gnd vdd FILL
XFILL_2__10318_ gnd vdd FILL
XFILL111720x65050 gnd vdd FILL
X_7672_ _7670_/Y _7672_/B _7672_/C gnd _7766_/D vdd OAI21X1
XFILL_2__13106_ gnd vdd FILL
XFILL_5__11478_ gnd vdd FILL
XFILL_3__15445_ gnd vdd FILL
XFILL_3__8842_ gnd vdd FILL
XFILL_3__12657_ gnd vdd FILL
XFILL_4__14996_ gnd vdd FILL
XFILL_2__14086_ gnd vdd FILL
XFILL_1__13836_ gnd vdd FILL
XFILL_2__11298_ gnd vdd FILL
XFILL_0__15265_ gnd vdd FILL
XFILL_5__13217_ gnd vdd FILL
XFILL_5__16005_ gnd vdd FILL
XFILL_0__12477_ gnd vdd FILL
XSFILL109000x35050 gnd vdd FILL
XFILL_5__9758_ gnd vdd FILL
X_9411_ _9411_/A _9425_/A _9411_/C gnd _9411_/Y vdd OAI21X1
XFILL_5__10429_ gnd vdd FILL
XFILL112360x31050 gnd vdd FILL
XFILL_6__12768_ gnd vdd FILL
XFILL_5__14197_ gnd vdd FILL
XSFILL64120x57050 gnd vdd FILL
XFILL_2__13037_ gnd vdd FILL
XFILL_3__11608_ gnd vdd FILL
XFILL_4__13947_ gnd vdd FILL
XFILL_2__10249_ gnd vdd FILL
XFILL_3__15376_ gnd vdd FILL
XFILL_0__14216_ gnd vdd FILL
XFILL_3__12588_ gnd vdd FILL
XFILL_6__7502_ gnd vdd FILL
XFILL_3__8773_ gnd vdd FILL
XFILL_5__8709_ gnd vdd FILL
XFILL_0__11428_ gnd vdd FILL
XFILL_1__10979_ gnd vdd FILL
XFILL_0__15196_ gnd vdd FILL
XFILL_1__13767_ gnd vdd FILL
XFILL_5__13148_ gnd vdd FILL
X_9342_ _9342_/A _9339_/B _9341_/Y gnd _9432_/D vdd OAI21X1
XFILL_3__14327_ gnd vdd FILL
XFILL_4__13878_ gnd vdd FILL
XFILL_0__8995_ gnd vdd FILL
XFILL_1__15506_ gnd vdd FILL
XFILL_3__7724_ gnd vdd FILL
XFILL_3__11539_ gnd vdd FILL
XFILL_1__12718_ gnd vdd FILL
XFILL_0__14147_ gnd vdd FILL
XFILL_1__13698_ gnd vdd FILL
XFILL_0__11359_ gnd vdd FILL
XSFILL43960x15050 gnd vdd FILL
XFILL_0__7946_ gnd vdd FILL
XSFILL3560x64050 gnd vdd FILL
XFILL_5__13079_ gnd vdd FILL
XFILL_4__15617_ gnd vdd FILL
X_9273_ _9301_/B _8889_/B gnd _9274_/C vdd NAND2X1
XFILL_4_BUFX2_insert307 gnd vdd FILL
XFILL_4__12829_ gnd vdd FILL
XFILL_3__14258_ gnd vdd FILL
XFILL_1__12649_ gnd vdd FILL
XFILL_4_BUFX2_insert318 gnd vdd FILL
XFILL_1__15437_ gnd vdd FILL
XFILL_2__14988_ gnd vdd FILL
XFILL_0__14078_ gnd vdd FILL
XFILL_4_BUFX2_insert329 gnd vdd FILL
X_8224_ _8292_/Q gnd _8224_/Y vdd INVX1
XFILL_3__13209_ gnd vdd FILL
XSFILL28760x76050 gnd vdd FILL
XFILL_4__15548_ gnd vdd FILL
XFILL_0__7877_ gnd vdd FILL
XFILL_3__14189_ gnd vdd FILL
XFILL_0__13029_ gnd vdd FILL
XFILL_2__13939_ gnd vdd FILL
XSFILL44040x24050 gnd vdd FILL
XFILL_1__15368_ gnd vdd FILL
XFILL_3__7586_ gnd vdd FILL
XFILL_0__9616_ gnd vdd FILL
X_8155_ _8069_/A _8663_/CLK _9944_/R vdd _8155_/D gnd vdd DFFSR
XFILL_4__15479_ gnd vdd FILL
XFILL_1__14319_ gnd vdd FILL
XFILL_1__15299_ gnd vdd FILL
X_7106_ _7061_/A _8642_/B gnd _7107_/C vdd NAND2X1
XFILL_0__9547_ gnd vdd FILL
XFILL_1__8340_ gnd vdd FILL
X_8086_ _8084_/Y _8082_/A _8086_/C gnd _8160_/D vdd OAI21X1
XFILL_2__15609_ gnd vdd FILL
XFILL_3__9256_ gnd vdd FILL
XFILL_1__8271_ gnd vdd FILL
X_7037_ _7061_/A _7037_/B gnd _7037_/Y vdd NAND2X1
XFILL_3__8207_ gnd vdd FILL
XFILL_0__9478_ gnd vdd FILL
XFILL112440x11050 gnd vdd FILL
XSFILL64200x37050 gnd vdd FILL
XFILL_1__7222_ gnd vdd FILL
XSFILL38920x5050 gnd vdd FILL
XFILL_3__8138_ gnd vdd FILL
XFILL_4__8951_ gnd vdd FILL
X_8988_ _8988_/A _8996_/A _8988_/C gnd _9058_/D vdd OAI21X1
XFILL_3__8069_ gnd vdd FILL
XFILL_1__7084_ gnd vdd FILL
X_7939_ _7970_/B _8195_/B gnd _7940_/C vdd NAND2X1
XFILL_4__8882_ gnd vdd FILL
XSFILL94280x32050 gnd vdd FILL
XFILL_0_BUFX2_insert908 gnd vdd FILL
XFILL_4__7833_ gnd vdd FILL
XFILL_0_BUFX2_insert919 gnd vdd FILL
X_11540_ _11660_/A _11535_/Y _11539_/Y gnd _11540_/Y vdd NAND3X1
X_9609_ _9615_/A _7177_/B gnd _9610_/C vdd NAND2X1
XFILL_4__7764_ gnd vdd FILL
X_11471_ _11490_/A _11433_/Y _11324_/Y gnd _11471_/Y vdd AOI21X1
XFILL_4__9503_ gnd vdd FILL
XFILL_1__7986_ gnd vdd FILL
X_10422_ _10423_/B _7990_/B gnd _10422_/Y vdd NAND2X1
X_13210_ _13246_/A _13215_/A gnd _13239_/B vdd NAND2X1
XFILL_4__7695_ gnd vdd FILL
X_14190_ _8933_/Q gnd _14190_/Y vdd INVX1
XFILL_1__9725_ gnd vdd FILL
XFILL_1__6937_ gnd vdd FILL
X_13141_ _13139_/Y _13134_/A _13141_/C gnd _13195_/D vdd OAI21X1
X_10353_ _10311_/A _7786_/CLK _8053_/R vdd _10353_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert830 gnd vdd FILL
XSFILL48600x71050 gnd vdd FILL
XFILL_1__9656_ gnd vdd FILL
XFILL_4_BUFX2_insert841 gnd vdd FILL
XFILL_4_BUFX2_insert852 gnd vdd FILL
XFILL_1__6868_ gnd vdd FILL
XSFILL89240x21050 gnd vdd FILL
XFILL_4__9365_ gnd vdd FILL
XFILL_4_BUFX2_insert863 gnd vdd FILL
X_13072_ _6895_/A _8815_/CLK _9056_/R vdd _13072_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert874 gnd vdd FILL
X_10284_ _10284_/A gnd _10284_/Y vdd INVX1
XFILL_1__8607_ gnd vdd FILL
XFILL_4_BUFX2_insert885 gnd vdd FILL
XFILL_2__8380_ gnd vdd FILL
XFILL_4_BUFX2_insert896 gnd vdd FILL
XFILL_4__8316_ gnd vdd FILL
X_12023_ _12031_/A _12023_/B _12031_/C gnd _12026_/A vdd NAND3X1
XFILL_4__9296_ gnd vdd FILL
XFILL_2__7331_ gnd vdd FILL
XSFILL28920x36050 gnd vdd FILL
XFILL_5__7040_ gnd vdd FILL
XFILL_4__8247_ gnd vdd FILL
XSFILL94360x12050 gnd vdd FILL
XSFILL68520x22050 gnd vdd FILL
XFILL_5__10780_ gnd vdd FILL
XSFILL69000x29050 gnd vdd FILL
XFILL_1__8469_ gnd vdd FILL
XSFILL79160x73050 gnd vdd FILL
XFILL_2__9001_ gnd vdd FILL
XFILL_3__10910_ gnd vdd FILL
XFILL_1__10000_ gnd vdd FILL
XFILL_4__11160_ gnd vdd FILL
X_13974_ _13974_/A _13974_/B gnd _13975_/A vdd NOR2X1
XFILL_2__7193_ gnd vdd FILL
XFILL_3__11890_ gnd vdd FILL
X_15713_ _14218_/Y _15924_/B _16000_/A _15713_/D gnd _15713_/Y vdd OAI22X1
XFILL_4__10111_ gnd vdd FILL
XFILL_5__12450_ gnd vdd FILL
X_12925_ _12841_/A _8161_/CLK _7140_/R vdd _12925_/D gnd vdd DFFSR
XFILL_5__8991_ gnd vdd FILL
XFILL_2__12270_ gnd vdd FILL
XFILL_4__11091_ gnd vdd FILL
XFILL_0__10661_ gnd vdd FILL
XSFILL18040x69050 gnd vdd FILL
XFILL_5__11401_ gnd vdd FILL
XFILL_5__7942_ gnd vdd FILL
XSFILL84280x64050 gnd vdd FILL
X_15644_ _15369_/A _14164_/B _15644_/C _15644_/D gnd _15645_/A vdd OAI22X1
XFILL_5__12381_ gnd vdd FILL
X_12856_ _12856_/A gnd _12856_/Y vdd INVX1
XFILL_4__10042_ gnd vdd FILL
XFILL_1_BUFX2_insert720 gnd vdd FILL
XFILL_2__11221_ gnd vdd FILL
XSFILL58440x74050 gnd vdd FILL
XFILL_1_BUFX2_insert731 gnd vdd FILL
XFILL_0__12400_ gnd vdd FILL
XFILL_3__13560_ gnd vdd FILL
XFILL_1__11951_ gnd vdd FILL
XFILL_1_BUFX2_insert742 gnd vdd FILL
XFILL_3__10772_ gnd vdd FILL
XFILL_0__13380_ gnd vdd FILL
XFILL_5__14120_ gnd vdd FILL
XFILL_1_BUFX2_insert753 gnd vdd FILL
XFILL_5__7873_ gnd vdd FILL
X_11807_ _11249_/Y _11768_/B _11806_/Y gnd _11808_/B vdd OAI21X1
XFILL_5__11332_ gnd vdd FILL
XFILL_1_BUFX2_insert764 gnd vdd FILL
XFILL_4__14850_ gnd vdd FILL
XFILL_3__12511_ gnd vdd FILL
XSFILL59080x40050 gnd vdd FILL
XFILL_2__9903_ gnd vdd FILL
X_15575_ _14078_/A _15175_/B _15087_/B _7581_/A gnd _15580_/B vdd AOI22X1
X_12787_ _12785_/Y _12789_/A _12787_/C gnd _12821_/D vdd OAI21X1
XFILL_1__10902_ gnd vdd FILL
XFILL_2__11152_ gnd vdd FILL
XFILL_1_BUFX2_insert775 gnd vdd FILL
XFILL_5__9612_ gnd vdd FILL
XFILL_1_BUFX2_insert786 gnd vdd FILL
XFILL_0__12331_ gnd vdd FILL
XFILL_3__13491_ gnd vdd FILL
XFILL_1__11882_ gnd vdd FILL
XFILL_1__14670_ gnd vdd FILL
XFILL_1_BUFX2_insert797 gnd vdd FILL
XFILL_4__13801_ gnd vdd FILL
X_14526_ _14526_/A _14525_/Y _14526_/C gnd _14527_/B vdd NAND3X1
XFILL_5__14051_ gnd vdd FILL
XFILL_3__15230_ gnd vdd FILL
XFILL_5__11263_ gnd vdd FILL
XFILL_2__10103_ gnd vdd FILL
X_11738_ _11731_/B _11079_/Y _11743_/A gnd _11739_/A vdd OAI21X1
XFILL_3__12442_ gnd vdd FILL
XFILL_4__14781_ gnd vdd FILL
XFILL_1__13621_ gnd vdd FILL
XFILL112280x46050 gnd vdd FILL
XFILL_0__15050_ gnd vdd FILL
XFILL_2__15960_ gnd vdd FILL
XFILL_4__11993_ gnd vdd FILL
XFILL_4_BUFX2_insert13 gnd vdd FILL
XFILL_2__11083_ gnd vdd FILL
XFILL_1__10833_ gnd vdd FILL
XFILL_5__9543_ gnd vdd FILL
XFILL_0__12262_ gnd vdd FILL
XFILL_4_BUFX2_insert24 gnd vdd FILL
XFILL_5__13002_ gnd vdd FILL
XFILL_4_BUFX2_insert35 gnd vdd FILL
X_14457_ _14453_/Y _14457_/B gnd _14460_/C vdd NOR2X1
XFILL_4__13732_ gnd vdd FILL
XFILL_4__10944_ gnd vdd FILL
XFILL_4_BUFX2_insert46 gnd vdd FILL
XFILL_0__14001_ gnd vdd FILL
X_11669_ _11060_/Y _11682_/B _11668_/Y gnd _11669_/Y vdd OAI21X1
XFILL_2__10034_ gnd vdd FILL
XFILL_3__15161_ gnd vdd FILL
XFILL_5__11194_ gnd vdd FILL
XFILL_2__14911_ gnd vdd FILL
XFILL_1__16340_ gnd vdd FILL
XFILL_4_BUFX2_insert57 gnd vdd FILL
XFILL_2__9765_ gnd vdd FILL
XFILL_3__12373_ gnd vdd FILL
XFILL_1__13552_ gnd vdd FILL
XFILL_0__11213_ gnd vdd FILL
XFILL_1__10764_ gnd vdd FILL
XFILL_4_BUFX2_insert68 gnd vdd FILL
XFILL_2__6977_ gnd vdd FILL
XFILL_2__15891_ gnd vdd FILL
XFILL_5__9474_ gnd vdd FILL
XFILL_4_BUFX2_insert79 gnd vdd FILL
X_13408_ _13407_/Y _13718_/A gnd _13876_/C vdd NAND2X1
XFILL_0__7800_ gnd vdd FILL
XFILL_0__12193_ gnd vdd FILL
XFILL_4__16451_ gnd vdd FILL
XFILL_6__12484_ gnd vdd FILL
XFILL_5__10145_ gnd vdd FILL
XFILL_3__14112_ gnd vdd FILL
XFILL_2__8716_ gnd vdd FILL
XFILL_1__12503_ gnd vdd FILL
XFILL_4__13663_ gnd vdd FILL
XFILL_0__8780_ gnd vdd FILL
X_14388_ _9193_/Q _14868_/D _13645_/C _9961_/Q gnd _14390_/A vdd AOI22X1
XFILL_3__11324_ gnd vdd FILL
XFILL_2__14842_ gnd vdd FILL
XSFILL79240x53050 gnd vdd FILL
XFILL_4__10875_ gnd vdd FILL
XFILL_3__15092_ gnd vdd FILL
XFILL_0__11144_ gnd vdd FILL
XFILL_1__13483_ gnd vdd FILL
XFILL_1__16271_ gnd vdd FILL
XFILL_4__15402_ gnd vdd FILL
XFILL_1__10695_ gnd vdd FILL
X_16127_ _16106_/A _16127_/B _15726_/A _16127_/D gnd _16127_/Y vdd OAI22X1
X_13339_ _13289_/B _13295_/A gnd _13339_/Y vdd NAND2X1
XFILL_4__12614_ gnd vdd FILL
XFILL_0__7731_ gnd vdd FILL
XFILL_4__16382_ gnd vdd FILL
XFILL_3__14043_ gnd vdd FILL
XFILL_5__14953_ gnd vdd FILL
XFILL_1__12434_ gnd vdd FILL
XFILL_3__7440_ gnd vdd FILL
XFILL_4__13594_ gnd vdd FILL
XFILL_1__15222_ gnd vdd FILL
XFILL_2__8647_ gnd vdd FILL
XFILL_3__11255_ gnd vdd FILL
XFILL_2__14773_ gnd vdd FILL
XFILL_5__8356_ gnd vdd FILL
XSFILL114440x62050 gnd vdd FILL
XFILL_2__11985_ gnd vdd FILL
XFILL_0__15952_ gnd vdd FILL
XSFILL43480x32050 gnd vdd FILL
XFILL_0__11075_ gnd vdd FILL
XFILL_4__15333_ gnd vdd FILL
XFILL_5__13904_ gnd vdd FILL
X_16058_ _16056_/Y _16058_/B gnd _16058_/Y vdd NOR2X1
XFILL_2_BUFX2_insert1007 gnd vdd FILL
XFILL_1__15153_ gnd vdd FILL
XFILL_3__11186_ gnd vdd FILL
XFILL_2__13724_ gnd vdd FILL
XFILL_5__14884_ gnd vdd FILL
XFILL_1__12365_ gnd vdd FILL
XFILL_2__10936_ gnd vdd FILL
XFILL_3__7371_ gnd vdd FILL
XFILL_5__7307_ gnd vdd FILL
XFILL_2__8578_ gnd vdd FILL
XFILL_2_BUFX2_insert1018 gnd vdd FILL
XSFILL84360x44050 gnd vdd FILL
XSFILL13560x2050 gnd vdd FILL
XFILL_0__14903_ gnd vdd FILL
XFILL_0__10026_ gnd vdd FILL
XFILL_2_BUFX2_insert1029 gnd vdd FILL
XFILL_6__13105_ gnd vdd FILL
X_15009_ _14989_/A _15061_/C _15636_/B gnd _15009_/Y vdd NAND3X1
XFILL_0__9401_ gnd vdd FILL
XFILL_0__15883_ gnd vdd FILL
XFILL_5__13835_ gnd vdd FILL
XFILL_0__7593_ gnd vdd FILL
XFILL_3__9110_ gnd vdd FILL
XSFILL53720x7050 gnd vdd FILL
XFILL_4__15264_ gnd vdd FILL
XFILL_1__14104_ gnd vdd FILL
XFILL_3__10137_ gnd vdd FILL
XFILL_4__12476_ gnd vdd FILL
XFILL_1__11316_ gnd vdd FILL
XFILL_3__15994_ gnd vdd FILL
XFILL_2__13655_ gnd vdd FILL
XFILL_1__15084_ gnd vdd FILL
XSFILL99400x66050 gnd vdd FILL
XFILL_0__14834_ gnd vdd FILL
XFILL_5__7238_ gnd vdd FILL
XFILL_1__12296_ gnd vdd FILL
XSFILL59160x20050 gnd vdd FILL
XFILL_6__10248_ gnd vdd FILL
XFILL_4__14215_ gnd vdd FILL
XFILL_4__11427_ gnd vdd FILL
XFILL_5__10978_ gnd vdd FILL
XFILL_4__15195_ gnd vdd FILL
XFILL_2__12606_ gnd vdd FILL
XFILL_5__13766_ gnd vdd FILL
XFILL_1__14035_ gnd vdd FILL
XFILL_3__10068_ gnd vdd FILL
XFILL_3__9041_ gnd vdd FILL
XFILL_3__14945_ gnd vdd FILL
X_9960_ _9960_/Q _7527_/CLK _8935_/R vdd _9902_/Y gnd vdd DFFSR
XFILL_2__16374_ gnd vdd FILL
XFILL_1__11247_ gnd vdd FILL
XFILL_2__13586_ gnd vdd FILL
XFILL_2__10798_ gnd vdd FILL
XFILL_0__14765_ gnd vdd FILL
XFILL_5__7169_ gnd vdd FILL
XFILL_5__15505_ gnd vdd FILL
XFILL_0__11977_ gnd vdd FILL
XSFILL38840x19050 gnd vdd FILL
X_8911_ _8909_/Y _8896_/B _8910_/Y gnd _8947_/D vdd OAI21X1
XFILL_5__12717_ gnd vdd FILL
XFILL_4__14146_ gnd vdd FILL
XFILL_0__9263_ gnd vdd FILL
XFILL112360x26050 gnd vdd FILL
XFILL_2__15325_ gnd vdd FILL
XFILL_5__13697_ gnd vdd FILL
XFILL_4__11358_ gnd vdd FILL
X_9891_ _9957_/Q gnd _9891_/Y vdd INVX1
XFILL_3__14876_ gnd vdd FILL
XFILL_0__13716_ gnd vdd FILL
XFILL_0__10928_ gnd vdd FILL
XFILL_0_BUFX2_insert1000 gnd vdd FILL
XFILL_1__11178_ gnd vdd FILL
XFILL_0_BUFX2_insert1011 gnd vdd FILL
XFILL_0__14696_ gnd vdd FILL
XFILL_0__8214_ gnd vdd FILL
XFILL_0_BUFX2_insert1022 gnd vdd FILL
XFILL_4__10309_ gnd vdd FILL
XFILL_5__15436_ gnd vdd FILL
XFILL_5__12648_ gnd vdd FILL
X_8842_ _8840_/Y _8823_/B _8842_/C gnd _8924_/D vdd OAI21X1
XFILL_3__13827_ gnd vdd FILL
XSFILL109400x51050 gnd vdd FILL
XFILL_4__14077_ gnd vdd FILL
XFILL_0_BUFX2_insert1033 gnd vdd FILL
XFILL_2__15256_ gnd vdd FILL
XFILL_4__11289_ gnd vdd FILL
XFILL_1__10129_ gnd vdd FILL
XFILL_0_BUFX2_insert1044 gnd vdd FILL
XFILL_0__13647_ gnd vdd FILL
XFILL_2__12468_ gnd vdd FILL
XFILL_6__9721_ gnd vdd FILL
XFILL_1__15986_ gnd vdd FILL
XFILL_0_BUFX2_insert1055 gnd vdd FILL
XSFILL49080x72050 gnd vdd FILL
XFILL_0_BUFX2_insert1066 gnd vdd FILL
XFILL_4__13028_ gnd vdd FILL
XFILL_0__8145_ gnd vdd FILL
XFILL_5__12579_ gnd vdd FILL
XFILL_5__15367_ gnd vdd FILL
XFILL_2__14207_ gnd vdd FILL
X_8773_ _8759_/B _8005_/B gnd _8774_/C vdd NAND2X1
XFILL_3__13758_ gnd vdd FILL
XFILL_6_BUFX2_insert914 gnd vdd FILL
XFILL_2__11419_ gnd vdd FILL
XFILL_2__15187_ gnd vdd FILL
XFILL_2__12399_ gnd vdd FILL
XFILL_0_BUFX2_insert1088 gnd vdd FILL
XFILL_1__14937_ gnd vdd FILL
XFILL_0__16366_ gnd vdd FILL
XFILL_6_BUFX2_insert925 gnd vdd FILL
XFILL_0__13578_ gnd vdd FILL
XFILL_0__8076_ gnd vdd FILL
XFILL_5__14318_ gnd vdd FILL
X_7724_ _7724_/A gnd _7724_/Y vdd INVX1
XFILL_3__12709_ gnd vdd FILL
XFILL_5__15298_ gnd vdd FILL
XFILL_2__14138_ gnd vdd FILL
XSFILL114520x42050 gnd vdd FILL
XFILL_0__15317_ gnd vdd FILL
XSFILL115000x49050 gnd vdd FILL
XFILL_0__12529_ gnd vdd FILL
XFILL_3__9874_ gnd vdd FILL
XFILL_3__13689_ gnd vdd FILL
XSFILL44040x19050 gnd vdd FILL
XFILL_1__14868_ gnd vdd FILL
XFILL_0__16297_ gnd vdd FILL
XFILL_6__15608_ gnd vdd FILL
XFILL_5__14249_ gnd vdd FILL
X_7655_ _7593_/A _7016_/CLK _9064_/R vdd _7655_/D gnd vdd DFFSR
XFILL_3__15428_ gnd vdd FILL
XFILL_3__8825_ gnd vdd FILL
XFILL_1__13819_ gnd vdd FILL
XFILL_0__15248_ gnd vdd FILL
XFILL_4__14979_ gnd vdd FILL
XFILL_2__14069_ gnd vdd FILL
XFILL_1__14799_ gnd vdd FILL
XFILL_1__7840_ gnd vdd FILL
XFILL_3__15359_ gnd vdd FILL
X_7586_ _7584_/Y _7606_/A _7586_/C gnd _7652_/D vdd OAI21X1
XFILL_3__8756_ gnd vdd FILL
XFILL_0__15179_ gnd vdd FILL
X_9325_ _9325_/Q _9453_/CLK _9453_/R vdd _9325_/D gnd vdd DFFSR
XFILL_3__7707_ gnd vdd FILL
XFILL_0__8978_ gnd vdd FILL
XFILL_4_BUFX2_insert104 gnd vdd FILL
XFILL_4__7480_ gnd vdd FILL
XFILL_1__9510_ gnd vdd FILL
X_9256_ _9254_/Y _9277_/B _9256_/C gnd _9318_/D vdd OAI21X1
XFILL_0__7929_ gnd vdd FILL
XSFILL23720x41050 gnd vdd FILL
X_8207_ _8208_/B _8207_/B gnd _8208_/C vdd NAND2X1
XSFILL89960x55050 gnd vdd FILL
X_9187_ _9117_/A _9077_/CLK _7665_/R vdd _9119_/Y gnd vdd DFFSR
XFILL_4__9150_ gnd vdd FILL
XFILL_3_BUFX2_insert804 gnd vdd FILL
XFILL_3__7569_ gnd vdd FILL
XSFILL3640x39050 gnd vdd FILL
XFILL_3_BUFX2_insert815 gnd vdd FILL
X_8138_ _8138_/A gnd _8140_/A vdd INVX1
XFILL_3_BUFX2_insert826 gnd vdd FILL
XFILL_1__9372_ gnd vdd FILL
XFILL_4__8101_ gnd vdd FILL
XFILL_3_BUFX2_insert837 gnd vdd FILL
XFILL_3_BUFX2_insert848 gnd vdd FILL
XFILL_6__9017_ gnd vdd FILL
XFILL_3_BUFX2_insert859 gnd vdd FILL
XFILL_4__9081_ gnd vdd FILL
XFILL_1__8323_ gnd vdd FILL
XSFILL94280x27050 gnd vdd FILL
XSFILL114600x22050 gnd vdd FILL
X_8069_ _8069_/A gnd _8071_/A vdd INVX1
XFILL_3__9239_ gnd vdd FILL
XFILL_1__8254_ gnd vdd FILL
XSFILL103640x46050 gnd vdd FILL
XFILL_1__7205_ gnd vdd FILL
X_10971_ _10965_/Y _10971_/B gnd _10971_/Y vdd NAND2X1
XFILL_1__8185_ gnd vdd FILL
XFILL_4__9983_ gnd vdd FILL
X_12710_ _12710_/A gnd _12710_/Y vdd INVX1
X_13690_ _7643_/Q _14290_/C _13690_/C gnd _13698_/B vdd AOI21X1
XSFILL33560x44050 gnd vdd FILL
X_12641_ _12639_/Y vdd _12641_/C gnd _12687_/D vdd OAI21X1
XSFILL23800x21050 gnd vdd FILL
XFILL_1__7067_ gnd vdd FILL
XSFILL59080x7050 gnd vdd FILL
XFILL_4__8865_ gnd vdd FILL
XFILL_0_CLKBUF1_insert120 gnd vdd FILL
XFILL_0_CLKBUF1_insert131 gnd vdd FILL
X_15360_ _10333_/Q _15178_/C _15359_/Y gnd _15361_/C vdd AOI21X1
XFILL_0_BUFX2_insert705 gnd vdd FILL
XFILL_0_CLKBUF1_insert142 gnd vdd FILL
X_12572_ _12570_/Y vdd _12572_/C gnd _12664_/D vdd OAI21X1
XFILL_0_BUFX2_insert716 gnd vdd FILL
XFILL_2__6900_ gnd vdd FILL
XFILL_0_BUFX2_insert727 gnd vdd FILL
XFILL_0_CLKBUF1_insert153 gnd vdd FILL
XFILL_4__7816_ gnd vdd FILL
XFILL_0_CLKBUF1_insert164 gnd vdd FILL
XFILL_0_BUFX2_insert738 gnd vdd FILL
XSFILL3720x19050 gnd vdd FILL
XFILL_2__7880_ gnd vdd FILL
XFILL_0_BUFX2_insert749 gnd vdd FILL
X_14311_ _14311_/A _14311_/B gnd _14312_/A vdd NOR2X1
X_11523_ _11159_/Y gnd _11542_/B vdd INVX1
XFILL_0_CLKBUF1_insert175 gnd vdd FILL
XFILL_0_CLKBUF1_insert186 gnd vdd FILL
X_15291_ _15291_/A _15581_/C _16314_/A _13711_/D gnd _15293_/A vdd OAI22X1
XFILL_0_CLKBUF1_insert197 gnd vdd FILL
XFILL_4__7747_ gnd vdd FILL
X_14242_ _14234_/Y _14242_/B gnd _14243_/B vdd NAND2X1
XSFILL74280x1050 gnd vdd FILL
X_11454_ _11454_/A _11318_/C _11325_/Y gnd _11454_/Y vdd OAI21X1
XFILL_2__9550_ gnd vdd FILL
XSFILL13720x73050 gnd vdd FILL
XFILL_1__7969_ gnd vdd FILL
X_10405_ _10405_/A _10405_/B _10404_/Y gnd _10405_/Y vdd OAI21X1
XFILL_4__7678_ gnd vdd FILL
XFILL_2__8501_ gnd vdd FILL
X_14173_ _10469_/Q gnd _15674_/A vdd INVX1
X_11385_ _11380_/Y _11382_/Y _11385_/C gnd _11385_/Y vdd AOI21X1
XFILL_4__10660_ gnd vdd FILL
XFILL_2__9481_ gnd vdd FILL
XFILL_4__9417_ gnd vdd FILL
XFILL_5__8210_ gnd vdd FILL
X_13124_ _13190_/Q gnd _13126_/A vdd INVX1
XFILL_5__11950_ gnd vdd FILL
XFILL_4_BUFX2_insert660 gnd vdd FILL
X_10336_ _15474_/A _7791_/CLK _9711_/R vdd _10336_/D gnd vdd DFFSR
XFILL_3__11040_ gnd vdd FILL
XFILL_1__9639_ gnd vdd FILL
XFILL_4_BUFX2_insert671 gnd vdd FILL
XSFILL29400x61050 gnd vdd FILL
XFILL_4_BUFX2_insert682 gnd vdd FILL
XFILL_5__8141_ gnd vdd FILL
XFILL_4__9348_ gnd vdd FILL
XFILL_2__11770_ gnd vdd FILL
XFILL_5__10901_ gnd vdd FILL
XFILL_4_BUFX2_insert693 gnd vdd FILL
X_13055_ _6878_/A _7406_/CLK _8430_/R vdd _13055_/D gnd vdd DFFSR
XSFILL84280x59050 gnd vdd FILL
XFILL_4__12330_ gnd vdd FILL
X_10267_ _10285_/A _8091_/B gnd _10267_/Y vdd NAND2X1
XFILL_5__11881_ gnd vdd FILL
XFILL_0__11900_ gnd vdd FILL
XFILL_1__12150_ gnd vdd FILL
XFILL_2__8363_ gnd vdd FILL
XFILL_4__9279_ gnd vdd FILL
XFILL_5__8072_ gnd vdd FILL
X_12006_ _12006_/A _12006_/B _12005_/Y gnd _13092_/B vdd NAND3X1
XFILL_0__12880_ gnd vdd FILL
XFILL_5__13620_ gnd vdd FILL
XFILL_5__10832_ gnd vdd FILL
X_10198_ _10198_/Q _7382_/CLK _8674_/R vdd _10198_/D gnd vdd DFFSR
XFILL_4__12261_ gnd vdd FILL
XFILL_1__11101_ gnd vdd FILL
XFILL_2__7314_ gnd vdd FILL
XFILL_2__13440_ gnd vdd FILL
XFILL_2__10652_ gnd vdd FILL
XFILL_1__12081_ gnd vdd FILL
XFILL_3__12991_ gnd vdd FILL
XFILL_0__11831_ gnd vdd FILL
XFILL_4__14000_ gnd vdd FILL
XSFILL99480x40050 gnd vdd FILL
XFILL_5__13551_ gnd vdd FILL
XFILL_4__11212_ gnd vdd FILL
XFILL_5__10763_ gnd vdd FILL
XFILL_3__14730_ gnd vdd FILL
XFILL_2__7245_ gnd vdd FILL
XFILL_3__11942_ gnd vdd FILL
XFILL_4__12192_ gnd vdd FILL
XFILL_1__11032_ gnd vdd FILL
XFILL_0__14550_ gnd vdd FILL
XFILL_2__13371_ gnd vdd FILL
XFILL_0__11762_ gnd vdd FILL
XFILL_5__12502_ gnd vdd FILL
XFILL_4__11143_ gnd vdd FILL
X_13957_ _8928_/Q gnd _13959_/A vdd INVX1
XFILL_5__13482_ gnd vdd FILL
XFILL_2__15110_ gnd vdd FILL
XFILL_5__16270_ gnd vdd FILL
XFILL_5__10694_ gnd vdd FILL
XFILL_2__12322_ gnd vdd FILL
XFILL_3__14661_ gnd vdd FILL
XFILL_0__13501_ gnd vdd FILL
XFILL_2__7176_ gnd vdd FILL
XFILL_3__11873_ gnd vdd FILL
XFILL_2__16090_ gnd vdd FILL
XFILL_1__15840_ gnd vdd FILL
XFILL_0__14481_ gnd vdd FILL
XFILL_5__8974_ gnd vdd FILL
X_12908_ vdd _12908_/B gnd _12909_/C vdd NAND2X1
XFILL_5__15221_ gnd vdd FILL
XFILL_3__16400_ gnd vdd FILL
XFILL_5__12433_ gnd vdd FILL
XFILL_0__11693_ gnd vdd FILL
XSFILL74200x9050 gnd vdd FILL
XFILL_3__13612_ gnd vdd FILL
XSFILL13800x53050 gnd vdd FILL
XFILL_0__16220_ gnd vdd FILL
XFILL_2__15041_ gnd vdd FILL
XFILL_4__15951_ gnd vdd FILL
XFILL_2__12253_ gnd vdd FILL
XFILL_4__11074_ gnd vdd FILL
X_13888_ _9951_/Q gnd _15423_/D vdd INVX1
XFILL_3__10824_ gnd vdd FILL
XFILL_3__14592_ gnd vdd FILL
XFILL_0__13432_ gnd vdd FILL
XSFILL79240x48050 gnd vdd FILL
XFILL_1__15771_ gnd vdd FILL
XFILL_0__10644_ gnd vdd FILL
X_15627_ _15622_/Y _15627_/B _15627_/C gnd _15628_/C vdd NOR3X1
XFILL_1__12983_ gnd vdd FILL
XFILL_6__10935_ gnd vdd FILL
XFILL_5__12364_ gnd vdd FILL
XFILL_3__16331_ gnd vdd FILL
X_12839_ vdd _12839_/B gnd _12840_/C vdd NAND2X1
XFILL_5__15152_ gnd vdd FILL
XFILL_1_BUFX2_insert550 gnd vdd FILL
XFILL_4__14902_ gnd vdd FILL
XFILL_4__10025_ gnd vdd FILL
XFILL_1_BUFX2_insert561 gnd vdd FILL
XFILL_2__11204_ gnd vdd FILL
XFILL_3__13543_ gnd vdd FILL
XFILL_1_BUFX2_insert572 gnd vdd FILL
XFILL_2__12184_ gnd vdd FILL
XFILL_3__10755_ gnd vdd FILL
XFILL_3__6940_ gnd vdd FILL
XFILL_1__14722_ gnd vdd FILL
XFILL_0__16151_ gnd vdd FILL
XFILL_4__15882_ gnd vdd FILL
XFILL_0__13363_ gnd vdd FILL
XFILL_1__11934_ gnd vdd FILL
XFILL_0__10575_ gnd vdd FILL
XFILL_1_BUFX2_insert583 gnd vdd FILL
XSFILL114440x57050 gnd vdd FILL
XFILL_5__7856_ gnd vdd FILL
XFILL_5__14103_ gnd vdd FILL
XFILL_5__11315_ gnd vdd FILL
XFILL_1_BUFX2_insert594 gnd vdd FILL
XFILL_6__13654_ gnd vdd FILL
XFILL_5__15083_ gnd vdd FILL
X_15558_ _15322_/A _14050_/Y _14033_/Y _15558_/D gnd _15558_/Y vdd OAI22X1
XFILL_4__14833_ gnd vdd FILL
XFILL_5__12295_ gnd vdd FILL
XFILL_2__11135_ gnd vdd FILL
XFILL_0__15102_ gnd vdd FILL
XFILL_3__16262_ gnd vdd FILL
XFILL_3__13474_ gnd vdd FILL
XFILL_0__12314_ gnd vdd FILL
XFILL_3__10686_ gnd vdd FILL
XSFILL84360x39050 gnd vdd FILL
XFILL_1__11865_ gnd vdd FILL
XFILL_3__6871_ gnd vdd FILL
XFILL_1__14653_ gnd vdd FILL
XFILL_0__16082_ gnd vdd FILL
XFILL_0__13294_ gnd vdd FILL
X_14509_ _14509_/A _14466_/C gnd _14510_/C vdd NOR2X1
XFILL_5__14034_ gnd vdd FILL
XFILL_0__8901_ gnd vdd FILL
X_7440_ _7440_/A _7425_/B _7439_/Y gnd _7440_/Y vdd OAI21X1
XFILL_3__15213_ gnd vdd FILL
XFILL_5__11246_ gnd vdd FILL
XFILL_3__12425_ gnd vdd FILL
XFILL_3__8610_ gnd vdd FILL
XFILL_0__9881_ gnd vdd FILL
X_15489_ _8212_/A gnd _15490_/D vdd INVX1
XFILL_4__14764_ gnd vdd FILL
XFILL_1__13604_ gnd vdd FILL
XFILL_4__11976_ gnd vdd FILL
XFILL_3__16193_ gnd vdd FILL
XFILL_0__15033_ gnd vdd FILL
XFILL_2__15943_ gnd vdd FILL
XFILL_2__11066_ gnd vdd FILL
XFILL_5__9526_ gnd vdd FILL
XFILL_1__10816_ gnd vdd FILL
XFILL_3__9590_ gnd vdd FILL
XFILL_0__12245_ gnd vdd FILL
XFILL_1__14584_ gnd vdd FILL
XFILL_1__11796_ gnd vdd FILL
XSFILL59160x15050 gnd vdd FILL
XFILL_0__8832_ gnd vdd FILL
X_7371_ _7297_/B _7499_/B gnd _7372_/C vdd NAND2X1
XFILL_4__10927_ gnd vdd FILL
XFILL_2__10017_ gnd vdd FILL
XFILL_4__13715_ gnd vdd FILL
XFILL_3__15144_ gnd vdd FILL
XFILL_5__11177_ gnd vdd FILL
XFILL_3__12356_ gnd vdd FILL
XFILL_1__16323_ gnd vdd FILL
XFILL_4__14695_ gnd vdd FILL
XFILL_2__9748_ gnd vdd FILL
XFILL_1__13535_ gnd vdd FILL
XFILL_1__10747_ gnd vdd FILL
XFILL_2__15874_ gnd vdd FILL
X_9110_ _9108_/Y _9170_/B _9110_/C gnd _9184_/D vdd OAI21X1
XFILL_0__12176_ gnd vdd FILL
XFILL_5__10128_ gnd vdd FILL
XFILL_6__15255_ gnd vdd FILL
XFILL111880x14050 gnd vdd FILL
XFILL_0__8763_ gnd vdd FILL
XFILL_4__13646_ gnd vdd FILL
XFILL_3__11307_ gnd vdd FILL
XFILL_5__15985_ gnd vdd FILL
XFILL_2__14825_ gnd vdd FILL
XFILL_3__15075_ gnd vdd FILL
XFILL_2__9679_ gnd vdd FILL
XFILL_3__8472_ gnd vdd FILL
XFILL_3__12287_ gnd vdd FILL
XFILL_0__11127_ gnd vdd FILL
XFILL_1__16254_ gnd vdd FILL
XFILL_1__10678_ gnd vdd FILL
XFILL_6__14206_ gnd vdd FILL
XFILL_1__13466_ gnd vdd FILL
XSFILL23640x56050 gnd vdd FILL
XFILL_0__7714_ gnd vdd FILL
XFILL_5__9388_ gnd vdd FILL
X_9041_ _9017_/A _9041_/B gnd _9041_/Y vdd NAND2X1
XFILL_5__10059_ gnd vdd FILL
XFILL_3__14026_ gnd vdd FILL
XFILL_5__14936_ gnd vdd FILL
XFILL_3__7423_ gnd vdd FILL
XFILL_1__15205_ gnd vdd FILL
XFILL_4__16365_ gnd vdd FILL
XSFILL109400x46050 gnd vdd FILL
XFILL_0__8694_ gnd vdd FILL
XFILL_4__13577_ gnd vdd FILL
XFILL_3__11238_ gnd vdd FILL
XFILL_4__10789_ gnd vdd FILL
XFILL_1__12417_ gnd vdd FILL
XFILL_2__14756_ gnd vdd FILL
XFILL_1__13397_ gnd vdd FILL
XFILL_1__16185_ gnd vdd FILL
XFILL_0__15935_ gnd vdd FILL
XFILL_2__11968_ gnd vdd FILL
XFILL_5__8339_ gnd vdd FILL
XFILL_0__11058_ gnd vdd FILL
XSFILL49080x67050 gnd vdd FILL
XFILL_4__15316_ gnd vdd FILL
XFILL_4__12528_ gnd vdd FILL
XSFILL79320x28050 gnd vdd FILL
XFILL_6__11349_ gnd vdd FILL
XFILL_5__14867_ gnd vdd FILL
XFILL_4__16296_ gnd vdd FILL
XFILL_2__13707_ gnd vdd FILL
XFILL_2__10919_ gnd vdd FILL
XFILL_0__10009_ gnd vdd FILL
XFILL_3__7354_ gnd vdd FILL
XFILL_1__12348_ gnd vdd FILL
XFILL_1__15136_ gnd vdd FILL
XFILL_3__11169_ gnd vdd FILL
XFILL_2__14687_ gnd vdd FILL
XFILL_2__11899_ gnd vdd FILL
XFILL_0__15866_ gnd vdd FILL
XCLKBUF1_insert1078 clk gnd CLKBUF1_insert216/A vdd CLKBUF1
XSFILL64120x70050 gnd vdd FILL
XFILL_5__13818_ gnd vdd FILL
XFILL_4__15247_ gnd vdd FILL
XFILL_6__14068_ gnd vdd FILL
XFILL_4__12459_ gnd vdd FILL
XFILL_0__7576_ gnd vdd FILL
XFILL_2__13638_ gnd vdd FILL
XFILL_5__14798_ gnd vdd FILL
XSFILL114520x37050 gnd vdd FILL
XFILL_3__15977_ gnd vdd FILL
XFILL_0__14817_ gnd vdd FILL
XFILL_1__15067_ gnd vdd FILL
XFILL_1__12279_ gnd vdd FILL
XFILL_0_BUFX2_insert11 gnd vdd FILL
XFILL_0__15797_ gnd vdd FILL
XFILL_4__15178_ gnd vdd FILL
XFILL_5__13749_ gnd vdd FILL
XFILL_3__9024_ gnd vdd FILL
X_9943_ _9849_/A _7515_/CLK _7515_/R vdd _9851_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert22 gnd vdd FILL
XFILL_1__14018_ gnd vdd FILL
XFILL_2__16357_ gnd vdd FILL
XFILL_0_BUFX2_insert33 gnd vdd FILL
XFILL_3__14928_ gnd vdd FILL
XFILL_2__13569_ gnd vdd FILL
XFILL_0_BUFX2_insert44 gnd vdd FILL
XFILL_0__14748_ gnd vdd FILL
XFILL_0_BUFX2_insert55 gnd vdd FILL
XFILL_4__14129_ gnd vdd FILL
XFILL_0__9246_ gnd vdd FILL
XFILL_2__15308_ gnd vdd FILL
XFILL_0_BUFX2_insert66 gnd vdd FILL
XSFILL69080x2050 gnd vdd FILL
XFILL_3__14859_ gnd vdd FILL
XFILL_0_BUFX2_insert77 gnd vdd FILL
X_9874_ _9937_/A _9362_/B gnd _9874_/Y vdd NAND2X1
XFILL_2__16288_ gnd vdd FILL
XSFILL84040x21050 gnd vdd FILL
XFILL_0_BUFX2_insert88 gnd vdd FILL
XFILL_0_BUFX2_insert99 gnd vdd FILL
XFILL_0__14679_ gnd vdd FILL
XFILL_5__15419_ gnd vdd FILL
X_8825_ _8919_/Q gnd _8827_/A vdd INVX1
XFILL_2__15239_ gnd vdd FILL
XFILL_5__16399_ gnd vdd FILL
XFILL_6_BUFX2_insert700 gnd vdd FILL
XFILL_1__15969_ gnd vdd FILL
XFILL_4__6980_ gnd vdd FILL
XFILL_0__8128_ gnd vdd FILL
XFILL_3__9926_ gnd vdd FILL
X_8756_ _8756_/A _8788_/A _8756_/C gnd _8810_/D vdd OAI21X1
XFILL_1__9990_ gnd vdd FILL
XSFILL23720x36050 gnd vdd FILL
XFILL_0__16349_ gnd vdd FILL
XFILL_6_BUFX2_insert766 gnd vdd FILL
XFILL_6__6847_ gnd vdd FILL
XSFILL33880x80050 gnd vdd FILL
X_7707_ _7672_/B _7451_/B gnd _7708_/C vdd NAND2X1
XFILL_0__8059_ gnd vdd FILL
XSFILL18840x4050 gnd vdd FILL
XFILL_3__9857_ gnd vdd FILL
XFILL_4__8650_ gnd vdd FILL
X_8687_ _8687_/Q _7651_/CLK _7665_/R vdd _8643_/Y gnd vdd DFFSR
XFILL_1__8872_ gnd vdd FILL
X_7638_ _7638_/Q _8818_/CLK _9430_/R vdd _7544_/Y gnd vdd DFFSR
XFILL_4__7601_ gnd vdd FILL
XSFILL39400x24050 gnd vdd FILL
XFILL_3__9788_ gnd vdd FILL
XSFILL64200x50050 gnd vdd FILL
XFILL_4__8581_ gnd vdd FILL
XFILL_1_CLKBUF1_insert204 gnd vdd FILL
XSFILL79000x10050 gnd vdd FILL
XFILL_1__7823_ gnd vdd FILL
XFILL_1_CLKBUF1_insert215 gnd vdd FILL
XSFILL114600x17050 gnd vdd FILL
X_7569_ _7647_/Q gnd _7569_/Y vdd INVX1
XFILL_3__8739_ gnd vdd FILL
X_9308_ _9224_/A _9436_/CLK _9454_/R vdd _9226_/Y gnd vdd DFFSR
XFILL_1__7754_ gnd vdd FILL
XFILL_4__7463_ gnd vdd FILL
X_11170_ _11480_/A gnd _11174_/C vdd INVX4
X_9239_ _9313_/Q gnd _9241_/A vdd INVX1
XFILL_1__7685_ gnd vdd FILL
X_10121_ _10127_/A _6921_/B gnd _10122_/C vdd NAND2X1
XFILL_3_BUFX2_insert601 gnd vdd FILL
XFILL_3_BUFX2_insert612 gnd vdd FILL
XFILL_1__9424_ gnd vdd FILL
XFILL_3_BUFX2_insert623 gnd vdd FILL
XFILL_4__9133_ gnd vdd FILL
XFILL_3_BUFX2_insert634 gnd vdd FILL
XSFILL104520x69050 gnd vdd FILL
X_10052_ _14734_/A gnd _10054_/A vdd INVX1
XFILL_3_BUFX2_insert645 gnd vdd FILL
XFILL_3_BUFX2_insert656 gnd vdd FILL
XSFILL8760x67050 gnd vdd FILL
XFILL_1__9355_ gnd vdd FILL
XFILL_3_BUFX2_insert667 gnd vdd FILL
XSFILL23800x16050 gnd vdd FILL
XFILL_3_BUFX2_insert678 gnd vdd FILL
XSFILL84200x4050 gnd vdd FILL
XFILL_3_BUFX2_insert689 gnd vdd FILL
X_14860_ _9075_/Q gnd _14860_/Y vdd INVX1
XFILL_4__8015_ gnd vdd FILL
XFILL_1__9286_ gnd vdd FILL
XSFILL49240x27050 gnd vdd FILL
X_13811_ _8925_/Q gnd _13811_/Y vdd INVX1
XFILL_2__7030_ gnd vdd FILL
XFILL_1__8237_ gnd vdd FILL
X_14791_ _14765_/Y _14790_/Y _14791_/C gnd _13033_/B vdd AOI21X1
X_13742_ _13864_/B _8668_/Q _10844_/Q _13884_/C gnd _13750_/B vdd AOI22X1
X_10954_ _10941_/Y _10954_/B gnd _10955_/C vdd NOR2X1
XFILL_1__7119_ gnd vdd FILL
X_13673_ _13669_/Y _13673_/B gnd _13674_/C vdd NOR2X1
X_10885_ _12704_/A _12701_/A gnd _10892_/C vdd OR2X2
XFILL_1__8099_ gnd vdd FILL
XFILL_2__8981_ gnd vdd FILL
XFILL_5__7710_ gnd vdd FILL
X_15412_ _15412_/A _15411_/Y _15399_/Y gnd _15413_/B vdd NAND3X1
XFILL_4__8917_ gnd vdd FILL
X_12624_ _12624_/A gnd _12626_/A vdd INVX1
XFILL_4__9897_ gnd vdd FILL
X_16392_ _16392_/A gnd _16392_/C gnd _16392_/Y vdd OAI21X1
XFILL_0_BUFX2_insert502 gnd vdd FILL
XFILL_3__10540_ gnd vdd FILL
XFILL_2__7932_ gnd vdd FILL
XFILL_0_BUFX2_insert513 gnd vdd FILL
XFILL_0_BUFX2_insert524 gnd vdd FILL
XFILL_4__8848_ gnd vdd FILL
XFILL_0__10360_ gnd vdd FILL
XFILL_5__11100_ gnd vdd FILL
XFILL_0_BUFX2_insert535 gnd vdd FILL
X_15343_ _15343_/A _15342_/Y _15341_/Y gnd _15343_/Y vdd NOR3X1
XFILL_5__12080_ gnd vdd FILL
XFILL_0_BUFX2_insert546 gnd vdd FILL
X_12555_ _12403_/A _13201_/CLK _13201_/R vdd _12555_/D gnd vdd DFFSR
XFILL_4__11830_ gnd vdd FILL
XFILL_6__10651_ gnd vdd FILL
XFILL_0_BUFX2_insert557 gnd vdd FILL
XFILL_2__7863_ gnd vdd FILL
XFILL_0_BUFX2_insert568 gnd vdd FILL
XFILL_1__11650_ gnd vdd FILL
XFILL_4__8779_ gnd vdd FILL
XFILL_0_BUFX2_insert579 gnd vdd FILL
XFILL_5__7572_ gnd vdd FILL
X_11506_ _11571_/A _11500_/C gnd _11507_/C vdd NAND2X1
XFILL_5__11031_ gnd vdd FILL
XFILL_0__10291_ gnd vdd FILL
XFILL_2__9602_ gnd vdd FILL
XFILL_3__12210_ gnd vdd FILL
X_15274_ _15274_/A _15274_/B gnd _15296_/A vdd NOR2X1
X_12486_ _12484_/Y vdd _12485_/Y gnd _12486_/Y vdd OAI21X1
XFILL_4__11761_ gnd vdd FILL
XFILL_0__12030_ gnd vdd FILL
XFILL_1__11581_ gnd vdd FILL
X_14225_ _7398_/Q _14626_/A _13864_/C _8550_/Q gnd _14227_/A vdd AOI22X1
XSFILL99480x35050 gnd vdd FILL
XFILL_6__12321_ gnd vdd FILL
XFILL_4__13500_ gnd vdd FILL
X_11437_ _11437_/A _11435_/A _11437_/C gnd _11437_/Y vdd OAI21X1
XFILL_2__9533_ gnd vdd FILL
XFILL_4__14480_ gnd vdd FILL
XFILL_3__12141_ gnd vdd FILL
XSFILL74120x33050 gnd vdd FILL
XFILL_1__13320_ gnd vdd FILL
XFILL_1__10532_ gnd vdd FILL
XFILL_4__11692_ gnd vdd FILL
XFILL_5__9242_ gnd vdd FILL
XFILL_2__12871_ gnd vdd FILL
XFILL_6__15040_ gnd vdd FILL
X_14156_ _14156_/A gnd _14157_/C vdd INVX1
XFILL_4__13431_ gnd vdd FILL
XFILL_2__14610_ gnd vdd FILL
XFILL_5__15770_ gnd vdd FILL
XFILL_4__10643_ gnd vdd FILL
X_11368_ _11201_/Y _11349_/B _11367_/Y gnd _11417_/C vdd OAI21X1
XFILL_1__13251_ gnd vdd FILL
XFILL_3__12072_ gnd vdd FILL
XFILL_2__9464_ gnd vdd FILL
XFILL_5__12982_ gnd vdd FILL
XFILL_2__11822_ gnd vdd FILL
XCLKBUF1_insert203 CLKBUF1_insert192/A gnd _8947_/CLK vdd CLKBUF1
XFILL_2__15590_ gnd vdd FILL
XCLKBUF1_insert214 CLKBUF1_insert206/A gnd _9818_/CLK vdd CLKBUF1
XFILL_0__13981_ gnd vdd FILL
X_13107_ _13108_/B _12026_/Y gnd _13107_/Y vdd NAND2X1
XFILL_5__9173_ gnd vdd FILL
X_10319_ _10317_/Y _10318_/A _10319_/C gnd _10319_/Y vdd OAI21X1
XFILL_5__14721_ gnd vdd FILL
XFILL_6__12183_ gnd vdd FILL
XFILL_4_BUFX2_insert490 gnd vdd FILL
XFILL_4__16150_ gnd vdd FILL
XFILL_4__13362_ gnd vdd FILL
XFILL_3__15900_ gnd vdd FILL
XFILL_5__11933_ gnd vdd FILL
XFILL_1__12202_ gnd vdd FILL
XSFILL13800x48050 gnd vdd FILL
X_14087_ _7197_/A gnd _14088_/A vdd INVX1
XFILL_3__11023_ gnd vdd FILL
XFILL_4__10574_ gnd vdd FILL
XFILL_2__14541_ gnd vdd FILL
XSFILL78760x36050 gnd vdd FILL
X_11299_ _11133_/Y gnd _11620_/B vdd INVX1
XFILL_5__8124_ gnd vdd FILL
XFILL_0__15720_ gnd vdd FILL
XFILL_2__9395_ gnd vdd FILL
XFILL_2__11753_ gnd vdd FILL
XFILL_1__10394_ gnd vdd FILL
XFILL_6__11134_ gnd vdd FILL
XFILL_4__15101_ gnd vdd FILL
X_13038_ _6899_/A gnd _13038_/Y vdd INVX1
XFILL_4__12313_ gnd vdd FILL
XFILL_0__7430_ gnd vdd FILL
XFILL_5__14652_ gnd vdd FILL
XFILL_4__16081_ gnd vdd FILL
XFILL_4__13293_ gnd vdd FILL
XFILL_1__12133_ gnd vdd FILL
XFILL_2__8346_ gnd vdd FILL
XFILL_3__15831_ gnd vdd FILL
XFILL_5__11864_ gnd vdd FILL
XFILL_2__10704_ gnd vdd FILL
XFILL_2__14472_ gnd vdd FILL
XFILL_5__8055_ gnd vdd FILL
XFILL_0__15651_ gnd vdd FILL
XFILL_2__11684_ gnd vdd FILL
XFILL_0__12863_ gnd vdd FILL
XFILL_5__13603_ gnd vdd FILL
XFILL_4__15032_ gnd vdd FILL
XFILL_5__10815_ gnd vdd FILL
XFILL_2__16211_ gnd vdd FILL
XFILL_4__12244_ gnd vdd FILL
XFILL_0__7361_ gnd vdd FILL
XFILL_5__14583_ gnd vdd FILL
XFILL_2__13423_ gnd vdd FILL
XFILL_3__15762_ gnd vdd FILL
XFILL_5__11795_ gnd vdd FILL
XFILL_2__10635_ gnd vdd FILL
XFILL_0__14602_ gnd vdd FILL
XFILL_3__12974_ gnd vdd FILL
XFILL_1__12064_ gnd vdd FILL
XFILL_2__8277_ gnd vdd FILL
XFILL_3__7070_ gnd vdd FILL
XFILL_0__11814_ gnd vdd FILL
XFILL_0__9100_ gnd vdd FILL
XFILL_6__10016_ gnd vdd FILL
XFILL_0__15582_ gnd vdd FILL
XFILL_5__16322_ gnd vdd FILL
X_6940_ _6940_/A _6948_/A _6939_/Y gnd _7010_/D vdd OAI21X1
XFILL_3__14713_ gnd vdd FILL
XFILL_5__10746_ gnd vdd FILL
XFILL_5__13534_ gnd vdd FILL
XFILL_0__7292_ gnd vdd FILL
XFILL_2__7228_ gnd vdd FILL
X_14989_ _14989_/A _14982_/Y _15061_/C gnd _14989_/Y vdd NAND3X1
XFILL_3__11925_ gnd vdd FILL
XFILL_4__12175_ gnd vdd FILL
XSFILL43880x43050 gnd vdd FILL
XFILL_2__16142_ gnd vdd FILL
XFILL_1__11015_ gnd vdd FILL
XFILL_2__13354_ gnd vdd FILL
XFILL_3__15693_ gnd vdd FILL
XFILL_0__14533_ gnd vdd FILL
XFILL_2__10566_ gnd vdd FILL
XFILL_0__11745_ gnd vdd FILL
XFILL_0__9031_ gnd vdd FILL
XFILL_3_CLKBUF1_insert170 gnd vdd FILL
XFILL_4__11126_ gnd vdd FILL
XFILL_5__16253_ gnd vdd FILL
XFILL_5__10677_ gnd vdd FILL
XFILL_3_CLKBUF1_insert181 gnd vdd FILL
XFILL_3__14644_ gnd vdd FILL
XFILL_5__13465_ gnd vdd FILL
XFILL_2__12305_ gnd vdd FILL
X_6871_ _6871_/A gnd memoryWriteData[1] vdd BUFX2
XFILL_3_CLKBUF1_insert192 gnd vdd FILL
XFILL_2__7159_ gnd vdd FILL
XFILL_1__15823_ gnd vdd FILL
XFILL_3__11856_ gnd vdd FILL
XFILL_2__16073_ gnd vdd FILL
XSFILL99560x15050 gnd vdd FILL
XFILL_2__13285_ gnd vdd FILL
XFILL_2__10497_ gnd vdd FILL
XFILL_0__14464_ gnd vdd FILL
XFILL_5__15204_ gnd vdd FILL
XFILL_0__11676_ gnd vdd FILL
XSFILL74200x13050 gnd vdd FILL
XFILL_5__12416_ gnd vdd FILL
X_8610_ _8610_/A _8609_/A _8610_/C gnd _8676_/D vdd OAI21X1
XFILL_5__8957_ gnd vdd FILL
XFILL_3__10807_ gnd vdd FILL
XFILL_5__16184_ gnd vdd FILL
XFILL_5__13396_ gnd vdd FILL
X_9590_ _9686_/Q gnd _9590_/Y vdd INVX1
XFILL_4__15934_ gnd vdd FILL
XFILL_2__15024_ gnd vdd FILL
XFILL_4__11057_ gnd vdd FILL
XFILL_3__14575_ gnd vdd FILL
XFILL_0__16203_ gnd vdd FILL
XFILL_0__13415_ gnd vdd FILL
XFILL_2__12236_ gnd vdd FILL
XFILL_3__7972_ gnd vdd FILL
XFILL_0__10627_ gnd vdd FILL
XFILL_3__11787_ gnd vdd FILL
XFILL_1__15754_ gnd vdd FILL
XFILL_0__14395_ gnd vdd FILL
XFILL_1__12966_ gnd vdd FILL
XFILL_5__12347_ gnd vdd FILL
XFILL_5__8888_ gnd vdd FILL
XFILL_4__10008_ gnd vdd FILL
XFILL_1_BUFX2_insert380 gnd vdd FILL
XFILL_3__16314_ gnd vdd FILL
XFILL_5__15135_ gnd vdd FILL
X_8541_ _8459_/A _8541_/CLK _8285_/R vdd _8461_/Y gnd vdd DFFSR
XFILL_1_BUFX2_insert391 gnd vdd FILL
XFILL_3__13526_ gnd vdd FILL
XFILL_3__6923_ gnd vdd FILL
XFILL_1__14705_ gnd vdd FILL
XFILL_4__15865_ gnd vdd FILL
XFILL_0__13346_ gnd vdd FILL
XFILL_6__9420_ gnd vdd FILL
XFILL_1__11917_ gnd vdd FILL
XFILL_2__12167_ gnd vdd FILL
XFILL_0__16134_ gnd vdd FILL
XFILL_0__10558_ gnd vdd FILL
XFILL_1__15685_ gnd vdd FILL
XFILL_5_BUFX2_insert707 gnd vdd FILL
XFILL_5__7839_ gnd vdd FILL
XFILL_0__9933_ gnd vdd FILL
XFILL_1__12897_ gnd vdd FILL
XFILL_5_BUFX2_insert718 gnd vdd FILL
XFILL111720x73050 gnd vdd FILL
X_8472_ _8503_/B _8472_/B gnd _8473_/C vdd NAND2X1
XFILL_5__15066_ gnd vdd FILL
XFILL_4__14816_ gnd vdd FILL
XFILL_5_BUFX2_insert729 gnd vdd FILL
XFILL_5__12278_ gnd vdd FILL
XFILL_3__16245_ gnd vdd FILL
XFILL_3__13457_ gnd vdd FILL
XFILL_2__11118_ gnd vdd FILL
XFILL_3__9642_ gnd vdd FILL
XFILL_1__14636_ gnd vdd FILL
XFILL_3__6854_ gnd vdd FILL
XFILL_2__12098_ gnd vdd FILL
XFILL_4__15796_ gnd vdd FILL
XFILL_3__10669_ gnd vdd FILL
XFILL_0__16065_ gnd vdd FILL
XFILL_0__13277_ gnd vdd FILL
XSFILL89480x67050 gnd vdd FILL
XFILL_1__11848_ gnd vdd FILL
X_7423_ _7513_/Q gnd _7425_/A vdd INVX1
XFILL_5__14017_ gnd vdd FILL
XFILL_0__10489_ gnd vdd FILL
XFILL_5__11229_ gnd vdd FILL
XFILL_3__12408_ gnd vdd FILL
XSFILL64120x65050 gnd vdd FILL
XFILL_0__9864_ gnd vdd FILL
XFILL_2__15926_ gnd vdd FILL
XFILL_4__11959_ gnd vdd FILL
XFILL_3__16176_ gnd vdd FILL
XFILL_4__14747_ gnd vdd FILL
XFILL_0__15016_ gnd vdd FILL
XFILL_2__11049_ gnd vdd FILL
XFILL_3__13388_ gnd vdd FILL
XFILL_0__12228_ gnd vdd FILL
XFILL_5__9509_ gnd vdd FILL
XFILL_1__14567_ gnd vdd FILL
XFILL_1__11779_ gnd vdd FILL
X_7354_ _7352_/Y _7354_/B _7353_/Y gnd _7354_/Y vdd OAI21X1
XFILL_3__15127_ gnd vdd FILL
XFILL_3__8524_ gnd vdd FILL
XFILL_3__12339_ gnd vdd FILL
XFILL_1__16306_ gnd vdd FILL
XFILL_0__9795_ gnd vdd FILL
XFILL_4__14678_ gnd vdd FILL
XFILL_1__13518_ gnd vdd FILL
XFILL_2__15857_ gnd vdd FILL
XFILL_0__12159_ gnd vdd FILL
XFILL_1__14498_ gnd vdd FILL
XSFILL43960x23050 gnd vdd FILL
XSFILL3560x72050 gnd vdd FILL
XFILL_0__8746_ gnd vdd FILL
XFILL_4__13629_ gnd vdd FILL
XFILL_2__14808_ gnd vdd FILL
XFILL_3__15058_ gnd vdd FILL
XFILL_5__15968_ gnd vdd FILL
X_7285_ _7251_/A _9447_/CLK _7285_/R vdd _7285_/D gnd vdd DFFSR
XFILL_1__16237_ gnd vdd FILL
XFILL_3__8455_ gnd vdd FILL
XFILL_1__13449_ gnd vdd FILL
XSFILL84840x35050 gnd vdd FILL
XFILL_2__15788_ gnd vdd FILL
X_9024_ _9022_/Y _8996_/A _9024_/C gnd _9024_/Y vdd OAI21X1
XFILL_3__14009_ gnd vdd FILL
XFILL_5__14919_ gnd vdd FILL
XSFILL83800x71050 gnd vdd FILL
XFILL_1__7470_ gnd vdd FILL
XFILL_4__16348_ gnd vdd FILL
XFILL_5__15899_ gnd vdd FILL
XFILL_2__14739_ gnd vdd FILL
XFILL_6__7115_ gnd vdd FILL
XFILL_0__15918_ gnd vdd FILL
XFILL_1__16168_ gnd vdd FILL
XFILL_3__8386_ gnd vdd FILL
XFILL_0__7628_ gnd vdd FILL
XFILL_3__7337_ gnd vdd FILL
XFILL_1__15119_ gnd vdd FILL
XFILL_4__16279_ gnd vdd FILL
XFILL_1__16099_ gnd vdd FILL
XFILL_0__15849_ gnd vdd FILL
XFILL_2_BUFX2_insert608 gnd vdd FILL
XFILL_1__9140_ gnd vdd FILL
XSFILL33880x75050 gnd vdd FILL
XFILL_2__16409_ gnd vdd FILL
XFILL_2_BUFX2_insert619 gnd vdd FILL
XFILL_0__7559_ gnd vdd FILL
XFILL111800x53050 gnd vdd FILL
XSFILL23320x33050 gnd vdd FILL
X_9926_ _9924_/Y _9868_/A _9925_/Y gnd _9968_/D vdd OAI21X1
XFILL_3__9007_ gnd vdd FILL
XSFILL89560x47050 gnd vdd FILL
XSFILL38920x12050 gnd vdd FILL
XSFILL64200x45050 gnd vdd FILL
XFILL_3__7199_ gnd vdd FILL
XFILL_0__9229_ gnd vdd FILL
X_9857_ _9857_/A _9920_/B _9857_/C gnd _9945_/D vdd OAI21X1
XFILL_6__8997_ gnd vdd FILL
XSFILL68680x4050 gnd vdd FILL
XSFILL39000x21050 gnd vdd FILL
XFILL_6__7948_ gnd vdd FILL
X_8808_ _8808_/Q _7016_/CLK _9704_/R vdd _8808_/D gnd vdd DFFSR
X_9788_ _9789_/B _9788_/B gnd _9788_/Y vdd NAND2X1
XFILL_4__9751_ gnd vdd FILL
XSFILL3640x52050 gnd vdd FILL
XFILL_6_BUFX2_insert541 gnd vdd FILL
XFILL_4__6963_ gnd vdd FILL
XBUFX2_insert607 BUFX2_insert607/A gnd _9061_/R vdd BUFX2
X_10670_ _10670_/A _10615_/B _10670_/C gnd _10728_/D vdd OAI21X1
XBUFX2_insert618 _13430_/Y gnd _14762_/B vdd BUFX2
X_8739_ _8805_/Q gnd _8741_/A vdd INVX1
XFILL_4__8702_ gnd vdd FILL
XFILL_3__9909_ gnd vdd FILL
XBUFX2_insert629 _13465_/Y gnd _14744_/B vdd BUFX2
XSFILL28040x45050 gnd vdd FILL
XFILL_4__9682_ gnd vdd FILL
XSFILL94280x40050 gnd vdd FILL
XFILL_4__6894_ gnd vdd FILL
XFILL_4__8633_ gnd vdd FILL
X_12340_ _12312_/A _12340_/B _12312_/C gnd _12342_/B vdd NAND3X1
XFILL_6__9549_ gnd vdd FILL
XFILL_1__8855_ gnd vdd FILL
X_12271_ _12255_/A gnd _12255_/C gnd _12271_/Y vdd NAND3X1
XFILL_1__7806_ gnd vdd FILL
XFILL_1__8786_ gnd vdd FILL
X_14010_ _14010_/A _13803_/A _14575_/C _14008_/Y gnd _14010_/Y vdd OAI22X1
XSFILL74040x48050 gnd vdd FILL
XFILL_4__8495_ gnd vdd FILL
X_11222_ _11218_/B _11227_/A gnd _11222_/Y vdd AND2X2
XFILL_1__7737_ gnd vdd FILL
XFILL_4__7446_ gnd vdd FILL
X_11153_ _12290_/Y _11153_/B gnd _11153_/Y vdd NOR2X1
XFILL_3_BUFX2_insert420 gnd vdd FILL
XFILL_3_BUFX2_insert431 gnd vdd FILL
X_10104_ _10104_/A _10140_/B _10103_/Y gnd _10198_/D vdd OAI21X1
XFILL_4__7377_ gnd vdd FILL
XFILL_1__9407_ gnd vdd FILL
XFILL_2__8200_ gnd vdd FILL
XFILL_3_BUFX2_insert442 gnd vdd FILL
X_15961_ _15646_/D _14532_/D _15899_/C _15961_/D gnd _15961_/Y vdd OAI22X1
X_11084_ _12262_/Y _11083_/Y gnd _11085_/C vdd NOR2X1
XFILL_3_BUFX2_insert453 gnd vdd FILL
XFILL_4__9116_ gnd vdd FILL
XSFILL3720x32050 gnd vdd FILL
XFILL_3_BUFX2_insert464 gnd vdd FILL
XFILL_1__7599_ gnd vdd FILL
XFILL_3_BUFX2_insert475 gnd vdd FILL
XSFILL94360x5050 gnd vdd FILL
X_10035_ _10054_/B _9011_/B gnd _10036_/C vdd NAND2X1
X_14912_ _14910_/Y _14506_/C _14718_/B _14911_/Y gnd _14916_/B vdd OAI22X1
XFILL_3_BUFX2_insert486 gnd vdd FILL
X_15892_ _9269_/A _15892_/B gnd _15892_/Y vdd NAND2X1
XFILL_3_BUFX2_insert497 gnd vdd FILL
XFILL_2__8131_ gnd vdd FILL
XFILL_1__9338_ gnd vdd FILL
XSFILL79560x79050 gnd vdd FILL
XFILL_4__10290_ gnd vdd FILL
XSFILL28120x25050 gnd vdd FILL
XSFILL94360x20050 gnd vdd FILL
X_14843_ _7027_/Q gnd _14843_/Y vdd INVX1
XFILL_5__11580_ gnd vdd FILL
XFILL_1__9269_ gnd vdd FILL
XFILL_2__10420_ gnd vdd FILL
XFILL_2__8062_ gnd vdd FILL
XFILL_5__10531_ gnd vdd FILL
XFILL_5__9860_ gnd vdd FILL
XFILL_3__11710_ gnd vdd FILL
X_14774_ _8433_/Q _14037_/B _14956_/D _14774_/D gnd _14774_/Y vdd AOI22X1
X_11986_ _12072_/A gnd _12072_/C gnd _11986_/Y vdd NAND3X1
XFILL_0_BUFX2_insert3 gnd vdd FILL
XFILL_0__11530_ gnd vdd FILL
XFILL_5__9791_ gnd vdd FILL
XFILL_5__13250_ gnd vdd FILL
X_13725_ _13725_/A _13868_/B _14456_/C _13725_/D gnd _13726_/B vdd OAI22X1
X_10937_ _12779_/A gnd _10957_/B vdd INVX2
XFILL_4_CLKBUF1_insert210 gnd vdd FILL
XSFILL74120x28050 gnd vdd FILL
XFILL_3__11641_ gnd vdd FILL
XFILL_4__13980_ gnd vdd FILL
XFILL_2__10282_ gnd vdd FILL
XFILL_5__8742_ gnd vdd FILL
XFILL_5__12201_ gnd vdd FILL
XFILL_4_CLKBUF1_insert221 gnd vdd FILL
XFILL_0__11461_ gnd vdd FILL
X_16444_ _14776_/A _6999_/CLK _7011_/R vdd _16404_/Y gnd vdd DFFSR
X_13656_ _8962_/A gnd _15211_/A vdd INVX1
XFILL_2__12021_ gnd vdd FILL
XFILL_5__10393_ gnd vdd FILL
XFILL_3__14360_ gnd vdd FILL
X_10868_ _14883_/A _8297_/CLK _7796_/R vdd _10868_/D gnd vdd DFFSR
XFILL_2__8964_ gnd vdd FILL
XFILL_0__10412_ gnd vdd FILL
XFILL_3__11572_ gnd vdd FILL
XFILL_1__12751_ gnd vdd FILL
XFILL_0__14180_ gnd vdd FILL
XFILL_0_BUFX2_insert310 gnd vdd FILL
XFILL_6__10703_ gnd vdd FILL
X_12607_ vdd memoryOutData[13] gnd _12608_/C vdd NAND2X1
XFILL_0_BUFX2_insert321 gnd vdd FILL
XFILL_0__11392_ gnd vdd FILL
XFILL_5__12132_ gnd vdd FILL
XFILL_3__13311_ gnd vdd FILL
X_16375_ _15787_/A gnd _16375_/Y vdd INVX1
XFILL_0_BUFX2_insert332 gnd vdd FILL
X_13587_ _13587_/A _13586_/Y _13587_/C _13587_/D gnd _13591_/A vdd OAI22X1
XFILL_4__15650_ gnd vdd FILL
XFILL_3__10523_ gnd vdd FILL
XFILL_0_BUFX2_insert343 gnd vdd FILL
XFILL_4__12862_ gnd vdd FILL
XFILL_0__13131_ gnd vdd FILL
X_10799_ _14358_/A gnd _10801_/A vdd INVX1
XFILL_3__14291_ gnd vdd FILL
XFILL_1__11702_ gnd vdd FILL
XSFILL109480x15050 gnd vdd FILL
XFILL_2__8895_ gnd vdd FILL
XFILL_0_BUFX2_insert354 gnd vdd FILL
XFILL_5__7624_ gnd vdd FILL
XFILL_1__15470_ gnd vdd FILL
X_15326_ _13767_/Y _15681_/B _15681_/C _13744_/Y gnd _15329_/B vdd OAI22X1
XFILL_0_BUFX2_insert365 gnd vdd FILL
XSFILL8760x6050 gnd vdd FILL
XFILL_4__14601_ gnd vdd FILL
X_12538_ _12352_/A _12538_/CLK _12795_/R vdd _12450_/Y gnd vdd DFFSR
XFILL_3__16030_ gnd vdd FILL
XFILL_5__12063_ gnd vdd FILL
XFILL_0_BUFX2_insert376 gnd vdd FILL
XFILL_0__6930_ gnd vdd FILL
XFILL_4__11813_ gnd vdd FILL
XFILL_3__13242_ gnd vdd FILL
XFILL_0_BUFX2_insert387 gnd vdd FILL
XSFILL54120x8050 gnd vdd FILL
XFILL_2__7846_ gnd vdd FILL
XFILL112280x54050 gnd vdd FILL
XSFILL93800x34050 gnd vdd FILL
XFILL_1__14421_ gnd vdd FILL
XFILL_4__15581_ gnd vdd FILL
XFILL_0_BUFX2_insert398 gnd vdd FILL
XFILL_1__11633_ gnd vdd FILL
XFILL_2__13972_ gnd vdd FILL
XFILL_5__7555_ gnd vdd FILL
XFILL_0__10274_ gnd vdd FILL
XFILL_5__11014_ gnd vdd FILL
X_15257_ _15250_/Y _15257_/B _15257_/C gnd _15258_/B vdd NAND3X1
XFILL_2__15711_ gnd vdd FILL
XFILL_0__6861_ gnd vdd FILL
XSFILL53800x50050 gnd vdd FILL
XFILL_4__14532_ gnd vdd FILL
X_12469_ _12027_/B gnd _12469_/Y vdd INVX1
XFILL_4__11744_ gnd vdd FILL
XFILL_0__12013_ gnd vdd FILL
XFILL_3__13173_ gnd vdd FILL
XFILL_1__14352_ gnd vdd FILL
XFILL_3__10385_ gnd vdd FILL
XFILL_1__11564_ gnd vdd FILL
X_14208_ _14208_/A _14643_/B _13467_/A _14207_/Y gnd _14208_/Y vdd OAI22X1
XFILL_0__8600_ gnd vdd FILL
XFILL_5__7486_ gnd vdd FILL
XFILL_5__15822_ gnd vdd FILL
XFILL_4__14463_ gnd vdd FILL
X_15188_ _13628_/Y _15972_/B _15392_/C _13629_/Y gnd _15192_/A vdd OAI22X1
XFILL_3__12124_ gnd vdd FILL
XFILL_2__9516_ gnd vdd FILL
XFILL_1__13303_ gnd vdd FILL
XSFILL79240x61050 gnd vdd FILL
XFILL_2__15642_ gnd vdd FILL
XSFILL43880x38050 gnd vdd FILL
XFILL_4__11675_ gnd vdd FILL
XFILL_1__10515_ gnd vdd FILL
XFILL_5__9225_ gnd vdd FILL
XFILL_2__12854_ gnd vdd FILL
XFILL_1__11495_ gnd vdd FILL
XFILL_1__14283_ gnd vdd FILL
XFILL_4__16202_ gnd vdd FILL
X_14139_ _8736_/A gnd _14141_/B vdd INVX1
XFILL_4__13414_ gnd vdd FILL
XFILL_0__8531_ gnd vdd FILL
XFILL_4__10626_ gnd vdd FILL
X_7070_ _7061_/A _8606_/B gnd _7071_/C vdd NAND2X1
XFILL_5__15753_ gnd vdd FILL
XFILL_1__16022_ gnd vdd FILL
XFILL_5__12965_ gnd vdd FILL
XFILL_3__12055_ gnd vdd FILL
XFILL_5_BUFX2_insert1000 gnd vdd FILL
XFILL_4__14394_ gnd vdd FILL
XFILL_3__8240_ gnd vdd FILL
XFILL_2__11805_ gnd vdd FILL
XFILL_1__10446_ gnd vdd FILL
XFILL_1__13234_ gnd vdd FILL
XFILL_5_BUFX2_insert1011 gnd vdd FILL
XFILL_2__15573_ gnd vdd FILL
XSFILL18680x14050 gnd vdd FILL
XFILL_2__12785_ gnd vdd FILL
XFILL_5__9156_ gnd vdd FILL
XSFILL8520x24050 gnd vdd FILL
XFILL_5_BUFX2_insert1022 gnd vdd FILL
XFILL_5__14704_ gnd vdd FILL
XFILL_0__13964_ gnd vdd FILL
XFILL_5_BUFX2_insert1033 gnd vdd FILL
XFILL_4__13345_ gnd vdd FILL
XFILL_0__8462_ gnd vdd FILL
XFILL_5__11916_ gnd vdd FILL
XFILL_3__11006_ gnd vdd FILL
XFILL_4__16133_ gnd vdd FILL
XFILL_5_BUFX2_insert1044 gnd vdd FILL
XFILL_5__15684_ gnd vdd FILL
XFILL_4__10557_ gnd vdd FILL
XFILL_2__14524_ gnd vdd FILL
XFILL_5__12896_ gnd vdd FILL
XFILL_0__15703_ gnd vdd FILL
XFILL_2__9378_ gnd vdd FILL
XFILL_1__13165_ gnd vdd FILL
XSFILL84360x52050 gnd vdd FILL
XFILL_5_BUFX2_insert1055 gnd vdd FILL
XFILL_2__11736_ gnd vdd FILL
XFILL_5__8107_ gnd vdd FILL
XFILL_1__10377_ gnd vdd FILL
XFILL_5_BUFX2_insert1066 gnd vdd FILL
XFILL_0__12915_ gnd vdd FILL
XFILL_5__9087_ gnd vdd FILL
XSFILL59000x69050 gnd vdd FILL
XFILL_5__14635_ gnd vdd FILL
XFILL_0__13895_ gnd vdd FILL
XFILL_4__16064_ gnd vdd FILL
XFILL_4__13276_ gnd vdd FILL
XFILL_2__8329_ gnd vdd FILL
XFILL_5_BUFX2_insert1088 gnd vdd FILL
XFILL_1__12116_ gnd vdd FILL
XFILL_3__15814_ gnd vdd FILL
XFILL_3__7122_ gnd vdd FILL
XFILL_5__11847_ gnd vdd FILL
XFILL_0__8393_ gnd vdd FILL
XFILL_2__14455_ gnd vdd FILL
XFILL_4__10488_ gnd vdd FILL
XFILL_0__15634_ gnd vdd FILL
XFILL_1__13096_ gnd vdd FILL
XFILL_2__11667_ gnd vdd FILL
XFILL_6__15925_ gnd vdd FILL
XFILL_0__12846_ gnd vdd FILL
XFILL_4__15015_ gnd vdd FILL
XFILL_4__12227_ gnd vdd FILL
XFILL_0__7344_ gnd vdd FILL
XFILL_5__14566_ gnd vdd FILL
XFILL_2__13406_ gnd vdd FILL
XFILL_3__7053_ gnd vdd FILL
X_7972_ _7972_/A _7972_/B gnd _7973_/C vdd NAND2X1
XFILL_1__12047_ gnd vdd FILL
XFILL_2__10618_ gnd vdd FILL
XFILL_3__12957_ gnd vdd FILL
XFILL_5__11778_ gnd vdd FILL
XFILL_3__15745_ gnd vdd FILL
XFILL_2__14386_ gnd vdd FILL
XFILL_0__12777_ gnd vdd FILL
XFILL_0__15565_ gnd vdd FILL
XFILL_5__16305_ gnd vdd FILL
XFILL_2__11598_ gnd vdd FILL
XFILL112360x34050 gnd vdd FILL
X_9711_ _9711_/Q _7651_/CLK _9711_/R vdd _9711_/D gnd vdd DFFSR
XFILL_5__13517_ gnd vdd FILL
X_6923_ _7005_/Q gnd _6923_/Y vdd INVX1
XFILL_3__11908_ gnd vdd FILL
XFILL_4__12158_ gnd vdd FILL
XFILL_2__16125_ gnd vdd FILL
XFILL_2__13337_ gnd vdd FILL
XFILL_3__15676_ gnd vdd FILL
XFILL_5__14497_ gnd vdd FILL
XFILL_2__10549_ gnd vdd FILL
XFILL_3__12888_ gnd vdd FILL
XFILL_0__14516_ gnd vdd FILL
XSFILL79720x39050 gnd vdd FILL
XFILL_0__11728_ gnd vdd FILL
XFILL_0__9014_ gnd vdd FILL
XFILL_5__16236_ gnd vdd FILL
XFILL_0__15496_ gnd vdd FILL
XFILL_4__11109_ gnd vdd FILL
XFILL_3__14627_ gnd vdd FILL
XFILL_5__13448_ gnd vdd FILL
XFILL_6__15787_ gnd vdd FILL
XFILL_5__9989_ gnd vdd FILL
X_9642_ _9628_/B _9898_/B gnd _9642_/Y vdd NAND2X1
X_6854_ _6854_/A gnd memoryAddress[16] vdd BUFX2
XFILL_4__12089_ gnd vdd FILL
XFILL_1__15806_ gnd vdd FILL
XFILL_3_BUFX2_insert1070 gnd vdd FILL
XFILL_2__16056_ gnd vdd FILL
XFILL_3__11839_ gnd vdd FILL
XFILL_2__13268_ gnd vdd FILL
XFILL_0__11659_ gnd vdd FILL
XFILL_0__14447_ gnd vdd FILL
XFILL_1__13998_ gnd vdd FILL
XSFILL79320x41050 gnd vdd FILL
XFILL_3_BUFX2_insert1092 gnd vdd FILL
XFILL_6__14738_ gnd vdd FILL
XSFILL43960x18050 gnd vdd FILL
XFILL_4__15917_ gnd vdd FILL
XFILL_5__16167_ gnd vdd FILL
XFILL_2__15007_ gnd vdd FILL
X_9573_ _9507_/A _7790_/CLK _9566_/R vdd _9573_/D gnd vdd DFFSR
XSFILL3560x67050 gnd vdd FILL
XFILL_3__14558_ gnd vdd FILL
XFILL_5__13379_ gnd vdd FILL
XFILL_2__12219_ gnd vdd FILL
XFILL_1__15737_ gnd vdd FILL
XFILL_3__7955_ gnd vdd FILL
XFILL_0__14378_ gnd vdd FILL
XFILL_5_BUFX2_insert504 gnd vdd FILL
XFILL_5__15118_ gnd vdd FILL
XSFILL28760x79050 gnd vdd FILL
X_8524_ _8524_/A _8440_/B _8524_/C gnd _8524_/Y vdd OAI21X1
XFILL_3__13509_ gnd vdd FILL
XFILL_5_BUFX2_insert515 gnd vdd FILL
XSFILL114520x50050 gnd vdd FILL
XFILL_1__6970_ gnd vdd FILL
XFILL_5__16098_ gnd vdd FILL
XFILL_4__15848_ gnd vdd FILL
XFILL_3__6906_ gnd vdd FILL
XFILL_0__13329_ gnd vdd FILL
XFILL_3__14489_ gnd vdd FILL
XFILL_0__16117_ gnd vdd FILL
XFILL_5_BUFX2_insert526 gnd vdd FILL
XFILL_3__7886_ gnd vdd FILL
XFILL_1__15668_ gnd vdd FILL
XFILL_5_BUFX2_insert537 gnd vdd FILL
XFILL_0__9916_ gnd vdd FILL
XFILL_5_BUFX2_insert548 gnd vdd FILL
XFILL_5_BUFX2_insert559 gnd vdd FILL
XFILL_5__15049_ gnd vdd FILL
XSFILL84440x32050 gnd vdd FILL
XFILL_3__16228_ gnd vdd FILL
XFILL_3__9625_ gnd vdd FILL
X_8455_ _8455_/A _8494_/B _8455_/C gnd _8539_/D vdd OAI21X1
XFILL_3__6837_ gnd vdd FILL
XFILL_1__14619_ gnd vdd FILL
XFILL_4__15779_ gnd vdd FILL
XFILL_3_BUFX2_insert7 gnd vdd FILL
XFILL_0__16048_ gnd vdd FILL
XFILL_6__16339_ gnd vdd FILL
XFILL_1__15599_ gnd vdd FILL
XSFILL103560x74050 gnd vdd FILL
XFILL_1__8640_ gnd vdd FILL
X_7406_ _7406_/Q _7406_/CLK _9692_/R vdd _7360_/Y gnd vdd DFFSR
XFILL_0__9847_ gnd vdd FILL
X_8386_ _8372_/B _7490_/B gnd _8387_/C vdd NAND2X1
XFILL_3__16159_ gnd vdd FILL
XFILL_2__15909_ gnd vdd FILL
XFILL_3__9556_ gnd vdd FILL
XFILL111800x48050 gnd vdd FILL
XFILL_6__9265_ gnd vdd FILL
X_7337_ _7337_/A gnd _7337_/Y vdd INVX1
XFILL_3__8507_ gnd vdd FILL
XFILL_4__7300_ gnd vdd FILL
XFILL_3_BUFX2_insert70 gnd vdd FILL
XFILL_1__8571_ gnd vdd FILL
XFILL_0__9778_ gnd vdd FILL
XFILL_3_BUFX2_insert81 gnd vdd FILL
XFILL_3__9487_ gnd vdd FILL
XFILL_3_BUFX2_insert92 gnd vdd FILL
XFILL_6__8216_ gnd vdd FILL
XFILL112440x14050 gnd vdd FILL
XFILL_0__8729_ gnd vdd FILL
X_7268_ _7268_/Q _7268_/CLK _8688_/R vdd _7268_/D gnd vdd DFFSR
XSFILL38920x8050 gnd vdd FILL
XFILL_2_CLKBUF1_insert118 gnd vdd FILL
XFILL_4__7231_ gnd vdd FILL
XFILL_3__8438_ gnd vdd FILL
XFILL_2_CLKBUF1_insert129 gnd vdd FILL
X_9007_ _9065_/Q gnd _9009_/A vdd INVX1
XSFILL39000x16050 gnd vdd FILL
XFILL_1__7453_ gnd vdd FILL
X_7199_ _7197_/Y _7166_/B _7199_/C gnd _7199_/Y vdd OAI21X1
XFILL_3__8369_ gnd vdd FILL
XFILL_4__7162_ gnd vdd FILL
XSFILL3640x47050 gnd vdd FILL
XFILL_2_BUFX2_insert405 gnd vdd FILL
XFILL_2_BUFX2_insert416 gnd vdd FILL
XFILL_4__7093_ gnd vdd FILL
XSFILL28840x59050 gnd vdd FILL
XFILL_2_BUFX2_insert427 gnd vdd FILL
XFILL_1__9123_ gnd vdd FILL
XFILL_2_BUFX2_insert438 gnd vdd FILL
XSFILL94280x35050 gnd vdd FILL
XSFILL114600x30050 gnd vdd FILL
XFILL_2_BUFX2_insert449 gnd vdd FILL
X_11840_ _11839_/Y _11762_/B _11836_/Y gnd _11840_/Y vdd OAI21X1
X_9909_ _9963_/Q gnd _9909_/Y vdd INVX1
XSFILL69080x11050 gnd vdd FILL
XSFILL103640x54050 gnd vdd FILL
XSFILL69320x73050 gnd vdd FILL
XFILL_1__8005_ gnd vdd FILL
X_11771_ _11245_/Y _11770_/B _11771_/C gnd _11772_/C vdd OAI21X1
XFILL_4__9803_ gnd vdd FILL
X_13510_ _13509_/Y _14237_/B _13876_/C _13510_/D gnd _13510_/Y vdd OAI22X1
XFILL_4__7995_ gnd vdd FILL
X_10722_ _15566_/A _7778_/CLK _8418_/R vdd _10652_/Y gnd vdd DFFSR
XSFILL64120x3050 gnd vdd FILL
X_14490_ _14486_/Y _14489_/Y gnd _14490_/Y vdd NOR2X1
XSFILL104520x82050 gnd vdd FILL
XBUFX2_insert404 _10920_/Y gnd _12422_/A vdd BUFX2
XBUFX2_insert415 _15050_/Y gnd _16036_/A vdd BUFX2
XFILL_4__6946_ gnd vdd FILL
XBUFX2_insert426 _15047_/Y gnd _15774_/C vdd BUFX2
XFILL_4__9734_ gnd vdd FILL
X_13441_ _9558_/Q gnd _13441_/Y vdd INVX1
XBUFX2_insert437 _13326_/Y gnd _8759_/B vdd BUFX2
XFILL_6_BUFX2_insert382 gnd vdd FILL
XSFILL8760x80050 gnd vdd FILL
X_10653_ _15590_/A gnd _10655_/A vdd INVX1
XFILL_6_BUFX2_insert393 gnd vdd FILL
XBUFX2_insert448 _13276_/Y gnd _7250_/B vdd BUFX2
XBUFX2_insert459 _13442_/Y gnd _14718_/B vdd BUFX2
XFILL_4__9665_ gnd vdd FILL
XFILL_4__6877_ gnd vdd FILL
X_16160_ _16247_/C _16160_/B _14760_/A _16314_/D gnd _16160_/Y vdd OAI22X1
X_13372_ _13372_/A _13398_/A _13423_/B gnd _13372_/Y vdd NAND3X1
XFILL_1__8907_ gnd vdd FILL
XFILL_2__7700_ gnd vdd FILL
X_10584_ _13552_/A _8152_/CLK _9944_/R vdd _10584_/D gnd vdd DFFSR
XFILL_4__8616_ gnd vdd FILL
XSFILL3720x27050 gnd vdd FILL
XFILL_1__9887_ gnd vdd FILL
X_15111_ _15544_/A _13524_/Y _13520_/Y _15756_/D gnd _15111_/Y vdd OAI22X1
X_12323_ _12327_/A gnd _12319_/C gnd _12326_/A vdd NAND3X1
XFILL_4__9596_ gnd vdd FILL
X_16091_ _9200_/Q gnd _16091_/Y vdd INVX1
XFILL_2__7631_ gnd vdd FILL
XFILL_1__8838_ gnd vdd FILL
XSFILL28920x39050 gnd vdd FILL
XFILL_5__7340_ gnd vdd FILL
XSFILL94360x15050 gnd vdd FILL
X_15042_ _15187_/A _13416_/Y _15187_/C gnd _15076_/A vdd NOR3X1
X_12254_ _12254_/A _12254_/B _12253_/Y gnd _12254_/Y vdd NAND3X1
XSFILL13720x81050 gnd vdd FILL
XFILL_2__7562_ gnd vdd FILL
XFILL_3__10170_ gnd vdd FILL
XFILL_1__8769_ gnd vdd FILL
XSFILL79160x76050 gnd vdd FILL
XFILL_4__8478_ gnd vdd FILL
X_11205_ _11204_/Y gnd _11334_/A vdd INVX2
XSFILL29000x48050 gnd vdd FILL
XFILL_2__9301_ gnd vdd FILL
XFILL_1__10300_ gnd vdd FILL
X_12185_ _12179_/A _12942_/Q gnd _12186_/C vdd NAND2X1
XFILL_4__11460_ gnd vdd FILL
XFILL_5__9010_ gnd vdd FILL
XFILL_2__7493_ gnd vdd FILL
XFILL_1__11280_ gnd vdd FILL
XFILL_4__7429_ gnd vdd FILL
XSFILL109400x3050 gnd vdd FILL
XFILL_4__10411_ gnd vdd FILL
X_11136_ _12282_/Y gnd _11617_/B vdd INVX1
XFILL_2__9232_ gnd vdd FILL
XFILL_5__12750_ gnd vdd FILL
XFILL_1__10231_ gnd vdd FILL
XSFILL8440x39050 gnd vdd FILL
XFILL_4__11391_ gnd vdd FILL
XFILL_2__12570_ gnd vdd FILL
XFILL_3_BUFX2_insert250 gnd vdd FILL
XFILL_0__10961_ gnd vdd FILL
XFILL_3_BUFX2_insert261 gnd vdd FILL
XSFILL84280x67050 gnd vdd FILL
XFILL_4__13130_ gnd vdd FILL
XFILL_5__11701_ gnd vdd FILL
XFILL_3_BUFX2_insert272 gnd vdd FILL
X_15944_ _15708_/A _14513_/Y _15708_/C gnd _15967_/B vdd NOR3X1
X_11067_ _11065_/Y _11066_/Y _11062_/Y gnd _11067_/Y vdd OAI21X1
XFILL_3__13860_ gnd vdd FILL
XFILL_2__9163_ gnd vdd FILL
XFILL_3_BUFX2_insert283 gnd vdd FILL
XFILL_2__11521_ gnd vdd FILL
XFILL_0__12700_ gnd vdd FILL
XFILL_3_BUFX2_insert294 gnd vdd FILL
XFILL_1__10162_ gnd vdd FILL
XFILL_0__13680_ gnd vdd FILL
X_10018_ _10018_/A _9996_/A _10017_/Y gnd _10084_/D vdd OAI21X1
XFILL_0__10892_ gnd vdd FILL
XFILL_5__14420_ gnd vdd FILL
XFILL_2__8114_ gnd vdd FILL
XFILL_5__11632_ gnd vdd FILL
XFILL_6__13971_ gnd vdd FILL
X_15875_ _15874_/Y _15239_/B _15524_/A _15875_/D gnd _15875_/Y vdd OAI22X1
XFILL_2__14240_ gnd vdd FILL
XFILL_4__10273_ gnd vdd FILL
XFILL_0__12631_ gnd vdd FILL
XFILL_3__13791_ gnd vdd FILL
XFILL_2_BUFX2_insert950 gnd vdd FILL
XFILL_2__11452_ gnd vdd FILL
XFILL_2__9094_ gnd vdd FILL
XFILL_6__15710_ gnd vdd FILL
XFILL_5__9912_ gnd vdd FILL
XFILL_1__14970_ gnd vdd FILL
X_14826_ _7370_/A gnd _14826_/Y vdd INVX1
XFILL_4__12012_ gnd vdd FILL
XFILL_2_BUFX2_insert961 gnd vdd FILL
XFILL_2_BUFX2_insert972 gnd vdd FILL
XFILL_3__15530_ gnd vdd FILL
XFILL_5__14351_ gnd vdd FILL
XFILL_5__11563_ gnd vdd FILL
XFILL_2_BUFX2_insert983 gnd vdd FILL
XFILL_2__10403_ gnd vdd FILL
XFILL_3__12742_ gnd vdd FILL
XFILL_2_BUFX2_insert994 gnd vdd FILL
XFILL_2__14171_ gnd vdd FILL
XFILL_1__13921_ gnd vdd FILL
XFILL_0__15350_ gnd vdd FILL
XFILL112280x49050 gnd vdd FILL
XFILL_2__11383_ gnd vdd FILL
XFILL_5__13302_ gnd vdd FILL
XFILL_5__10514_ gnd vdd FILL
X_14757_ _14757_/A _13879_/B _13479_/C _14756_/Y gnd _14757_/Y vdd OAI22X1
XFILL_0__7060_ gnd vdd FILL
XFILL_2__13122_ gnd vdd FILL
X_11969_ _11969_/A _11969_/B gnd _11970_/C vdd NAND2X1
XFILL_5__11494_ gnd vdd FILL
XFILL_3__15461_ gnd vdd FILL
XFILL_5__14282_ gnd vdd FILL
XFILL_0__14301_ gnd vdd FILL
XFILL_0__11513_ gnd vdd FILL
XFILL_1__13852_ gnd vdd FILL
XFILL_0__15281_ gnd vdd FILL
XFILL_5__16021_ gnd vdd FILL
XFILL_0__12493_ gnd vdd FILL
XSFILL99160x1050 gnd vdd FILL
X_13708_ _13708_/A _14068_/C _14342_/B _13708_/D gnd _13712_/B vdd OAI22X1
XFILL_6__11804_ gnd vdd FILL
XFILL_5__13233_ gnd vdd FILL
XFILL_5__10445_ gnd vdd FILL
XFILL_5__6986_ gnd vdd FILL
XSFILL13800x61050 gnd vdd FILL
XFILL_6__15572_ gnd vdd FILL
XFILL_5__9774_ gnd vdd FILL
XFILL_3__14412_ gnd vdd FILL
XFILL_6__12784_ gnd vdd FILL
XFILL_3__11624_ gnd vdd FILL
X_14688_ _16071_/A _14358_/B _14739_/C _16072_/A gnd _14690_/A vdd AOI22X1
XFILL_0__14232_ gnd vdd FILL
XFILL_3__15392_ gnd vdd FILL
XSFILL79240x56050 gnd vdd FILL
XFILL_2__10265_ gnd vdd FILL
XFILL_4__13963_ gnd vdd FILL
XFILL_2__9996_ gnd vdd FILL
XFILL_0__11444_ gnd vdd FILL
XFILL_1__13783_ gnd vdd FILL
XFILL_6__14523_ gnd vdd FILL
XFILL_5__8725_ gnd vdd FILL
XFILL_4__15702_ gnd vdd FILL
X_13639_ _9562_/Q gnd _13640_/D vdd INVX1
XFILL_5__13164_ gnd vdd FILL
X_16427_ _15482_/A _7535_/CLK _7648_/R vdd _16353_/Y gnd vdd DFFSR
XFILL_1__10995_ gnd vdd FILL
XFILL_5__10376_ gnd vdd FILL
XFILL_2__12004_ gnd vdd FILL
XFILL_3__14343_ gnd vdd FILL
XFILL_4__12914_ gnd vdd FILL
XFILL_3__7740_ gnd vdd FILL
XFILL_1__15522_ gnd vdd FILL
XFILL_3__11555_ gnd vdd FILL
XFILL_1__12734_ gnd vdd FILL
XFILL_0__14163_ gnd vdd FILL
XFILL_2__10196_ gnd vdd FILL
XFILL_4__13894_ gnd vdd FILL
XBUFX2_insert960 _13361_/Y gnd _10363_/B vdd BUFX2
XFILL_5__8656_ gnd vdd FILL
XSFILL8520x19050 gnd vdd FILL
XFILL_0__11375_ gnd vdd FILL
XFILL_5__12115_ gnd vdd FILL
XBUFX2_insert971 _16451_/Y gnd _13149_/A vdd BUFX2
X_16358_ gnd gnd gnd _16358_/Y vdd NAND2X1
XFILL_3__10506_ gnd vdd FILL
XFILL_4__15633_ gnd vdd FILL
XBUFX2_insert982 _13455_/Y gnd _14496_/A vdd BUFX2
XFILL_0__7962_ gnd vdd FILL
XFILL_5__13095_ gnd vdd FILL
XFILL_6__11666_ gnd vdd FILL
XFILL_4__12845_ gnd vdd FILL
XFILL_0__13114_ gnd vdd FILL
XFILL_3__14274_ gnd vdd FILL
XBUFX2_insert993 _12408_/Y gnd _9782_/B vdd BUFX2
XFILL_3__7671_ gnd vdd FILL
XSFILL84360x47050 gnd vdd FILL
XFILL_2__8878_ gnd vdd FILL
XFILL_3__11486_ gnd vdd FILL
XFILL_1__15453_ gnd vdd FILL
XFILL_5__7607_ gnd vdd FILL
X_15309_ _15309_/A _15305_/Y _15309_/C gnd _15310_/A vdd NAND3X1
XSFILL13560x5050 gnd vdd FILL
XFILL_0__14094_ gnd vdd FILL
XFILL_0__6913_ gnd vdd FILL
XFILL_5__8587_ gnd vdd FILL
XFILL_3__16013_ gnd vdd FILL
XFILL_5__12046_ gnd vdd FILL
X_8240_ _8216_/A _8624_/B gnd _8241_/C vdd NAND2X1
XSFILL48920x3050 gnd vdd FILL
XFILL_3__13225_ gnd vdd FILL
X_16289_ _16014_/C _8275_/A _8659_/A _16212_/A gnd _16289_/Y vdd AOI22X1
XFILL_6__14385_ gnd vdd FILL
XFILL_3__9410_ gnd vdd FILL
XFILL_4__12776_ gnd vdd FILL
XFILL_3__10437_ gnd vdd FILL
XFILL_4__15564_ gnd vdd FILL
XFILL_0__7893_ gnd vdd FILL
XFILL_2__7829_ gnd vdd FILL
XFILL_1__14404_ gnd vdd FILL
XFILL_0__13045_ gnd vdd FILL
XFILL_1__11616_ gnd vdd FILL
XFILL_2__13955_ gnd vdd FILL
XSFILL99400x69050 gnd vdd FILL
XFILL_1__15384_ gnd vdd FILL
XFILL_0__10257_ gnd vdd FILL
XFILL_6__13336_ gnd vdd FILL
XFILL_1__12596_ gnd vdd FILL
XFILL_0__9632_ gnd vdd FILL
X_8171_ _8171_/Q _8171_/CLK _8171_/R vdd _8171_/D gnd vdd DFFSR
XFILL_0__6844_ gnd vdd FILL
XFILL_4__14515_ gnd vdd FILL
XFILL_6__10548_ gnd vdd FILL
XFILL_3__13156_ gnd vdd FILL
XFILL_2__12906_ gnd vdd FILL
XFILL_4__11727_ gnd vdd FILL
XFILL_3__9341_ gnd vdd FILL
XFILL_3__10368_ gnd vdd FILL
XFILL_1__14335_ gnd vdd FILL
XFILL_4__15495_ gnd vdd FILL
XFILL_2__13886_ gnd vdd FILL
XFILL_1__11547_ gnd vdd FILL
XFILL_0__10188_ gnd vdd FILL
XFILL_5__15805_ gnd vdd FILL
XFILL_5__7469_ gnd vdd FILL
X_7122_ _7122_/A _7064_/A _7122_/C gnd _7156_/D vdd OAI21X1
XFILL111880x22050 gnd vdd FILL
XFILL_3__12107_ gnd vdd FILL
XFILL_2__15625_ gnd vdd FILL
XFILL112360x29050 gnd vdd FILL
XFILL_4__11658_ gnd vdd FILL
XFILL_4__14446_ gnd vdd FILL
XFILL_2__12837_ gnd vdd FILL
XFILL_3__13087_ gnd vdd FILL
XFILL_3__9272_ gnd vdd FILL
XFILL_5__13997_ gnd vdd FILL
XFILL_3__10299_ gnd vdd FILL
XFILL_5__9208_ gnd vdd FILL
XFILL_1__11478_ gnd vdd FILL
XFILL_1__14266_ gnd vdd FILL
XFILL_6__12218_ gnd vdd FILL
XFILL_0__8514_ gnd vdd FILL
X_7053_ _7051_/Y _7095_/B _7053_/C gnd _7133_/D vdd OAI21X1
XFILL_0__14996_ gnd vdd FILL
XFILL_5__15736_ gnd vdd FILL
XFILL_1__16005_ gnd vdd FILL
XFILL_3__12038_ gnd vdd FILL
XFILL_0__9494_ gnd vdd FILL
XFILL_3__8223_ gnd vdd FILL
XFILL_1__13217_ gnd vdd FILL
XFILL_2__15556_ gnd vdd FILL
XFILL_4__14377_ gnd vdd FILL
XFILL_4__11589_ gnd vdd FILL
XFILL_1__10429_ gnd vdd FILL
XFILL_2__12768_ gnd vdd FILL
XFILL_5__9139_ gnd vdd FILL
XFILL_1__14197_ gnd vdd FILL
XFILL_0__13947_ gnd vdd FILL
XSFILL49080x75050 gnd vdd FILL
XFILL_4__16116_ gnd vdd FILL
XFILL_0__8445_ gnd vdd FILL
XFILL_4__13328_ gnd vdd FILL
XFILL_5__15667_ gnd vdd FILL
XFILL_2__14507_ gnd vdd FILL
XFILL_5__12879_ gnd vdd FILL
XFILL_2__11719_ gnd vdd FILL
XFILL_1__13148_ gnd vdd FILL
XFILL_2__15487_ gnd vdd FILL
XFILL_2__12699_ gnd vdd FILL
XFILL_0__13878_ gnd vdd FILL
XFILL_5__14618_ gnd vdd FILL
XFILL_4__13259_ gnd vdd FILL
XFILL_0__8376_ gnd vdd FILL
XFILL_3__7105_ gnd vdd FILL
XSFILL109560x9050 gnd vdd FILL
XFILL_4__16047_ gnd vdd FILL
XSFILL114520x45050 gnd vdd FILL
XFILL_5__15598_ gnd vdd FILL
XFILL_2__14438_ gnd vdd FILL
XFILL_0__15617_ gnd vdd FILL
XFILL_3__8085_ gnd vdd FILL
XFILL_1__13079_ gnd vdd FILL
XFILL_3__13989_ gnd vdd FILL
XFILL_6__8903_ gnd vdd FILL
XFILL_0__12829_ gnd vdd FILL
XFILL_0__7327_ gnd vdd FILL
XFILL_5__14549_ gnd vdd FILL
XFILL_3__15728_ gnd vdd FILL
XFILL_3__7036_ gnd vdd FILL
X_7955_ _7955_/A _7955_/B _7954_/Y gnd _8031_/D vdd OAI21X1
XFILL_2__14369_ gnd vdd FILL
XFILL_0__15548_ gnd vdd FILL
XFILL_2__16108_ gnd vdd FILL
X_6906_ _6955_/B _6906_/B gnd _6907_/C vdd NAND2X1
X_7886_ _7887_/B _8014_/B gnd _7887_/C vdd NAND2X1
XFILL_3__15659_ gnd vdd FILL
XFILL_5__16219_ gnd vdd FILL
XFILL_0__15479_ gnd vdd FILL
X_9625_ _9623_/Y _9625_/B _9625_/C gnd _9697_/D vdd OAI21X1
X_6837_ _6837_/A gnd MemWrite vdd BUFX2
XFILL_2__16039_ gnd vdd FILL
XFILL_0__7189_ gnd vdd FILL
XFILL_3__8987_ gnd vdd FILL
XFILL_1__9810_ gnd vdd FILL
XFILL_5_BUFX2_insert301 gnd vdd FILL
X_9556_ _9466_/A _9556_/B gnd _9557_/C vdd NAND2X1
XFILL_3__7938_ gnd vdd FILL
XFILL_5_BUFX2_insert312 gnd vdd FILL
XFILL_5_BUFX2_insert323 gnd vdd FILL
XSFILL89160x39050 gnd vdd FILL
XFILL_5_BUFX2_insert334 gnd vdd FILL
XBUFX2_insert13 _14989_/Y gnd _16099_/C vdd BUFX2
X_8507_ _8507_/A gnd _8507_/Y vdd INVX1
XFILL_1__9741_ gnd vdd FILL
XFILL112040x11050 gnd vdd FILL
XBUFX2_insert24 _11344_/Y gnd _11571_/A vdd BUFX2
XFILL_5_BUFX2_insert345 gnd vdd FILL
XFILL_1__6953_ gnd vdd FILL
X_9487_ _9548_/B _9487_/B gnd _9488_/C vdd NAND2X1
XBUFX2_insert35 _13265_/Y gnd _6988_/B vdd BUFX2
XFILL_5_BUFX2_insert356 gnd vdd FILL
XFILL_3__7869_ gnd vdd FILL
XBUFX2_insert46 _14986_/Y gnd _15677_/A vdd BUFX2
XFILL_5_BUFX2_insert367 gnd vdd FILL
XBUFX2_insert57 _13309_/Y gnd _8079_/A vdd BUFX2
XFILL_5_BUFX2_insert378 gnd vdd FILL
XBUFX2_insert68 _13393_/Y gnd _14317_/C vdd BUFX2
XFILL_5_BUFX2_insert389 gnd vdd FILL
X_8438_ _8438_/A gnd _8438_/Y vdd INVX1
XFILL_1__9672_ gnd vdd FILL
XFILL_4__8401_ gnd vdd FILL
XFILL_3__9608_ gnd vdd FILL
XBUFX2_insert79 _15015_/Y gnd _15407_/C vdd BUFX2
XFILL_1__6884_ gnd vdd FILL
XFILL_4__9381_ gnd vdd FILL
XFILL_1__8623_ gnd vdd FILL
XSFILL114600x25050 gnd vdd FILL
XFILL_4__8332_ gnd vdd FILL
X_8369_ _8369_/A _8345_/B _8369_/C gnd _8369_/Y vdd OAI21X1
XFILL_3__9539_ gnd vdd FILL
XFILL_4__8263_ gnd vdd FILL
XFILL_1__7505_ gnd vdd FILL
XFILL_1__8485_ gnd vdd FILL
XFILL_4__7214_ gnd vdd FILL
XFILL_4__8194_ gnd vdd FILL
XFILL_1__7436_ gnd vdd FILL
X_13990_ _9623_/A gnd _13990_/Y vdd INVX1
X_12941_ _12889_/A _7532_/CLK _8816_/R vdd _12941_/D gnd vdd DFFSR
XSFILL8760x75050 gnd vdd FILL
XSFILL23800x24050 gnd vdd FILL
XFILL_1__7367_ gnd vdd FILL
XFILL_2_BUFX2_insert235 gnd vdd FILL
XFILL_2_BUFX2_insert246 gnd vdd FILL
XSFILL89240x19050 gnd vdd FILL
XFILL_4__7076_ gnd vdd FILL
XFILL_2_BUFX2_insert257 gnd vdd FILL
X_15660_ _15660_/A _15659_/Y _15658_/Y gnd _15660_/Y vdd NAND3X1
XFILL_1__9106_ gnd vdd FILL
XFILL_2_BUFX2_insert268 gnd vdd FILL
X_12872_ vdd _12872_/B gnd _12873_/C vdd NAND2X1
XFILL_2_BUFX2_insert279 gnd vdd FILL
XFILL_1__7298_ gnd vdd FILL
X_14611_ _10430_/A gnd _14611_/Y vdd INVX1
XFILL_1_BUFX2_insert902 gnd vdd FILL
XFILL_1_BUFX2_insert913 gnd vdd FILL
X_11823_ _11821_/Y _11809_/C _11822_/Y gnd _11829_/A vdd AOI21X1
XFILL_1__9037_ gnd vdd FILL
XFILL_1_BUFX2_insert924 gnd vdd FILL
X_15591_ _7011_/Q gnd _15591_/Y vdd INVX1
XFILL_1_BUFX2_insert935 gnd vdd FILL
XFILL_1_BUFX2_insert946 gnd vdd FILL
XFILL_5__6840_ gnd vdd FILL
X_14542_ _14540_/Y _13836_/B _13467_/A _14541_/Y gnd _14546_/A vdd OAI22X1
XFILL_1_BUFX2_insert957 gnd vdd FILL
XFILL_1_BUFX2_insert968 gnd vdd FILL
X_11754_ _11754_/A gnd _12021_/A vdd INVX1
XSFILL74280x4050 gnd vdd FILL
XFILL_1_BUFX2_insert979 gnd vdd FILL
XFILL_2__9850_ gnd vdd FILL
XSFILL113880x4050 gnd vdd FILL
XSFILL13720x76050 gnd vdd FILL
XSFILL54360x26050 gnd vdd FILL
XFILL_5__10230_ gnd vdd FILL
X_10705_ _10676_/B _8273_/B gnd _10705_/Y vdd NAND2X1
XFILL_4__7978_ gnd vdd FILL
X_14473_ _14473_/A _14473_/B gnd _14500_/B vdd NOR2X1
XSFILL94760x31050 gnd vdd FILL
XFILL_4__10960_ gnd vdd FILL
XBUFX2_insert234 _12348_/Y gnd _8314_/B vdd BUFX2
XFILL_2__10050_ gnd vdd FILL
X_11685_ _12266_/Y _11064_/Y _11045_/Y gnd _11686_/A vdd OAI21X1
XFILL_2__9781_ gnd vdd FILL
XFILL_5__8510_ gnd vdd FILL
XBUFX2_insert245 _13460_/Y gnd _13795_/B vdd BUFX2
XSFILL68920x41050 gnd vdd FILL
XSFILL103720x29050 gnd vdd FILL
X_16212_ _16212_/A _8653_/A _9677_/A _15652_/D gnd _16219_/B vdd AOI22X1
XFILL_1__10780_ gnd vdd FILL
XBUFX2_insert256 _12423_/Y gnd _9797_/B vdd BUFX2
XFILL_2__6993_ gnd vdd FILL
XSFILL94200x74050 gnd vdd FILL
X_13424_ _13381_/A _13381_/B _13418_/A gnd _13424_/Y vdd NAND3X1
XFILL_4__6929_ gnd vdd FILL
XFILL_5__9490_ gnd vdd FILL
X_10636_ _10678_/A _9100_/B gnd _10637_/C vdd NAND2X1
XBUFX2_insert267 _15024_/Y gnd _15410_/D vdd BUFX2
XFILL_5__10161_ gnd vdd FILL
XBUFX2_insert278 _13419_/Y gnd _14479_/B vdd BUFX2
XFILL_2__8732_ gnd vdd FILL
XFILL_3__11340_ gnd vdd FILL
XBUFX2_insert289 _15059_/Y gnd _16099_/B vdd BUFX2
XFILL_4__10891_ gnd vdd FILL
XFILL_1__9939_ gnd vdd FILL
XFILL_5_CLKBUF1_insert113 gnd vdd FILL
XFILL_5_CLKBUF1_insert124 gnd vdd FILL
XFILL_0__11160_ gnd vdd FILL
XFILL_5__8441_ gnd vdd FILL
XFILL_4__9648_ gnd vdd FILL
XFILL_5_CLKBUF1_insert135 gnd vdd FILL
X_16143_ _15760_/A _14743_/Y _16143_/C gnd _16147_/A vdd OAI21X1
XFILL_4__12630_ gnd vdd FILL
X_13355_ _13225_/D _13220_/A _13219_/B gnd _13355_/Y vdd OAI21X1
XFILL_5_CLKBUF1_insert146 gnd vdd FILL
XFILL_6__11451_ gnd vdd FILL
XSFILL104600x57050 gnd vdd FILL
X_10567_ _14763_/B gnd _10569_/A vdd INVX1
XFILL_5_CLKBUF1_insert157 gnd vdd FILL
XFILL_0__10111_ gnd vdd FILL
XFILL_3__11271_ gnd vdd FILL
XFILL_5_CLKBUF1_insert168 gnd vdd FILL
XFILL_5_BUFX2_insert890 gnd vdd FILL
XFILL_1__12450_ gnd vdd FILL
XFILL_5_CLKBUF1_insert179 gnd vdd FILL
XSFILL74520x39050 gnd vdd FILL
X_12306_ _12306_/A _12306_/B _12306_/C gnd _12306_/Y vdd NAND3X1
XFILL_0__11091_ gnd vdd FILL
XFILL_5__8372_ gnd vdd FILL
XSFILL98840x77050 gnd vdd FILL
XFILL_6__14170_ gnd vdd FILL
XFILL_3__13010_ gnd vdd FILL
X_16074_ _14689_/B _15916_/B _16074_/C gnd _16075_/B vdd AOI21X1
XFILL_5__13920_ gnd vdd FILL
X_13286_ _13297_/A _13286_/B gnd _13287_/B vdd OR2X2
XFILL_2__7614_ gnd vdd FILL
X_10498_ _13682_/B gnd _10500_/A vdd INVX1
XFILL_2__13740_ gnd vdd FILL
XFILL_1__11401_ gnd vdd FILL
XFILL_2__10952_ gnd vdd FILL
XFILL_1__12381_ gnd vdd FILL
XFILL_5__7323_ gnd vdd FILL
XFILL_0__10042_ gnd vdd FILL
XFILL_2__8594_ gnd vdd FILL
X_15025_ _13395_/Y _15025_/B _16018_/C _13469_/Y gnd _15025_/Y vdd OAI22X1
X_12237_ _6875_/A _12237_/B _12269_/C _12704_/A gnd _12237_/Y vdd AOI22X1
XFILL_4__14300_ gnd vdd FILL
XFILL_4__11512_ gnd vdd FILL
XFILL_5__13851_ gnd vdd FILL
XSFILL74120x41050 gnd vdd FILL
XFILL_4__15280_ gnd vdd FILL
XFILL_4__12492_ gnd vdd FILL
XFILL_3__10153_ gnd vdd FILL
XFILL_2__7545_ gnd vdd FILL
XFILL_1__14120_ gnd vdd FILL
XFILL_1__11332_ gnd vdd FILL
XFILL_2__13671_ gnd vdd FILL
XFILL_0__14850_ gnd vdd FILL
XFILL_2__10883_ gnd vdd FILL
XFILL_2__15410_ gnd vdd FILL
XFILL_4__14231_ gnd vdd FILL
XFILL_6__10264_ gnd vdd FILL
X_12168_ _12168_/A _12117_/B _12168_/C gnd _12168_/Y vdd OAI21X1
XFILL_4__11443_ gnd vdd FILL
XFILL_2__12622_ gnd vdd FILL
XFILL_5__13782_ gnd vdd FILL
XFILL_2__16390_ gnd vdd FILL
XFILL_0__13801_ gnd vdd FILL
XSFILL108840x62050 gnd vdd FILL
XFILL_1__14051_ gnd vdd FILL
XFILL_3__14961_ gnd vdd FILL
XFILL_1__11263_ gnd vdd FILL
XFILL_2__7476_ gnd vdd FILL
XFILL_5__10994_ gnd vdd FILL
XFILL_5__15521_ gnd vdd FILL
XFILL_0__11993_ gnd vdd FILL
X_11119_ _11118_/Y _11143_/A gnd _11141_/A vdd AND2X2
XFILL_5__7185_ gnd vdd FILL
XFILL_0__14781_ gnd vdd FILL
XFILL_2__9215_ gnd vdd FILL
XFILL_5__12733_ gnd vdd FILL
XSFILL13800x56050 gnd vdd FILL
XFILL_4__14162_ gnd vdd FILL
XFILL_2__15341_ gnd vdd FILL
X_12099_ _12047_/A _12427_/A _12011_/C gnd _12102_/A vdd NAND3X1
XFILL_3__13912_ gnd vdd FILL
XFILL_4__11374_ gnd vdd FILL
XFILL_1__13002_ gnd vdd FILL
XFILL_3__14892_ gnd vdd FILL
XFILL_0__10944_ gnd vdd FILL
XFILL_0__13732_ gnd vdd FILL
XFILL_1__11194_ gnd vdd FILL
XFILL_0__8230_ gnd vdd FILL
XFILL_4__13113_ gnd vdd FILL
X_15927_ _15923_/Y _15927_/B _15927_/C gnd _15928_/B vdd NAND3X1
XFILL_5__15452_ gnd vdd FILL
XFILL_4__10325_ gnd vdd FILL
XFILL_2__9146_ gnd vdd FILL
XFILL_4__14093_ gnd vdd FILL
XFILL_2__11504_ gnd vdd FILL
XFILL_3__13843_ gnd vdd FILL
XFILL_1__10145_ gnd vdd FILL
XFILL_2__15272_ gnd vdd FILL
XFILL_0__16451_ gnd vdd FILL
XFILL_2__12484_ gnd vdd FILL
XFILL_0__13663_ gnd vdd FILL
XFILL_0__10875_ gnd vdd FILL
XFILL_5__14403_ gnd vdd FILL
XFILL_4__13044_ gnd vdd FILL
XFILL_5__11615_ gnd vdd FILL
XFILL_4__10256_ gnd vdd FILL
XFILL_5__15383_ gnd vdd FILL
XFILL_2__14223_ gnd vdd FILL
X_15858_ _7914_/Q _16204_/B gnd _15860_/A vdd NAND2X1
XFILL_3__13774_ gnd vdd FILL
XFILL_0__15402_ gnd vdd FILL
XFILL_5__12595_ gnd vdd FILL
XFILL_2__11435_ gnd vdd FILL
XFILL_0__12614_ gnd vdd FILL
XFILL_2_BUFX2_insert780 gnd vdd FILL
XFILL_1__14953_ gnd vdd FILL
XFILL_0__16382_ gnd vdd FILL
XFILL_0__13594_ gnd vdd FILL
XFILL_0__7112_ gnd vdd FILL
XFILL_2_BUFX2_insert791 gnd vdd FILL
X_14809_ _13871_/A _14809_/B _13850_/B _14808_/Y gnd _14810_/B vdd OAI22X1
XFILL_5__14334_ gnd vdd FILL
XFILL_0__8092_ gnd vdd FILL
X_7740_ _7744_/B _9788_/B gnd _7741_/C vdd NAND2X1
XFILL_3__12725_ gnd vdd FILL
XSFILL43880x51050 gnd vdd FILL
XFILL_3__15513_ gnd vdd FILL
XFILL_5__11546_ gnd vdd FILL
XFILL_3__8910_ gnd vdd FILL
XFILL_4__10187_ gnd vdd FILL
XFILL_2__14154_ gnd vdd FILL
X_15789_ _7400_/Q _15789_/B _15794_/B gnd _15789_/Y vdd NAND3X1
XFILL_1__13904_ gnd vdd FILL
XFILL_0__15333_ gnd vdd FILL
XFILL_3__9890_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1075 gnd vdd FILL
XFILL_2__11366_ gnd vdd FILL
XSFILL59160x18050 gnd vdd FILL
XFILL_1__14884_ gnd vdd FILL
XFILL_0__7043_ gnd vdd FILL
XFILL_6__12836_ gnd vdd FILL
XFILL_5__14265_ gnd vdd FILL
XFILL_2__13105_ gnd vdd FILL
XFILL_3__12656_ gnd vdd FILL
XFILL_3__8841_ gnd vdd FILL
XFILL_2__10317_ gnd vdd FILL
X_7671_ _8823_/A _7690_/B gnd _7672_/C vdd NAND2X1
XFILL_5__11477_ gnd vdd FILL
XFILL_3__15444_ gnd vdd FILL
XFILL_1__13835_ gnd vdd FILL
XFILL_4__14995_ gnd vdd FILL
XFILL_2__14085_ gnd vdd FILL
XFILL_5__16004_ gnd vdd FILL
XFILL_0__12476_ gnd vdd FILL
XFILL_2__11297_ gnd vdd FILL
XFILL_0__15264_ gnd vdd FILL
XSFILL74200x21050 gnd vdd FILL
XFILL_5__13216_ gnd vdd FILL
XFILL_5__9757_ gnd vdd FILL
X_9410_ _9425_/A _9282_/B gnd _9411_/C vdd NAND2X1
XFILL_5__10428_ gnd vdd FILL
XFILL_5__6969_ gnd vdd FILL
XFILL_3__11607_ gnd vdd FILL
XFILL_3__15375_ gnd vdd FILL
XFILL_5__14196_ gnd vdd FILL
XFILL_2__13036_ gnd vdd FILL
XFILL_4__13946_ gnd vdd FILL
XFILL_2__10248_ gnd vdd FILL
XFILL_3__12587_ gnd vdd FILL
XFILL_0__14215_ gnd vdd FILL
XFILL_3__8772_ gnd vdd FILL
XFILL_0__11427_ gnd vdd FILL
XFILL_5__8708_ gnd vdd FILL
XFILL_1__13766_ gnd vdd FILL
XFILL_2__9979_ gnd vdd FILL
XSFILL59000x82050 gnd vdd FILL
XFILL_1__10978_ gnd vdd FILL
XFILL_0__15195_ gnd vdd FILL
XFILL_5__10359_ gnd vdd FILL
XFILL_5__13147_ gnd vdd FILL
XFILL_3__14326_ gnd vdd FILL
X_9341_ _9339_/B _8701_/B gnd _9341_/Y vdd NAND2X1
XFILL_0__8994_ gnd vdd FILL
XFILL_1__15505_ gnd vdd FILL
XFILL_3__11538_ gnd vdd FILL
XFILL_3__7723_ gnd vdd FILL
XFILL_1__12717_ gnd vdd FILL
XFILL_4__13877_ gnd vdd FILL
XSFILL109400x49050 gnd vdd FILL
XFILL_0__14146_ gnd vdd FILL
XFILL_2__10179_ gnd vdd FILL
XFILL_0__11358_ gnd vdd FILL
XBUFX2_insert790 _15052_/Y gnd _16155_/D vdd BUFX2
XFILL_5__8639_ gnd vdd FILL
XFILL_1__13697_ gnd vdd FILL
XFILL_0__7945_ gnd vdd FILL
XFILL_4__15616_ gnd vdd FILL
XFILL_3__14257_ gnd vdd FILL
X_9272_ _9272_/A gnd _9272_/Y vdd INVX1
XFILL_4__12828_ gnd vdd FILL
XFILL_4_BUFX2_insert308 gnd vdd FILL
XFILL_0__10309_ gnd vdd FILL
XFILL_1__15436_ gnd vdd FILL
XFILL_3__11469_ gnd vdd FILL
XFILL_1__12648_ gnd vdd FILL
XFILL_2__14987_ gnd vdd FILL
XFILL_4_BUFX2_insert319 gnd vdd FILL
XFILL_0__14077_ gnd vdd FILL
XFILL_0__11289_ gnd vdd FILL
XFILL_6__7363_ gnd vdd FILL
XFILL_3__13208_ gnd vdd FILL
XSFILL64120x73050 gnd vdd FILL
XFILL_5__12029_ gnd vdd FILL
X_8223_ _8223_/A _8244_/B _8222_/Y gnd _8223_/Y vdd OAI21X1
XFILL_4__15547_ gnd vdd FILL
XFILL_0__7876_ gnd vdd FILL
XFILL_4__12759_ gnd vdd FILL
XFILL_3__14188_ gnd vdd FILL
XFILL_2__13938_ gnd vdd FILL
XFILL_0__13028_ gnd vdd FILL
XFILL_1__15367_ gnd vdd FILL
XFILL_3__7585_ gnd vdd FILL
XFILL_0__9615_ gnd vdd FILL
XFILL_1__12579_ gnd vdd FILL
X_8154_ _8066_/A _8541_/CLK _8285_/R vdd _8068_/Y gnd vdd DFFSR
XFILL_3__13139_ gnd vdd FILL
XFILL_1__14318_ gnd vdd FILL
XFILL_4__15478_ gnd vdd FILL
XFILL_2__13869_ gnd vdd FILL
XFILL_6__16038_ gnd vdd FILL
XFILL_1__15298_ gnd vdd FILL
XSFILL43960x31050 gnd vdd FILL
XFILL_0__9546_ gnd vdd FILL
X_7105_ _7105_/A gnd _7105_/Y vdd INVX1
XSFILL3560x80050 gnd vdd FILL
X_8085_ _8082_/A _7445_/B gnd _8086_/C vdd NAND2X1
XFILL_4__14429_ gnd vdd FILL
XFILL_3__9255_ gnd vdd FILL
XSFILL18600x48050 gnd vdd FILL
XSFILL69080x5050 gnd vdd FILL
XFILL_2__15608_ gnd vdd FILL
XFILL_1__14249_ gnd vdd FILL
XFILL_5__15719_ gnd vdd FILL
XFILL_0__14979_ gnd vdd FILL
X_7036_ _7128_/Q gnd _7038_/A vdd INVX1
XFILL_3__8206_ gnd vdd FILL
XFILL_1__8270_ gnd vdd FILL
XFILL_0__9477_ gnd vdd FILL
XFILL_2__15539_ gnd vdd FILL
XSFILL44040x40050 gnd vdd FILL
XFILL_1__7221_ gnd vdd FILL
XFILL_3__8137_ gnd vdd FILL
XSFILL23720x39050 gnd vdd FILL
XSFILL33880x83050 gnd vdd FILL
XFILL_0__8359_ gnd vdd FILL
XFILL_3__8068_ gnd vdd FILL
X_8987_ _8996_/A _8987_/B gnd _8988_/C vdd NAND2X1
XSFILL18840x7050 gnd vdd FILL
XFILL_4__8950_ gnd vdd FILL
XFILL111800x61050 gnd vdd FILL
X_7938_ _7938_/A gnd _7938_/Y vdd INVX1
XFILL_1__7083_ gnd vdd FILL
XSFILL38920x20050 gnd vdd FILL
XFILL_4__8881_ gnd vdd FILL
XSFILL79000x13050 gnd vdd FILL
XFILL_6__9797_ gnd vdd FILL
X_7869_ _7867_/Y _7872_/B _7868_/Y gnd _7917_/D vdd OAI21X1
XFILL_4__7832_ gnd vdd FILL
XFILL_0_BUFX2_insert909 gnd vdd FILL
X_9608_ _9608_/A gnd _9608_/Y vdd INVX1
XFILL_6__8748_ gnd vdd FILL
XFILL_4__7763_ gnd vdd FILL
XSFILL3640x60050 gnd vdd FILL
X_11470_ _11467_/Y _11469_/Y _11470_/C gnd _11479_/B vdd AOI21X1
X_9539_ _9537_/Y _9554_/B _9539_/C gnd _9583_/D vdd OAI21X1
XFILL_1__7985_ gnd vdd FILL
XFILL_4__9502_ gnd vdd FILL
XSFILL28840x72050 gnd vdd FILL
X_10421_ _10475_/Q gnd _10423_/A vdd INVX1
XFILL_4__7694_ gnd vdd FILL
XFILL_1__9724_ gnd vdd FILL
XFILL_1__6936_ gnd vdd FILL
X_13140_ _13134_/A _13140_/B gnd _13141_/C vdd NAND2X1
X_10352_ _14703_/A _7268_/CLK _7649_/R vdd _10352_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert820 gnd vdd FILL
XFILL_1__9655_ gnd vdd FILL
XSFILL44040x2050 gnd vdd FILL
XFILL_1__6867_ gnd vdd FILL
XFILL_4_BUFX2_insert831 gnd vdd FILL
XFILL_4_BUFX2_insert842 gnd vdd FILL
XFILL_4__9364_ gnd vdd FILL
XFILL_4_BUFX2_insert853 gnd vdd FILL
XFILL_6_CLKBUF1_insert208 gnd vdd FILL
X_13071_ _6894_/A _9060_/CLK _9060_/R vdd _13071_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert864 gnd vdd FILL
XFILL_1__8606_ gnd vdd FILL
XFILL_6_CLKBUF1_insert219 gnd vdd FILL
XFILL_4_BUFX2_insert875 gnd vdd FILL
X_10283_ _10281_/Y _10285_/A _10282_/Y gnd _10343_/D vdd OAI21X1
XFILL_4__8315_ gnd vdd FILL
XFILL_4_BUFX2_insert886 gnd vdd FILL
XFILL_4__9295_ gnd vdd FILL
XFILL_4_BUFX2_insert897 gnd vdd FILL
X_12022_ _12019_/Y _12022_/B _12022_/C gnd _12022_/Y vdd NAND3X1
XFILL_2__7330_ gnd vdd FILL
XFILL_4__8246_ gnd vdd FILL
XSFILL49640x51050 gnd vdd FILL
XFILL_1__8468_ gnd vdd FILL
XFILL_2__9000_ gnd vdd FILL
X_13973_ _13971_/Y _13973_/B _13973_/C gnd _13974_/A vdd NAND3X1
XFILL_1__7419_ gnd vdd FILL
XSFILL3720x40050 gnd vdd FILL
XFILL_1__8399_ gnd vdd FILL
XFILL_2__7192_ gnd vdd FILL
X_15712_ _8230_/A gnd _15713_/D vdd INVX1
XFILL_4__10110_ gnd vdd FILL
X_12924_ _12131_/B _9823_/CLK _9823_/R vdd _12924_/D gnd vdd DFFSR
XFILL_5__8990_ gnd vdd FILL
XSFILL28920x52050 gnd vdd FILL
XFILL_4__11090_ gnd vdd FILL
XFILL_0__10660_ gnd vdd FILL
XFILL_4__7059_ gnd vdd FILL
XFILL_5__7941_ gnd vdd FILL
XFILL_5__11400_ gnd vdd FILL
XFILL_6__10951_ gnd vdd FILL
X_15643_ _8292_/Q gnd _15644_/C vdd INVX1
XFILL_1_BUFX2_insert710 gnd vdd FILL
XFILL_4__10041_ gnd vdd FILL
X_12855_ _12853_/Y vdd _12855_/C gnd _12855_/Y vdd OAI21X1
XFILL_5__12380_ gnd vdd FILL
XFILL_1_BUFX2_insert721 gnd vdd FILL
XFILL_2__11220_ gnd vdd FILL
XFILL_3__10771_ gnd vdd FILL
XFILL_1__11950_ gnd vdd FILL
XFILL_1_BUFX2_insert732 gnd vdd FILL
XFILL_5__7872_ gnd vdd FILL
XFILL_1_BUFX2_insert743 gnd vdd FILL
X_11806_ _11249_/Y _11768_/B _11835_/C gnd _11806_/Y vdd AOI21X1
XFILL_3__12510_ gnd vdd FILL
XFILL_5__11331_ gnd vdd FILL
X_15574_ _8733_/A _15821_/B _15978_/C _8477_/A gnd _15580_/A vdd AOI22X1
XFILL_1_BUFX2_insert754 gnd vdd FILL
X_12786_ _12789_/A memoryOutData[30] gnd _12787_/C vdd NAND2X1
XFILL_1_BUFX2_insert765 gnd vdd FILL
XFILL_2__9902_ gnd vdd FILL
XFILL_1__10901_ gnd vdd FILL
XFILL_3__13490_ gnd vdd FILL
XFILL_0__12330_ gnd vdd FILL
XFILL_2__11151_ gnd vdd FILL
XFILL_5__9611_ gnd vdd FILL
XFILL_1_BUFX2_insert776 gnd vdd FILL
XFILL_1__11881_ gnd vdd FILL
X_14525_ _8760_/A _13853_/B _14525_/C gnd _14525_/Y vdd AOI21X1
XFILL_1_BUFX2_insert787 gnd vdd FILL
XFILL_4__13800_ gnd vdd FILL
XFILL_1_BUFX2_insert798 gnd vdd FILL
XFILL_5__14050_ gnd vdd FILL
XSFILL99480x38050 gnd vdd FILL
XFILL_5__11262_ gnd vdd FILL
X_11737_ _11731_/B _11079_/Y _11737_/C gnd _11740_/B vdd NAND3X1
XFILL_3__12441_ gnd vdd FILL
XFILL_2__10102_ gnd vdd FILL
XFILL_1__13620_ gnd vdd FILL
XFILL_4__14780_ gnd vdd FILL
XFILL_4__11992_ gnd vdd FILL
XFILL_0__12261_ gnd vdd FILL
XFILL_2__11082_ gnd vdd FILL
XFILL_1__10832_ gnd vdd FILL
XSFILL84280x80050 gnd vdd FILL
XFILL_4_BUFX2_insert14 gnd vdd FILL
XFILL_5__9542_ gnd vdd FILL
XFILL_5__13001_ gnd vdd FILL
X_14456_ _14456_/A _13587_/C _14456_/C _14454_/Y gnd _14457_/B vdd OAI22X1
XFILL_4_BUFX2_insert25 gnd vdd FILL
XFILL_4_BUFX2_insert36 gnd vdd FILL
X_11668_ _11059_/Y _11681_/B gnd _11668_/Y vdd NAND2X1
XFILL_4__13731_ gnd vdd FILL
XFILL_3__15160_ gnd vdd FILL
XFILL_5__11193_ gnd vdd FILL
XFILL_2__9764_ gnd vdd FILL
XFILL_4__10943_ gnd vdd FILL
XFILL_3__12372_ gnd vdd FILL
XFILL_0__14000_ gnd vdd FILL
XFILL_2__10033_ gnd vdd FILL
XFILL_4_BUFX2_insert47 gnd vdd FILL
XFILL_2__14910_ gnd vdd FILL
XFILL_0__11212_ gnd vdd FILL
XFILL_2__6976_ gnd vdd FILL
XFILL_1__13551_ gnd vdd FILL
XFILL_2__15890_ gnd vdd FILL
XFILL_1__10763_ gnd vdd FILL
X_13407_ _12809_/Q _13406_/Y gnd _13407_/Y vdd NOR2X1
XFILL_4_BUFX2_insert58 gnd vdd FILL
XFILL_0__12192_ gnd vdd FILL
XFILL_5__9473_ gnd vdd FILL
XFILL_5__10144_ gnd vdd FILL
XFILL_4_BUFX2_insert69 gnd vdd FILL
X_10619_ _10617_/Y _10619_/B _10618_/Y gnd _10619_/Y vdd OAI21X1
XFILL_3__14111_ gnd vdd FILL
XFILL_4__16450_ gnd vdd FILL
X_14387_ _14387_/A _14387_/B gnd _14387_/Y vdd NOR2X1
XFILL_3__11323_ gnd vdd FILL
XFILL_2__14841_ gnd vdd FILL
XFILL_2__8715_ gnd vdd FILL
XFILL_1__12502_ gnd vdd FILL
XFILL_4__13662_ gnd vdd FILL
XFILL_4__10874_ gnd vdd FILL
X_11599_ _11660_/A _11598_/Y _11599_/C gnd _11599_/Y vdd NAND3X1
XFILL_3__15091_ gnd vdd FILL
XFILL_0__11143_ gnd vdd FILL
XFILL_1__16270_ gnd vdd FILL
XSFILL109480x23050 gnd vdd FILL
X_16126_ _14768_/B _15569_/C _15687_/A _16126_/D gnd _16128_/A vdd OAI22X1
XFILL_1__13482_ gnd vdd FILL
X_13338_ _13337_/Y _13335_/Y gnd _13338_/Y vdd NOR2X1
XFILL_4__15401_ gnd vdd FILL
XFILL_1__10694_ gnd vdd FILL
XFILL_0__7730_ gnd vdd FILL
XFILL_4__12613_ gnd vdd FILL
XFILL_3__14042_ gnd vdd FILL
XFILL_5__14952_ gnd vdd FILL
XFILL_1__15221_ gnd vdd FILL
XFILL_2__8646_ gnd vdd FILL
XFILL_4__16381_ gnd vdd FILL
XFILL_3__11254_ gnd vdd FILL
XFILL112280x62050 gnd vdd FILL
XFILL_4__13593_ gnd vdd FILL
XFILL_1__12433_ gnd vdd FILL
XFILL_2__14772_ gnd vdd FILL
XFILL_5__8355_ gnd vdd FILL
XFILL_2__11984_ gnd vdd FILL
XFILL_0__15951_ gnd vdd FILL
XFILL_0__11074_ gnd vdd FILL
XFILL_5__13903_ gnd vdd FILL
X_16057_ _16261_/A _14675_/D _14675_/A _16261_/D gnd _16058_/B vdd OAI22X1
X_13269_ _13297_/C _13269_/B gnd _13269_/Y vdd NOR2X1
XFILL_4__15332_ gnd vdd FILL
XFILL_2__13723_ gnd vdd FILL
XFILL_5__14883_ gnd vdd FILL
XFILL_2__8577_ gnd vdd FILL
XFILL_2__10935_ gnd vdd FILL
XFILL_3__7370_ gnd vdd FILL
XFILL_5__7306_ gnd vdd FILL
XFILL_2_BUFX2_insert1008 gnd vdd FILL
XFILL_3__11185_ gnd vdd FILL
XFILL_1__15152_ gnd vdd FILL
XFILL_0__14902_ gnd vdd FILL
XFILL_0__10025_ gnd vdd FILL
XFILL_1__12364_ gnd vdd FILL
X_15008_ _15008_/A _15008_/B _15008_/C gnd _15028_/B vdd NAND3X1
XFILL_0__9400_ gnd vdd FILL
XFILL_2_BUFX2_insert1019 gnd vdd FILL
XFILL_0__15882_ gnd vdd FILL
XFILL_5__13834_ gnd vdd FILL
XFILL_0__7592_ gnd vdd FILL
XFILL_3__10136_ gnd vdd FILL
XFILL_4__12475_ gnd vdd FILL
XFILL_1__14103_ gnd vdd FILL
XFILL_4__15263_ gnd vdd FILL
XFILL_2__13654_ gnd vdd FILL
XFILL_1__11315_ gnd vdd FILL
XFILL_3__15993_ gnd vdd FILL
XFILL_0__14833_ gnd vdd FILL
XFILL_5__7237_ gnd vdd FILL
XFILL_1__15083_ gnd vdd FILL
XFILL_1__12295_ gnd vdd FILL
XFILL_4__14214_ gnd vdd FILL
XFILL_4__11426_ gnd vdd FILL
XFILL_2__12605_ gnd vdd FILL
XFILL_5__13765_ gnd vdd FILL
XFILL_3__9040_ gnd vdd FILL
XSFILL28840x2050 gnd vdd FILL
XFILL_5__10977_ gnd vdd FILL
XFILL_4__15194_ gnd vdd FILL
XFILL_2__7459_ gnd vdd FILL
XFILL_1__14034_ gnd vdd FILL
XFILL_3__10067_ gnd vdd FILL
XFILL_3__14944_ gnd vdd FILL
XFILL_2__16373_ gnd vdd FILL
XSFILL18680x22050 gnd vdd FILL
XFILL_2__13585_ gnd vdd FILL
XFILL_1__11246_ gnd vdd FILL
XFILL_5__7168_ gnd vdd FILL
XFILL_5__15504_ gnd vdd FILL
XFILL_2__10797_ gnd vdd FILL
XSFILL74200x16050 gnd vdd FILL
XFILL_0__14764_ gnd vdd FILL
X_8910_ _8896_/B _8910_/B gnd _8910_/Y vdd NAND2X1
XFILL_5__12716_ gnd vdd FILL
XFILL_0__11976_ gnd vdd FILL
XFILL_0__9262_ gnd vdd FILL
XFILL_2__15324_ gnd vdd FILL
XFILL_4__14145_ gnd vdd FILL
XFILL_4__11357_ gnd vdd FILL
X_9890_ _9890_/A _9868_/A _9890_/C gnd _9890_/Y vdd OAI21X1
XFILL_5__13696_ gnd vdd FILL
XFILL_3__14875_ gnd vdd FILL
XFILL_0__13715_ gnd vdd FILL
XFILL_1__11177_ gnd vdd FILL
XFILL_0__10927_ gnd vdd FILL
XFILL_0__8213_ gnd vdd FILL
XFILL_5__7099_ gnd vdd FILL
XSFILL59000x77050 gnd vdd FILL
XFILL_0_BUFX2_insert1001 gnd vdd FILL
XFILL_4__10308_ gnd vdd FILL
XFILL_0__14695_ gnd vdd FILL
XFILL_5__15435_ gnd vdd FILL
X_8841_ _8823_/B _7177_/B gnd _8842_/C vdd NAND2X1
XFILL_5__12647_ gnd vdd FILL
XFILL_0_BUFX2_insert1012 gnd vdd FILL
XFILL_4__14076_ gnd vdd FILL
XFILL_2__9129_ gnd vdd FILL
XFILL_1__10128_ gnd vdd FILL
XFILL_3__13826_ gnd vdd FILL
XFILL_2__15255_ gnd vdd FILL
XFILL_4__11288_ gnd vdd FILL
XFILL_0_BUFX2_insert1023 gnd vdd FILL
XSFILL99400x82050 gnd vdd FILL
XFILL_2__12467_ gnd vdd FILL
XFILL_0_BUFX2_insert1034 gnd vdd FILL
XFILL_1__15985_ gnd vdd FILL
XFILL_0__13646_ gnd vdd FILL
XFILL_4__13027_ gnd vdd FILL
XFILL_0__8144_ gnd vdd FILL
XFILL_0_BUFX2_insert1045 gnd vdd FILL
XFILL_4__10239_ gnd vdd FILL
XFILL_5__15366_ gnd vdd FILL
XFILL_2__14206_ gnd vdd FILL
XFILL_0_BUFX2_insert1056 gnd vdd FILL
XFILL_5__12578_ gnd vdd FILL
X_8772_ _8772_/A gnd _8772_/Y vdd INVX1
XFILL_0_BUFX2_insert1067 gnd vdd FILL
XFILL_2__11418_ gnd vdd FILL
XFILL_3__10969_ gnd vdd FILL
XFILL_6_BUFX2_insert904 gnd vdd FILL
XFILL_2__15186_ gnd vdd FILL
XFILL_1__10059_ gnd vdd FILL
XFILL_3__13757_ gnd vdd FILL
XFILL_1__14936_ gnd vdd FILL
XFILL_0_BUFX2_insert1089 gnd vdd FILL
XFILL_2__12398_ gnd vdd FILL
XFILL_0__16365_ gnd vdd FILL
XSFILL38840x35050 gnd vdd FILL
XFILL_0__10789_ gnd vdd FILL
XFILL112360x42050 gnd vdd FILL
XFILL_5__14317_ gnd vdd FILL
XFILL_0__13577_ gnd vdd FILL
XFILL_6__13868_ gnd vdd FILL
XSFILL64120x68050 gnd vdd FILL
XFILL_0__8075_ gnd vdd FILL
XFILL_6__6863_ gnd vdd FILL
XFILL_5__11529_ gnd vdd FILL
X_7723_ _7723_/A _7723_/B _7722_/Y gnd _7783_/D vdd OAI21X1
XFILL_3__12708_ gnd vdd FILL
XFILL_5__15297_ gnd vdd FILL
XFILL_2__14137_ gnd vdd FILL
XFILL_0__15316_ gnd vdd FILL
XFILL_3__13688_ gnd vdd FILL
XFILL_2__11349_ gnd vdd FILL
XFILL_1__14867_ gnd vdd FILL
XFILL_0__12528_ gnd vdd FILL
XFILL_3__9873_ gnd vdd FILL
XFILL_5__9809_ gnd vdd FILL
XFILL_0__16296_ gnd vdd FILL
XFILL_5__14248_ gnd vdd FILL
X_7654_ _7590_/A _8038_/CLK _8038_/R vdd _7592_/Y gnd vdd DFFSR
XFILL_3__12639_ gnd vdd FILL
XFILL_3__15427_ gnd vdd FILL
XFILL_1__13818_ gnd vdd FILL
XFILL_3__8824_ gnd vdd FILL
XFILL_2__14068_ gnd vdd FILL
XFILL_4__14978_ gnd vdd FILL
XFILL_0__15247_ gnd vdd FILL
XFILL_0__12459_ gnd vdd FILL
XFILL_1__14798_ gnd vdd FILL
XSFILL3560x75050 gnd vdd FILL
XFILL_5__14179_ gnd vdd FILL
XFILL_2__13019_ gnd vdd FILL
XFILL_4__13929_ gnd vdd FILL
XFILL_3__15358_ gnd vdd FILL
X_7585_ _7606_/A _9633_/B gnd _7586_/C vdd NAND2X1
XSFILL94200x2050 gnd vdd FILL
XFILL_1__13749_ gnd vdd FILL
XFILL_3__8755_ gnd vdd FILL
XFILL_0__15178_ gnd vdd FILL
XFILL_6__8464_ gnd vdd FILL
X_9324_ _9272_/A _9958_/CLK _9580_/R vdd _9324_/D gnd vdd DFFSR
XFILL_3__14309_ gnd vdd FILL
XFILL_0__8977_ gnd vdd FILL
XSFILL8600x12050 gnd vdd FILL
XFILL_3__7706_ gnd vdd FILL
XSFILL44040x35050 gnd vdd FILL
XFILL_3__15289_ gnd vdd FILL
XFILL_4_BUFX2_insert105 gnd vdd FILL
XFILL_0__14129_ gnd vdd FILL
XFILL_6__7415_ gnd vdd FILL
XFILL_0__7928_ gnd vdd FILL
X_9255_ _9277_/B _9895_/B gnd _9256_/C vdd NAND2X1
XFILL_3__7637_ gnd vdd FILL
XFILL_1__15419_ gnd vdd FILL
XFILL_1__16399_ gnd vdd FILL
X_8206_ _8206_/A gnd _8208_/A vdd INVX1
XFILL_0__7859_ gnd vdd FILL
XSFILL33880x78050 gnd vdd FILL
X_9186_ _9186_/Q _7382_/CLK _8674_/R vdd _9116_/Y gnd vdd DFFSR
XFILL_3__7568_ gnd vdd FILL
XFILL_3_BUFX2_insert805 gnd vdd FILL
XFILL_3_BUFX2_insert816 gnd vdd FILL
XFILL_4__8100_ gnd vdd FILL
XFILL_3_BUFX2_insert827 gnd vdd FILL
XFILL_1__9371_ gnd vdd FILL
X_8137_ _8137_/A _8098_/B _8136_/Y gnd _8137_/Y vdd OAI21X1
XFILL_3_BUFX2_insert838 gnd vdd FILL
XFILL_4__9080_ gnd vdd FILL
XFILL112440x22050 gnd vdd FILL
XFILL_3__7499_ gnd vdd FILL
XSFILL64200x48050 gnd vdd FILL
XFILL_3_BUFX2_insert849 gnd vdd FILL
XFILL_1__8322_ gnd vdd FILL
XFILL_0__9529_ gnd vdd FILL
X_8068_ _8066_/Y _8118_/A _8068_/C gnd _8068_/Y vdd OAI21X1
XFILL_3__9238_ gnd vdd FILL
XFILL_1__8253_ gnd vdd FILL
X_7019_ _7019_/Q _7147_/CLK _7531_/R vdd _6967_/Y gnd vdd DFFSR
XFILL_3__9169_ gnd vdd FILL
XFILL_1__7204_ gnd vdd FILL
XSFILL3640x55050 gnd vdd FILL
X_10970_ _10970_/A _10970_/B _10936_/B gnd _10971_/B vdd OAI21X1
XFILL_1__8184_ gnd vdd FILL
XSFILL28840x67050 gnd vdd FILL
XSFILL94280x43050 gnd vdd FILL
XFILL_4__9982_ gnd vdd FILL
X_12640_ vdd memoryOutData[24] gnd _12641_/C vdd NAND2X1
XFILL_1__7066_ gnd vdd FILL
XFILL_4__8864_ gnd vdd FILL
XFILL_0_CLKBUF1_insert121 gnd vdd FILL
X_12571_ vdd memoryOutData[1] gnd _12572_/C vdd NAND2X1
XSFILL33960x58050 gnd vdd FILL
XFILL_0_BUFX2_insert706 gnd vdd FILL
XFILL_0_CLKBUF1_insert132 gnd vdd FILL
XFILL_0_BUFX2_insert717 gnd vdd FILL
XFILL_0_CLKBUF1_insert143 gnd vdd FILL
XFILL_0_BUFX2_insert728 gnd vdd FILL
X_14310_ _14306_/Y _14310_/B _14310_/C gnd _14311_/B vdd NAND3X1
XFILL_4__7815_ gnd vdd FILL
XFILL_0_CLKBUF1_insert154 gnd vdd FILL
XFILL_0_BUFX2_insert739 gnd vdd FILL
X_11522_ _11107_/B _11517_/Y _11543_/C gnd _11522_/Y vdd NAND3X1
XFILL_0_CLKBUF1_insert165 gnd vdd FILL
XFILL_0_CLKBUF1_insert176 gnd vdd FILL
X_15290_ _7813_/A gnd _15291_/A vdd INVX1
XFILL_0_CLKBUF1_insert187 gnd vdd FILL
XSFILL33560x60050 gnd vdd FILL
XFILL_0_CLKBUF1_insert198 gnd vdd FILL
XSFILL48360x20050 gnd vdd FILL
X_14241_ _14237_/Y _14241_/B gnd _14242_/B vdd NOR2X1
XFILL_4__7746_ gnd vdd FILL
X_11453_ _11289_/C _11449_/Y _11452_/Y gnd _11454_/A vdd AOI21X1
XFILL_1__7968_ gnd vdd FILL
XSFILL89240x32050 gnd vdd FILL
X_10404_ _10405_/B _7972_/B gnd _10404_/Y vdd NAND2X1
XFILL_4__7677_ gnd vdd FILL
X_14172_ _16432_/Q gnd _14174_/D vdd INVX1
XFILL_2__8500_ gnd vdd FILL
XFILL_1__6919_ gnd vdd FILL
X_11384_ _11384_/A _11038_/Y _11383_/Y gnd _11385_/C vdd OAI21X1
XFILL_2__9480_ gnd vdd FILL
XSFILL3720x35050 gnd vdd FILL
XFILL_4__9416_ gnd vdd FILL
X_13123_ _13123_/A _13099_/B _13122_/Y gnd _13123_/Y vdd OAI21X1
XSFILL94360x8050 gnd vdd FILL
XSFILL13320x68050 gnd vdd FILL
XFILL_4_BUFX2_insert650 gnd vdd FILL
X_10335_ _13920_/A _7274_/CLK _7274_/R vdd _10335_/D gnd vdd DFFSR
XFILL_1__9638_ gnd vdd FILL
XSFILL28920x47050 gnd vdd FILL
XFILL_4_BUFX2_insert661 gnd vdd FILL
XFILL_4_BUFX2_insert672 gnd vdd FILL
XFILL_5__8140_ gnd vdd FILL
XSFILL94360x23050 gnd vdd FILL
XFILL_4__9347_ gnd vdd FILL
XFILL_4_BUFX2_insert683 gnd vdd FILL
XFILL_5__10900_ gnd vdd FILL
X_13054_ _6877_/A _12669_/CLK _12795_/R vdd _13054_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert694 gnd vdd FILL
X_10266_ _15537_/B gnd _10268_/A vdd INVX1
XFILL_5__11880_ gnd vdd FILL
XFILL_2__8362_ gnd vdd FILL
XFILL_4__9278_ gnd vdd FILL
X_12005_ _12005_/A _12093_/B _12061_/C gnd gnd _12005_/Y vdd AOI22X1
XFILL_5__8071_ gnd vdd FILL
XFILL_5__10831_ gnd vdd FILL
XFILL_4__12260_ gnd vdd FILL
XFILL_2__7313_ gnd vdd FILL
XSFILL103720x42050 gnd vdd FILL
X_10197_ _10197_/A _10160_/A _10196_/Y gnd _10197_/Y vdd OAI21X1
XFILL_1__11100_ gnd vdd FILL
XFILL_4__8229_ gnd vdd FILL
XFILL_1__12080_ gnd vdd FILL
XFILL_2__10651_ gnd vdd FILL
XFILL_3__12990_ gnd vdd FILL
XFILL_0__11830_ gnd vdd FILL
XFILL_4__11211_ gnd vdd FILL
XFILL_5__13550_ gnd vdd FILL
XFILL_2__7244_ gnd vdd FILL
XFILL_5__10762_ gnd vdd FILL
XFILL_3__11941_ gnd vdd FILL
XFILL_4__12191_ gnd vdd FILL
XFILL_1__11031_ gnd vdd FILL
XFILL_2__13370_ gnd vdd FILL
XFILL_6__14840_ gnd vdd FILL
XFILL_5__12501_ gnd vdd FILL
XSFILL33640x40050 gnd vdd FILL
XFILL_0__11761_ gnd vdd FILL
XSFILL84280x75050 gnd vdd FILL
XFILL_4__11142_ gnd vdd FILL
XFILL_2__12321_ gnd vdd FILL
X_13956_ _13956_/A _14725_/A _14949_/C _13956_/D gnd _13960_/B vdd OAI22X1
XFILL_5__13481_ gnd vdd FILL
XFILL_3__11872_ gnd vdd FILL
XFILL_5__10693_ gnd vdd FILL
XFILL_3__14660_ gnd vdd FILL
XFILL_0__13500_ gnd vdd FILL
XFILL_2__7175_ gnd vdd FILL
XSFILL74520x52050 gnd vdd FILL
XFILL_0__14480_ gnd vdd FILL
XFILL_5__15220_ gnd vdd FILL
XFILL_0__11692_ gnd vdd FILL
XFILL_5__12432_ gnd vdd FILL
XFILL_5__8973_ gnd vdd FILL
XSFILL59080x51050 gnd vdd FILL
X_12907_ _12907_/A gnd _12907_/Y vdd INVX1
XSFILL89320x12050 gnd vdd FILL
X_13887_ _13863_/Y _13886_/Y _14265_/C gnd _12976_/B vdd AOI21X1
XFILL_3__13611_ gnd vdd FILL
XFILL_6__11983_ gnd vdd FILL
XFILL_2__15040_ gnd vdd FILL
XFILL_4__15950_ gnd vdd FILL
XFILL_4__11073_ gnd vdd FILL
XFILL_3__10823_ gnd vdd FILL
XFILL_3__14591_ gnd vdd FILL
XFILL_2__12252_ gnd vdd FILL
XFILL_0__13431_ gnd vdd FILL
XFILL_1__15770_ gnd vdd FILL
XFILL_0__10643_ gnd vdd FILL
XSFILL109480x18050 gnd vdd FILL
XFILL_1__12982_ gnd vdd FILL
XFILL_4__10024_ gnd vdd FILL
X_15626_ _15626_/A _15899_/A gnd _15627_/C vdd NOR2X1
XSFILL8760x9050 gnd vdd FILL
X_12838_ _12131_/B gnd _12838_/Y vdd INVX1
XFILL_5__15151_ gnd vdd FILL
XFILL_4__14901_ gnd vdd FILL
XFILL_1_BUFX2_insert540 gnd vdd FILL
XFILL_5__12363_ gnd vdd FILL
XFILL_3__16330_ gnd vdd FILL
XFILL_3__13542_ gnd vdd FILL
XFILL_2__11203_ gnd vdd FILL
XFILL_3__10754_ gnd vdd FILL
XFILL_1__14721_ gnd vdd FILL
XFILL_1_BUFX2_insert551 gnd vdd FILL
XFILL_4__15881_ gnd vdd FILL
XFILL_1_BUFX2_insert562 gnd vdd FILL
XFILL112280x57050 gnd vdd FILL
XFILL_1__11933_ gnd vdd FILL
XFILL_2__12183_ gnd vdd FILL
XFILL_0__16150_ gnd vdd FILL
XFILL_0__10574_ gnd vdd FILL
XFILL_0__13362_ gnd vdd FILL
XFILL_1_BUFX2_insert573 gnd vdd FILL
XFILL_5__14102_ gnd vdd FILL
XFILL_1_BUFX2_insert584 gnd vdd FILL
XFILL_5__7855_ gnd vdd FILL
XFILL_5__11314_ gnd vdd FILL
X_12769_ _12767_/Y _12723_/A _12769_/C gnd _12815_/D vdd OAI21X1
XFILL_4__14832_ gnd vdd FILL
X_15557_ _14058_/A _15378_/B _15556_/Y gnd _15559_/A vdd OAI21X1
XFILL_5__15082_ gnd vdd FILL
XFILL_1_BUFX2_insert595 gnd vdd FILL
XFILL_3__13473_ gnd vdd FILL
XFILL_5__12294_ gnd vdd FILL
XFILL_2__11134_ gnd vdd FILL
XFILL_0__15101_ gnd vdd FILL
XFILL_3__16261_ gnd vdd FILL
XFILL_3__10685_ gnd vdd FILL
XFILL_0__12313_ gnd vdd FILL
XFILL_3__6870_ gnd vdd FILL
XFILL_1__14652_ gnd vdd FILL
XFILL_0__13293_ gnd vdd FILL
XFILL_1__11864_ gnd vdd FILL
XFILL_0__16081_ gnd vdd FILL
X_14508_ _10220_/Q gnd _14509_/A vdd INVX1
XFILL_5__14033_ gnd vdd FILL
XFILL_0__8900_ gnd vdd FILL
XFILL_0__9880_ gnd vdd FILL
XFILL_3__15212_ gnd vdd FILL
XFILL_3__12424_ gnd vdd FILL
X_15488_ _8340_/A gnd _15488_/Y vdd INVX1
XFILL_5__11245_ gnd vdd FILL
XFILL_1__13603_ gnd vdd FILL
XFILL_3__16192_ gnd vdd FILL
XFILL_6__10796_ gnd vdd FILL
XFILL_4__14763_ gnd vdd FILL
XFILL_1__10815_ gnd vdd FILL
XFILL_4__11975_ gnd vdd FILL
XFILL_0__15032_ gnd vdd FILL
XFILL_2__15942_ gnd vdd FILL
XFILL_0__12244_ gnd vdd FILL
XFILL_2__11065_ gnd vdd FILL
XFILL_5__9525_ gnd vdd FILL
XFILL_1__14583_ gnd vdd FILL
XFILL_0__8831_ gnd vdd FILL
XFILL_1__11795_ gnd vdd FILL
XFILL_3__15143_ gnd vdd FILL
XFILL_5__11176_ gnd vdd FILL
XFILL_4__13714_ gnd vdd FILL
X_14439_ _10418_/A gnd _15870_/A vdd INVX1
X_7370_ _7370_/A gnd _7372_/A vdd INVX1
XFILL_4__10926_ gnd vdd FILL
XFILL_2__10016_ gnd vdd FILL
XFILL_1__16322_ gnd vdd FILL
XFILL_3__12355_ gnd vdd FILL
XFILL_2__6959_ gnd vdd FILL
XFILL_4__14694_ gnd vdd FILL
XFILL_2__9747_ gnd vdd FILL
XFILL_1__13534_ gnd vdd FILL
XFILL_0__12175_ gnd vdd FILL
XFILL_2__15873_ gnd vdd FILL
XFILL_1__10746_ gnd vdd FILL
XSFILL18680x17050 gnd vdd FILL
XSFILL114440x73050 gnd vdd FILL
XSFILL8520x27050 gnd vdd FILL
XFILL_5__10127_ gnd vdd FILL
XFILL_0__8762_ gnd vdd FILL
XFILL_3__11306_ gnd vdd FILL
XFILL_5__15984_ gnd vdd FILL
XFILL_4__13645_ gnd vdd FILL
XFILL_3__15074_ gnd vdd FILL
XFILL_3__8471_ gnd vdd FILL
XFILL_2__14824_ gnd vdd FILL
XFILL_0__11126_ gnd vdd FILL
XFILL_1__16253_ gnd vdd FILL
XFILL_3__12286_ gnd vdd FILL
XFILL_2__9678_ gnd vdd FILL
XSFILL84360x55050 gnd vdd FILL
XFILL_1__13465_ gnd vdd FILL
XFILL_1__10677_ gnd vdd FILL
XFILL_0__7713_ gnd vdd FILL
X_16109_ _16107_/Y _15239_/B _15953_/A _16108_/Y gnd _16109_/Y vdd OAI22X1
XFILL_5__10058_ gnd vdd FILL
XFILL_3__14025_ gnd vdd FILL
X_9040_ _9040_/A gnd _9042_/A vdd INVX1
XFILL_5__14935_ gnd vdd FILL
XFILL_5__9387_ gnd vdd FILL
XFILL_1__15204_ gnd vdd FILL
XFILL_4__16364_ gnd vdd FILL
XFILL_6__12397_ gnd vdd FILL
XFILL_3__7422_ gnd vdd FILL
XFILL_3__11237_ gnd vdd FILL
XFILL_4__10788_ gnd vdd FILL
XFILL_2__8629_ gnd vdd FILL
XFILL_1__12416_ gnd vdd FILL
XFILL_4__13576_ gnd vdd FILL
XFILL_2__14755_ gnd vdd FILL
XFILL_1__16184_ gnd vdd FILL
XFILL_2__11967_ gnd vdd FILL
XFILL_0__15934_ gnd vdd FILL
XSFILL59160x31050 gnd vdd FILL
XFILL_0__11057_ gnd vdd FILL
XFILL_1__13396_ gnd vdd FILL
XFILL_5__8338_ gnd vdd FILL
XFILL_4__15315_ gnd vdd FILL
XFILL_5__14866_ gnd vdd FILL
XFILL_4__12527_ gnd vdd FILL
XFILL_2__13706_ gnd vdd FILL
XFILL_2__10918_ gnd vdd FILL
XFILL_0__10008_ gnd vdd FILL
XFILL_3__7353_ gnd vdd FILL
XFILL_4__16295_ gnd vdd FILL
XFILL_1__15135_ gnd vdd FILL
XFILL_3__11168_ gnd vdd FILL
XFILL_1__12347_ gnd vdd FILL
XFILL_2__14686_ gnd vdd FILL
XFILL_5__8269_ gnd vdd FILL
XFILL_2__11898_ gnd vdd FILL
XFILL_0__15865_ gnd vdd FILL
XFILL_5__13817_ gnd vdd FILL
XFILL_4__15246_ gnd vdd FILL
XFILL_0__7575_ gnd vdd FILL
XFILL112360x37050 gnd vdd FILL
XFILL_3__10119_ gnd vdd FILL
XFILL_2__13637_ gnd vdd FILL
XFILL_5__14797_ gnd vdd FILL
XFILL_4__12458_ gnd vdd FILL
XCLKBUF1_insert1079 clk gnd CLKBUF1_insert193/A vdd CLKBUF1
XFILL_3__15976_ gnd vdd FILL
XFILL_1__15066_ gnd vdd FILL
XFILL_0__14816_ gnd vdd FILL
XFILL_3__11099_ gnd vdd FILL
XFILL_1__12278_ gnd vdd FILL
XFILL_0__15796_ gnd vdd FILL
XFILL_3__9023_ gnd vdd FILL
XFILL_5__13748_ gnd vdd FILL
X_9942_ _9942_/Q _6998_/CLK _7644_/R vdd _9942_/D gnd vdd DFFSR
XFILL_4__11409_ gnd vdd FILL
XFILL_4__15177_ gnd vdd FILL
XFILL_4__12389_ gnd vdd FILL
XFILL_1__14017_ gnd vdd FILL
XFILL_2__16356_ gnd vdd FILL
XFILL_0_BUFX2_insert12 gnd vdd FILL
XFILL_3__14927_ gnd vdd FILL
XFILL_2__13568_ gnd vdd FILL
XFILL_0_BUFX2_insert23 gnd vdd FILL
XFILL_1__11229_ gnd vdd FILL
XFILL_0_BUFX2_insert34 gnd vdd FILL
XFILL_0__14747_ gnd vdd FILL
XFILL_0__11959_ gnd vdd FILL
XSFILL79320x44050 gnd vdd FILL
XFILL_0_BUFX2_insert45 gnd vdd FILL
XFILL_0__9245_ gnd vdd FILL
XSFILL49080x83050 gnd vdd FILL
XFILL_4__14128_ gnd vdd FILL
XFILL_0_BUFX2_insert56 gnd vdd FILL
XFILL_2__15307_ gnd vdd FILL
XFILL_5__13679_ gnd vdd FILL
XFILL_2__12519_ gnd vdd FILL
X_9873_ _9951_/Q gnd _9875_/A vdd INVX1
XFILL_3__14858_ gnd vdd FILL
XFILL_2__16287_ gnd vdd FILL
XFILL_0_BUFX2_insert67 gnd vdd FILL
XFILL_0_BUFX2_insert78 gnd vdd FILL
XFILL_2__13499_ gnd vdd FILL
XFILL_0_BUFX2_insert89 gnd vdd FILL
XFILL_0__14678_ gnd vdd FILL
XFILL_5__15418_ gnd vdd FILL
X_8824_ _8822_/Y _8823_/B _8823_/Y gnd _8918_/D vdd OAI21X1
XFILL_3__13809_ gnd vdd FILL
XFILL_2__15238_ gnd vdd FILL
XFILL_4__14059_ gnd vdd FILL
XFILL_5__16398_ gnd vdd FILL
XSFILL114520x53050 gnd vdd FILL
XFILL_0__13629_ gnd vdd FILL
XFILL_1__15968_ gnd vdd FILL
XFILL_3__14789_ gnd vdd FILL
XFILL_0__8127_ gnd vdd FILL
XFILL_5__15349_ gnd vdd FILL
X_8755_ _8788_/A _8243_/B gnd _8756_/C vdd NAND2X1
XFILL_2__15169_ gnd vdd FILL
XFILL_3__9925_ gnd vdd FILL
XFILL_0__16348_ gnd vdd FILL
XFILL_1__14919_ gnd vdd FILL
XFILL_1__15899_ gnd vdd FILL
XFILL_6_BUFX2_insert756 gnd vdd FILL
X_7706_ _7706_/A gnd _7708_/A vdd INVX1
XFILL_0__8058_ gnd vdd FILL
XSFILL59240x11050 gnd vdd FILL
X_8686_ _8638_/A _8046_/CLK _9692_/R vdd _8686_/D gnd vdd DFFSR
XFILL_3__9856_ gnd vdd FILL
XFILL_0__16279_ gnd vdd FILL
XFILL_1__8871_ gnd vdd FILL
X_7637_ _7637_/A _7598_/B _7637_/C gnd _7669_/D vdd OAI21X1
XFILL111960x10050 gnd vdd FILL
XFILL_4__7600_ gnd vdd FILL
XFILL_4__8580_ gnd vdd FILL
XFILL_3__9787_ gnd vdd FILL
XFILL_6__8516_ gnd vdd FILL
XFILL112440x17050 gnd vdd FILL
XFILL_1__7822_ gnd vdd FILL
XSFILL73880x80050 gnd vdd FILL
XFILL_1_CLKBUF1_insert205 gnd vdd FILL
XFILL_1_CLKBUF1_insert216 gnd vdd FILL
X_7568_ _7566_/Y _7568_/B _7567_/Y gnd _7568_/Y vdd OAI21X1
XSFILL23720x52050 gnd vdd FILL
XFILL_3__8738_ gnd vdd FILL
XSFILL39000x19050 gnd vdd FILL
X_9307_ _9221_/A _7143_/CLK _7015_/R vdd _9223_/Y gnd vdd DFFSR
XFILL_1__7753_ gnd vdd FILL
XFILL_4__7462_ gnd vdd FILL
X_7499_ _7460_/A _7499_/B gnd _7499_/Y vdd NAND2X1
X_9238_ _9238_/A _9238_/B _9238_/C gnd _9312_/D vdd OAI21X1
XFILL_1__7684_ gnd vdd FILL
X_10120_ _10120_/A gnd _10122_/A vdd INVX1
XFILL_1__9423_ gnd vdd FILL
XFILL_3_BUFX2_insert602 gnd vdd FILL
XSFILL94280x38050 gnd vdd FILL
XSFILL114600x33050 gnd vdd FILL
XFILL_3_BUFX2_insert613 gnd vdd FILL
XFILL_4__9132_ gnd vdd FILL
X_9169_ _9112_/A _8401_/B gnd _9170_/C vdd NAND2X1
XFILL_3_BUFX2_insert624 gnd vdd FILL
XFILL_3_BUFX2_insert635 gnd vdd FILL
XFILL_3_BUFX2_insert646 gnd vdd FILL
X_10051_ _10051_/A _10054_/B _10050_/Y gnd _10095_/D vdd OAI21X1
XFILL_1__9354_ gnd vdd FILL
XSFILL69080x14050 gnd vdd FILL
XFILL_3_BUFX2_insert657 gnd vdd FILL
XFILL_3_BUFX2_insert668 gnd vdd FILL
XFILL_3_BUFX2_insert679 gnd vdd FILL
XFILL_4__8014_ gnd vdd FILL
XFILL_1__9285_ gnd vdd FILL
XSFILL104280x23050 gnd vdd FILL
X_13810_ _13808_/Y _14466_/C _14555_/C _13809_/Y gnd _13814_/B vdd OAI22X1
XFILL_1__8236_ gnd vdd FILL
X_14790_ _14789_/Y _14790_/B gnd _14790_/Y vdd NOR2X1
XSFILL33560x55050 gnd vdd FILL
X_13741_ _13854_/B _9224_/A _8328_/A _13848_/B gnd _13741_/Y vdd AOI22X1
XSFILL8760x83050 gnd vdd FILL
X_10953_ _10952_/Y gnd _10954_/B vdd INVX1
XFILL_1__7118_ gnd vdd FILL
X_13672_ _15233_/C _14466_/C _14555_/C _13671_/Y gnd _13673_/B vdd OAI22X1
X_10884_ _12695_/A _10883_/Y gnd _10887_/C vdd NOR2X1
XFILL_1__8098_ gnd vdd FILL
XSFILL59800x5050 gnd vdd FILL
XFILL_2__8980_ gnd vdd FILL
XFILL_4__8916_ gnd vdd FILL
X_12623_ _12621_/Y vdd _12623_/C gnd _12681_/D vdd OAI21X1
X_15411_ _15411_/A _15410_/Y gnd _15411_/Y vdd NOR2X1
XFILL_4__9896_ gnd vdd FILL
X_16391_ gnd gnd gnd _16392_/C vdd NAND2X1
XFILL_1__7049_ gnd vdd FILL
XFILL_0_BUFX2_insert503 gnd vdd FILL
XFILL_2__7931_ gnd vdd FILL
XFILL_0_BUFX2_insert514 gnd vdd FILL
XFILL_4__8847_ gnd vdd FILL
X_15342_ _13801_/Y _15342_/B gnd _15342_/Y vdd NOR2X1
XFILL_0_BUFX2_insert525 gnd vdd FILL
XSFILL94360x18050 gnd vdd FILL
X_12554_ _12496_/A _13201_/CLK _13201_/R vdd _12554_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert536 gnd vdd FILL
XFILL_2__7862_ gnd vdd FILL
XFILL_0_BUFX2_insert547 gnd vdd FILL
XFILL_0_BUFX2_insert558 gnd vdd FILL
XFILL_0_BUFX2_insert569 gnd vdd FILL
XSFILL28520x44050 gnd vdd FILL
X_11505_ _11185_/B _11185_/A gnd _11505_/Y vdd NOR2X1
XFILL_5__7571_ gnd vdd FILL
XFILL_5__11030_ gnd vdd FILL
XFILL_0__10290_ gnd vdd FILL
XFILL_4__8778_ gnd vdd FILL
X_15273_ _15273_/A _15273_/B _15273_/C gnd _15274_/A vdd NAND3X1
XFILL_2__9601_ gnd vdd FILL
X_12485_ vdd _12485_/B gnd _12485_/Y vdd NAND2X1
XFILL_4__11760_ gnd vdd FILL
XSFILL69400x56050 gnd vdd FILL
XSFILL94200x82050 gnd vdd FILL
X_14224_ _14223_/Y _14224_/B gnd _14224_/Y vdd NOR2X1
XFILL_1__11580_ gnd vdd FILL
XFILL_4__7729_ gnd vdd FILL
XSFILL109400x6050 gnd vdd FILL
X_11436_ _11312_/Y gnd _11437_/A vdd INVX2
XFILL_3__12140_ gnd vdd FILL
XFILL_2__9532_ gnd vdd FILL
XFILL_4__11691_ gnd vdd FILL
XFILL_1__10531_ gnd vdd FILL
XFILL_2__12870_ gnd vdd FILL
XFILL_5__9241_ gnd vdd FILL
X_14155_ _10656_/A gnd _15633_/B vdd INVX1
XFILL_4__13430_ gnd vdd FILL
XFILL_4__10642_ gnd vdd FILL
X_11367_ _11414_/A _11764_/A _11366_/Y gnd _11367_/Y vdd AOI21X1
XFILL_3__12071_ gnd vdd FILL
XFILL_2__9463_ gnd vdd FILL
XFILL_5__12981_ gnd vdd FILL
XFILL_2__11821_ gnd vdd FILL
XFILL_1__13250_ gnd vdd FILL
X_13106_ _11914_/A gnd _13108_/A vdd INVX1
XCLKBUF1_insert204 CLKBUF1_insert182/A gnd _7007_/CLK vdd CLKBUF1
XFILL_5__9172_ gnd vdd FILL
X_10318_ _10318_/A _8654_/B gnd _10319_/C vdd NAND2X1
XCLKBUF1_insert215 CLKBUF1_insert218/A gnd _7147_/CLK vdd CLKBUF1
XFILL_0__13980_ gnd vdd FILL
XFILL_5__14720_ gnd vdd FILL
XFILL_5__11932_ gnd vdd FILL
XFILL_4_BUFX2_insert480 gnd vdd FILL
X_14086_ _9757_/A gnd _14088_/D vdd INVX1
XFILL_3__11022_ gnd vdd FILL
XFILL_4__10573_ gnd vdd FILL
XFILL_4__13361_ gnd vdd FILL
XFILL_2__14540_ gnd vdd FILL
XFILL_1__12201_ gnd vdd FILL
X_11298_ _11297_/Y gnd _11298_/Y vdd INVX1
XFILL_4_BUFX2_insert491 gnd vdd FILL
XFILL_5__8123_ gnd vdd FILL
XFILL_2__9394_ gnd vdd FILL
XFILL_2__11752_ gnd vdd FILL
XSFILL99480x51050 gnd vdd FILL
XFILL_1__10393_ gnd vdd FILL
XFILL_4__15100_ gnd vdd FILL
X_13037_ _13035_/Y vdd _13037_/C gnd _13075_/D vdd OAI21X1
X_10249_ _10304_/B _7177_/B gnd _10250_/C vdd NAND2X1
XFILL_4__12312_ gnd vdd FILL
XFILL_5__14651_ gnd vdd FILL
XFILL_4__13292_ gnd vdd FILL
XFILL_2__10703_ gnd vdd FILL
XFILL_2__8345_ gnd vdd FILL
XFILL_3__15830_ gnd vdd FILL
XFILL_5__11863_ gnd vdd FILL
XFILL_4__16080_ gnd vdd FILL
XFILL_2__14471_ gnd vdd FILL
XFILL_1__12132_ gnd vdd FILL
XFILL_0__15650_ gnd vdd FILL
XFILL_2__11683_ gnd vdd FILL
XFILL_5__8054_ gnd vdd FILL
XFILL_5__13602_ gnd vdd FILL
XFILL_0__12862_ gnd vdd FILL
XFILL_5__10814_ gnd vdd FILL
XFILL_2__16210_ gnd vdd FILL
XFILL_0__7360_ gnd vdd FILL
XFILL_4__15031_ gnd vdd FILL
XFILL_4__12243_ gnd vdd FILL
XFILL_5__14582_ gnd vdd FILL
XFILL_2__13422_ gnd vdd FILL
XSFILL53800x48050 gnd vdd FILL
XFILL_0__14601_ gnd vdd FILL
XFILL_2__10634_ gnd vdd FILL
XFILL_2__8276_ gnd vdd FILL
XFILL_5__11794_ gnd vdd FILL
XFILL_3__15761_ gnd vdd FILL
XFILL_3__12973_ gnd vdd FILL
XFILL_1__12063_ gnd vdd FILL
XFILL_0__11813_ gnd vdd FILL
XSFILL109320x77050 gnd vdd FILL
XFILL_5__16321_ gnd vdd FILL
XFILL_0__15581_ gnd vdd FILL
XFILL_5__13533_ gnd vdd FILL
XFILL_2__7227_ gnd vdd FILL
XFILL_3__14712_ gnd vdd FILL
XFILL_4__12174_ gnd vdd FILL
XFILL_5__10745_ gnd vdd FILL
XFILL_2__16141_ gnd vdd FILL
XFILL_0__7291_ gnd vdd FILL
XFILL_2__13353_ gnd vdd FILL
X_14988_ _12813_/Q _12812_/Q gnd _15061_/C vdd AND2X2
XFILL_3__11924_ gnd vdd FILL
XFILL_1__11014_ gnd vdd FILL
XSFILL28600x24050 gnd vdd FILL
XFILL_3__15692_ gnd vdd FILL
XFILL_0__14532_ gnd vdd FILL
XFILL_2__10565_ gnd vdd FILL
XFILL_0__9030_ gnd vdd FILL
XFILL_0__11744_ gnd vdd FILL
XFILL_3_CLKBUF1_insert160 gnd vdd FILL
XFILL_4__11125_ gnd vdd FILL
XFILL_5__16252_ gnd vdd FILL
XFILL_5__13464_ gnd vdd FILL
XFILL_2__12304_ gnd vdd FILL
XFILL_3_CLKBUF1_insert171 gnd vdd FILL
X_13939_ _7520_/Q gnd _13940_/D vdd INVX1
XFILL_3__14643_ gnd vdd FILL
XFILL_2__7158_ gnd vdd FILL
X_6870_ _6870_/A gnd memoryWriteData[0] vdd BUFX2
XFILL_1__15822_ gnd vdd FILL
XFILL_2__16072_ gnd vdd FILL
XFILL_5__10676_ gnd vdd FILL
XFILL_3__11855_ gnd vdd FILL
XFILL_2__13284_ gnd vdd FILL
XFILL_3_CLKBUF1_insert182 gnd vdd FILL
XFILL_3_CLKBUF1_insert193 gnd vdd FILL
XFILL_2__10496_ gnd vdd FILL
XFILL_0__14463_ gnd vdd FILL
XFILL_5__15203_ gnd vdd FILL
XSFILL114440x68050 gnd vdd FILL
XFILL_5__12415_ gnd vdd FILL
XFILL_5__8956_ gnd vdd FILL
XFILL_0__11675_ gnd vdd FILL
XFILL_5__16183_ gnd vdd FILL
XFILL_4__15933_ gnd vdd FILL
XFILL_2__15023_ gnd vdd FILL
XFILL_4__11056_ gnd vdd FILL
XFILL_3__10806_ gnd vdd FILL
XFILL_0__16202_ gnd vdd FILL
XFILL_5__13395_ gnd vdd FILL
XFILL_2__12235_ gnd vdd FILL
XFILL_3__14574_ gnd vdd FILL
XFILL_0__13414_ gnd vdd FILL
XFILL_2__7089_ gnd vdd FILL
XSFILL33720x15050 gnd vdd FILL
XFILL_3__11786_ gnd vdd FILL
XFILL_1__15753_ gnd vdd FILL
XFILL_3__7971_ gnd vdd FILL
XFILL_0__10626_ gnd vdd FILL
XFILL_1__12965_ gnd vdd FILL
XSFILL115080x34050 gnd vdd FILL
XFILL_4__10007_ gnd vdd FILL
XFILL_0__14394_ gnd vdd FILL
XSFILL48920x6050 gnd vdd FILL
X_15609_ _15609_/A _15609_/B _15609_/C gnd _15610_/B vdd NOR3X1
XFILL_5__15134_ gnd vdd FILL
XFILL_6__13705_ gnd vdd FILL
XFILL_5__8887_ gnd vdd FILL
X_8540_ _8540_/Q _7534_/CLK _8156_/R vdd _8540_/D gnd vdd DFFSR
XFILL_5__12346_ gnd vdd FILL
XFILL_1_BUFX2_insert370 gnd vdd FILL
XFILL_3__16313_ gnd vdd FILL
XFILL_1_BUFX2_insert381 gnd vdd FILL
XFILL_1__14704_ gnd vdd FILL
XFILL_4__15864_ gnd vdd FILL
XFILL_3__13525_ gnd vdd FILL
XFILL_3__6922_ gnd vdd FILL
XFILL_1_BUFX2_insert392 gnd vdd FILL
XFILL_1__11916_ gnd vdd FILL
XFILL_2__12166_ gnd vdd FILL
XFILL_0__16133_ gnd vdd FILL
XFILL_0__13345_ gnd vdd FILL
XFILL_1__15684_ gnd vdd FILL
XFILL_1__12896_ gnd vdd FILL
XFILL_0__10557_ gnd vdd FILL
XFILL_5_BUFX2_insert708 gnd vdd FILL
XFILL_5__7838_ gnd vdd FILL
XSFILL59160x26050 gnd vdd FILL
XFILL_4__14815_ gnd vdd FILL
XFILL_0__9932_ gnd vdd FILL
XFILL_5__15065_ gnd vdd FILL
XFILL_3__16244_ gnd vdd FILL
X_8471_ _8545_/Q gnd _8471_/Y vdd INVX1
XFILL_5_BUFX2_insert719 gnd vdd FILL
XFILL_5__12277_ gnd vdd FILL
XFILL_2__11117_ gnd vdd FILL
XFILL_1__14635_ gnd vdd FILL
XFILL_3__6853_ gnd vdd FILL
XFILL_3__13456_ gnd vdd FILL
XFILL_4__15795_ gnd vdd FILL
XFILL_3__10668_ gnd vdd FILL
XFILL_3__9641_ gnd vdd FILL
XFILL_2__12097_ gnd vdd FILL
XFILL_0__16064_ gnd vdd FILL
XFILL_1__11847_ gnd vdd FILL
XFILL_0__13276_ gnd vdd FILL
XFILL_0__10488_ gnd vdd FILL
XFILL_5__14016_ gnd vdd FILL
XFILL_6__16355_ gnd vdd FILL
XFILL_6__13567_ gnd vdd FILL
X_7422_ _7422_/A _7470_/B _7421_/Y gnd _7512_/D vdd OAI21X1
XFILL_5__11228_ gnd vdd FILL
XFILL111880x25050 gnd vdd FILL
XFILL_3__12407_ gnd vdd FILL
XFILL_0__9863_ gnd vdd FILL
XFILL_4__14746_ gnd vdd FILL
XFILL_2__15925_ gnd vdd FILL
XFILL_3__16175_ gnd vdd FILL
XFILL_4__11958_ gnd vdd FILL
XFILL_3__13387_ gnd vdd FILL
XFILL_0__15015_ gnd vdd FILL
XFILL_2__11048_ gnd vdd FILL
XFILL_5__9508_ gnd vdd FILL
XFILL_1__14566_ gnd vdd FILL
XFILL_0__12227_ gnd vdd FILL
XFILL_6__15306_ gnd vdd FILL
XFILL_1__11778_ gnd vdd FILL
XFILL_6__9281_ gnd vdd FILL
XFILL_4__10909_ gnd vdd FILL
X_7353_ _7354_/B _9657_/B gnd _7353_/Y vdd NAND2X1
XFILL_1__16305_ gnd vdd FILL
XFILL_3__12338_ gnd vdd FILL
XFILL_0__9794_ gnd vdd FILL
XFILL_5__11159_ gnd vdd FILL
XFILL_3__15126_ gnd vdd FILL
XSFILL109400x57050 gnd vdd FILL
XFILL_3__8523_ gnd vdd FILL
XFILL_4__14677_ gnd vdd FILL
XFILL_1__13517_ gnd vdd FILL
XFILL_4__11889_ gnd vdd FILL
XFILL_2__15856_ gnd vdd FILL
XFILL_1__14497_ gnd vdd FILL
XFILL_6__8232_ gnd vdd FILL
XFILL_0__12158_ gnd vdd FILL
XFILL_6__12449_ gnd vdd FILL
XFILL_4__16416_ gnd vdd FILL
XFILL_0__8745_ gnd vdd FILL
XSFILL49080x78050 gnd vdd FILL
XFILL_4__13628_ gnd vdd FILL
XFILL_1__16236_ gnd vdd FILL
XFILL_2__14807_ gnd vdd FILL
XFILL_3__15057_ gnd vdd FILL
XFILL_5__15967_ gnd vdd FILL
XFILL_3__12269_ gnd vdd FILL
XFILL_3__8454_ gnd vdd FILL
X_7284_ _7248_/A _9194_/CLK _7775_/R vdd _7284_/D gnd vdd DFFSR
XFILL_1__13448_ gnd vdd FILL
XFILL_0__11109_ gnd vdd FILL
XFILL_0__12089_ gnd vdd FILL
XFILL_2__12999_ gnd vdd FILL
XFILL_2__15787_ gnd vdd FILL
XSFILL64120x81050 gnd vdd FILL
XFILL_6__15168_ gnd vdd FILL
X_9023_ _8996_/A _8511_/B gnd _9024_/C vdd NAND2X1
XFILL_4__16347_ gnd vdd FILL
XFILL_3__14008_ gnd vdd FILL
XFILL_5__14918_ gnd vdd FILL
XFILL_5__15898_ gnd vdd FILL
XSFILL104440x50 gnd vdd FILL
XFILL_4__13559_ gnd vdd FILL
XFILL_0__15917_ gnd vdd FILL
XFILL_1__16167_ gnd vdd FILL
XSFILL114520x48050 gnd vdd FILL
XFILL_2__14738_ gnd vdd FILL
XFILL_3__8385_ gnd vdd FILL
XSFILL74120x1050 gnd vdd FILL
XFILL_1__13379_ gnd vdd FILL
XFILL_6__14119_ gnd vdd FILL
XFILL_0__7627_ gnd vdd FILL
XFILL_5__14849_ gnd vdd FILL
XFILL_3__7336_ gnd vdd FILL
XFILL_1__15118_ gnd vdd FILL
XFILL_4__16278_ gnd vdd FILL
XFILL_1__16098_ gnd vdd FILL
XFILL_0__15848_ gnd vdd FILL
XFILL_2__14669_ gnd vdd FILL
XFILL_4__15229_ gnd vdd FILL
XFILL_0__7558_ gnd vdd FILL
XFILL_2__16408_ gnd vdd FILL
XFILL_2_BUFX2_insert609 gnd vdd FILL
XFILL_1__15049_ gnd vdd FILL
XFILL_3__15959_ gnd vdd FILL
XFILL_0__15779_ gnd vdd FILL
X_9925_ _9868_/A _9413_/B gnd _9925_/Y vdd NAND2X1
XFILL_3__9006_ gnd vdd FILL
XFILL_0__7489_ gnd vdd FILL
XFILL_2__16339_ gnd vdd FILL
XFILL_3__7198_ gnd vdd FILL
XFILL_0__9228_ gnd vdd FILL
XFILL_1__8021_ gnd vdd FILL
X_9856_ _9917_/B _9600_/B gnd _9857_/C vdd NAND2X1
XSFILL23720x47050 gnd vdd FILL
XFILL_0__9159_ gnd vdd FILL
X_8807_ _8745_/A _8551_/CLK _9064_/R vdd _8807_/D gnd vdd DFFSR
XFILL112040x14050 gnd vdd FILL
X_9787_ _9837_/Q gnd _9787_/Y vdd INVX1
XSFILL64600x59050 gnd vdd FILL
X_6999_ _6999_/Q _6999_/CLK _7000_/R vdd _6999_/D gnd vdd DFFSR
XFILL_6_BUFX2_insert531 gnd vdd FILL
XFILL_4__9750_ gnd vdd FILL
XFILL_4__6962_ gnd vdd FILL
X_8738_ _8736_/Y _8759_/B _8738_/C gnd _8804_/D vdd OAI21X1
XBUFX2_insert608 _15035_/Y gnd _15708_/A vdd BUFX2
XFILL_3__9908_ gnd vdd FILL
XBUFX2_insert619 _13430_/Y gnd _14458_/C vdd BUFX2
XFILL_4__8701_ gnd vdd FILL
XFILL_4__6893_ gnd vdd FILL
XFILL_6__9617_ gnd vdd FILL
XFILL_4__9681_ gnd vdd FILL
XSFILL79000x21050 gnd vdd FILL
XFILL_6_BUFX2_insert597 gnd vdd FILL
X_8669_ _8669_/Q _7915_/CLK _8669_/R vdd _8589_/Y gnd vdd DFFSR
XFILL_4__8632_ gnd vdd FILL
XFILL_1__8854_ gnd vdd FILL
X_12270_ _12267_/Y _12270_/B _12270_/C gnd _12270_/Y vdd NAND3X1
XFILL_1__7805_ gnd vdd FILL
XFILL_1__8785_ gnd vdd FILL
XSFILL28840x80050 gnd vdd FILL
XFILL_4__8494_ gnd vdd FILL
X_11221_ _10889_/Y _10882_/Y gnd _11227_/A vdd NOR2X1
XFILL_1__7736_ gnd vdd FILL
XFILL_4__7445_ gnd vdd FILL
X_11152_ _12171_/Y gnd _11153_/B vdd INVX1
XSFILL8760x78050 gnd vdd FILL
XSFILL23800x27050 gnd vdd FILL
XFILL_3_BUFX2_insert410 gnd vdd FILL
XFILL_3_BUFX2_insert421 gnd vdd FILL
X_10103_ _8951_/A _10140_/B gnd _10103_/Y vdd NAND2X1
XFILL_4__7376_ gnd vdd FILL
XSFILL33960x71050 gnd vdd FILL
XFILL_1__9406_ gnd vdd FILL
X_15960_ _9964_/Q gnd _15961_/D vdd INVX1
X_11083_ _12150_/Y gnd _11083_/Y vdd INVX2
XFILL_3_BUFX2_insert432 gnd vdd FILL
XFILL_3_BUFX2_insert443 gnd vdd FILL
XFILL_3_BUFX2_insert454 gnd vdd FILL
XFILL_4__9115_ gnd vdd FILL
XFILL_1__7598_ gnd vdd FILL
XFILL_3_BUFX2_insert465 gnd vdd FILL
X_10034_ _14442_/A gnd _10034_/Y vdd INVX1
X_14911_ _9552_/A gnd _14911_/Y vdd INVX1
XFILL_3_BUFX2_insert476 gnd vdd FILL
XFILL_2__8130_ gnd vdd FILL
XFILL_3_BUFX2_insert487 gnd vdd FILL
XFILL_1__9337_ gnd vdd FILL
X_15891_ _15891_/A _15891_/B _14402_/C gnd _12884_/B vdd AOI21X1
XFILL_3_BUFX2_insert498 gnd vdd FILL
X_14842_ _10483_/Q gnd _14842_/Y vdd INVX1
XSFILL74280x7050 gnd vdd FILL
XFILL_1__9268_ gnd vdd FILL
XFILL_2__8061_ gnd vdd FILL
XSFILL58920x1050 gnd vdd FILL
XFILL_5__10530_ gnd vdd FILL
XFILL_1__8219_ gnd vdd FILL
X_11985_ _12047_/A gnd _11985_/Y vdd INVX8
X_14773_ _7367_/A _14353_/A _14847_/C _7153_/Q gnd _14775_/A vdd AOI22X1
XFILL_0_BUFX2_insert4 gnd vdd FILL
XFILL_5__9790_ gnd vdd FILL
X_10936_ _12773_/A _10936_/B _10936_/C gnd _10945_/C vdd NAND3X1
X_13724_ _8283_/Q gnd _13725_/A vdd INVX1
XSFILL28920x60050 gnd vdd FILL
XFILL_3__11640_ gnd vdd FILL
XFILL_4_CLKBUF1_insert200 gnd vdd FILL
XFILL_4_CLKBUF1_insert211 gnd vdd FILL
XFILL_2__10281_ gnd vdd FILL
XFILL_0__11460_ gnd vdd FILL
XFILL_5__8741_ gnd vdd FILL
XFILL_5__12200_ gnd vdd FILL
XFILL_4_CLKBUF1_insert222 gnd vdd FILL
X_16443_ _14713_/A _8289_/CLK _8688_/R vdd _16443_/D gnd vdd DFFSR
X_10867_ _10867_/Q _8051_/CLK _7789_/R vdd _10831_/Y gnd vdd DFFSR
X_13655_ _13651_/Y _13655_/B gnd _13663_/B vdd NOR2X1
XFILL_2__12020_ gnd vdd FILL
XFILL_5__10392_ gnd vdd FILL
XFILL_3__11571_ gnd vdd FILL
XFILL_1__12750_ gnd vdd FILL
XFILL_0_BUFX2_insert300 gnd vdd FILL
XFILL_2__8963_ gnd vdd FILL
XFILL_0__10411_ gnd vdd FILL
XFILL_0__11391_ gnd vdd FILL
XFILL_0_BUFX2_insert311 gnd vdd FILL
X_12606_ _12676_/Q gnd _12606_/Y vdd INVX1
XFILL_4__9879_ gnd vdd FILL
XFILL_5__12131_ gnd vdd FILL
X_13586_ _7769_/Q gnd _13586_/Y vdd INVX1
XFILL_3__13310_ gnd vdd FILL
XFILL_0_BUFX2_insert322 gnd vdd FILL
XFILL_3__10522_ gnd vdd FILL
X_16374_ _16374_/A gnd _16374_/C gnd _16434_/D vdd OAI21X1
XFILL_4__12861_ gnd vdd FILL
X_10798_ _10798_/A _10797_/A _10798_/C gnd _10798_/Y vdd OAI21X1
XFILL_3__14290_ gnd vdd FILL
XFILL_1__11701_ gnd vdd FILL
XFILL_0_BUFX2_insert333 gnd vdd FILL
XFILL_0__13130_ gnd vdd FILL
XFILL_0_BUFX2_insert344 gnd vdd FILL
XFILL_2__8894_ gnd vdd FILL
XFILL_0_BUFX2_insert355 gnd vdd FILL
XFILL_5__7623_ gnd vdd FILL
XFILL_4__14600_ gnd vdd FILL
X_15325_ _16339_/A _15680_/B _15680_/C gnd _15336_/C vdd NAND3X1
X_12537_ _12349_/A _12537_/CLK _9060_/R vdd _12447_/Y gnd vdd DFFSR
XSFILL99480x46050 gnd vdd FILL
XFILL_0_BUFX2_insert366 gnd vdd FILL
XFILL_3__13241_ gnd vdd FILL
XFILL_5__12062_ gnd vdd FILL
XSFILL74120x44050 gnd vdd FILL
XFILL_4__11812_ gnd vdd FILL
XFILL_3__10453_ gnd vdd FILL
XFILL_0_BUFX2_insert377 gnd vdd FILL
XFILL_1__14420_ gnd vdd FILL
XFILL_4__15580_ gnd vdd FILL
XFILL_0_BUFX2_insert388 gnd vdd FILL
XFILL_2__7845_ gnd vdd FILL
XFILL_1__11632_ gnd vdd FILL
XFILL_2__13971_ gnd vdd FILL
XFILL_0__10273_ gnd vdd FILL
XFILL_0_BUFX2_insert399 gnd vdd FILL
XFILL_6__16140_ gnd vdd FILL
XFILL_6__13352_ gnd vdd FILL
XFILL_5__7554_ gnd vdd FILL
XFILL_5__11013_ gnd vdd FILL
X_15256_ _15253_/Y _15256_/B gnd _15257_/B vdd NOR2X1
XFILL_0__6860_ gnd vdd FILL
X_12468_ _12468_/A vdd _12467_/Y gnd _12468_/Y vdd OAI21X1
XFILL_4__14531_ gnd vdd FILL
XFILL_2__15710_ gnd vdd FILL
XFILL_3__13172_ gnd vdd FILL
XFILL_4__11743_ gnd vdd FILL
XFILL_3__10384_ gnd vdd FILL
XFILL_0__12012_ gnd vdd FILL
XFILL_1__14351_ gnd vdd FILL
XSFILL108840x65050 gnd vdd FILL
XFILL_1__11563_ gnd vdd FILL
XFILL_5__7485_ gnd vdd FILL
X_14207_ _8549_/Q gnd _14207_/Y vdd INVX1
X_11419_ _11419_/A _11204_/Y _11207_/B gnd _11419_/Y vdd NAND3X1
X_15187_ _15187_/A _15187_/B _15187_/C gnd _15187_/Y vdd NOR3X1
XFILL_5__15821_ gnd vdd FILL
XFILL_3__12123_ gnd vdd FILL
XFILL_1__13302_ gnd vdd FILL
XFILL_4__14462_ gnd vdd FILL
X_12399_ _12397_/Y _12359_/A _12399_/C gnd _12399_/Y vdd OAI21X1
XFILL_2__9515_ gnd vdd FILL
XFILL_2__15641_ gnd vdd FILL
XFILL_4__11674_ gnd vdd FILL
XFILL_2__12853_ gnd vdd FILL
XFILL_1__10514_ gnd vdd FILL
XFILL_5__9224_ gnd vdd FILL
XFILL_1__14282_ gnd vdd FILL
XFILL_4__16201_ gnd vdd FILL
X_14138_ _14138_/A _14479_/B _14555_/C _14137_/Y gnd _14138_/Y vdd OAI22X1
XFILL_6__12234_ gnd vdd FILL
XFILL_1__11494_ gnd vdd FILL
XFILL_0__8530_ gnd vdd FILL
XFILL_4__13413_ gnd vdd FILL
XFILL_5__15752_ gnd vdd FILL
XFILL_4__10625_ gnd vdd FILL
XFILL_1__16021_ gnd vdd FILL
XFILL_5__12964_ gnd vdd FILL
XFILL_3__12054_ gnd vdd FILL
XFILL_2__11804_ gnd vdd FILL
XFILL_1__13233_ gnd vdd FILL
XFILL_4__14393_ gnd vdd FILL
XSFILL54040x11050 gnd vdd FILL
XFILL_2__12784_ gnd vdd FILL
XFILL_1__10445_ gnd vdd FILL
XFILL_5_BUFX2_insert1001 gnd vdd FILL
XFILL_2__15572_ gnd vdd FILL
XFILL_5_BUFX2_insert1012 gnd vdd FILL
XFILL_5__14703_ gnd vdd FILL
XFILL_5__9155_ gnd vdd FILL
XFILL_0__13963_ gnd vdd FILL
XFILL_0__8461_ gnd vdd FILL
XFILL_5__11915_ gnd vdd FILL
X_14069_ _15547_/A gnd _14069_/Y vdd INVX1
XFILL_5_BUFX2_insert1023 gnd vdd FILL
XFILL_3__11005_ gnd vdd FILL
XFILL_4__16132_ gnd vdd FILL
XFILL_4__13344_ gnd vdd FILL
XFILL_5__15683_ gnd vdd FILL
XFILL_5_BUFX2_insert1034 gnd vdd FILL
XFILL_0__15702_ gnd vdd FILL
XFILL_5__12895_ gnd vdd FILL
XFILL_4__10556_ gnd vdd FILL
XFILL_2__14523_ gnd vdd FILL
XFILL_2__11735_ gnd vdd FILL
XFILL_2__9377_ gnd vdd FILL
XFILL_1__13164_ gnd vdd FILL
XFILL_0__12914_ gnd vdd FILL
XFILL_5__8106_ gnd vdd FILL
XFILL_5_BUFX2_insert1045 gnd vdd FILL
XFILL_1__10376_ gnd vdd FILL
XFILL_5_BUFX2_insert1056 gnd vdd FILL
XFILL_5__14634_ gnd vdd FILL
XFILL_5_BUFX2_insert1067 gnd vdd FILL
XFILL_0__13894_ gnd vdd FILL
XFILL_5__9086_ gnd vdd FILL
XFILL_6__12096_ gnd vdd FILL
XFILL_3__15813_ gnd vdd FILL
XFILL_4__16063_ gnd vdd FILL
XFILL_3__7121_ gnd vdd FILL
XFILL_0__8392_ gnd vdd FILL
XFILL_5__11846_ gnd vdd FILL
XFILL_5_BUFX2_insert1089 gnd vdd FILL
XFILL_4__13275_ gnd vdd FILL
XFILL_2__14454_ gnd vdd FILL
XSFILL114040x65050 gnd vdd FILL
XFILL_2__8328_ gnd vdd FILL
XFILL_1__12115_ gnd vdd FILL
XSFILL43880x54050 gnd vdd FILL
XFILL_4__10487_ gnd vdd FILL
XFILL_0__15633_ gnd vdd FILL
XFILL_2__11666_ gnd vdd FILL
XFILL_0__12845_ gnd vdd FILL
XFILL_1__13095_ gnd vdd FILL
XFILL_4__15014_ gnd vdd FILL
XFILL_0__7343_ gnd vdd FILL
XFILL_6__11047_ gnd vdd FILL
XFILL_5__14565_ gnd vdd FILL
XFILL_2__13405_ gnd vdd FILL
XFILL_4__12226_ gnd vdd FILL
XFILL_3__7052_ gnd vdd FILL
X_7971_ _7971_/A gnd _7973_/A vdd INVX1
XSFILL58120x57050 gnd vdd FILL
XSFILL18680x30050 gnd vdd FILL
XFILL_2__8259_ gnd vdd FILL
XFILL_2__10617_ gnd vdd FILL
XFILL_5__11777_ gnd vdd FILL
XFILL_3__15744_ gnd vdd FILL
XSFILL58920x76050 gnd vdd FILL
XFILL_1__12046_ gnd vdd FILL
XFILL_2__14385_ gnd vdd FILL
XFILL_3__12956_ gnd vdd FILL
XFILL_0__15564_ gnd vdd FILL
XFILL_5__16304_ gnd vdd FILL
XFILL_2__11597_ gnd vdd FILL
XSFILL74200x24050 gnd vdd FILL
XFILL_0__12776_ gnd vdd FILL
X_9710_ _9710_/Q _8046_/CLK _9061_/R vdd _9710_/D gnd vdd DFFSR
XFILL_5__13516_ gnd vdd FILL
X_6922_ _6920_/Y _6988_/B _6922_/C gnd _7004_/D vdd OAI21X1
XFILL_2__13336_ gnd vdd FILL
XFILL_5__14496_ gnd vdd FILL
XFILL_3__11907_ gnd vdd FILL
XFILL_4__12157_ gnd vdd FILL
XFILL_2__16124_ gnd vdd FILL
XFILL_3__15675_ gnd vdd FILL
XFILL_0__14515_ gnd vdd FILL
XFILL_2__10548_ gnd vdd FILL
XFILL_0__9013_ gnd vdd FILL
XFILL_3__12887_ gnd vdd FILL
XFILL_0__11727_ gnd vdd FILL
XFILL_5__16235_ gnd vdd FILL
XFILL_0__15495_ gnd vdd FILL
XFILL_5__9988_ gnd vdd FILL
XFILL_5__13447_ gnd vdd FILL
XFILL_4__11108_ gnd vdd FILL
X_9641_ _9641_/A gnd _9641_/Y vdd INVX1
XFILL_5__10659_ gnd vdd FILL
XFILL_3__14626_ gnd vdd FILL
X_6853_ _6853_/A gnd memoryAddress[15] vdd BUFX2
XFILL_4__12088_ gnd vdd FILL
XFILL_2__16055_ gnd vdd FILL
XFILL_2__13267_ gnd vdd FILL
XFILL_3_BUFX2_insert1060 gnd vdd FILL
XFILL_1__15805_ gnd vdd FILL
XFILL_3__11838_ gnd vdd FILL
XFILL_3_BUFX2_insert1071 gnd vdd FILL
XFILL_0__14446_ gnd vdd FILL
XFILL_1__13997_ gnd vdd FILL
XFILL_0__11658_ gnd vdd FILL
XFILL_4__15916_ gnd vdd FILL
XFILL_5__16166_ gnd vdd FILL
XFILL_2__15006_ gnd vdd FILL
XFILL_3_BUFX2_insert1093 gnd vdd FILL
XFILL_4__11039_ gnd vdd FILL
X_9572_ _9572_/Q _9707_/CLK _8801_/R vdd _9572_/D gnd vdd DFFSR
XFILL_5__13378_ gnd vdd FILL
XFILL_2__12218_ gnd vdd FILL
XFILL_3__14557_ gnd vdd FILL
XFILL_3__7954_ gnd vdd FILL
XFILL_3__11769_ gnd vdd FILL
XFILL_1__15736_ gnd vdd FILL
XFILL_0__14377_ gnd vdd FILL
XFILL_5__15117_ gnd vdd FILL
XFILL112360x50050 gnd vdd FILL
X_8523_ _8440_/B _8011_/B gnd _8524_/C vdd NAND2X1
XFILL_5__12329_ gnd vdd FILL
XFILL_0__11589_ gnd vdd FILL
XSFILL89960x50 gnd vdd FILL
XSFILL64120x76050 gnd vdd FILL
XFILL_5_BUFX2_insert505 gnd vdd FILL
XFILL_5__16097_ gnd vdd FILL
XFILL_4__15847_ gnd vdd FILL
XFILL_3__13508_ gnd vdd FILL
XFILL_0__16116_ gnd vdd FILL
XFILL_5_BUFX2_insert516 gnd vdd FILL
XFILL_2__12149_ gnd vdd FILL
XFILL_3__6905_ gnd vdd FILL
XFILL_0__13328_ gnd vdd FILL
XFILL_3__14488_ gnd vdd FILL
XFILL_1__15667_ gnd vdd FILL
XFILL_5_BUFX2_insert527 gnd vdd FILL
XFILL_3__7885_ gnd vdd FILL
XFILL_1__12879_ gnd vdd FILL
XFILL_0__9915_ gnd vdd FILL
XFILL_5__15048_ gnd vdd FILL
XFILL_5_BUFX2_insert538 gnd vdd FILL
XFILL_5_BUFX2_insert549 gnd vdd FILL
XFILL_3__16227_ gnd vdd FILL
X_8454_ _8494_/B _8582_/B gnd _8455_/C vdd NAND2X1
XFILL_1__14618_ gnd vdd FILL
XFILL_3__9624_ gnd vdd FILL
XFILL_3__13439_ gnd vdd FILL
XFILL_4__15778_ gnd vdd FILL
XFILL_3__6836_ gnd vdd FILL
XFILL_0__16047_ gnd vdd FILL
XFILL_0__13259_ gnd vdd FILL
XFILL_3_BUFX2_insert8 gnd vdd FILL
XFILL_1__15598_ gnd vdd FILL
X_7405_ _7355_/A _7411_/CLK _7411_/R vdd _7405_/D gnd vdd DFFSR
XSFILL43960x34050 gnd vdd FILL
XSFILL3560x83050 gnd vdd FILL
XFILL_0__9846_ gnd vdd FILL
XFILL_4__14729_ gnd vdd FILL
XSFILL68760x79050 gnd vdd FILL
XFILL_2__15908_ gnd vdd FILL
X_8385_ _8385_/A gnd _8385_/Y vdd INVX1
XSFILL69080x8050 gnd vdd FILL
XFILL_3__16158_ gnd vdd FILL
XFILL_1__14549_ gnd vdd FILL
XFILL_3__9555_ gnd vdd FILL
XSFILL108680x8050 gnd vdd FILL
XSFILL18760x10050 gnd vdd FILL
X_7336_ _7334_/Y _7336_/B _7336_/C gnd _7336_/Y vdd OAI21X1
XFILL_3_BUFX2_insert60 gnd vdd FILL
XFILL_1__8570_ gnd vdd FILL
XFILL_3__15109_ gnd vdd FILL
XFILL_0__6989_ gnd vdd FILL
XFILL_3__8506_ gnd vdd FILL
XFILL_0__9777_ gnd vdd FILL
XSFILL8600x20050 gnd vdd FILL
XSFILL68360x81050 gnd vdd FILL
XSFILL44040x43050 gnd vdd FILL
XFILL_3__16089_ gnd vdd FILL
XFILL_3_BUFX2_insert71 gnd vdd FILL
XFILL_2__15839_ gnd vdd FILL
XFILL_3__9486_ gnd vdd FILL
XFILL_3_BUFX2_insert82 gnd vdd FILL
XFILL_3_BUFX2_insert93 gnd vdd FILL
XFILL_0__8728_ gnd vdd FILL
XFILL_4__7230_ gnd vdd FILL
XFILL_2_CLKBUF1_insert119 gnd vdd FILL
XFILL_1__16219_ gnd vdd FILL
X_7267_ _7197_/A _9077_/CLK _7515_/R vdd _7199_/Y gnd vdd DFFSR
XSFILL84280x2050 gnd vdd FILL
X_9006_ _9004_/Y _9005_/A _9006_/C gnd _9064_/D vdd OAI21X1
XFILL_1__7452_ gnd vdd FILL
XFILL_0__8659_ gnd vdd FILL
X_7198_ _7166_/B _7326_/B gnd _7199_/C vdd NAND2X1
XFILL_4__7161_ gnd vdd FILL
XFILL_3__8368_ gnd vdd FILL
XFILL111800x64050 gnd vdd FILL
XFILL_6__8077_ gnd vdd FILL
XFILL_2_BUFX2_insert406 gnd vdd FILL
XFILL_3__7319_ gnd vdd FILL
XFILL112440x30050 gnd vdd FILL
XFILL_4__7092_ gnd vdd FILL
XFILL_2_BUFX2_insert417 gnd vdd FILL
XFILL_1__9122_ gnd vdd FILL
XSFILL64200x56050 gnd vdd FILL
XFILL_2_BUFX2_insert428 gnd vdd FILL
XSFILL79000x16050 gnd vdd FILL
XSFILL49560x74050 gnd vdd FILL
XFILL_2_BUFX2_insert439 gnd vdd FILL
X_9908_ _9908_/A _9896_/B _9907_/Y gnd _9908_/Y vdd OAI21X1
XSFILL3640x63050 gnd vdd FILL
XFILL_1__8004_ gnd vdd FILL
X_11770_ _11245_/Y _11770_/B _11835_/C gnd _11771_/C vdd AOI21X1
X_9839_ _9839_/Q _7647_/CLK _9823_/R vdd _9839_/D gnd vdd DFFSR
XFILL_4__9802_ gnd vdd FILL
XSFILL28840x75050 gnd vdd FILL
X_10721_ _10647_/A _9953_/CLK _9580_/R vdd _10721_/D gnd vdd DFFSR
XSFILL94280x51050 gnd vdd FILL
XFILL_4__7994_ gnd vdd FILL
XBUFX2_insert405 _10920_/Y gnd _12395_/A vdd BUFX2
XFILL_4__9733_ gnd vdd FILL
XBUFX2_insert416 _15050_/Y gnd _15899_/A vdd BUFX2
XFILL_4__6945_ gnd vdd FILL
X_13440_ _9686_/Q gnd _13444_/A vdd INVX1
XFILL_6_BUFX2_insert372 gnd vdd FILL
X_10652_ _10650_/Y _10615_/B _10652_/C gnd _10652_/Y vdd OAI21X1
XBUFX2_insert427 _15047_/Y gnd _15813_/C vdd BUFX2
XBUFX2_insert438 _15086_/Y gnd _15383_/A vdd BUFX2
XSFILL44040x5050 gnd vdd FILL
XBUFX2_insert449 _13276_/Y gnd _7207_/A vdd BUFX2
XFILL_4__9664_ gnd vdd FILL
X_13371_ _12807_/Q _13371_/B gnd _13423_/B vdd NOR2X1
XFILL_4__6876_ gnd vdd FILL
XFILL_1__8906_ gnd vdd FILL
X_10583_ _15122_/A _8152_/CLK _8664_/R vdd _10583_/D gnd vdd DFFSR
XFILL_4__8615_ gnd vdd FILL
XFILL_1__9886_ gnd vdd FILL
X_12322_ _12322_/A _12320_/Y _12322_/C gnd _12322_/Y vdd NAND3X1
X_15110_ _15802_/A _13499_/Y _15110_/C _15774_/C gnd _15110_/Y vdd OAI22X1
X_16090_ _16090_/A _15342_/B gnd _16093_/B vdd NOR2X1
XFILL_4__9595_ gnd vdd FILL
XFILL_2__7630_ gnd vdd FILL
XFILL_1__8837_ gnd vdd FILL
XSFILL88600x74050 gnd vdd FILL
X_15041_ _15040_/Y _15245_/B gnd _15041_/Y vdd OR2X2
X_12253_ _6879_/A _12237_/B _12269_/C _12716_/A gnd _12253_/Y vdd AOI22X1
XFILL_2__7561_ gnd vdd FILL
XSFILL89240x40050 gnd vdd FILL
XFILL_1__8768_ gnd vdd FILL
XSFILL53880x17050 gnd vdd FILL
X_11204_ _11203_/Y _11202_/Y gnd _11204_/Y vdd NOR2X1
XFILL_4__8477_ gnd vdd FILL
X_12184_ _12184_/A gnd _12184_/Y vdd INVX1
XFILL_2__9300_ gnd vdd FILL
XFILL_1__7719_ gnd vdd FILL
XSFILL3720x43050 gnd vdd FILL
XFILL_2__7492_ gnd vdd FILL
XFILL_4__7428_ gnd vdd FILL
XFILL_1__8699_ gnd vdd FILL
X_11135_ _12165_/Y gnd _11617_/A vdd INVX2
XFILL_4__10410_ gnd vdd FILL
XFILL_2__9231_ gnd vdd FILL
XFILL_4__11390_ gnd vdd FILL
XSFILL28920x55050 gnd vdd FILL
XFILL_3_BUFX2_insert240 gnd vdd FILL
XFILL_1__10230_ gnd vdd FILL
XFILL_0__10960_ gnd vdd FILL
XFILL_4__7359_ gnd vdd FILL
XFILL_5__11700_ gnd vdd FILL
XFILL_3_BUFX2_insert251 gnd vdd FILL
X_15943_ _15943_/A _15943_/B gnd _15968_/A vdd NOR2X1
XFILL_3_BUFX2_insert262 gnd vdd FILL
X_11066_ _12266_/Y _12153_/Y gnd _11066_/Y vdd NOR2X1
XFILL_3_BUFX2_insert273 gnd vdd FILL
XFILL_2__9162_ gnd vdd FILL
XFILL_2__11520_ gnd vdd FILL
XFILL_3_BUFX2_insert284 gnd vdd FILL
XFILL_3_BUFX2_insert295 gnd vdd FILL
XFILL_1__10161_ gnd vdd FILL
X_10017_ _9996_/A _9889_/B gnd _10017_/Y vdd NAND2X1
XSFILL29000x64050 gnd vdd FILL
XFILL_0__10891_ gnd vdd FILL
XFILL_2__8113_ gnd vdd FILL
XFILL_5__11631_ gnd vdd FILL
XFILL_4__10272_ gnd vdd FILL
X_15874_ _10802_/A gnd _15874_/Y vdd INVX1
XFILL_2__9093_ gnd vdd FILL
XFILL_2__11451_ gnd vdd FILL
XFILL_0__12630_ gnd vdd FILL
XFILL_5__9911_ gnd vdd FILL
XFILL_3__13790_ gnd vdd FILL
XFILL_4__9029_ gnd vdd FILL
XFILL_2_BUFX2_insert940 gnd vdd FILL
XFILL_2_BUFX2_insert951 gnd vdd FILL
XFILL_2_BUFX2_insert962 gnd vdd FILL
X_14825_ _7922_/Q gnd _14825_/Y vdd INVX1
XFILL_4__12011_ gnd vdd FILL
XFILL_5__14350_ gnd vdd FILL
XFILL_2__10402_ gnd vdd FILL
XFILL_5__11562_ gnd vdd FILL
XFILL_3__12741_ gnd vdd FILL
XFILL_2__14170_ gnd vdd FILL
XFILL_2_BUFX2_insert973 gnd vdd FILL
XFILL_1__13920_ gnd vdd FILL
XFILL_2__11382_ gnd vdd FILL
XFILL_2_BUFX2_insert984 gnd vdd FILL
XFILL_5__13301_ gnd vdd FILL
XFILL_2_BUFX2_insert995 gnd vdd FILL
XSFILL84280x83050 gnd vdd FILL
XFILL_6__12852_ gnd vdd FILL
XFILL_5__10513_ gnd vdd FILL
XFILL_2__13121_ gnd vdd FILL
X_14756_ _9031_/A gnd _14756_/Y vdd INVX1
XFILL_5__14281_ gnd vdd FILL
X_11968_ _13202_/Q gnd _11970_/A vdd INVX1
XFILL_0__14300_ gnd vdd FILL
XFILL_5__11493_ gnd vdd FILL
XFILL_3__15460_ gnd vdd FILL
XFILL_1__13851_ gnd vdd FILL
XFILL_0__11512_ gnd vdd FILL
XFILL_5__16020_ gnd vdd FILL
XFILL_0__15280_ gnd vdd FILL
XFILL_5__13232_ gnd vdd FILL
XFILL_0__12492_ gnd vdd FILL
XFILL_5__9773_ gnd vdd FILL
X_13707_ _8795_/Q gnd _13708_/A vdd INVX1
XFILL_5__10444_ gnd vdd FILL
X_10919_ _10924_/A _10906_/Y gnd _11874_/B vdd NOR2X1
XFILL_3__14411_ gnd vdd FILL
XFILL_5__6985_ gnd vdd FILL
X_11899_ _12127_/A gnd _11901_/A vdd INVX1
XFILL_3__11623_ gnd vdd FILL
XFILL_4__13962_ gnd vdd FILL
X_14687_ _14687_/A _14687_/B gnd _14687_/Y vdd NOR2X1
XFILL_3__15391_ gnd vdd FILL
XFILL_0__14231_ gnd vdd FILL
XFILL_2__10264_ gnd vdd FILL
XFILL_2__9995_ gnd vdd FILL
XFILL_1__13782_ gnd vdd FILL
XFILL_5__8724_ gnd vdd FILL
XFILL_0__11443_ gnd vdd FILL
XFILL_4__15701_ gnd vdd FILL
X_16426_ _13909_/A _7156_/CLK _9823_/R vdd _16426_/D gnd vdd DFFSR
XFILL_1__10994_ gnd vdd FILL
X_13638_ _9602_/A gnd _13640_/A vdd INVX1
XFILL_5__13163_ gnd vdd FILL
XFILL_2__12003_ gnd vdd FILL
XFILL_4__12913_ gnd vdd FILL
XSFILL38760x58050 gnd vdd FILL
XSFILL93800x45050 gnd vdd FILL
XFILL_1__15521_ gnd vdd FILL
XFILL_3__14342_ gnd vdd FILL
XFILL_5__10375_ gnd vdd FILL
XFILL_3__11554_ gnd vdd FILL
XFILL_1__12733_ gnd vdd FILL
XFILL112280x65050 gnd vdd FILL
XFILL_4__13893_ gnd vdd FILL
XFILL_0__14162_ gnd vdd FILL
XFILL_2__10195_ gnd vdd FILL
XBUFX2_insert950 _13365_/Y gnd _10809_/A vdd BUFX2
XFILL_5__8655_ gnd vdd FILL
XFILL_5__12114_ gnd vdd FILL
XFILL_0__11374_ gnd vdd FILL
XFILL_3__10505_ gnd vdd FILL
XFILL_4__15632_ gnd vdd FILL
XFILL_0__7961_ gnd vdd FILL
X_16357_ _14043_/A gnd _16357_/Y vdd INVX1
XBUFX2_insert961 _13361_/Y gnd _10395_/A vdd BUFX2
XSFILL68520x4050 gnd vdd FILL
XSFILL94440x11050 gnd vdd FILL
XFILL_4__12844_ gnd vdd FILL
XBUFX2_insert972 _16451_/Y gnd _13168_/B vdd BUFX2
X_13569_ _13876_/C gnd _13569_/Y vdd INVX8
XFILL_5__13094_ gnd vdd FILL
XBUFX2_insert983 _13351_/Y gnd _9996_/A vdd BUFX2
XFILL_3__7670_ gnd vdd FILL
XFILL_0__13113_ gnd vdd FILL
XFILL_3__14273_ gnd vdd FILL
XFILL_1__15452_ gnd vdd FILL
XFILL_3__11485_ gnd vdd FILL
XBUFX2_insert994 _12408_/Y gnd _8630_/B vdd BUFX2
XFILL_5__7606_ gnd vdd FILL
XFILL_2__8877_ gnd vdd FILL
XFILL_0__10325_ gnd vdd FILL
XFILL_0__6912_ gnd vdd FILL
X_15308_ _15307_/Y _15308_/B gnd _15309_/C vdd NOR2X1
XFILL_6__10616_ gnd vdd FILL
XFILL_0__14093_ gnd vdd FILL
XFILL_5__8586_ gnd vdd FILL
XFILL_3__16012_ gnd vdd FILL
XFILL_5__12045_ gnd vdd FILL
XFILL_3__13224_ gnd vdd FILL
XFILL_3__10436_ gnd vdd FILL
XFILL_4__15563_ gnd vdd FILL
X_16288_ _8531_/A _15978_/C gnd _16290_/B vdd NAND2X1
XFILL_1__14403_ gnd vdd FILL
XFILL_0__7892_ gnd vdd FILL
XFILL_4__12775_ gnd vdd FILL
XSFILL79240x72050 gnd vdd FILL
XFILL_2__7828_ gnd vdd FILL
XFILL_1__11615_ gnd vdd FILL
XFILL_0__10256_ gnd vdd FILL
XFILL_1__15383_ gnd vdd FILL
XFILL_0__13044_ gnd vdd FILL
XFILL_2__13954_ gnd vdd FILL
XFILL_1__12595_ gnd vdd FILL
XFILL_4__14514_ gnd vdd FILL
X_15239_ _15239_/A _15239_/B _15915_/C _15238_/Y gnd _15239_/Y vdd OAI22X1
XFILL_0__6843_ gnd vdd FILL
XFILL_0__9631_ gnd vdd FILL
XFILL_3__13155_ gnd vdd FILL
X_8170_ _8170_/Q _9328_/CLK _7920_/R vdd _8116_/Y gnd vdd DFFSR
XFILL_4__11726_ gnd vdd FILL
XSFILL28840x5050 gnd vdd FILL
XFILL_3__10367_ gnd vdd FILL
XFILL_1__14334_ gnd vdd FILL
XFILL_3__9340_ gnd vdd FILL
XFILL_4__15494_ gnd vdd FILL
XFILL_2__12905_ gnd vdd FILL
XFILL_2__7759_ gnd vdd FILL
XFILL_1__11546_ gnd vdd FILL
XSFILL18680x25050 gnd vdd FILL
XSFILL114440x81050 gnd vdd FILL
XFILL_2__13885_ gnd vdd FILL
XFILL_0__10187_ gnd vdd FILL
XFILL_3__12106_ gnd vdd FILL
XFILL_5__15804_ gnd vdd FILL
XFILL_5__7468_ gnd vdd FILL
XSFILL74200x19050 gnd vdd FILL
X_7121_ _7064_/A _8273_/B gnd _7122_/C vdd NAND2X1
XFILL_4__14445_ gnd vdd FILL
XFILL_2__15624_ gnd vdd FILL
XFILL_3__13086_ gnd vdd FILL
XFILL_5__13996_ gnd vdd FILL
XFILL_4__11657_ gnd vdd FILL
XFILL_3__9271_ gnd vdd FILL
XSFILL84360x63050 gnd vdd FILL
XFILL_1__14265_ gnd vdd FILL
XFILL_2__12836_ gnd vdd FILL
XFILL_5__9207_ gnd vdd FILL
XFILL_3__10298_ gnd vdd FILL
XFILL_1__11477_ gnd vdd FILL
XFILL_0__14995_ gnd vdd FILL
XFILL_0__8513_ gnd vdd FILL
X_7052_ _7095_/B _7180_/B gnd _7053_/C vdd NAND2X1
XFILL_1__16004_ gnd vdd FILL
XFILL_3__12037_ gnd vdd FILL
XFILL_0__9493_ gnd vdd FILL
XFILL_5__15735_ gnd vdd FILL
XFILL_1__13216_ gnd vdd FILL
XFILL_2__9429_ gnd vdd FILL
XFILL_4__14376_ gnd vdd FILL
XFILL_3__8222_ gnd vdd FILL
XFILL_1__10428_ gnd vdd FILL
XFILL_2__12767_ gnd vdd FILL
XFILL_2__15555_ gnd vdd FILL
XFILL_4__11588_ gnd vdd FILL
XFILL_1__14196_ gnd vdd FILL
XFILL_5__9138_ gnd vdd FILL
XFILL_0__13946_ gnd vdd FILL
XFILL_4__16115_ gnd vdd FILL
XFILL_0__8444_ gnd vdd FILL
XFILL_4__13327_ gnd vdd FILL
XFILL_5__15666_ gnd vdd FILL
XFILL_4__10539_ gnd vdd FILL
XFILL_2__14506_ gnd vdd FILL
XFILL_5__12878_ gnd vdd FILL
XFILL_2__11718_ gnd vdd FILL
XFILL_1__13147_ gnd vdd FILL
XFILL_2__12698_ gnd vdd FILL
XFILL_1__10359_ gnd vdd FILL
XFILL_2__15486_ gnd vdd FILL
XFILL_0__13877_ gnd vdd FILL
XSFILL109800x68050 gnd vdd FILL
XFILL_5__14617_ gnd vdd FILL
XSFILL38840x38050 gnd vdd FILL
XFILL_0__8375_ gnd vdd FILL
XFILL_3__7104_ gnd vdd FILL
XFILL_4__16046_ gnd vdd FILL
XFILL_5__11829_ gnd vdd FILL
XFILL_4__13258_ gnd vdd FILL
XFILL_5__15597_ gnd vdd FILL
XFILL_0__15616_ gnd vdd FILL
XFILL_2__11649_ gnd vdd FILL
XFILL_3__8084_ gnd vdd FILL
XFILL_2__14437_ gnd vdd FILL
XFILL_3__13988_ gnd vdd FILL
XFILL_0__12828_ gnd vdd FILL
XSFILL23640x80050 gnd vdd FILL
XFILL_0__7326_ gnd vdd FILL
XFILL_5__14548_ gnd vdd FILL
XSFILL38440x40050 gnd vdd FILL
XFILL_4__12209_ gnd vdd FILL
XFILL_3__15727_ gnd vdd FILL
XFILL_3__7035_ gnd vdd FILL
X_7954_ _7955_/B _7954_/B gnd _7954_/Y vdd NAND2X1
XFILL_1__12029_ gnd vdd FILL
XFILL_2__14368_ gnd vdd FILL
XFILL_0__15547_ gnd vdd FILL
XFILL_0__12759_ gnd vdd FILL
XSFILL79320x52050 gnd vdd FILL
XFILL_6__15838_ gnd vdd FILL
XSFILL43960x29050 gnd vdd FILL
X_6905_ _6999_/Q gnd _6905_/Y vdd INVX1
XFILL_5__14479_ gnd vdd FILL
XFILL_2__16107_ gnd vdd FILL
X_7885_ _7885_/A gnd _7887_/A vdd INVX1
XFILL_2__13319_ gnd vdd FILL
XFILL_3__15658_ gnd vdd FILL
XSFILL94200x5050 gnd vdd FILL
XFILL_2__14299_ gnd vdd FILL
XFILL_0__15478_ gnd vdd FILL
XFILL_6__8764_ gnd vdd FILL
XFILL_5__16218_ gnd vdd FILL
X_9624_ _9625_/B _9624_/B gnd _9625_/C vdd NAND2X1
X_6836_ gnd gnd MemRead vdd BUFX2
XFILL_3__14609_ gnd vdd FILL
XFILL_0__7188_ gnd vdd FILL
XFILL_2__16038_ gnd vdd FILL
XSFILL114520x61050 gnd vdd FILL
XSFILL8600x15050 gnd vdd FILL
XSFILL44040x38050 gnd vdd FILL
XFILL_3__15589_ gnd vdd FILL
XFILL_0__14429_ gnd vdd FILL
XFILL_6__7715_ gnd vdd FILL
XFILL_3__8986_ gnd vdd FILL
XFILL_5__16149_ gnd vdd FILL
X_9555_ _9555_/A gnd _9555_/Y vdd INVX1
XFILL_5_BUFX2_insert302 gnd vdd FILL
XFILL_3__7937_ gnd vdd FILL
XFILL_1__15719_ gnd vdd FILL
XFILL_5_BUFX2_insert313 gnd vdd FILL
X_8506_ _8504_/Y _8503_/B _8506_/C gnd _8506_/Y vdd OAI21X1
XFILL_5_BUFX2_insert324 gnd vdd FILL
XFILL_1__6952_ gnd vdd FILL
XFILL_1__9740_ gnd vdd FILL
XBUFX2_insert14 _14989_/Y gnd _15569_/C vdd BUFX2
XFILL_5_BUFX2_insert335 gnd vdd FILL
X_9486_ _9566_/Q gnd _9488_/A vdd INVX1
XBUFX2_insert25 _11344_/Y gnd _11802_/A vdd BUFX2
XFILL_5_BUFX2_insert346 gnd vdd FILL
XBUFX2_insert36 _13265_/Y gnd _6948_/A vdd BUFX2
XFILL_3__7868_ gnd vdd FILL
XFILL_5_BUFX2_insert357 gnd vdd FILL
XBUFX2_insert47 _13381_/Y gnd _14441_/B vdd BUFX2
XFILL_5_BUFX2_insert368 gnd vdd FILL
XFILL_5_BUFX2_insert379 gnd vdd FILL
X_8437_ _8437_/Q _9589_/CLK _7285_/R vdd _8437_/D gnd vdd DFFSR
XBUFX2_insert58 _13309_/Y gnd _8107_/B vdd BUFX2
XBUFX2_insert69 _13393_/Y gnd _13803_/A vdd BUFX2
XFILL_1__9671_ gnd vdd FILL
XFILL_3__9607_ gnd vdd FILL
XFILL_1__6883_ gnd vdd FILL
XFILL_4__8400_ gnd vdd FILL
XSFILL38920x18050 gnd vdd FILL
XFILL_4__9380_ gnd vdd FILL
XFILL112440x25050 gnd vdd FILL
XFILL_3__7799_ gnd vdd FILL
XFILL_1__8622_ gnd vdd FILL
X_8368_ _8345_/B _7856_/B gnd _8369_/C vdd NAND2X1
XFILL_4__8331_ gnd vdd FILL
XFILL_3__9538_ gnd vdd FILL
XSFILL24200x67050 gnd vdd FILL
X_7319_ _7319_/A gnd _7319_/Y vdd INVX1
X_8299_ _8299_/Q _7147_/CLK _7133_/R vdd _8299_/D gnd vdd DFFSR
XSFILL8600x6050 gnd vdd FILL
XFILL_4__8262_ gnd vdd FILL
XFILL_3__9469_ gnd vdd FILL
XFILL_1__7504_ gnd vdd FILL
XFILL_1__8484_ gnd vdd FILL
XFILL_4__7213_ gnd vdd FILL
XFILL_4__8193_ gnd vdd FILL
XFILL_1__7435_ gnd vdd FILL
XSFILL94280x46050 gnd vdd FILL
XSFILL84520x23050 gnd vdd FILL
X_12940_ _12886_/A _12669_/CLK _9050_/R vdd _12940_/D gnd vdd DFFSR
XFILL_2_BUFX2_insert225 gnd vdd FILL
XFILL_1__7366_ gnd vdd FILL
XFILL_2_BUFX2_insert236 gnd vdd FILL
XFILL_4__7075_ gnd vdd FILL
XFILL_2_BUFX2_insert247 gnd vdd FILL
XFILL_2_BUFX2_insert258 gnd vdd FILL
XFILL_1__9105_ gnd vdd FILL
X_12871_ _12871_/A gnd _12871_/Y vdd INVX1
XFILL_2_BUFX2_insert269 gnd vdd FILL
XFILL_1__7297_ gnd vdd FILL
XFILL_1_BUFX2_insert903 gnd vdd FILL
X_14610_ _16393_/A gnd _14610_/Y vdd INVX1
XFILL_1__9036_ gnd vdd FILL
XFILL_1_BUFX2_insert914 gnd vdd FILL
X_11822_ _11821_/Y _11809_/C _11802_/A gnd _11822_/Y vdd OAI21X1
X_15590_ _15590_/A gnd _15590_/Y vdd INVX1
XSFILL33560x63050 gnd vdd FILL
XFILL_1_BUFX2_insert925 gnd vdd FILL
XFILL_1_BUFX2_insert936 gnd vdd FILL
XFILL_1_BUFX2_insert947 gnd vdd FILL
X_14541_ _8556_/Q gnd _14541_/Y vdd INVX1
XFILL_1_BUFX2_insert958 gnd vdd FILL
X_11753_ _11753_/A _11753_/B gnd _11754_/A vdd NOR2X1
XFILL_1_BUFX2_insert969 gnd vdd FILL
XSFILL89240x35050 gnd vdd FILL
X_10704_ _14882_/A gnd _10706_/A vdd INVX1
XFILL_4__7977_ gnd vdd FILL
X_14472_ _14472_/A _14472_/B _14467_/Y gnd _14473_/A vdd NAND3X1
X_11684_ _11046_/Y _11684_/B gnd _11684_/Y vdd NOR2X1
XBUFX2_insert235 _12348_/Y gnd _9978_/B vdd BUFX2
XFILL_2__6992_ gnd vdd FILL
XFILL_2__9780_ gnd vdd FILL
XFILL_4__6928_ gnd vdd FILL
X_16211_ _7155_/Q _16293_/A gnd _16219_/A vdd NAND2X1
XBUFX2_insert246 _13460_/Y gnd _13876_/B vdd BUFX2
X_10635_ _10717_/Q gnd _10635_/Y vdd INVX1
XSFILL12840x64050 gnd vdd FILL
X_13423_ _13423_/A _13423_/B _13407_/Y gnd _13423_/Y vdd NAND3X1
XBUFX2_insert257 _12423_/Y gnd _6981_/B vdd BUFX2
XFILL_5__10160_ gnd vdd FILL
XBUFX2_insert268 _15024_/Y gnd _15756_/D vdd BUFX2
XFILL_2__8731_ gnd vdd FILL
XBUFX2_insert279 _13419_/Y gnd _14901_/B vdd BUFX2
XFILL_1__9938_ gnd vdd FILL
XFILL_5_CLKBUF1_insert114 gnd vdd FILL
XFILL_4__10890_ gnd vdd FILL
XFILL_5__8440_ gnd vdd FILL
XFILL_4__9647_ gnd vdd FILL
XSFILL94360x26050 gnd vdd FILL
X_13354_ _13354_/A _13312_/A gnd _13356_/B vdd OR2X2
XFILL_4__6859_ gnd vdd FILL
X_16142_ _7367_/A _15789_/B _15794_/B gnd _16143_/C vdd NAND3X1
XFILL_5_CLKBUF1_insert125 gnd vdd FILL
XFILL_5_CLKBUF1_insert136 gnd vdd FILL
X_10566_ _10566_/A _10500_/B _10566_/C gnd _10566_/Y vdd OAI21X1
XFILL_0__10110_ gnd vdd FILL
XFILL_5_CLKBUF1_insert147 gnd vdd FILL
XFILL_3__11270_ gnd vdd FILL
XFILL_1__9869_ gnd vdd FILL
XFILL_5_CLKBUF1_insert158 gnd vdd FILL
XFILL_5_BUFX2_insert880 gnd vdd FILL
XFILL_5_BUFX2_insert891 gnd vdd FILL
X_12305_ _6892_/A _12301_/B _12301_/C _12313_/D gnd _12306_/C vdd AOI22X1
XFILL_0__11090_ gnd vdd FILL
XFILL_5_CLKBUF1_insert169 gnd vdd FILL
XFILL_5__8371_ gnd vdd FILL
X_13285_ _13291_/A _13285_/B _13284_/Y gnd _13286_/B vdd NAND3X1
X_16073_ _16071_/Y _16151_/B _16247_/C _16072_/Y gnd _16074_/C vdd OAI22X1
X_10497_ _10495_/Y _10511_/A _10497_/C gnd _10585_/D vdd OAI21X1
XFILL_2__7613_ gnd vdd FILL
XFILL_1__11400_ gnd vdd FILL
XFILL_2__10951_ gnd vdd FILL
XFILL_0__10041_ gnd vdd FILL
XFILL_1__12380_ gnd vdd FILL
XFILL_5__7322_ gnd vdd FILL
XFILL_6__13120_ gnd vdd FILL
XFILL_2__8593_ gnd vdd FILL
XFILL_4__8529_ gnd vdd FILL
X_15024_ _14983_/A _14982_/Y _15024_/C gnd _15024_/Y vdd NAND3X1
X_12236_ _12248_/A _12710_/A _12248_/C gnd _12238_/B vdd NAND3X1
XFILL_5__13850_ gnd vdd FILL
XFILL_4__11511_ gnd vdd FILL
XFILL_3__10152_ gnd vdd FILL
XSFILL104360x11050 gnd vdd FILL
XFILL_2__13670_ gnd vdd FILL
XFILL_2__7544_ gnd vdd FILL
XFILL_4__12491_ gnd vdd FILL
XFILL_1__11331_ gnd vdd FILL
XFILL_2__10882_ gnd vdd FILL
XFILL_5__7253_ gnd vdd FILL
XSFILL84280x78050 gnd vdd FILL
XFILL_4__14230_ gnd vdd FILL
X_12167_ _12117_/B _12936_/Q gnd _12168_/C vdd NAND2X1
XFILL_2__12621_ gnd vdd FILL
XFILL_5__13781_ gnd vdd FILL
XFILL_4__11442_ gnd vdd FILL
XFILL_0__13800_ gnd vdd FILL
XFILL_1__14050_ gnd vdd FILL
XFILL_3__14960_ gnd vdd FILL
XFILL_5__10993_ gnd vdd FILL
XFILL_2__7475_ gnd vdd FILL
XFILL_1__11262_ gnd vdd FILL
XFILL_5__7184_ gnd vdd FILL
XFILL_5__15520_ gnd vdd FILL
X_11118_ _11553_/B _11117_/Y gnd _11118_/Y vdd NOR2X1
XFILL_0__14780_ gnd vdd FILL
XFILL_5__12732_ gnd vdd FILL
XFILL_0__11992_ gnd vdd FILL
XFILL_4__14161_ gnd vdd FILL
X_12098_ _12098_/A _12098_/B _12097_/Y gnd _13161_/B vdd NAND3X1
XFILL_1__13001_ gnd vdd FILL
XFILL_3__13911_ gnd vdd FILL
XSFILL89320x15050 gnd vdd FILL
XFILL_2__9214_ gnd vdd FILL
XFILL_2__15340_ gnd vdd FILL
XFILL_4__11373_ gnd vdd FILL
XFILL_0__13731_ gnd vdd FILL
XFILL_3__14891_ gnd vdd FILL
XFILL_0__10943_ gnd vdd FILL
XFILL_1__11193_ gnd vdd FILL
XSFILL19080x70050 gnd vdd FILL
X_15926_ _15926_/A _15926_/B gnd _15927_/B vdd NOR2X1
XFILL_4__13112_ gnd vdd FILL
X_11049_ _12254_/Y _12144_/Y gnd _11731_/B vdd XOR2X1
XFILL_5__15451_ gnd vdd FILL
XFILL_2__11503_ gnd vdd FILL
XFILL_4__10324_ gnd vdd FILL
XFILL_3__13842_ gnd vdd FILL
XFILL_2__9145_ gnd vdd FILL
XFILL_4__14092_ gnd vdd FILL
XFILL_2__15271_ gnd vdd FILL
XFILL_0__16450_ gnd vdd FILL
XFILL_1__10144_ gnd vdd FILL
XFILL_2__12483_ gnd vdd FILL
XFILL_0__13662_ gnd vdd FILL
XFILL_5__14402_ gnd vdd FILL
XFILL_0__10874_ gnd vdd FILL
XFILL_5__11614_ gnd vdd FILL
XFILL_2__14222_ gnd vdd FILL
XFILL_4__10255_ gnd vdd FILL
XFILL_5__15382_ gnd vdd FILL
X_15857_ _15978_/C _8498_/A _8242_/A _16014_/C gnd _15860_/C vdd AOI22X1
XFILL_4__13043_ gnd vdd FILL
XFILL_0__15401_ gnd vdd FILL
XFILL_5__12594_ gnd vdd FILL
XFILL_2__11434_ gnd vdd FILL
XFILL_3__13773_ gnd vdd FILL
XFILL_0__12613_ gnd vdd FILL
XFILL_2_BUFX2_insert770 gnd vdd FILL
XFILL_1__14952_ gnd vdd FILL
XFILL_0__7111_ gnd vdd FILL
XFILL_0__16381_ gnd vdd FILL
XFILL_2_BUFX2_insert781 gnd vdd FILL
X_14808_ _7538_/Q gnd _14808_/Y vdd INVX1
XFILL_0__13593_ gnd vdd FILL
XFILL_2_BUFX2_insert792 gnd vdd FILL
XFILL_5__14333_ gnd vdd FILL
XSFILL13800x72050 gnd vdd FILL
XFILL_3__15512_ gnd vdd FILL
XFILL_0__8091_ gnd vdd FILL
XFILL_5__11545_ gnd vdd FILL
XFILL_6__13884_ gnd vdd FILL
XFILL_3__12724_ gnd vdd FILL
XFILL_4__10186_ gnd vdd FILL
XFILL_2__14153_ gnd vdd FILL
X_15788_ _15550_/A _15787_/Y _15550_/C gnd _15788_/Y vdd NOR3X1
XSFILL79240x67050 gnd vdd FILL
XFILL_0__15332_ gnd vdd FILL
XFILL_1__13903_ gnd vdd FILL
XFILL_2__11365_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1076 gnd vdd FILL
XFILL_1__14883_ gnd vdd FILL
XFILL_6__15623_ gnd vdd FILL
XFILL_0__7042_ gnd vdd FILL
XFILL_5__14264_ gnd vdd FILL
XFILL_2__13104_ gnd vdd FILL
X_14739_ _9200_/Q _14868_/D _14739_/C _10608_/Q gnd _14740_/B vdd AOI22X1
XFILL_2__10316_ gnd vdd FILL
X_7670_ _7766_/Q gnd _7670_/Y vdd INVX1
XFILL_5__11476_ gnd vdd FILL
XFILL_3__15443_ gnd vdd FILL
XFILL_3__12655_ gnd vdd FILL
XFILL_3__8840_ gnd vdd FILL
XFILL_1__13834_ gnd vdd FILL
XFILL_4__14994_ gnd vdd FILL
XFILL_2__14084_ gnd vdd FILL
XFILL_5__16003_ gnd vdd FILL
XFILL_2__11296_ gnd vdd FILL
XFILL_0__15263_ gnd vdd FILL
XFILL_5__13215_ gnd vdd FILL
XFILL_5__9756_ gnd vdd FILL
XFILL_0__12475_ gnd vdd FILL
XFILL_5__10427_ gnd vdd FILL
XFILL_5__6968_ gnd vdd FILL
XFILL_5__14195_ gnd vdd FILL
XFILL_2__13035_ gnd vdd FILL
XFILL_3__11606_ gnd vdd FILL
XFILL_4__13945_ gnd vdd FILL
XFILL_3__15374_ gnd vdd FILL
XFILL_0__14214_ gnd vdd FILL
XFILL_2__10247_ gnd vdd FILL
XFILL_3__12586_ gnd vdd FILL
XFILL_5__8707_ gnd vdd FILL
XSFILL84360x58050 gnd vdd FILL
XFILL_1__13765_ gnd vdd FILL
XFILL_3__8771_ gnd vdd FILL
XFILL_2__9978_ gnd vdd FILL
XFILL_0__11426_ gnd vdd FILL
XFILL_1__10977_ gnd vdd FILL
XFILL_0__15194_ gnd vdd FILL
X_16409_ gnd gnd gnd _16410_/C vdd NAND2X1
XFILL_5__13146_ gnd vdd FILL
XFILL_6__8480_ gnd vdd FILL
X_9340_ _9340_/A gnd _9342_/A vdd INVX1
XFILL_6__11717_ gnd vdd FILL
XFILL_6__12697_ gnd vdd FILL
XFILL_5__10358_ gnd vdd FILL
XFILL_5__6899_ gnd vdd FILL
XFILL_3__14325_ gnd vdd FILL
XFILL_6__15485_ gnd vdd FILL
XFILL_1__12716_ gnd vdd FILL
XFILL_4__13876_ gnd vdd FILL
XFILL_0__8993_ gnd vdd FILL
XFILL_1__15504_ gnd vdd FILL
XFILL_3__11537_ gnd vdd FILL
XFILL_3__7722_ gnd vdd FILL
XFILL_0__14145_ gnd vdd FILL
XFILL_2__10178_ gnd vdd FILL
XFILL_5__8638_ gnd vdd FILL
XBUFX2_insert780 _10911_/Y gnd _12134_/A vdd BUFX2
XFILL_6__7431_ gnd vdd FILL
XFILL_1__13696_ gnd vdd FILL
XFILL_0__11357_ gnd vdd FILL
XFILL_4__15615_ gnd vdd FILL
XBUFX2_insert791 _15052_/Y gnd _15801_/C vdd BUFX2
XFILL_6__14436_ gnd vdd FILL
XFILL_0__7944_ gnd vdd FILL
X_9271_ _9271_/A _9228_/A _9270_/Y gnd _9323_/D vdd OAI21X1
XSFILL34600x51050 gnd vdd FILL
XFILL_4__12827_ gnd vdd FILL
XFILL_3__14256_ gnd vdd FILL
XFILL_5__10289_ gnd vdd FILL
XFILL_1__15435_ gnd vdd FILL
XFILL_1__12647_ gnd vdd FILL
XFILL_0__10308_ gnd vdd FILL
XFILL_3__11468_ gnd vdd FILL
XFILL_2__14986_ gnd vdd FILL
XFILL_0__14076_ gnd vdd FILL
XFILL_4_BUFX2_insert309 gnd vdd FILL
XFILL_5__12028_ gnd vdd FILL
XFILL_0__11288_ gnd vdd FILL
X_8222_ _8244_/B _9246_/B gnd _8222_/Y vdd NAND2X1
XFILL_5__8569_ gnd vdd FILL
XFILL_3__13207_ gnd vdd FILL
XFILL_4__15546_ gnd vdd FILL
XFILL_6__11579_ gnd vdd FILL
XFILL_4__12758_ gnd vdd FILL
XFILL_3__10419_ gnd vdd FILL
XFILL_0__7875_ gnd vdd FILL
XFILL_3__14187_ gnd vdd FILL
XFILL_1__15366_ gnd vdd FILL
XFILL_0__13027_ gnd vdd FILL
XFILL_3__11399_ gnd vdd FILL
XFILL_2__13937_ gnd vdd FILL
XFILL_1__12578_ gnd vdd FILL
XFILL_0__10239_ gnd vdd FILL
XFILL_3__7584_ gnd vdd FILL
XSFILL23640x75050 gnd vdd FILL
XFILL_0__9614_ gnd vdd FILL
X_8153_ _8153_/Q _9817_/CLK _8542_/R vdd _8065_/Y gnd vdd DFFSR
XFILL_6__14298_ gnd vdd FILL
XFILL_4__11709_ gnd vdd FILL
XFILL_3__13138_ gnd vdd FILL
XFILL_1__14317_ gnd vdd FILL
XFILL_4__15477_ gnd vdd FILL
XFILL_1__11529_ gnd vdd FILL
XFILL_2__13868_ gnd vdd FILL
XFILL_1__15297_ gnd vdd FILL
XFILL_6__9032_ gnd vdd FILL
XFILL_6__13249_ gnd vdd FILL
X_7104_ _7102_/Y _7055_/A _7104_/C gnd _7104_/Y vdd OAI21X1
XSFILL79320x47050 gnd vdd FILL
XFILL_0__9545_ gnd vdd FILL
XFILL_4__14428_ gnd vdd FILL
X_8084_ _8160_/Q gnd _8084_/Y vdd INVX1
XFILL_2__15607_ gnd vdd FILL
XFILL_1__14248_ gnd vdd FILL
XFILL_3__9254_ gnd vdd FILL
XFILL_5__13979_ gnd vdd FILL
XFILL_2__13799_ gnd vdd FILL
XFILL_0__14978_ gnd vdd FILL
XFILL_5__15718_ gnd vdd FILL
X_7035_ _7035_/A _7061_/A _7034_/Y gnd _7127_/D vdd OAI21X1
XFILL_0__9476_ gnd vdd FILL
XFILL_3__8205_ gnd vdd FILL
XFILL_4__14359_ gnd vdd FILL
XFILL_2__15538_ gnd vdd FILL
XFILL_1__14179_ gnd vdd FILL
XFILL_0__13929_ gnd vdd FILL
XFILL_1__7220_ gnd vdd FILL
XFILL_5__15649_ gnd vdd FILL
XSFILL84440x38050 gnd vdd FILL
XFILL_3__8136_ gnd vdd FILL
XFILL_2__15469_ gnd vdd FILL
XFILL_0__8358_ gnd vdd FILL
XFILL_4__16029_ gnd vdd FILL
XFILL_3__8067_ gnd vdd FILL
X_8986_ _8986_/A gnd _8988_/A vdd INVX1
XFILL_0__7309_ gnd vdd FILL
XFILL_6__9865_ gnd vdd FILL
X_7937_ _7935_/Y _7937_/B _7936_/Y gnd _8025_/D vdd OAI21X1
XFILL_1__7082_ gnd vdd FILL
XFILL111960x13050 gnd vdd FILL
XFILL_4__8880_ gnd vdd FILL
X_7868_ _7887_/B _7868_/B gnd _7868_/Y vdd NAND2X1
XSFILL23720x55050 gnd vdd FILL
XFILL_4__7831_ gnd vdd FILL
X_9607_ _9605_/Y _9597_/A _9607_/C gnd _9691_/D vdd OAI21X1
XFILL112040x22050 gnd vdd FILL
X_7799_ _8823_/A _7824_/B gnd _7800_/C vdd NAND2X1
XFILL_3__8969_ gnd vdd FILL
XSFILL79400x27050 gnd vdd FILL
XFILL_4__7762_ gnd vdd FILL
XFILL_5_BUFX2_insert110 gnd vdd FILL
X_9538_ _9554_/B _8642_/B gnd _9539_/C vdd NAND2X1
XFILL_4__9501_ gnd vdd FILL
XSFILL39400x43050 gnd vdd FILL
XFILL_1__7984_ gnd vdd FILL
X_10420_ _10420_/A _10426_/B _10419_/Y gnd _10474_/D vdd OAI21X1
XFILL_4__7693_ gnd vdd FILL
XSFILL114600x36050 gnd vdd FILL
XFILL_1__9723_ gnd vdd FILL
XFILL_1__6935_ gnd vdd FILL
X_9469_ _9514_/A _9597_/B gnd _9469_/Y vdd NAND2X1
X_10351_ _10305_/A _9716_/CLK _8431_/R vdd _10307_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert810 gnd vdd FILL
XFILL_1__9654_ gnd vdd FILL
XFILL_4_BUFX2_insert821 gnd vdd FILL
XSFILL69080x17050 gnd vdd FILL
XFILL_1__6866_ gnd vdd FILL
XFILL_4_BUFX2_insert832 gnd vdd FILL
XFILL_4_BUFX2_insert843 gnd vdd FILL
XFILL_4__9363_ gnd vdd FILL
X_13070_ _6893_/A _7005_/CLK _7133_/R vdd _13070_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert854 gnd vdd FILL
X_10282_ _10285_/A _8874_/B gnd _10282_/Y vdd NAND2X1
XSFILL109480x1050 gnd vdd FILL
XFILL_1__8605_ gnd vdd FILL
XFILL_4_BUFX2_insert865 gnd vdd FILL
XFILL_4_BUFX2_insert876 gnd vdd FILL
XFILL_4__8314_ gnd vdd FILL
XFILL_4_BUFX2_insert887 gnd vdd FILL
X_12021_ _12021_/A _12105_/B _12001_/C gnd gnd _12022_/C vdd AOI22X1
XFILL_4__9294_ gnd vdd FILL
XFILL_4_BUFX2_insert898 gnd vdd FILL
XFILL_4__8245_ gnd vdd FILL
XSFILL23800x35050 gnd vdd FILL
XFILL_1__8467_ gnd vdd FILL
X_13972_ _13972_/A _14389_/B _14358_/B _10848_/Q gnd _13973_/B vdd AOI22X1
XFILL_1__7418_ gnd vdd FILL
XFILL_1__8398_ gnd vdd FILL
XFILL_2__7191_ gnd vdd FILL
X_15711_ _15711_/A _15683_/B _15683_/C _15711_/D gnd _15714_/A vdd OAI22X1
X_12923_ _12923_/Q _9060_/CLK _7140_/R vdd _12837_/Y gnd vdd DFFSR
XFILL_1__7349_ gnd vdd FILL
XFILL_5__7940_ gnd vdd FILL
XFILL_4__7058_ gnd vdd FILL
X_15642_ _14138_/A _15981_/B _15351_/A _15642_/D gnd _15642_/Y vdd OAI22X1
XFILL_4__10040_ gnd vdd FILL
XFILL_1_BUFX2_insert700 gnd vdd FILL
X_12854_ vdd _12854_/B gnd _12855_/C vdd NAND2X1
XFILL_1_BUFX2_insert711 gnd vdd FILL
XFILL_3__10770_ gnd vdd FILL
XFILL_1_BUFX2_insert722 gnd vdd FILL
XFILL_1_BUFX2_insert733 gnd vdd FILL
XFILL_5__7871_ gnd vdd FILL
XFILL_5__11330_ gnd vdd FILL
X_11805_ _11794_/Y _11846_/C _11805_/C gnd _11808_/A vdd AOI21X1
XFILL_1__9019_ gnd vdd FILL
XFILL_1_BUFX2_insert744 gnd vdd FILL
X_15573_ _15573_/A _15572_/Y _15338_/C gnd _12860_/B vdd AOI21X1
XFILL_2__9901_ gnd vdd FILL
X_12785_ _12785_/A gnd _12785_/Y vdd INVX1
XFILL_1__10900_ gnd vdd FILL
XFILL_1_BUFX2_insert755 gnd vdd FILL
XFILL_2__11150_ gnd vdd FILL
XFILL_5__9610_ gnd vdd FILL
XFILL_1_BUFX2_insert766 gnd vdd FILL
XFILL_1__11880_ gnd vdd FILL
XSFILL69400x59050 gnd vdd FILL
XFILL_1_BUFX2_insert777 gnd vdd FILL
XFILL_1_BUFX2_insert788 gnd vdd FILL
X_14524_ _14524_/A _14815_/C gnd _14525_/C vdd NOR2X1
XSFILL109400x9050 gnd vdd FILL
XFILL_5__11261_ gnd vdd FILL
X_11736_ _11028_/Y _11041_/Y _11386_/Y gnd _11737_/C vdd OAI21X1
XFILL_1_BUFX2_insert799 gnd vdd FILL
XFILL_3__12440_ gnd vdd FILL
XFILL_1__10831_ gnd vdd FILL
XFILL_4__11991_ gnd vdd FILL
XFILL_2__11081_ gnd vdd FILL
XFILL_5__13000_ gnd vdd FILL
XFILL_5__9541_ gnd vdd FILL
XFILL_0__12260_ gnd vdd FILL
XFILL_4_BUFX2_insert15 gnd vdd FILL
X_14455_ _7605_/A gnd _14456_/A vdd INVX1
XFILL_4__13730_ gnd vdd FILL
XFILL_4__10942_ gnd vdd FILL
XFILL_4_BUFX2_insert26 gnd vdd FILL
XFILL_3__12371_ gnd vdd FILL
XFILL_2__10032_ gnd vdd FILL
X_11667_ _11649_/Y _11748_/A _11666_/Y gnd _11670_/B vdd OAI21X1
XFILL_5__11192_ gnd vdd FILL
XFILL_2__9763_ gnd vdd FILL
XFILL_4_BUFX2_insert37 gnd vdd FILL
XFILL_1__13550_ gnd vdd FILL
XFILL_0__11211_ gnd vdd FILL
XFILL_2__6975_ gnd vdd FILL
XFILL_1__10762_ gnd vdd FILL
XFILL_4_BUFX2_insert48 gnd vdd FILL
XFILL_6__11502_ gnd vdd FILL
XFILL_5__9472_ gnd vdd FILL
X_13406_ _11881_/A gnd _13406_/Y vdd INVX1
XFILL_4_BUFX2_insert59 gnd vdd FILL
XFILL_6__15270_ gnd vdd FILL
XFILL_0__12191_ gnd vdd FILL
X_10618_ _10619_/B _6906_/B gnd _10618_/Y vdd NAND2X1
XFILL_3__14110_ gnd vdd FILL
XFILL_5__10143_ gnd vdd FILL
XFILL_4__13661_ gnd vdd FILL
XFILL_2__8714_ gnd vdd FILL
XFILL_1__12501_ gnd vdd FILL
X_14386_ _15820_/A _14697_/B _14725_/A _14386_/D gnd _14387_/A vdd OAI22X1
X_11598_ _11597_/Y _11130_/B _11146_/B gnd _11598_/Y vdd OAI21X1
XFILL_3__11322_ gnd vdd FILL
XFILL_2__14840_ gnd vdd FILL
XFILL_3__15090_ gnd vdd FILL
XFILL_4__10873_ gnd vdd FILL
XFILL_0__11142_ gnd vdd FILL
XFILL_1__13481_ gnd vdd FILL
XFILL_4__15400_ gnd vdd FILL
XSFILL99480x54050 gnd vdd FILL
XFILL_6__14221_ gnd vdd FILL
XFILL_1__10693_ gnd vdd FILL
X_16125_ _8519_/A gnd _16126_/D vdd INVX1
X_13337_ _13337_/A _13337_/B _13337_/C gnd _13337_/Y vdd NAND3X1
X_10549_ _14454_/A gnd _10551_/A vdd INVX1
XFILL_4__12612_ gnd vdd FILL
XFILL_1__15220_ gnd vdd FILL
XFILL_3__14041_ gnd vdd FILL
XFILL_5__14951_ gnd vdd FILL
XFILL_4__16380_ gnd vdd FILL
XFILL_3__11253_ gnd vdd FILL
XFILL_1__12432_ gnd vdd FILL
XFILL_4__13592_ gnd vdd FILL
XFILL_2__8645_ gnd vdd FILL
XFILL_2__11983_ gnd vdd FILL
XFILL_0__15950_ gnd vdd FILL
XFILL_0__11073_ gnd vdd FILL
XFILL_2__14771_ gnd vdd FILL
XFILL_5__8354_ gnd vdd FILL
XFILL_4__15331_ gnd vdd FILL
XFILL_5__13902_ gnd vdd FILL
X_16056_ _15172_/A _16055_/Y _16155_/D _16056_/D gnd _16056_/Y vdd OAI22X1
XFILL_6__11364_ gnd vdd FILL
X_13268_ _13297_/A _13268_/B gnd _13269_/B vdd OR2X2
XFILL_5__14882_ gnd vdd FILL
XFILL_3__11184_ gnd vdd FILL
XFILL_1__15151_ gnd vdd FILL
XFILL_2__13722_ gnd vdd FILL
XFILL_0__14901_ gnd vdd FILL
XFILL_2__10934_ gnd vdd FILL
XFILL_2__8576_ gnd vdd FILL
XFILL_1__12363_ gnd vdd FILL
XFILL_5__7305_ gnd vdd FILL
XFILL_0__10024_ gnd vdd FILL
XFILL_6__10315_ gnd vdd FILL
X_15007_ _15356_/C _10486_/A _10198_/Q _15695_/D gnd _15008_/B vdd AOI22X1
XFILL_2_BUFX2_insert1009 gnd vdd FILL
XFILL_0__15881_ gnd vdd FILL
XSFILL53960x10050 gnd vdd FILL
XFILL_6__14083_ gnd vdd FILL
X_12219_ _12227_/A gnd _12307_/C gnd _12219_/Y vdd NAND3X1
XFILL_0__7591_ gnd vdd FILL
XSFILL13800x67050 gnd vdd FILL
XFILL_5__13833_ gnd vdd FILL
X_13199_ _11959_/A _12538_/CLK _13199_/R vdd _13199_/D gnd vdd DFFSR
XFILL_3__10135_ gnd vdd FILL
XFILL_1__14102_ gnd vdd FILL
XFILL_4__15262_ gnd vdd FILL
XFILL_4__12474_ gnd vdd FILL
XFILL_1__11314_ gnd vdd FILL
XFILL_2__13653_ gnd vdd FILL
XFILL_3__15992_ gnd vdd FILL
XFILL_0__14832_ gnd vdd FILL
XFILL_1__15082_ gnd vdd FILL
XFILL_5__7236_ gnd vdd FILL
XFILL_1__12294_ gnd vdd FILL
XFILL_4__14213_ gnd vdd FILL
XFILL_5__13764_ gnd vdd FILL
XFILL_4__11425_ gnd vdd FILL
XSFILL39240x78050 gnd vdd FILL
XFILL_5__10976_ gnd vdd FILL
XFILL_2__12604_ gnd vdd FILL
XFILL_4__15193_ gnd vdd FILL
XFILL_1__14033_ gnd vdd FILL
XFILL_3__14943_ gnd vdd FILL
XFILL_3__10066_ gnd vdd FILL
XFILL_2__7458_ gnd vdd FILL
XFILL_2__16372_ gnd vdd FILL
XFILL_2__13584_ gnd vdd FILL
XFILL_1__11245_ gnd vdd FILL
XFILL_2__10796_ gnd vdd FILL
XFILL_0__14763_ gnd vdd FILL
XFILL_5__7167_ gnd vdd FILL
XFILL_5__12715_ gnd vdd FILL
XFILL_0__11975_ gnd vdd FILL
XFILL_5__15503_ gnd vdd FILL
XFILL_0__9261_ gnd vdd FILL
XFILL_4__14144_ gnd vdd FILL
XFILL_2__15323_ gnd vdd FILL
XFILL_4__11356_ gnd vdd FILL
XFILL_5__13695_ gnd vdd FILL
XFILL_3__14874_ gnd vdd FILL
XSFILL83880x46050 gnd vdd FILL
XFILL_0__13714_ gnd vdd FILL
XFILL_0__10926_ gnd vdd FILL
XFILL_0__8212_ gnd vdd FILL
XFILL_1__11176_ gnd vdd FILL
X_15909_ _15903_/Y _15909_/B _15908_/Y gnd _15910_/A vdd NAND3X1
XFILL_0__14694_ gnd vdd FILL
X_8840_ _8924_/Q gnd _8840_/Y vdd INVX1
XFILL_5__12646_ gnd vdd FILL
XFILL_5__7098_ gnd vdd FILL
XFILL_0_BUFX2_insert1002 gnd vdd FILL
XFILL_4__10307_ gnd vdd FILL
XFILL_5__15434_ gnd vdd FILL
XFILL_3__13825_ gnd vdd FILL
XSFILL43880x62050 gnd vdd FILL
XFILL_2__9128_ gnd vdd FILL
XFILL_4__14075_ gnd vdd FILL
XFILL_1__10127_ gnd vdd FILL
XFILL_2__15254_ gnd vdd FILL
XFILL_2__12466_ gnd vdd FILL
XFILL_0_BUFX2_insert1013 gnd vdd FILL
XFILL_4__11287_ gnd vdd FILL
XFILL_0__13645_ gnd vdd FILL
XFILL_0_BUFX2_insert1024 gnd vdd FILL
XFILL_0_BUFX2_insert1035 gnd vdd FILL
XFILL_0__8143_ gnd vdd FILL
XFILL_1__15984_ gnd vdd FILL
XSFILL59160x29050 gnd vdd FILL
XFILL_5__15365_ gnd vdd FILL
XFILL_4__13026_ gnd vdd FILL
XFILL_0_BUFX2_insert1046 gnd vdd FILL
XFILL_5__12577_ gnd vdd FILL
XFILL_2__14205_ gnd vdd FILL
XFILL_0_BUFX2_insert1057 gnd vdd FILL
X_8771_ _8771_/A _8753_/B _8771_/C gnd _8815_/D vdd OAI21X1
XFILL_4__10238_ gnd vdd FILL
XFILL_2__11417_ gnd vdd FILL
XFILL_3__13756_ gnd vdd FILL
XFILL_3__9941_ gnd vdd FILL
XFILL_3__10968_ gnd vdd FILL
XFILL_2__15185_ gnd vdd FILL
XFILL_1__10058_ gnd vdd FILL
XFILL_0__16364_ gnd vdd FILL
XFILL_0_BUFX2_insert1068 gnd vdd FILL
XFILL_2__12397_ gnd vdd FILL
XFILL_1__14935_ gnd vdd FILL
XFILL_5__14316_ gnd vdd FILL
XSFILL74200x32050 gnd vdd FILL
XFILL_0__13576_ gnd vdd FILL
XFILL_0__10788_ gnd vdd FILL
XFILL_0__8074_ gnd vdd FILL
XFILL_5__11528_ gnd vdd FILL
X_7722_ _7723_/B _9898_/B gnd _7722_/Y vdd NAND2X1
XSFILL99000x77050 gnd vdd FILL
XFILL_3__12707_ gnd vdd FILL
XFILL_5__15296_ gnd vdd FILL
XFILL_0__15315_ gnd vdd FILL
XFILL_2__14136_ gnd vdd FILL
XFILL_4__10169_ gnd vdd FILL
XFILL_2__11348_ gnd vdd FILL
XFILL_3__9872_ gnd vdd FILL
XFILL_0__12527_ gnd vdd FILL
XFILL_3__13687_ gnd vdd FILL
XFILL_5__9808_ gnd vdd FILL
XFILL_1__14866_ gnd vdd FILL
XFILL_3__10899_ gnd vdd FILL
XFILL_0__16295_ gnd vdd FILL
XFILL_5__14247_ gnd vdd FILL
X_7653_ _7653_/Q _7406_/CLK _8430_/R vdd _7589_/Y gnd vdd DFFSR
XFILL_5__11459_ gnd vdd FILL
XFILL_3__15426_ gnd vdd FILL
XSFILL37960x23050 gnd vdd FILL
XFILL_3__12638_ gnd vdd FILL
XFILL_3__8823_ gnd vdd FILL
XFILL_2__14067_ gnd vdd FILL
XFILL_4__14977_ gnd vdd FILL
XFILL_1__13817_ gnd vdd FILL
XFILL_0__15246_ gnd vdd FILL
XFILL112440x2050 gnd vdd FILL
XFILL_2__11279_ gnd vdd FILL
XFILL_5__9739_ gnd vdd FILL
XFILL_0__12458_ gnd vdd FILL
XFILL_1__14797_ gnd vdd FILL
XSFILL78840x35050 gnd vdd FILL
XFILL_5__14178_ gnd vdd FILL
XFILL_2__13018_ gnd vdd FILL
XFILL_4__13928_ gnd vdd FILL
XSFILL23240x72050 gnd vdd FILL
XFILL_3__15357_ gnd vdd FILL
X_7584_ _7584_/A gnd _7584_/Y vdd INVX1
XFILL_3__12569_ gnd vdd FILL
XFILL_3__8754_ gnd vdd FILL
XFILL_0__11409_ gnd vdd FILL
XSFILL109800x81050 gnd vdd FILL
XFILL_0__15177_ gnd vdd FILL
XSFILL109000x62050 gnd vdd FILL
XFILL_1__13748_ gnd vdd FILL
X_9323_ _9269_/A _7389_/CLK _7531_/R vdd _9323_/D gnd vdd DFFSR
XFILL_0__12389_ gnd vdd FILL
XFILL_5__13129_ gnd vdd FILL
XFILL_3__14308_ gnd vdd FILL
XFILL_4__13859_ gnd vdd FILL
XFILL_0__8976_ gnd vdd FILL
XFILL_3__7705_ gnd vdd FILL
XFILL_0__14128_ gnd vdd FILL
XFILL_3__15288_ gnd vdd FILL
XFILL_1__13679_ gnd vdd FILL
XSFILL74120x4050 gnd vdd FILL
XFILL_4_BUFX2_insert106 gnd vdd FILL
XSFILL113720x4050 gnd vdd FILL
X_9254_ _9318_/Q gnd _9254_/Y vdd INVX1
XFILL_0__7927_ gnd vdd FILL
XFILL_3__14239_ gnd vdd FILL
XFILL_3__7636_ gnd vdd FILL
XFILL_1__15418_ gnd vdd FILL
XFILL_0__14059_ gnd vdd FILL
XFILL_2__14969_ gnd vdd FILL
X_8205_ _8205_/A _8246_/A _8204_/Y gnd _8205_/Y vdd OAI21X1
XSFILL43960x42050 gnd vdd FILL
XFILL_1__16398_ gnd vdd FILL
XFILL_4__15529_ gnd vdd FILL
X_9185_ _9185_/Q _7916_/CLK _7276_/R vdd _9185_/D gnd vdd DFFSR
XFILL_0__7858_ gnd vdd FILL
XFILL_3__7567_ gnd vdd FILL
XFILL_1__15349_ gnd vdd FILL
XFILL_3_BUFX2_insert806 gnd vdd FILL
X_8136_ _8098_/B _8136_/B gnd _8136_/Y vdd NAND2X1
XFILL_1__9370_ gnd vdd FILL
XFILL_3_BUFX2_insert817 gnd vdd FILL
XFILL_3_BUFX2_insert828 gnd vdd FILL
XSFILL44040x51050 gnd vdd FILL
XFILL_3_BUFX2_insert839 gnd vdd FILL
XFILL_3__7498_ gnd vdd FILL
XFILL_1__8321_ gnd vdd FILL
XFILL_0__9528_ gnd vdd FILL
X_8067_ _8118_/A _8195_/B gnd _8068_/C vdd NAND2X1
XFILL_3__9237_ gnd vdd FILL
XFILL_1__8252_ gnd vdd FILL
X_7018_ _6962_/A _7530_/CLK _7523_/R vdd _6964_/Y gnd vdd DFFSR
XSFILL78920x15050 gnd vdd FILL
XFILL_3__9168_ gnd vdd FILL
XFILL_1__7203_ gnd vdd FILL
XFILL_1__8183_ gnd vdd FILL
XFILL_3__8119_ gnd vdd FILL
XFILL_3__9099_ gnd vdd FILL
XSFILL64200x64050 gnd vdd FILL
XFILL_4__9981_ gnd vdd FILL
X_8969_ _8969_/A _9353_/B gnd _8969_/Y vdd NAND2X1
XFILL_1__7065_ gnd vdd FILL
XSFILL3640x71050 gnd vdd FILL
XFILL_4__8863_ gnd vdd FILL
X_12570_ _12570_/A gnd _12570_/Y vdd INVX1
XFILL_0_CLKBUF1_insert111 gnd vdd FILL
XFILL_0_CLKBUF1_insert122 gnd vdd FILL
XFILL_0_CLKBUF1_insert133 gnd vdd FILL
XFILL_0_BUFX2_insert707 gnd vdd FILL
XFILL_0_CLKBUF1_insert144 gnd vdd FILL
XFILL_0_BUFX2_insert718 gnd vdd FILL
XFILL_4__7814_ gnd vdd FILL
XSFILL28840x83050 gnd vdd FILL
XFILL_0_BUFX2_insert729 gnd vdd FILL
XFILL_0_CLKBUF1_insert155 gnd vdd FILL
X_11521_ _11521_/A _11159_/Y _11521_/C gnd _11543_/C vdd OAI21X1
XFILL_0_CLKBUF1_insert166 gnd vdd FILL
XFILL_0_CLKBUF1_insert177 gnd vdd FILL
XFILL_0_CLKBUF1_insert188 gnd vdd FILL
XFILL_0_CLKBUF1_insert199 gnd vdd FILL
XFILL_4__7745_ gnd vdd FILL
X_14240_ _14238_/Y _14203_/B _14489_/C _14240_/D gnd _14241_/B vdd OAI22X1
X_11452_ _11435_/Y _11550_/A gnd _11452_/Y vdd NAND2X1
XFILL_1__7967_ gnd vdd FILL
X_10403_ _10469_/Q gnd _10405_/A vdd INVX1
XSFILL33960x74050 gnd vdd FILL
X_14171_ _14171_/A _14171_/B _15651_/C gnd _12994_/B vdd AOI21X1
XFILL_4__7676_ gnd vdd FILL
X_11383_ _11383_/A _11018_/Y _11037_/Y gnd _11383_/Y vdd OAI21X1
XFILL_1__6918_ gnd vdd FILL
XFILL_4__9415_ gnd vdd FILL
XSFILL74040x67050 gnd vdd FILL
X_10334_ _10334_/Q _7781_/CLK _8670_/R vdd _10256_/Y gnd vdd DFFSR
X_13122_ _13099_/B _13122_/B gnd _13122_/Y vdd NAND2X1
XFILL_4_BUFX2_insert640 gnd vdd FILL
XFILL_1__9637_ gnd vdd FILL
XFILL_4_BUFX2_insert651 gnd vdd FILL
XSFILL34040x83050 gnd vdd FILL
XFILL_1__6849_ gnd vdd FILL
XFILL_4_BUFX2_insert662 gnd vdd FILL
XFILL_4__9346_ gnd vdd FILL
XFILL_4_BUFX2_insert673 gnd vdd FILL
X_13053_ _6876_/A _13184_/CLK _8176_/R vdd _13053_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert684 gnd vdd FILL
X_10265_ _10265_/A _10264_/A _10265_/C gnd _10265_/Y vdd OAI21X1
XFILL_4_BUFX2_insert695 gnd vdd FILL
XFILL_2__8361_ gnd vdd FILL
X_12004_ _12012_/A _12701_/A _11996_/C gnd _12006_/B vdd NAND3X1
XFILL_4__9277_ gnd vdd FILL
XFILL_5__8070_ gnd vdd FILL
XFILL_5__10830_ gnd vdd FILL
XFILL_2__7312_ gnd vdd FILL
XFILL_1__8519_ gnd vdd FILL
X_10196_ _10160_/A _9940_/B gnd _10196_/Y vdd NAND2X1
XSFILL33880x50 gnd vdd FILL
XFILL_2__10650_ gnd vdd FILL
XFILL_4__8228_ gnd vdd FILL
XFILL_1__9499_ gnd vdd FILL
XFILL_6__10031_ gnd vdd FILL
XFILL_4__11210_ gnd vdd FILL
XFILL_2__7243_ gnd vdd FILL
XFILL_5__10761_ gnd vdd FILL
XSFILL28920x63050 gnd vdd FILL
XFILL_3__11940_ gnd vdd FILL
XFILL_1__11030_ gnd vdd FILL
XFILL_4__12190_ gnd vdd FILL
XFILL_2__10581_ gnd vdd FILL
XFILL_5__12500_ gnd vdd FILL
XFILL_0__11760_ gnd vdd FILL
XFILL_2__12320_ gnd vdd FILL
XFILL_5__13480_ gnd vdd FILL
XFILL_4__11141_ gnd vdd FILL
X_13955_ _7956_/A gnd _13956_/D vdd INVX1
XFILL_5__10692_ gnd vdd FILL
XFILL_2__7174_ gnd vdd FILL
XFILL_3__11871_ gnd vdd FILL
XFILL_5__12431_ gnd vdd FILL
XFILL_5__8972_ gnd vdd FILL
X_12906_ _12904_/Y vdd _12905_/Y gnd _12906_/Y vdd OAI21X1
XFILL_0__11691_ gnd vdd FILL
XFILL_3__13610_ gnd vdd FILL
X_13886_ _13873_/Y _13885_/Y gnd _13886_/Y vdd NOR2X1
XFILL_3__10822_ gnd vdd FILL
XFILL_2__12251_ gnd vdd FILL
XFILL_4__11072_ gnd vdd FILL
XFILL_3__14590_ gnd vdd FILL
XFILL_0__13430_ gnd vdd FILL
XFILL_1__12981_ gnd vdd FILL
XFILL_0__10642_ gnd vdd FILL
X_15625_ _9760_/A gnd _15626_/A vdd INVX1
XSFILL99480x49050 gnd vdd FILL
XFILL_5__15150_ gnd vdd FILL
XFILL_5__12362_ gnd vdd FILL
XFILL_4__10023_ gnd vdd FILL
X_12837_ _12837_/A vdd _12837_/C gnd _12837_/Y vdd OAI21X1
XFILL_1_BUFX2_insert530 gnd vdd FILL
XFILL_4__14900_ gnd vdd FILL
XFILL_2__11202_ gnd vdd FILL
XSFILL74120x47050 gnd vdd FILL
XFILL_3__13541_ gnd vdd FILL
XFILL_1_BUFX2_insert541 gnd vdd FILL
XFILL_4__15880_ gnd vdd FILL
XFILL_3__10753_ gnd vdd FILL
XFILL_1__11932_ gnd vdd FILL
XFILL_1__14720_ gnd vdd FILL
XFILL_2__12182_ gnd vdd FILL
XFILL_1_BUFX2_insert552 gnd vdd FILL
XFILL_0__13361_ gnd vdd FILL
XFILL_1_BUFX2_insert563 gnd vdd FILL
XSFILL89720x26050 gnd vdd FILL
XFILL_5__14101_ gnd vdd FILL
XFILL_0__10573_ gnd vdd FILL
XFILL_5__7854_ gnd vdd FILL
XFILL_5__11313_ gnd vdd FILL
XFILL_4__14831_ gnd vdd FILL
X_15556_ _9442_/Q _15044_/C _15071_/C gnd _15556_/Y vdd NAND3X1
XFILL_5__15081_ gnd vdd FILL
XFILL_1_BUFX2_insert574 gnd vdd FILL
X_12768_ _12768_/A memoryOutData[24] gnd _12769_/C vdd NAND2X1
XFILL_0__15100_ gnd vdd FILL
XFILL_1_BUFX2_insert585 gnd vdd FILL
XFILL_5__12293_ gnd vdd FILL
XFILL_2__11133_ gnd vdd FILL
XFILL_3__16260_ gnd vdd FILL
XFILL_3__13472_ gnd vdd FILL
XFILL_1_BUFX2_insert596 gnd vdd FILL
XFILL_0__12312_ gnd vdd FILL
XFILL_3__10684_ gnd vdd FILL
XFILL_1__11863_ gnd vdd FILL
XFILL_1__14651_ gnd vdd FILL
XFILL_0__16080_ gnd vdd FILL
XFILL_0__13292_ gnd vdd FILL
XFILL_6__12603_ gnd vdd FILL
X_14507_ _14507_/A _14506_/Y gnd _14512_/C vdd NOR2X1
XFILL_5__14032_ gnd vdd FILL
XFILL_3__15211_ gnd vdd FILL
X_11719_ _11392_/Y _11739_/B gnd _11720_/B vdd NOR2X1
XFILL_5__11244_ gnd vdd FILL
XFILL_3__12423_ gnd vdd FILL
X_15487_ _15486_/Y _15487_/B gnd _15495_/A vdd NOR2X1
XFILL_4__14762_ gnd vdd FILL
XFILL_1__10814_ gnd vdd FILL
X_12699_ _12721_/B memoryOutData[1] gnd _12700_/C vdd NAND2X1
XFILL_1__13602_ gnd vdd FILL
XFILL_4__11974_ gnd vdd FILL
XFILL_3__16191_ gnd vdd FILL
XFILL_0__15031_ gnd vdd FILL
XFILL_2__15941_ gnd vdd FILL
XSFILL109480x34050 gnd vdd FILL
XFILL_2__11064_ gnd vdd FILL
XFILL_1__14582_ gnd vdd FILL
XFILL_0__12243_ gnd vdd FILL
XFILL_5__9524_ gnd vdd FILL
XFILL_1__11794_ gnd vdd FILL
XFILL_0__8830_ gnd vdd FILL
XFILL_4__13713_ gnd vdd FILL
X_14438_ _14438_/A _14430_/Y gnd _14449_/A vdd NAND2X1
XFILL_4__10925_ gnd vdd FILL
XFILL_2__10015_ gnd vdd FILL
XFILL_3__15142_ gnd vdd FILL
XFILL_5__11175_ gnd vdd FILL
XFILL_3__12354_ gnd vdd FILL
XFILL112280x73050 gnd vdd FILL
XFILL_1__16321_ gnd vdd FILL
XFILL_4__14693_ gnd vdd FILL
XFILL_2__9746_ gnd vdd FILL
XFILL_1__13533_ gnd vdd FILL
XFILL_2__6958_ gnd vdd FILL
XFILL_2__15872_ gnd vdd FILL
XFILL_1__10745_ gnd vdd FILL
XSFILL54040x14050 gnd vdd FILL
XFILL_0__12174_ gnd vdd FILL
XFILL_5__10126_ gnd vdd FILL
XFILL_4__13644_ gnd vdd FILL
XFILL_0__8761_ gnd vdd FILL
X_14369_ _7273_/Q gnd _14370_/A vdd INVX1
XFILL_3__11305_ gnd vdd FILL
XFILL_5__15983_ gnd vdd FILL
XFILL_2__14823_ gnd vdd FILL
XFILL_3__15073_ gnd vdd FILL
XFILL_2__9677_ gnd vdd FILL
XFILL_1__13464_ gnd vdd FILL
XFILL_0__11125_ gnd vdd FILL
XFILL_3__8470_ gnd vdd FILL
XFILL_1__16252_ gnd vdd FILL
XFILL_3__12285_ gnd vdd FILL
X_16108_ _10608_/Q gnd _16108_/Y vdd INVX1
XFILL_2__6889_ gnd vdd FILL
XFILL_1__10676_ gnd vdd FILL
XFILL_0__7712_ gnd vdd FILL
XFILL_5__9386_ gnd vdd FILL
XFILL_4__16363_ gnd vdd FILL
XFILL_3__14024_ gnd vdd FILL
XFILL_5__14934_ gnd vdd FILL
XFILL_5__10057_ gnd vdd FILL
XSFILL79240x80050 gnd vdd FILL
XFILL_1__12415_ gnd vdd FILL
XFILL_1__15203_ gnd vdd FILL
XSFILL43880x57050 gnd vdd FILL
XFILL_3__7421_ gnd vdd FILL
XFILL_4__13575_ gnd vdd FILL
XFILL_2__8628_ gnd vdd FILL
XFILL_3__11236_ gnd vdd FILL
XFILL_4__10787_ gnd vdd FILL
XFILL_1__16183_ gnd vdd FILL
XFILL_2__14754_ gnd vdd FILL
XFILL_2__11966_ gnd vdd FILL
XFILL_0__15933_ gnd vdd FILL
XFILL_1__13395_ gnd vdd FILL
XFILL_5__8337_ gnd vdd FILL
XFILL_0__11056_ gnd vdd FILL
X_16039_ _16036_/Y _16039_/B gnd _16044_/A vdd NOR2X1
XFILL_4__15314_ gnd vdd FILL
XFILL_4__12526_ gnd vdd FILL
XFILL_5__14865_ gnd vdd FILL
XFILL_1__15134_ gnd vdd FILL
XFILL_2__13705_ gnd vdd FILL
XFILL_3__11167_ gnd vdd FILL
XFILL_4__16294_ gnd vdd FILL
XFILL_2__10917_ gnd vdd FILL
XFILL_0__10007_ gnd vdd FILL
XFILL_3__7352_ gnd vdd FILL
XFILL_1__12346_ gnd vdd FILL
XSFILL18680x33050 gnd vdd FILL
XFILL_2__14685_ gnd vdd FILL
XFILL_5__8268_ gnd vdd FILL
XFILL_2__11897_ gnd vdd FILL
XFILL_0__15864_ gnd vdd FILL
XSFILL74200x27050 gnd vdd FILL
XFILL_5__13816_ gnd vdd FILL
XFILL_4__15245_ gnd vdd FILL
XFILL_3__10118_ gnd vdd FILL
XFILL_0__7574_ gnd vdd FILL
XFILL_4__12457_ gnd vdd FILL
XFILL_2__13636_ gnd vdd FILL
XFILL_3__15975_ gnd vdd FILL
XFILL_5__14796_ gnd vdd FILL
XFILL_1__15065_ gnd vdd FILL
XFILL_3__11098_ gnd vdd FILL
XFILL_0__14815_ gnd vdd FILL
XFILL_6__13017_ gnd vdd FILL
XFILL_1__12277_ gnd vdd FILL
XFILL_5__7219_ gnd vdd FILL
XFILL_0__15795_ gnd vdd FILL
XFILL_4__11408_ gnd vdd FILL
XFILL_5__8199_ gnd vdd FILL
XFILL_5__10959_ gnd vdd FILL
XFILL_4__15176_ gnd vdd FILL
XFILL_5__13747_ gnd vdd FILL
XFILL_1__14016_ gnd vdd FILL
XFILL_3__10049_ gnd vdd FILL
XFILL_3__9022_ gnd vdd FILL
XFILL_3__14926_ gnd vdd FILL
X_9941_ _9941_/A _9941_/B _9940_/Y gnd _9973_/D vdd OAI21X1
XFILL_4__12388_ gnd vdd FILL
XFILL_2__16355_ gnd vdd FILL
XFILL_0_BUFX2_insert13 gnd vdd FILL
XFILL_1__11228_ gnd vdd FILL
XFILL_2__10779_ gnd vdd FILL
XFILL_0_BUFX2_insert24 gnd vdd FILL
XFILL_2__13567_ gnd vdd FILL
XFILL_0__14746_ gnd vdd FILL
XFILL_0__11958_ gnd vdd FILL
XFILL_0_BUFX2_insert35 gnd vdd FILL
XFILL_4__14127_ gnd vdd FILL
XFILL_0__9244_ gnd vdd FILL
XFILL_2__15306_ gnd vdd FILL
XFILL_0_BUFX2_insert46 gnd vdd FILL
XFILL_5__13678_ gnd vdd FILL
XFILL_4__11339_ gnd vdd FILL
XFILL_0_BUFX2_insert57 gnd vdd FILL
X_9872_ _9870_/Y _9920_/B _9872_/C gnd _9950_/D vdd OAI21X1
XFILL_3__14857_ gnd vdd FILL
XFILL_2__12518_ gnd vdd FILL
XFILL_0__10909_ gnd vdd FILL
XFILL_2__16286_ gnd vdd FILL
XFILL_0_BUFX2_insert68 gnd vdd FILL
XFILL_1__11159_ gnd vdd FILL
XSFILL38840x46050 gnd vdd FILL
XFILL_0__14677_ gnd vdd FILL
XFILL_2__13498_ gnd vdd FILL
XFILL_5__12629_ gnd vdd FILL
XFILL_0__11889_ gnd vdd FILL
XFILL_0_BUFX2_insert79 gnd vdd FILL
XFILL112360x53050 gnd vdd FILL
XFILL_6__7963_ gnd vdd FILL
XFILL_5__15417_ gnd vdd FILL
XSFILL64120x79050 gnd vdd FILL
XFILL_3__13808_ gnd vdd FILL
X_8823_ _8823_/A _8823_/B gnd _8823_/Y vdd NAND2X1
XFILL_4__14058_ gnd vdd FILL
XFILL_6__14968_ gnd vdd FILL
XFILL_2__15237_ gnd vdd FILL
XFILL_5__16397_ gnd vdd FILL
XFILL_0__13628_ gnd vdd FILL
XFILL_2__12449_ gnd vdd FILL
XFILL_0__16416_ gnd vdd FILL
XFILL_3__14788_ gnd vdd FILL
XFILL_6__6914_ gnd vdd FILL
XFILL_1__15967_ gnd vdd FILL
XFILL_0__8126_ gnd vdd FILL
XFILL_4__13009_ gnd vdd FILL
XFILL_5__15348_ gnd vdd FILL
X_8754_ _8810_/Q gnd _8756_/A vdd INVX1
XFILL_3__9924_ gnd vdd FILL
XFILL_3__13739_ gnd vdd FILL
XFILL_2__15168_ gnd vdd FILL
XFILL_0__16347_ gnd vdd FILL
XFILL_1__14918_ gnd vdd FILL
XFILL_0__13559_ gnd vdd FILL
XFILL_6_BUFX2_insert735 gnd vdd FILL
XFILL_1__15898_ gnd vdd FILL
X_7705_ _7705_/A _7684_/B _7705_/C gnd _7777_/D vdd OAI21X1
XFILL_6_BUFX2_insert746 gnd vdd FILL
XFILL_0__8057_ gnd vdd FILL
XFILL_5__15279_ gnd vdd FILL
X_8685_ _8685_/Q _7021_/CLK _9062_/R vdd _8637_/Y gnd vdd DFFSR
XFILL_2__14119_ gnd vdd FILL
XFILL_3__9855_ gnd vdd FILL
XFILL_1__14849_ gnd vdd FILL
XFILL_2__15099_ gnd vdd FILL
XFILL_0__16278_ gnd vdd FILL
XFILL_3__15409_ gnd vdd FILL
X_7636_ _7598_/B _7380_/B gnd _7637_/C vdd NAND2X1
XSFILL18760x13050 gnd vdd FILL
XFILL_1__8870_ gnd vdd FILL
XSFILL8600x23050 gnd vdd FILL
XFILL_3__16389_ gnd vdd FILL
XFILL_0__15229_ gnd vdd FILL
XFILL_3__9786_ gnd vdd FILL
XFILL_1__7821_ gnd vdd FILL
X_7567_ _7568_/B _7439_/B gnd _7567_/Y vdd NAND2X1
XFILL_1_CLKBUF1_insert206 gnd vdd FILL
XFILL_1_CLKBUF1_insert217 gnd vdd FILL
XFILL_3__8737_ gnd vdd FILL
X_9306_ _9306_/Q _9306_/CLK _9306_/R vdd _9220_/Y gnd vdd DFFSR
XSFILL84280x5050 gnd vdd FILL
XFILL_0__8959_ gnd vdd FILL
XFILL_1__7752_ gnd vdd FILL
X_7498_ _7538_/Q gnd _7498_/Y vdd INVX1
XFILL_4__7461_ gnd vdd FILL
X_9237_ _9238_/B _7061_/B gnd _9238_/C vdd NAND2X1
XFILL_1__7683_ gnd vdd FILL
XFILL_3__7619_ gnd vdd FILL
XSFILL38920x26050 gnd vdd FILL
XFILL112440x33050 gnd vdd FILL
XFILL_3__8599_ gnd vdd FILL
XFILL_1__9422_ gnd vdd FILL
XFILL_3_BUFX2_insert603 gnd vdd FILL
XSFILL49560x77050 gnd vdd FILL
X_9168_ _9204_/Q gnd _9170_/A vdd INVX1
XFILL_3_BUFX2_insert614 gnd vdd FILL
XFILL_4__9131_ gnd vdd FILL
XSFILL89160x63050 gnd vdd FILL
XFILL_3_BUFX2_insert625 gnd vdd FILL
X_10050_ _10054_/B _6978_/B gnd _10050_/Y vdd NAND2X1
XFILL_3_BUFX2_insert636 gnd vdd FILL
X_8119_ _8117_/Y _8118_/A _8119_/C gnd _8171_/D vdd OAI21X1
XFILL_1__9353_ gnd vdd FILL
XFILL_3_BUFX2_insert647 gnd vdd FILL
X_9099_ _9099_/A gnd _9101_/A vdd INVX1
XFILL_3_BUFX2_insert658 gnd vdd FILL
XFILL_3_BUFX2_insert669 gnd vdd FILL
XSFILL79400x40050 gnd vdd FILL
XSFILL3640x66050 gnd vdd FILL
XFILL_4__8013_ gnd vdd FILL
XFILL_1__9284_ gnd vdd FILL
XSFILL28840x78050 gnd vdd FILL
XSFILL94280x54050 gnd vdd FILL
XFILL_1__8235_ gnd vdd FILL
X_13740_ _14697_/C gnd _13854_/B vdd INVX8
X_10952_ _12779_/A _12782_/A gnd _10952_/Y vdd NOR2X1
XSFILL69080x30050 gnd vdd FILL
XSFILL44040x8050 gnd vdd FILL
XSFILL33960x69050 gnd vdd FILL
XFILL_1__7117_ gnd vdd FILL
X_13671_ _7002_/Q gnd _13671_/Y vdd INVX1
XFILL_1__8097_ gnd vdd FILL
X_10883_ _12792_/Q gnd _10883_/Y vdd INVX1
XFILL_4__8915_ gnd vdd FILL
X_15410_ _15180_/C _15409_/Y _15410_/C _15410_/D gnd _15410_/Y vdd OAI22X1
X_12622_ vdd memoryOutData[18] gnd _12623_/C vdd NAND2X1
XFILL_4__9895_ gnd vdd FILL
X_16390_ _16390_/A gnd _16392_/A vdd INVX1
XFILL_1__7048_ gnd vdd FILL
XFILL_2__7930_ gnd vdd FILL
XFILL_0_BUFX2_insert504 gnd vdd FILL
XFILL_4__8846_ gnd vdd FILL
XFILL_0_BUFX2_insert515 gnd vdd FILL
X_15341_ _15341_/A _15646_/D gnd _15341_/Y vdd NOR2X1
X_12553_ _12553_/Q _13175_/CLK _12536_/R vdd _12495_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert526 gnd vdd FILL
XFILL_0_BUFX2_insert537 gnd vdd FILL
XFILL_2__7861_ gnd vdd FILL
XFILL_0_BUFX2_insert548 gnd vdd FILL
XSFILL89240x43050 gnd vdd FILL
XFILL_0_BUFX2_insert559 gnd vdd FILL
X_11504_ _11492_/Y _11493_/Y _11504_/C gnd _12089_/A vdd OAI21X1
XFILL_5__7570_ gnd vdd FILL
XFILL_4__8777_ gnd vdd FILL
XFILL_2__9600_ gnd vdd FILL
X_15272_ _15269_/Y _15272_/B gnd _15273_/C vdd NOR2X1
X_12484_ _12388_/A gnd _12484_/Y vdd INVX1
XFILL_1__8999_ gnd vdd FILL
XFILL_4__7728_ gnd vdd FILL
X_14223_ _14222_/Y _13860_/B _13871_/D _14223_/D gnd _14223_/Y vdd OAI22X1
XSFILL13320x79050 gnd vdd FILL
X_11435_ _11435_/A _11294_/Y gnd _11435_/Y vdd NOR2X1
XFILL_2__9531_ gnd vdd FILL
XFILL_1__10530_ gnd vdd FILL
XFILL_4__11690_ gnd vdd FILL
XFILL_5__9240_ gnd vdd FILL
X_14154_ _14145_/Y _14146_/Y _14154_/C gnd _14170_/B vdd NAND3X1
XSFILL68520x44050 gnd vdd FILL
X_11366_ _11362_/Y _11366_/B _11366_/C gnd _11366_/Y vdd OAI21X1
XFILL_3__12070_ gnd vdd FILL
XFILL_5__12980_ gnd vdd FILL
XFILL_4__10641_ gnd vdd FILL
XFILL_2__9462_ gnd vdd FILL
XFILL_2__11820_ gnd vdd FILL
X_10317_ _10355_/Q gnd _10317_/Y vdd INVX1
X_13105_ _13105_/A _13168_/B _13104_/Y gnd _13183_/D vdd OAI21X1
XFILL_5__9171_ gnd vdd FILL
XSFILL69160x10050 gnd vdd FILL
XCLKBUF1_insert205 CLKBUF1_insert218/A gnd _9963_/CLK vdd CLKBUF1
XFILL_5__11931_ gnd vdd FILL
XFILL_4_BUFX2_insert470 gnd vdd FILL
XFILL_3__11021_ gnd vdd FILL
XCLKBUF1_insert216 CLKBUF1_insert216/A gnd _8025_/CLK vdd CLKBUF1
XFILL_4__13360_ gnd vdd FILL
XFILL_4_BUFX2_insert481 gnd vdd FILL
XFILL_1__12200_ gnd vdd FILL
X_11297_ _11582_/C _11146_/B gnd _11297_/Y vdd NAND2X1
X_14085_ _14085_/A _14085_/B _14085_/C gnd _14096_/B vdd NAND3X1
XFILL_4__10572_ gnd vdd FILL
XFILL_4_BUFX2_insert492 gnd vdd FILL
XFILL_5__8122_ gnd vdd FILL
XFILL_2__9393_ gnd vdd FILL
XFILL_2__11751_ gnd vdd FILL
XFILL_1__10392_ gnd vdd FILL
X_10248_ _10332_/Q gnd _10248_/Y vdd INVX1
X_13036_ vdd _13036_/B gnd _13037_/C vdd NAND2X1
XFILL_4__12311_ gnd vdd FILL
XFILL_5__14650_ gnd vdd FILL
XFILL_5__11862_ gnd vdd FILL
XFILL_4__13291_ gnd vdd FILL
XFILL_2__10702_ gnd vdd FILL
XFILL_2__8344_ gnd vdd FILL
XFILL_1__12131_ gnd vdd FILL
XFILL_2__14470_ gnd vdd FILL
XSFILL104520x2050 gnd vdd FILL
XFILL_2__11682_ gnd vdd FILL
XFILL_0__12861_ gnd vdd FILL
XFILL_5__10813_ gnd vdd FILL
XFILL_5__13601_ gnd vdd FILL
XFILL_4__15030_ gnd vdd FILL
XFILL_6__15940_ gnd vdd FILL
XFILL_5__14581_ gnd vdd FILL
XFILL_4__12242_ gnd vdd FILL
X_10179_ _10179_/A _10193_/A _10179_/C gnd _10223_/D vdd OAI21X1
XFILL_0__14600_ gnd vdd FILL
XFILL_2__13421_ gnd vdd FILL
XFILL_2__10633_ gnd vdd FILL
XFILL_3__15760_ gnd vdd FILL
XFILL_5__11793_ gnd vdd FILL
XFILL_3__12972_ gnd vdd FILL
XFILL_1__12062_ gnd vdd FILL
XFILL_2__8275_ gnd vdd FILL
XFILL_0__11812_ gnd vdd FILL
XFILL_0__15580_ gnd vdd FILL
XFILL_5__16320_ gnd vdd FILL
XFILL_5__13532_ gnd vdd FILL
XFILL_5__10744_ gnd vdd FILL
XFILL_3__14711_ gnd vdd FILL
XFILL_0__7290_ gnd vdd FILL
X_14987_ _15687_/A _14987_/B _16199_/C _13453_/Y gnd _14987_/Y vdd OAI22X1
XFILL_3__11923_ gnd vdd FILL
XFILL_2__7226_ gnd vdd FILL
XFILL_4__12173_ gnd vdd FILL
XFILL_1__11013_ gnd vdd FILL
XFILL_2__16140_ gnd vdd FILL
XFILL_2__13352_ gnd vdd FILL
XFILL_3__15691_ gnd vdd FILL
XFILL_0__14531_ gnd vdd FILL
XFILL_2__10564_ gnd vdd FILL
XSFILL109480x29050 gnd vdd FILL
XFILL_0__11743_ gnd vdd FILL
XFILL_5__13463_ gnd vdd FILL
XFILL_3_CLKBUF1_insert150 gnd vdd FILL
X_13938_ _7828_/A gnd _13940_/A vdd INVX1
XFILL_4__11124_ gnd vdd FILL
XFILL_5__16251_ gnd vdd FILL
XFILL_3__14642_ gnd vdd FILL
XFILL_2__12303_ gnd vdd FILL
XFILL_3_CLKBUF1_insert161 gnd vdd FILL
XFILL_5__10675_ gnd vdd FILL
XFILL_2__13283_ gnd vdd FILL
XFILL_1__15821_ gnd vdd FILL
XFILL_3_CLKBUF1_insert172 gnd vdd FILL
XFILL_2__16071_ gnd vdd FILL
XFILL_3__11854_ gnd vdd FILL
XFILL_2__10495_ gnd vdd FILL
XFILL112280x68050 gnd vdd FILL
XFILL_0__14462_ gnd vdd FILL
XFILL_3_CLKBUF1_insert183 gnd vdd FILL
XFILL_3_CLKBUF1_insert194 gnd vdd FILL
XFILL_5__12414_ gnd vdd FILL
XFILL_5__15202_ gnd vdd FILL
XFILL_0__11674_ gnd vdd FILL
XFILL_5__8955_ gnd vdd FILL
XFILL_5__16182_ gnd vdd FILL
XFILL_6__14753_ gnd vdd FILL
X_13869_ _10638_/A gnd _13869_/Y vdd INVX1
XFILL_3__10805_ gnd vdd FILL
XFILL_0__16201_ gnd vdd FILL
XFILL_4__15932_ gnd vdd FILL
XFILL_2__15022_ gnd vdd FILL
XFILL_5__13394_ gnd vdd FILL
XFILL_2__12234_ gnd vdd FILL
XFILL_4__11055_ gnd vdd FILL
XFILL_3__14573_ gnd vdd FILL
XFILL_0__13413_ gnd vdd FILL
XFILL_2__7088_ gnd vdd FILL
XFILL_0__10625_ gnd vdd FILL
XFILL_3__7970_ gnd vdd FILL
XFILL_3__11785_ gnd vdd FILL
XFILL_1__15752_ gnd vdd FILL
XFILL_1__12964_ gnd vdd FILL
XFILL_0__14393_ gnd vdd FILL
XFILL_5__15133_ gnd vdd FILL
X_15608_ _15608_/A _15607_/Y gnd _15609_/C vdd NAND2X1
XFILL_5__8886_ gnd vdd FILL
XFILL_5__12345_ gnd vdd FILL
XFILL_3__16312_ gnd vdd FILL
XFILL_1_BUFX2_insert360 gnd vdd FILL
XFILL_4__10006_ gnd vdd FILL
XFILL_3__13524_ gnd vdd FILL
XFILL_1_BUFX2_insert371 gnd vdd FILL
XSFILL79240x75050 gnd vdd FILL
XFILL_3__6921_ gnd vdd FILL
XFILL_6__11896_ gnd vdd FILL
XFILL_1__14703_ gnd vdd FILL
XFILL_2__12165_ gnd vdd FILL
XFILL_0__16132_ gnd vdd FILL
XFILL_1_BUFX2_insert382 gnd vdd FILL
XFILL_4__15863_ gnd vdd FILL
XFILL_0__13344_ gnd vdd FILL
XFILL_1__11915_ gnd vdd FILL
XFILL_1__15683_ gnd vdd FILL
XFILL_1__12895_ gnd vdd FILL
XFILL_0__10556_ gnd vdd FILL
XFILL_1_BUFX2_insert393 gnd vdd FILL
XFILL_5__7837_ gnd vdd FILL
XFILL_0__9931_ gnd vdd FILL
X_15539_ _16036_/A _14052_/Y _14060_/Y _15376_/B gnd _15541_/A vdd OAI22X1
XFILL_5__15064_ gnd vdd FILL
XFILL_3__16243_ gnd vdd FILL
XFILL_4__14814_ gnd vdd FILL
XFILL_5_BUFX2_insert709 gnd vdd FILL
XFILL_5__12276_ gnd vdd FILL
X_8470_ _8470_/A _8469_/A _8470_/C gnd _8544_/D vdd OAI21X1
XFILL_2__11116_ gnd vdd FILL
XFILL_3__9640_ gnd vdd FILL
XFILL_3__13455_ gnd vdd FILL
XFILL_4__15794_ gnd vdd FILL
XSFILL28840x8050 gnd vdd FILL
XFILL_1__14634_ gnd vdd FILL
XFILL_3__6852_ gnd vdd FILL
XFILL_2__12096_ gnd vdd FILL
XFILL_3__10667_ gnd vdd FILL
XSFILL18680x28050 gnd vdd FILL
XFILL_0__16063_ gnd vdd FILL
XFILL_1__11846_ gnd vdd FILL
XFILL_0__13275_ gnd vdd FILL
XFILL_5__14015_ gnd vdd FILL
XSFILL8520x38050 gnd vdd FILL
XFILL_0__10487_ gnd vdd FILL
X_7421_ _7470_/B _9981_/B gnd _7421_/Y vdd NAND2X1
XFILL_5__11227_ gnd vdd FILL
XFILL_3__12406_ gnd vdd FILL
XFILL_0__9862_ gnd vdd FILL
XFILL_4__14745_ gnd vdd FILL
XFILL_2__15924_ gnd vdd FILL
XFILL_3__16174_ gnd vdd FILL
XFILL_4__11957_ gnd vdd FILL
XFILL_0__15014_ gnd vdd FILL
XFILL_2__11047_ gnd vdd FILL
XFILL_5__9507_ gnd vdd FILL
XSFILL84360x66050 gnd vdd FILL
XFILL_3__13386_ gnd vdd FILL
XFILL_0__12226_ gnd vdd FILL
XFILL_1__14565_ gnd vdd FILL
XFILL_1__11777_ gnd vdd FILL
XFILL_4__10908_ gnd vdd FILL
X_7352_ _7404_/Q gnd _7352_/Y vdd INVX1
XFILL_5__11158_ gnd vdd FILL
XFILL_3__15125_ gnd vdd FILL
XFILL_5__7699_ gnd vdd FILL
XFILL_2__9729_ gnd vdd FILL
XFILL_3__8522_ gnd vdd FILL
XFILL_1__16304_ gnd vdd FILL
XFILL_4__14676_ gnd vdd FILL
XFILL_0__9793_ gnd vdd FILL
XFILL_3__12337_ gnd vdd FILL
XFILL_4__11888_ gnd vdd FILL
XFILL_2__15855_ gnd vdd FILL
XFILL_1__13516_ gnd vdd FILL
XFILL_1__14496_ gnd vdd FILL
XFILL_0__12157_ gnd vdd FILL
XSFILL59160x42050 gnd vdd FILL
XFILL_5__10109_ gnd vdd FILL
XFILL_4__13627_ gnd vdd FILL
XFILL_0__8744_ gnd vdd FILL
XFILL_4__16415_ gnd vdd FILL
X_7283_ _7245_/A _8429_/CLK _9203_/R vdd _7283_/D gnd vdd DFFSR
XFILL_2__14806_ gnd vdd FILL
XFILL_3__15056_ gnd vdd FILL
XFILL_5__15966_ gnd vdd FILL
XFILL_5__11089_ gnd vdd FILL
XFILL_1__16235_ gnd vdd FILL
XFILL_1__13447_ gnd vdd FILL
XFILL_3__12268_ gnd vdd FILL
XFILL_3__8453_ gnd vdd FILL
XFILL_0__11108_ gnd vdd FILL
XFILL_1__10659_ gnd vdd FILL
XFILL_2__15786_ gnd vdd FILL
XFILL_2__12998_ gnd vdd FILL
XFILL_5__9369_ gnd vdd FILL
XFILL_0__12088_ gnd vdd FILL
X_9022_ _9022_/A gnd _9022_/Y vdd INVX1
XFILL_4__16346_ gnd vdd FILL
XFILL_3__14007_ gnd vdd FILL
XFILL112360x48050 gnd vdd FILL
XFILL_5__14917_ gnd vdd FILL
XFILL_4__13558_ gnd vdd FILL
XFILL_3__11219_ gnd vdd FILL
XFILL_5__15897_ gnd vdd FILL
XFILL_2__14737_ gnd vdd FILL
XFILL_0__15916_ gnd vdd FILL
XFILL_3__8384_ gnd vdd FILL
XFILL_1__13378_ gnd vdd FILL
XFILL_1__16166_ gnd vdd FILL
XFILL_2__11949_ gnd vdd FILL
XFILL_3__12199_ gnd vdd FILL
XFILL_0__11039_ gnd vdd FILL
XFILL_4__12509_ gnd vdd FILL
XFILL_0__7626_ gnd vdd FILL
XFILL_5__14848_ gnd vdd FILL
XSFILL109400x73050 gnd vdd FILL
XFILL_4__16277_ gnd vdd FILL
XFILL_3__7335_ gnd vdd FILL
XFILL_1__12329_ gnd vdd FILL
XFILL_1__15117_ gnd vdd FILL
XFILL_4__13489_ gnd vdd FILL
XFILL_1__16097_ gnd vdd FILL
XSFILL8680x1050 gnd vdd FILL
XFILL_2__14668_ gnd vdd FILL
XFILL_0__15847_ gnd vdd FILL
XFILL_4__15228_ gnd vdd FILL
XFILL_2__16407_ gnd vdd FILL
XSFILL89400x1050 gnd vdd FILL
XFILL_0__7557_ gnd vdd FILL
XFILL_2__13619_ gnd vdd FILL
XFILL_3__15958_ gnd vdd FILL
XFILL_5__14779_ gnd vdd FILL
XFILL_1__15048_ gnd vdd FILL
XFILL_2__14599_ gnd vdd FILL
XFILL_0__15778_ gnd vdd FILL
X_9924_ _9924_/A gnd _9924_/Y vdd INVX1
XFILL_3__9005_ gnd vdd FILL
XFILL_4__15159_ gnd vdd FILL
XSFILL114520x64050 gnd vdd FILL
XFILL_0__7488_ gnd vdd FILL
XFILL_2__16338_ gnd vdd FILL
XSFILL8600x18050 gnd vdd FILL
XFILL_3__14909_ gnd vdd FILL
XFILL_3__15889_ gnd vdd FILL
XFILL_0__14729_ gnd vdd FILL
XFILL_3__7197_ gnd vdd FILL
XFILL_0__9227_ gnd vdd FILL
XFILL_1__8020_ gnd vdd FILL
XFILL_5__16449_ gnd vdd FILL
XSFILL33800x11050 gnd vdd FILL
X_9855_ _9945_/Q gnd _9857_/A vdd INVX1
XFILL_2__16269_ gnd vdd FILL
X_8806_ _8806_/Q _7282_/CLK _8166_/R vdd _8744_/Y gnd vdd DFFSR
XFILL_0__9158_ gnd vdd FILL
XFILL_6_BUFX2_insert510 gnd vdd FILL
X_6998_ _6998_/Q _6998_/CLK _7644_/R vdd _6998_/D gnd vdd DFFSR
X_9786_ _9786_/A _9785_/A _9786_/C gnd _9836_/D vdd OAI21X1
XFILL_6_BUFX2_insert521 gnd vdd FILL
XFILL_4__6961_ gnd vdd FILL
XFILL_0__8109_ gnd vdd FILL
XFILL_0__9089_ gnd vdd FILL
X_8737_ _8759_/B _8225_/B gnd _8738_/C vdd NAND2X1
XFILL_3__9907_ gnd vdd FILL
XFILL_4__8700_ gnd vdd FILL
XBUFX2_insert609 _15035_/Y gnd _16141_/A vdd BUFX2
XFILL111960x21050 gnd vdd FILL
XFILL112440x28050 gnd vdd FILL
XFILL_4__9680_ gnd vdd FILL
XFILL_4__6892_ gnd vdd FILL
XFILL_6_BUFX2_insert587 gnd vdd FILL
X_8668_ _8668_/Q _8046_/CLK _8670_/R vdd _8668_/D gnd vdd DFFSR
XFILL_4__8631_ gnd vdd FILL
XFILL112040x30050 gnd vdd FILL
XFILL_1__8853_ gnd vdd FILL
X_7619_ _7619_/A _7570_/A _7619_/C gnd _7663_/D vdd OAI21X1
X_8599_ _8599_/A gnd _8601_/A vdd INVX1
XSFILL8600x9050 gnd vdd FILL
XFILL_3__9769_ gnd vdd FILL
XFILL_6__9478_ gnd vdd FILL
XFILL_1__7804_ gnd vdd FILL
XFILL_1__8784_ gnd vdd FILL
X_11220_ _11220_/A _11220_/B _11219_/Y gnd _11342_/C vdd OAI21X1
XFILL_4__8493_ gnd vdd FILL
XSFILL94280x49050 gnd vdd FILL
XFILL_1__7735_ gnd vdd FILL
XFILL_4__7444_ gnd vdd FILL
X_11151_ _11150_/Y _11403_/A gnd _11156_/A vdd NAND2X1
XSFILL69080x25050 gnd vdd FILL
X_10102_ _10198_/Q gnd _10104_/A vdd INVX1
XFILL_3_BUFX2_insert400 gnd vdd FILL
XFILL_4__7375_ gnd vdd FILL
XFILL_3_BUFX2_insert411 gnd vdd FILL
XFILL_1__9405_ gnd vdd FILL
XFILL_3_BUFX2_insert422 gnd vdd FILL
X_11082_ _12258_/Y _11071_/Y gnd _11393_/A vdd NOR2X1
XFILL_3_BUFX2_insert433 gnd vdd FILL
XSFILL7880x66050 gnd vdd FILL
XFILL_3_BUFX2_insert444 gnd vdd FILL
XFILL_4__9114_ gnd vdd FILL
XFILL_1__7597_ gnd vdd FILL
XFILL_3_BUFX2_insert455 gnd vdd FILL
X_10033_ _10031_/Y _10024_/B _10033_/C gnd _10089_/D vdd OAI21X1
X_14910_ _9680_/A gnd _14910_/Y vdd INVX1
XFILL_3_BUFX2_insert466 gnd vdd FILL
XFILL_1__9336_ gnd vdd FILL
XFILL_3_BUFX2_insert477 gnd vdd FILL
X_15890_ _15890_/A _15890_/B _15889_/Y gnd _15891_/B vdd NOR3X1
XFILL_3_BUFX2_insert488 gnd vdd FILL
XFILL_4__9045_ gnd vdd FILL
XFILL_3_BUFX2_insert499 gnd vdd FILL
X_14841_ _14839_/Y _13846_/A _14575_/C _14840_/Y gnd _14841_/Y vdd OAI22X1
XSFILL105160x62050 gnd vdd FILL
XFILL_1__9267_ gnd vdd FILL
XFILL_2__8060_ gnd vdd FILL
XFILL112120x10050 gnd vdd FILL
XFILL_1__8218_ gnd vdd FILL
X_14772_ _14772_/A _14771_/Y gnd _14772_/Y vdd NOR2X1
X_11984_ _11999_/A _12343_/A _11999_/C gnd _11990_/A vdd NAND3X1
XFILL_0_BUFX2_insert5 gnd vdd FILL
X_13723_ _10501_/A gnd _13725_/D vdd INVX1
X_10935_ _10935_/A _10934_/Y gnd _10936_/C vdd NOR2X1
XFILL_1__8149_ gnd vdd FILL
XFILL_4_CLKBUF1_insert201 gnd vdd FILL
XFILL_2__10280_ gnd vdd FILL
XSFILL53720x79050 gnd vdd FILL
XFILL_5__8740_ gnd vdd FILL
XSFILL94360x29050 gnd vdd FILL
XFILL_4_CLKBUF1_insert212 gnd vdd FILL
X_16442_ _16076_/A _7535_/CLK _7648_/R vdd _16398_/Y gnd vdd DFFSR
XFILL_4_CLKBUF1_insert223 gnd vdd FILL
X_13654_ _13653_/Y _13795_/B _14489_/C _15213_/A gnd _13655_/B vdd OAI22X1
X_10866_ _14793_/C _7662_/CLK _9454_/R vdd _10828_/Y gnd vdd DFFSR
XFILL_5__10391_ gnd vdd FILL
XFILL_2__8962_ gnd vdd FILL
XFILL_0__10410_ gnd vdd FILL
XFILL_3__11570_ gnd vdd FILL
XFILL_0_BUFX2_insert301 gnd vdd FILL
X_12605_ _12605_/A vdd _12604_/Y gnd _12675_/D vdd OAI21X1
XFILL_5__12130_ gnd vdd FILL
XFILL_4__9878_ gnd vdd FILL
XFILL_0__11390_ gnd vdd FILL
X_16373_ gnd gnd gnd _16374_/C vdd NAND2X1
XFILL_6__11681_ gnd vdd FILL
XFILL_0_BUFX2_insert312 gnd vdd FILL
X_13585_ _7641_/Q gnd _13587_/D vdd INVX1
XFILL_3__10521_ gnd vdd FILL
XFILL_4__12860_ gnd vdd FILL
XFILL_1__11700_ gnd vdd FILL
XFILL_0_BUFX2_insert323 gnd vdd FILL
XSFILL68920x60050 gnd vdd FILL
XFILL_0_BUFX2_insert334 gnd vdd FILL
X_10797_ _10797_/A _7853_/B gnd _10798_/C vdd NAND2X1
XFILL_2__8893_ gnd vdd FILL
XFILL_5__7622_ gnd vdd FILL
XFILL_4__8829_ gnd vdd FILL
X_15324_ _15324_/A _15318_/Y _15323_/Y gnd _15324_/Y vdd NAND3X1
XFILL_0_BUFX2_insert345 gnd vdd FILL
XFILL_0_BUFX2_insert356 gnd vdd FILL
XFILL_5__12061_ gnd vdd FILL
X_12536_ _11991_/B _12537_/CLK _12536_/R vdd _12444_/Y gnd vdd DFFSR
XFILL_4__11811_ gnd vdd FILL
XFILL_3__13240_ gnd vdd FILL
XFILL_0_BUFX2_insert367 gnd vdd FILL
XSFILL104360x14050 gnd vdd FILL
XFILL_2__7844_ gnd vdd FILL
XFILL_3__10452_ gnd vdd FILL
XFILL_0_BUFX2_insert378 gnd vdd FILL
XFILL_1__11631_ gnd vdd FILL
XFILL_2__13970_ gnd vdd FILL
XFILL_5__7553_ gnd vdd FILL
XFILL_0__10272_ gnd vdd FILL
XFILL_0_BUFX2_insert389 gnd vdd FILL
XFILL_5__11012_ gnd vdd FILL
X_15255_ _15369_/A _15255_/B _15255_/C _15369_/D gnd _15256_/B vdd OAI22X1
XFILL_4__14530_ gnd vdd FILL
XFILL_6__10563_ gnd vdd FILL
X_12467_ vdd _12467_/B gnd _12467_/Y vdd NAND2X1
XFILL_4__11742_ gnd vdd FILL
XFILL_3__10383_ gnd vdd FILL
XFILL_0__12011_ gnd vdd FILL
XFILL_3__13171_ gnd vdd FILL
XFILL_1__14350_ gnd vdd FILL
XFILL_1__11562_ gnd vdd FILL
X_14206_ _8611_/A gnd _14208_/A vdd INVX1
XFILL_5__7484_ gnd vdd FILL
XFILL_5__15820_ gnd vdd FILL
X_11418_ _11359_/Y _11360_/Y _11417_/Y gnd _12105_/A vdd OAI21X1
XFILL_1__13301_ gnd vdd FILL
XFILL_4__14461_ gnd vdd FILL
X_15186_ _13594_/A gnd _15187_/B vdd INVX1
XFILL_3__12122_ gnd vdd FILL
XSFILL89320x18050 gnd vdd FILL
XFILL_2__9514_ gnd vdd FILL
X_12398_ _12380_/A _12621_/A gnd _12399_/C vdd NAND2X1
XFILL_2__15640_ gnd vdd FILL
XFILL_4__11673_ gnd vdd FILL
XFILL_1__10513_ gnd vdd FILL
XFILL_2__12852_ gnd vdd FILL
XFILL_5__9223_ gnd vdd FILL
XFILL_1__14281_ gnd vdd FILL
XSFILL99480x62050 gnd vdd FILL
XFILL_4__16200_ gnd vdd FILL
XFILL_1__11493_ gnd vdd FILL
XFILL_4__13412_ gnd vdd FILL
X_14137_ _7012_/Q gnd _14137_/Y vdd INVX1
XFILL_4__10624_ gnd vdd FILL
XSFILL74120x60050 gnd vdd FILL
XFILL_5__15751_ gnd vdd FILL
X_11349_ _10996_/Y _11349_/B _11231_/Y _11484_/B gnd _11350_/A vdd OAI22X1
XFILL_1__13232_ gnd vdd FILL
XFILL_1__16020_ gnd vdd FILL
XFILL_5__12963_ gnd vdd FILL
XFILL_3__12053_ gnd vdd FILL
XFILL_4__14392_ gnd vdd FILL
XFILL_2__11803_ gnd vdd FILL
XFILL_1__10444_ gnd vdd FILL
XFILL_2__15571_ gnd vdd FILL
XFILL_2__12783_ gnd vdd FILL
XFILL_5_BUFX2_insert1002 gnd vdd FILL
XFILL_5__9154_ gnd vdd FILL
XFILL_0__13962_ gnd vdd FILL
XFILL_5__14702_ gnd vdd FILL
XFILL_4__16131_ gnd vdd FILL
XFILL_4__13343_ gnd vdd FILL
XFILL_0__8460_ gnd vdd FILL
XFILL_5__11914_ gnd vdd FILL
XFILL_5_BUFX2_insert1013 gnd vdd FILL
X_14068_ _14068_/A _13775_/B _14068_/C _14067_/Y gnd _14068_/Y vdd OAI22X1
XFILL_3__11004_ gnd vdd FILL
XFILL_5__15682_ gnd vdd FILL
XFILL_5__12894_ gnd vdd FILL
XFILL_4__10555_ gnd vdd FILL
XFILL_2__14522_ gnd vdd FILL
XFILL_5_BUFX2_insert1024 gnd vdd FILL
XFILL_5_BUFX2_insert1035 gnd vdd FILL
XFILL_0__15701_ gnd vdd FILL
XFILL_2__9376_ gnd vdd FILL
XFILL_1__13163_ gnd vdd FILL
XFILL_0__12913_ gnd vdd FILL
XFILL_2__11734_ gnd vdd FILL
XFILL_5__8105_ gnd vdd FILL
XFILL_1__10375_ gnd vdd FILL
XFILL_5_BUFX2_insert1046 gnd vdd FILL
XFILL_5_BUFX2_insert1057 gnd vdd FILL
X_13019_ _13017_/Y vdd _13019_/C gnd _13069_/D vdd OAI21X1
XFILL_0__13893_ gnd vdd FILL
XFILL_5__9085_ gnd vdd FILL
XSFILL13800x75050 gnd vdd FILL
XFILL_5__14633_ gnd vdd FILL
XFILL_3__15812_ gnd vdd FILL
XFILL_4__16062_ gnd vdd FILL
XFILL_4__13274_ gnd vdd FILL
XFILL_5_BUFX2_insert1068 gnd vdd FILL
XFILL_1__12114_ gnd vdd FILL
XFILL_2__8327_ gnd vdd FILL
XFILL_3__7120_ gnd vdd FILL
XFILL_0__8391_ gnd vdd FILL
XFILL_5__11845_ gnd vdd FILL
XFILL_2__14453_ gnd vdd FILL
XFILL_4__10486_ gnd vdd FILL
XFILL_0__12844_ gnd vdd FILL
XFILL_0__15632_ gnd vdd FILL
XFILL_1__13094_ gnd vdd FILL
XFILL_2__11665_ gnd vdd FILL
XFILL_4__15013_ gnd vdd FILL
XFILL_0__7342_ gnd vdd FILL
XFILL_4__12225_ gnd vdd FILL
XFILL_5__14564_ gnd vdd FILL
XFILL_2__13404_ gnd vdd FILL
X_7970_ _7970_/A _7970_/B _7970_/C gnd _8036_/D vdd OAI21X1
XFILL_5__11776_ gnd vdd FILL
XFILL_3__15743_ gnd vdd FILL
XFILL_3__7051_ gnd vdd FILL
XFILL_2__10616_ gnd vdd FILL
XFILL_1__12045_ gnd vdd FILL
XFILL_2__8258_ gnd vdd FILL
XFILL_3__12955_ gnd vdd FILL
XFILL_0__15563_ gnd vdd FILL
XFILL_2__14384_ gnd vdd FILL
XFILL_2__11596_ gnd vdd FILL
XFILL_0__12775_ gnd vdd FILL
XFILL_5__16303_ gnd vdd FILL
XSFILL114440x79050 gnd vdd FILL
X_6921_ _6988_/B _6921_/B gnd _6922_/C vdd NAND2X1
XFILL_5__13515_ gnd vdd FILL
XFILL_5__14495_ gnd vdd FILL
XFILL_3__11906_ gnd vdd FILL
XFILL_2__16123_ gnd vdd FILL
XFILL_4__12156_ gnd vdd FILL
XFILL_2__7209_ gnd vdd FILL
XFILL_2__13335_ gnd vdd FILL
XFILL_3__15674_ gnd vdd FILL
XFILL_0__14514_ gnd vdd FILL
XFILL_3__12886_ gnd vdd FILL
XFILL_0__11726_ gnd vdd FILL
XFILL_2__8189_ gnd vdd FILL
XFILL_2__10547_ gnd vdd FILL
XFILL_6__14805_ gnd vdd FILL
XFILL_0__15494_ gnd vdd FILL
XFILL_0__9012_ gnd vdd FILL
XFILL_5__16234_ gnd vdd FILL
XFILL_5__9987_ gnd vdd FILL
XFILL_4__11107_ gnd vdd FILL
X_9640_ _9640_/A _9639_/A _9640_/C gnd _9702_/D vdd OAI21X1
XSFILL43880x70050 gnd vdd FILL
XFILL_3__14625_ gnd vdd FILL
XFILL_5__10658_ gnd vdd FILL
XFILL_5__13446_ gnd vdd FILL
X_6852_ _6852_/A gnd memoryAddress[14] vdd BUFX2
XFILL_4__12087_ gnd vdd FILL
XFILL_1__15804_ gnd vdd FILL
XFILL_3_BUFX2_insert1050 gnd vdd FILL
XFILL_2__16054_ gnd vdd FILL
XFILL_3__11837_ gnd vdd FILL
XFILL_2__13266_ gnd vdd FILL
XSFILL98920x76050 gnd vdd FILL
XFILL_3_BUFX2_insert1061 gnd vdd FILL
XFILL_0__14445_ gnd vdd FILL
XSFILL59160x37050 gnd vdd FILL
XFILL_0__11657_ gnd vdd FILL
XFILL_3_BUFX2_insert1072 gnd vdd FILL
XFILL_1__13996_ gnd vdd FILL
XFILL_4__15915_ gnd vdd FILL
XFILL_5__13377_ gnd vdd FILL
XFILL_5__16165_ gnd vdd FILL
XFILL_2__15005_ gnd vdd FILL
X_9571_ _9501_/A _6999_/CLK _7000_/R vdd _9503_/Y gnd vdd DFFSR
XFILL_4__11038_ gnd vdd FILL
XFILL_3__14556_ gnd vdd FILL
XFILL_2__12217_ gnd vdd FILL
XFILL_3__7953_ gnd vdd FILL
XFILL_3__11768_ gnd vdd FILL
XFILL_1__15735_ gnd vdd FILL
XSFILL74200x40050 gnd vdd FILL
XFILL_0__14376_ gnd vdd FILL
XFILL_5__8869_ gnd vdd FILL
X_8522_ _8522_/A gnd _8524_/A vdd INVX1
XFILL_5__12328_ gnd vdd FILL
XFILL_0__11588_ gnd vdd FILL
XFILL_5__15116_ gnd vdd FILL
XFILL_6__14667_ gnd vdd FILL
XFILL_3__13507_ gnd vdd FILL
XFILL_3__6904_ gnd vdd FILL
XFILL_5__16096_ gnd vdd FILL
XFILL_4__15846_ gnd vdd FILL
XFILL_5_BUFX2_insert506 gnd vdd FILL
XFILL_0__13327_ gnd vdd FILL
XFILL_3__14487_ gnd vdd FILL
XFILL_2__12148_ gnd vdd FILL
XFILL_0__16115_ gnd vdd FILL
XFILL_1__15666_ gnd vdd FILL
XFILL_3__7884_ gnd vdd FILL
XFILL_0__10539_ gnd vdd FILL
XFILL_6__16406_ gnd vdd FILL
XFILL_5_BUFX2_insert517 gnd vdd FILL
XFILL_3__11699_ gnd vdd FILL
XFILL_6__13618_ gnd vdd FILL
XFILL_5_BUFX2_insert528 gnd vdd FILL
XFILL_0__9914_ gnd vdd FILL
XFILL_1__12878_ gnd vdd FILL
XFILL_3__16226_ gnd vdd FILL
XFILL_5_BUFX2_insert539 gnd vdd FILL
XFILL_5__15047_ gnd vdd FILL
XFILL_5__12259_ gnd vdd FILL
X_8453_ _8453_/A gnd _8455_/A vdd INVX1
XFILL_3__9623_ gnd vdd FILL
XFILL_3__13438_ gnd vdd FILL
XFILL_1__14617_ gnd vdd FILL
XFILL_0__16046_ gnd vdd FILL
XFILL_2__12079_ gnd vdd FILL
XFILL_4__12989_ gnd vdd FILL
XFILL_4__15777_ gnd vdd FILL
XFILL_0__13258_ gnd vdd FILL
XFILL_1__11829_ gnd vdd FILL
X_7404_ _7404_/Q _7916_/CLK _9580_/R vdd _7354_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert9 gnd vdd FILL
XFILL_1__15597_ gnd vdd FILL
XFILL_0_BUFX2_insert890 gnd vdd FILL
XFILL_2__15907_ gnd vdd FILL
X_8384_ _8384_/A _8321_/B _8384_/C gnd _8384_/Y vdd OAI21X1
XFILL_4__14728_ gnd vdd FILL
XFILL_3__16157_ gnd vdd FILL
XFILL_3__13369_ gnd vdd FILL
XFILL_0__12209_ gnd vdd FILL
XFILL_3__9554_ gnd vdd FILL
XSFILL109000x70050 gnd vdd FILL
XFILL_1__14548_ gnd vdd FILL
X_7335_ _7297_/B _9383_/B gnd _7336_/C vdd NAND2X1
XFILL_6__16268_ gnd vdd FILL
XFILL_3__15108_ gnd vdd FILL
XFILL_3__8505_ gnd vdd FILL
XFILL_3_BUFX2_insert50 gnd vdd FILL
XFILL_0__9776_ gnd vdd FILL
XFILL_0__6988_ gnd vdd FILL
XFILL_3_BUFX2_insert61 gnd vdd FILL
XFILL_3__16088_ gnd vdd FILL
XFILL_2__15838_ gnd vdd FILL
XFILL_4__14659_ gnd vdd FILL
XFILL_3__9485_ gnd vdd FILL
XFILL_3_BUFX2_insert72 gnd vdd FILL
XFILL_1__14479_ gnd vdd FILL
XFILL_6__15219_ gnd vdd FILL
XFILL_3_BUFX2_insert83 gnd vdd FILL
XFILL_0__8727_ gnd vdd FILL
XFILL_3__15039_ gnd vdd FILL
XFILL_5__15949_ gnd vdd FILL
X_7266_ _7194_/A _7778_/CLK _8424_/R vdd _7266_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert94 gnd vdd FILL
XFILL_1__16218_ gnd vdd FILL
XFILL_2__15769_ gnd vdd FILL
XSFILL43960x50050 gnd vdd FILL
X_9005_ _9005_/A _9005_/B gnd _9006_/C vdd NAND2X1
XFILL_1__7451_ gnd vdd FILL
XFILL_4__16329_ gnd vdd FILL
XFILL_0__8658_ gnd vdd FILL
X_7197_ _7197_/A gnd _7197_/Y vdd INVX1
XFILL_4__7160_ gnd vdd FILL
XFILL_1__16149_ gnd vdd FILL
XFILL_3__8367_ gnd vdd FILL
XFILL_0__7609_ gnd vdd FILL
XFILL_0__8589_ gnd vdd FILL
XSFILL99560x2050 gnd vdd FILL
XFILL_3__7318_ gnd vdd FILL
XFILL_2_BUFX2_insert407 gnd vdd FILL
XFILL_4__7091_ gnd vdd FILL
XFILL_1__9121_ gnd vdd FILL
XFILL_2_BUFX2_insert418 gnd vdd FILL
XFILL_2_BUFX2_insert429 gnd vdd FILL
XFILL_3__7249_ gnd vdd FILL
X_9907_ _9896_/B _9907_/B gnd _9907_/Y vdd NAND2X1
XFILL112040x25050 gnd vdd FILL
XFILL_1__8003_ gnd vdd FILL
X_9838_ _9838_/Q _8942_/CLK _8942_/R vdd _9838_/D gnd vdd DFFSR
XFILL_4__9801_ gnd vdd FILL
XFILL_4__7993_ gnd vdd FILL
X_10720_ _10720_/Q _9834_/CLK _7793_/R vdd _10646_/Y gnd vdd DFFSR
XFILL_4__9732_ gnd vdd FILL
X_9769_ _9831_/Q gnd _9771_/A vdd INVX1
XBUFX2_insert406 _10920_/Y gnd _12371_/A vdd BUFX2
XFILL_4__6944_ gnd vdd FILL
XFILL_6_BUFX2_insert362 gnd vdd FILL
XBUFX2_insert417 _15050_/Y gnd _15172_/A vdd BUFX2
XBUFX2_insert428 _15047_/Y gnd _15972_/C vdd BUFX2
X_10651_ _10615_/B _7451_/B gnd _10652_/C vdd NAND2X1
XBUFX2_insert439 _15086_/Y gnd _15662_/A vdd BUFX2
XFILL_4__9663_ gnd vdd FILL
XFILL_4__6875_ gnd vdd FILL
X_10582_ _10486_/A _6998_/CLK _7644_/R vdd _10582_/D gnd vdd DFFSR
X_13370_ _14456_/C gnd _13370_/Y vdd INVX8
XFILL_1__8905_ gnd vdd FILL
XFILL_4__8614_ gnd vdd FILL
XFILL_1__9885_ gnd vdd FILL
X_12321_ _6896_/A _12301_/B _12301_/C _12313_/D gnd _12322_/C vdd AOI22X1
XFILL_4__9594_ gnd vdd FILL
XFILL_1__8836_ gnd vdd FILL
X_15040_ _15715_/C _15036_/A _15920_/B gnd _15040_/Y vdd OAI21X1
X_12252_ _12248_/A _12800_/Q _12248_/C gnd _12254_/B vdd NAND3X1
XFILL_1__8767_ gnd vdd FILL
XFILL_2__7560_ gnd vdd FILL
XSFILL33960x82050 gnd vdd FILL
XFILL_4__8476_ gnd vdd FILL
X_11203_ _12201_/Y _12330_/Y gnd _11203_/Y vdd NOR2X1
X_12183_ _12183_/A _12201_/B _12183_/C gnd _12183_/Y vdd OAI21X1
XFILL_1__7718_ gnd vdd FILL
XFILL_4__7427_ gnd vdd FILL
XFILL_2__7491_ gnd vdd FILL
XFILL_1__8698_ gnd vdd FILL
X_11134_ _12165_/Y _12282_/Y gnd _11634_/A vdd NAND2X1
XFILL_2__9230_ gnd vdd FILL
XFILL_3_BUFX2_insert230 gnd vdd FILL
XSFILL49640x70050 gnd vdd FILL
XFILL_4__7358_ gnd vdd FILL
XFILL_3_BUFX2_insert241 gnd vdd FILL
XFILL_3_BUFX2_insert252 gnd vdd FILL
X_15942_ _15939_/Y _15941_/Y _15942_/C gnd _15943_/B vdd NAND3X1
X_11065_ _11063_/Y _11064_/Y gnd _11065_/Y vdd NOR2X1
XFILL_3_BUFX2_insert263 gnd vdd FILL
XFILL_2__9161_ gnd vdd FILL
XFILL_3_BUFX2_insert274 gnd vdd FILL
XFILL_1__10160_ gnd vdd FILL
X_10016_ _10016_/A gnd _10018_/A vdd INVX1
XFILL_3_BUFX2_insert285 gnd vdd FILL
XFILL_3_BUFX2_insert296 gnd vdd FILL
XFILL_0__10890_ gnd vdd FILL
XFILL_5__11630_ gnd vdd FILL
XFILL_4__7289_ gnd vdd FILL
XFILL_2__8112_ gnd vdd FILL
X_15873_ _14407_/D _15595_/B _15873_/C gnd _15876_/A vdd OAI21X1
XFILL_4__10271_ gnd vdd FILL
XFILL_2__11450_ gnd vdd FILL
XFILL_2__9092_ gnd vdd FILL
XFILL_4__9028_ gnd vdd FILL
XFILL_2_BUFX2_insert930 gnd vdd FILL
XFILL_5__9910_ gnd vdd FILL
X_14824_ _7282_/Q _13619_/B _14214_/C _10098_/Q gnd _14824_/Y vdd AOI22X1
XFILL_4__12010_ gnd vdd FILL
XFILL_2_BUFX2_insert941 gnd vdd FILL
XFILL_5__11561_ gnd vdd FILL
XFILL_2_BUFX2_insert952 gnd vdd FILL
XSFILL28920x71050 gnd vdd FILL
XFILL_3__12740_ gnd vdd FILL
XFILL_2_BUFX2_insert963 gnd vdd FILL
XFILL_2__10401_ gnd vdd FILL
XFILL_2_BUFX2_insert974 gnd vdd FILL
XFILL_2__11381_ gnd vdd FILL
XFILL_2_BUFX2_insert985 gnd vdd FILL
XFILL_5__13300_ gnd vdd FILL
XFILL_5__10512_ gnd vdd FILL
XFILL_2_BUFX2_insert996 gnd vdd FILL
X_14755_ _9841_/Q gnd _14757_/A vdd INVX1
XFILL_5__14280_ gnd vdd FILL
X_11967_ _11967_/A _11955_/B _11967_/C gnd _6864_/A vdd OAI21X1
XFILL_2__13120_ gnd vdd FILL
XFILL_5__11492_ gnd vdd FILL
XFILL_0__11511_ gnd vdd FILL
XFILL_1__13850_ gnd vdd FILL
XFILL_5__9772_ gnd vdd FILL
XFILL_5__13231_ gnd vdd FILL
XSFILL8840x69050 gnd vdd FILL
XFILL_0__12491_ gnd vdd FILL
X_13706_ _9477_/A gnd _13708_/D vdd INVX1
XFILL_5__10443_ gnd vdd FILL
X_10918_ _10911_/A _10984_/Q gnd _10924_/A vdd NAND2X1
XFILL_3__14410_ gnd vdd FILL
XFILL_5__6984_ gnd vdd FILL
X_14686_ _14030_/A _16083_/C _14949_/C _14686_/D gnd _14687_/B vdd OAI22X1
XFILL_3__11622_ gnd vdd FILL
XFILL_4__13961_ gnd vdd FILL
XFILL_3__15390_ gnd vdd FILL
XFILL_0__14230_ gnd vdd FILL
X_11898_ _11896_/Y _11975_/A _11897_/Y gnd _6841_/A vdd OAI21X1
XFILL_2__10263_ gnd vdd FILL
XFILL_2__9994_ gnd vdd FILL
XFILL_5__8723_ gnd vdd FILL
XFILL_0__11442_ gnd vdd FILL
X_16425_ _16425_/Q _7406_/CLK _9692_/R vdd _16425_/D gnd vdd DFFSR
XSFILL99480x57050 gnd vdd FILL
XFILL_1__13781_ gnd vdd FILL
XFILL_1__10993_ gnd vdd FILL
X_13637_ _13637_/A _13637_/B _14265_/C gnd _12961_/B vdd AOI21X1
XFILL_4__15700_ gnd vdd FILL
XFILL_5__13162_ gnd vdd FILL
XFILL_4__12912_ gnd vdd FILL
XFILL_2__12002_ gnd vdd FILL
XSFILL74120x55050 gnd vdd FILL
X_10849_ _15509_/A _9953_/CLK _9580_/R vdd _10777_/Y gnd vdd DFFSR
XFILL_3__14341_ gnd vdd FILL
XFILL_5__10374_ gnd vdd FILL
XFILL_1__15520_ gnd vdd FILL
XFILL_4__13892_ gnd vdd FILL
XFILL_3__11553_ gnd vdd FILL
XFILL_1__12732_ gnd vdd FILL
XFILL_0__14161_ gnd vdd FILL
XFILL_2__10194_ gnd vdd FILL
XFILL_5__8654_ gnd vdd FILL
XFILL_5__12113_ gnd vdd FILL
XBUFX2_insert940 _12426_/Y gnd _7496_/B vdd BUFX2
XFILL_0__11373_ gnd vdd FILL
XFILL_6__14452_ gnd vdd FILL
XBUFX2_insert951 _13365_/Y gnd _10762_/B vdd BUFX2
X_16356_ _16356_/A gnd _16356_/C gnd _16428_/D vdd OAI21X1
XBUFX2_insert962 _13361_/Y gnd _10423_/B vdd BUFX2
XFILL_3__10504_ gnd vdd FILL
XFILL_4__15631_ gnd vdd FILL
XFILL_4__12843_ gnd vdd FILL
XFILL_0__7960_ gnd vdd FILL
XFILL_5__13093_ gnd vdd FILL
X_13568_ _14868_/A _15130_/B _13568_/C _14956_/D gnd _13571_/A vdd AOI22X1
XBUFX2_insert973 _16451_/Y gnd _13134_/A vdd BUFX2
XFILL_0__13112_ gnd vdd FILL
XFILL_3__14272_ gnd vdd FILL
XFILL_5__7605_ gnd vdd FILL
XFILL_2__8876_ gnd vdd FILL
XFILL_1__15451_ gnd vdd FILL
XFILL_3__11484_ gnd vdd FILL
XFILL_0__10324_ gnd vdd FILL
X_15307_ _13773_/Y _15386_/B _15386_/C _15307_/D gnd _15307_/Y vdd OAI22X1
XFILL_6__13403_ gnd vdd FILL
XFILL_0__14092_ gnd vdd FILL
XBUFX2_insert984 _13351_/Y gnd _10066_/B vdd BUFX2
XFILL_0__6911_ gnd vdd FILL
XBUFX2_insert995 _12408_/Y gnd _7990_/B vdd BUFX2
XFILL_5__8585_ gnd vdd FILL
XFILL_3__16011_ gnd vdd FILL
X_12519_ _12519_/A vdd _12518_/Y gnd _12519_/Y vdd OAI21X1
XFILL_5__12044_ gnd vdd FILL
XSFILL53960x13050 gnd vdd FILL
XFILL_3__13223_ gnd vdd FILL
X_16287_ _7925_/Q _16204_/B gnd _16287_/Y vdd NAND2X1
XFILL_4__12774_ gnd vdd FILL
XFILL_4__15562_ gnd vdd FILL
XFILL_0__7891_ gnd vdd FILL
XFILL_1__14402_ gnd vdd FILL
XFILL_3__10435_ gnd vdd FILL
XFILL_2__7827_ gnd vdd FILL
X_13499_ _9465_/A gnd _13499_/Y vdd INVX1
XSFILL109480x42050 gnd vdd FILL
XFILL_2__13953_ gnd vdd FILL
XFILL_1__11614_ gnd vdd FILL
XFILL_0__13043_ gnd vdd FILL
XFILL_0__10255_ gnd vdd FILL
XFILL_1__15382_ gnd vdd FILL
XFILL_1__12594_ gnd vdd FILL
X_15238_ _13682_/B gnd _15238_/Y vdd INVX1
XFILL_0__9630_ gnd vdd FILL
XFILL_4__14513_ gnd vdd FILL
XFILL_0__6842_ gnd vdd FILL
XFILL_4__11725_ gnd vdd FILL
XFILL112280x81050 gnd vdd FILL
XFILL_3__13154_ gnd vdd FILL
XFILL_2__12904_ gnd vdd FILL
XFILL_4__15493_ gnd vdd FILL
XFILL_2__7758_ gnd vdd FILL
XFILL_1__14333_ gnd vdd FILL
XFILL_1__11545_ gnd vdd FILL
XFILL_3__10366_ gnd vdd FILL
XSFILL54040x22050 gnd vdd FILL
XFILL_2__13884_ gnd vdd FILL
XFILL_0__10186_ gnd vdd FILL
XFILL_5__15803_ gnd vdd FILL
XFILL_5__7467_ gnd vdd FILL
XFILL_6__16053_ gnd vdd FILL
X_7120_ _7156_/Q gnd _7122_/A vdd INVX1
XFILL_6__13265_ gnd vdd FILL
X_15169_ _15169_/A _13623_/Y _15169_/C _15169_/D gnd _15169_/Y vdd OAI22X1
XFILL_3__12105_ gnd vdd FILL
XFILL_4__14444_ gnd vdd FILL
XFILL_2__15623_ gnd vdd FILL
XFILL_4__11656_ gnd vdd FILL
XFILL_3__9270_ gnd vdd FILL
XFILL_2__12835_ gnd vdd FILL
XFILL_3__13085_ gnd vdd FILL
XFILL_5__9206_ gnd vdd FILL
XFILL_5__13995_ gnd vdd FILL
XFILL_2__7689_ gnd vdd FILL
XFILL_1__14264_ gnd vdd FILL
XFILL_3__10297_ gnd vdd FILL
XFILL_1__11476_ gnd vdd FILL
XFILL_6__15004_ gnd vdd FILL
XFILL_0__8512_ gnd vdd FILL
X_7051_ _7133_/Q gnd _7051_/Y vdd INVX1
XFILL_0__14994_ gnd vdd FILL
XFILL_5__15734_ gnd vdd FILL
XFILL_1__16003_ gnd vdd FILL
XFILL_3__12036_ gnd vdd FILL
XFILL_2__9428_ gnd vdd FILL
XFILL_4__14375_ gnd vdd FILL
XFILL_0__9492_ gnd vdd FILL
XFILL_3__8221_ gnd vdd FILL
XFILL_1__13215_ gnd vdd FILL
XFILL_1__10427_ gnd vdd FILL
XFILL_2__15554_ gnd vdd FILL
XFILL_4__11587_ gnd vdd FILL
XFILL_2__12766_ gnd vdd FILL
XFILL_1__14195_ gnd vdd FILL
XFILL_5__9137_ gnd vdd FILL
XFILL_0__13945_ gnd vdd FILL
XFILL_4__13326_ gnd vdd FILL
XFILL_4__16114_ gnd vdd FILL
XFILL_6__12147_ gnd vdd FILL
XFILL_0__8443_ gnd vdd FILL
XFILL_5__15665_ gnd vdd FILL
XFILL_2__14505_ gnd vdd FILL
XFILL_4__10538_ gnd vdd FILL
XFILL_2__9359_ gnd vdd FILL
XFILL_1__13146_ gnd vdd FILL
XSFILL18680x41050 gnd vdd FILL
XFILL_5__12877_ gnd vdd FILL
XFILL_2__11717_ gnd vdd FILL
XFILL_1__10358_ gnd vdd FILL
XFILL_2__15485_ gnd vdd FILL
XFILL_2__12697_ gnd vdd FILL
XSFILL74200x35050 gnd vdd FILL
XFILL_0__13876_ gnd vdd FILL
XFILL_4__16045_ gnd vdd FILL
XFILL_5__14616_ gnd vdd FILL
XFILL_4__13257_ gnd vdd FILL
XFILL_0__8374_ gnd vdd FILL
XFILL_3__7103_ gnd vdd FILL
XFILL_5__11828_ gnd vdd FILL
XFILL_5__15596_ gnd vdd FILL
XFILL_2__14436_ gnd vdd FILL
XFILL_0__15615_ gnd vdd FILL
XFILL_3__13987_ gnd vdd FILL
XFILL_5__8019_ gnd vdd FILL
XFILL_2__11648_ gnd vdd FILL
XFILL_3__8083_ gnd vdd FILL
XFILL_1__10289_ gnd vdd FILL
XFILL_0__12827_ gnd vdd FILL
XFILL_6__9881_ gnd vdd FILL
XFILL_4__12208_ gnd vdd FILL
XSFILL49000x11050 gnd vdd FILL
XFILL_0__7325_ gnd vdd FILL
XFILL_5__14547_ gnd vdd FILL
XFILL_3__15726_ gnd vdd FILL
XFILL_1__12028_ gnd vdd FILL
XFILL_3__7034_ gnd vdd FILL
X_7953_ _7953_/A gnd _7955_/A vdd INVX1
XFILL_5__11759_ gnd vdd FILL
XFILL_2__14367_ gnd vdd FILL
XFILL112440x5050 gnd vdd FILL
XFILL_0__12758_ gnd vdd FILL
XFILL_0__15546_ gnd vdd FILL
XFILL_2__11579_ gnd vdd FILL
XFILL_6__8832_ gnd vdd FILL
XFILL_4__12139_ gnd vdd FILL
X_6904_ _6902_/Y _6948_/A _6904_/C gnd _6998_/D vdd OAI21X1
XFILL_2__16106_ gnd vdd FILL
XFILL_5__14478_ gnd vdd FILL
XFILL_2__13318_ gnd vdd FILL
XFILL_3__15657_ gnd vdd FILL
X_7884_ _7882_/Y _7824_/B _7884_/C gnd _7922_/D vdd OAI21X1
XFILL_3__12869_ gnd vdd FILL
XFILL_0__11709_ gnd vdd FILL
XFILL_2__14298_ gnd vdd FILL
XFILL_5__16217_ gnd vdd FILL
XFILL112360x61050 gnd vdd FILL
XFILL_0__15477_ gnd vdd FILL
XFILL_3__14608_ gnd vdd FILL
X_9623_ _9623_/A gnd _9623_/Y vdd INVX1
XFILL_5__13429_ gnd vdd FILL
XFILL_0__7187_ gnd vdd FILL
XFILL_2__16037_ gnd vdd FILL
XFILL_2__13249_ gnd vdd FILL
XFILL_3__15588_ gnd vdd FILL
XFILL_3__8985_ gnd vdd FILL
XSFILL74120x7050 gnd vdd FILL
XFILL_0__14428_ gnd vdd FILL
XFILL_1__13979_ gnd vdd FILL
XFILL_5__16148_ gnd vdd FILL
XFILL_3__14539_ gnd vdd FILL
X_9554_ _9554_/A _9554_/B _9553_/Y gnd _9588_/D vdd OAI21X1
XFILL_3__7936_ gnd vdd FILL
XFILL_1__15718_ gnd vdd FILL
XFILL_5_BUFX2_insert303 gnd vdd FILL
XFILL_0__14359_ gnd vdd FILL
XSFILL43960x45050 gnd vdd FILL
XFILL_5_BUFX2_insert314 gnd vdd FILL
X_8505_ _8503_/B _8377_/B gnd _8506_/C vdd NAND2X1
XFILL_1__6951_ gnd vdd FILL
XBUFX2_insert15 _14989_/Y gnd _15386_/C vdd BUFX2
XFILL_4__15829_ gnd vdd FILL
XFILL_5__16079_ gnd vdd FILL
XFILL_5_BUFX2_insert325 gnd vdd FILL
X_9485_ _9485_/A _9551_/B _9484_/Y gnd _9485_/Y vdd OAI21X1
XFILL_5_BUFX2_insert336 gnd vdd FILL
XFILL_3__7867_ gnd vdd FILL
XBUFX2_insert26 _13320_/Y gnd _8508_/A vdd BUFX2
XFILL_1__15649_ gnd vdd FILL
XFILL_5_BUFX2_insert347 gnd vdd FILL
XFILL_5_BUFX2_insert358 gnd vdd FILL
XBUFX2_insert37 _13265_/Y gnd _6982_/B vdd BUFX2
XFILL_3__16209_ gnd vdd FILL
XBUFX2_insert48 _13381_/Y gnd _14583_/B vdd BUFX2
XFILL_5_BUFX2_insert369 gnd vdd FILL
XSFILL18760x21050 gnd vdd FILL
XBUFX2_insert59 _14983_/Y gnd _15180_/C vdd BUFX2
XFILL_1__9670_ gnd vdd FILL
XFILL_3__9606_ gnd vdd FILL
X_8436_ _8436_/Q _9194_/CLK _7914_/R vdd _8436_/D gnd vdd DFFSR
XFILL_1__6882_ gnd vdd FILL
XFILL_0__16029_ gnd vdd FILL
XFILL_3__7798_ gnd vdd FILL
XFILL_1__8621_ gnd vdd FILL
X_8367_ _8367_/A gnd _8369_/A vdd INVX1
XFILL_4__8330_ gnd vdd FILL
XFILL_3__9537_ gnd vdd FILL
XSFILL54040x50 gnd vdd FILL
X_7318_ _7318_/A _7354_/B _7317_/Y gnd _7392_/D vdd OAI21X1
XFILL_0__9759_ gnd vdd FILL
XSFILL23880x12050 gnd vdd FILL
X_8298_ _8242_/A _9578_/CLK _9460_/R vdd _8244_/Y gnd vdd DFFSR
XFILL_4__8261_ gnd vdd FILL
XFILL_3__9468_ gnd vdd FILL
XFILL111800x75050 gnd vdd FILL
XFILL_1__7503_ gnd vdd FILL
X_7249_ _7250_/B _7889_/B gnd _7249_/Y vdd NAND2X1
XFILL_1__8483_ gnd vdd FILL
XFILL_4__7212_ gnd vdd FILL
XSFILL38920x34050 gnd vdd FILL
XFILL112440x41050 gnd vdd FILL
XFILL_4__8192_ gnd vdd FILL
XFILL_6__8128_ gnd vdd FILL
XSFILL64200x67050 gnd vdd FILL
XFILL_3__9399_ gnd vdd FILL
XFILL_1__7434_ gnd vdd FILL
XSFILL27960x58050 gnd vdd FILL
XFILL_1__7365_ gnd vdd FILL
XFILL_2_BUFX2_insert226 gnd vdd FILL
XFILL_4__7074_ gnd vdd FILL
XFILL_2_BUFX2_insert237 gnd vdd FILL
XSFILL3640x74050 gnd vdd FILL
XFILL_1__9104_ gnd vdd FILL
XFILL_2_BUFX2_insert248 gnd vdd FILL
XSFILL95000x1050 gnd vdd FILL
X_12870_ _12868_/Y vdd _12870_/C gnd _12934_/D vdd OAI21X1
XFILL_2_BUFX2_insert259 gnd vdd FILL
XSFILL3720x2050 gnd vdd FILL
XSFILL84120x18050 gnd vdd FILL
XFILL_1__7296_ gnd vdd FILL
XSFILL94280x62050 gnd vdd FILL
X_11821_ _12222_/Y _11007_/Y _11839_/A gnd _11821_/Y vdd OAI21X1
XFILL_1_BUFX2_insert904 gnd vdd FILL
XFILL_1__9035_ gnd vdd FILL
XSFILL68440x72050 gnd vdd FILL
XFILL_1_BUFX2_insert915 gnd vdd FILL
XFILL_1_BUFX2_insert926 gnd vdd FILL
XFILL_1_BUFX2_insert937 gnd vdd FILL
X_14540_ _8632_/A gnd _14540_/Y vdd INVX1
XFILL_1_BUFX2_insert948 gnd vdd FILL
X_11752_ _11750_/Y _11752_/B _11752_/C gnd _11753_/A vdd OAI21X1
XFILL_1_BUFX2_insert959 gnd vdd FILL
XFILL_4__7976_ gnd vdd FILL
X_10703_ _10701_/Y _10678_/A _10703_/C gnd _10739_/D vdd OAI21X1
XSFILL33960x77050 gnd vdd FILL
X_14471_ _10475_/Q _14389_/B _14867_/C _9963_/Q gnd _14472_/B vdd AOI22X1
X_11683_ _11680_/Y _11683_/B gnd _11683_/Y vdd NOR2X1
XBUFX2_insert225 _12432_/Y gnd _8910_/B vdd BUFX2
XFILL_2__6991_ gnd vdd FILL
XFILL_4__6927_ gnd vdd FILL
X_16210_ _16210_/A _16210_/B _16210_/C gnd _16220_/B vdd NAND3X1
XBUFX2_insert236 _12348_/Y gnd _9082_/B vdd BUFX2
X_13422_ _8150_/Q gnd _13422_/Y vdd INVX1
XBUFX2_insert247 _10922_/Y gnd _15651_/C vdd BUFX2
X_10634_ _10632_/Y _10700_/B _10634_/C gnd _10634_/Y vdd OAI21X1
XFILL_2__8730_ gnd vdd FILL
XBUFX2_insert258 _12423_/Y gnd _8005_/B vdd BUFX2
XFILL_1__9937_ gnd vdd FILL
XBUFX2_insert269 _13364_/Y gnd _10676_/B vdd BUFX2
XFILL_4__9646_ gnd vdd FILL
XFILL_4__6858_ gnd vdd FILL
X_16141_ _16141_/A _14778_/A _16141_/C gnd _16141_/Y vdd NOR3X1
XFILL_5_CLKBUF1_insert115 gnd vdd FILL
X_13353_ _13246_/A _13337_/B _13359_/A gnd _13354_/A vdd NAND3X1
XFILL_5_CLKBUF1_insert126 gnd vdd FILL
X_10565_ _10500_/B _6981_/B gnd _10566_/C vdd NAND2X1
XFILL_5_CLKBUF1_insert137 gnd vdd FILL
XFILL_1__9868_ gnd vdd FILL
XSFILL89240x51050 gnd vdd FILL
XSFILL18760x2050 gnd vdd FILL
XFILL_2__8661_ gnd vdd FILL
XFILL_5_BUFX2_insert870 gnd vdd FILL
XFILL_5_CLKBUF1_insert148 gnd vdd FILL
XFILL_5_BUFX2_insert881 gnd vdd FILL
X_12304_ _12312_/A _12340_/B _12312_/C gnd _12306_/B vdd NAND3X1
XFILL_5_CLKBUF1_insert159 gnd vdd FILL
XFILL_5__8370_ gnd vdd FILL
XFILL_5_BUFX2_insert892 gnd vdd FILL
X_16072_ _16072_/A gnd _16072_/Y vdd INVX1
X_13284_ _13295_/A _13284_/B _13295_/C gnd _13284_/Y vdd OAI21X1
XFILL_2__7612_ gnd vdd FILL
X_10496_ _10511_/A _8576_/B gnd _10497_/C vdd NAND2X1
XFILL_2__8592_ gnd vdd FILL
XFILL_2__10950_ gnd vdd FILL
XFILL_5__7321_ gnd vdd FILL
XFILL_0__10040_ gnd vdd FILL
XFILL_4__8528_ gnd vdd FILL
XFILL_1__9799_ gnd vdd FILL
X_15023_ _14982_/Y _16232_/B gnd _15023_/Y vdd NAND2X1
XSFILL73960x50 gnd vdd FILL
X_12235_ _12255_/A gnd _12255_/C gnd _12238_/A vdd NAND3X1
XFILL_4__11510_ gnd vdd FILL
XFILL_3__10151_ gnd vdd FILL
XSFILL28920x66050 gnd vdd FILL
XFILL_2__7543_ gnd vdd FILL
XFILL_4__12490_ gnd vdd FILL
XFILL_1__11330_ gnd vdd FILL
XSFILL94360x42050 gnd vdd FILL
XFILL_4__8459_ gnd vdd FILL
XFILL_2__10881_ gnd vdd FILL
XFILL_5__7252_ gnd vdd FILL
X_12166_ _13192_/Q gnd _12168_/A vdd INVX1
XFILL_4__11441_ gnd vdd FILL
XFILL_2__12620_ gnd vdd FILL
XFILL_5__13780_ gnd vdd FILL
XFILL_5__10992_ gnd vdd FILL
XFILL_1__11261_ gnd vdd FILL
XFILL_2__7474_ gnd vdd FILL
XFILL_5__7183_ gnd vdd FILL
XFILL_0__11991_ gnd vdd FILL
X_11117_ _11116_/Y _11115_/Y gnd _11117_/Y vdd NOR2X1
XFILL_5__12731_ gnd vdd FILL
XFILL_1__13000_ gnd vdd FILL
XFILL_4__14160_ gnd vdd FILL
XFILL_2__9213_ gnd vdd FILL
XFILL_3__13910_ gnd vdd FILL
X_12097_ _12521_/B _12113_/B _12113_/C gnd gnd _12097_/Y vdd AOI22X1
XSFILL108520x8050 gnd vdd FILL
XFILL_4__11372_ gnd vdd FILL
XFILL_3__14890_ gnd vdd FILL
XFILL_0__10942_ gnd vdd FILL
XFILL_0__13730_ gnd vdd FILL
XFILL_1__11192_ gnd vdd FILL
XFILL_4__13111_ gnd vdd FILL
X_15925_ _15180_/C _14452_/Y _14451_/Y _15410_/D gnd _15926_/B vdd OAI22X1
X_11048_ _11048_/A _11640_/C gnd _11056_/A vdd NAND2X1
XFILL_5__15450_ gnd vdd FILL
XFILL_4__10323_ gnd vdd FILL
XFILL_5__12662_ gnd vdd FILL
XFILL_3__13841_ gnd vdd FILL
XFILL_2__9144_ gnd vdd FILL
XFILL_4__14091_ gnd vdd FILL
XFILL_2__11502_ gnd vdd FILL
XFILL_1__10143_ gnd vdd FILL
XFILL_2__15270_ gnd vdd FILL
XFILL_0__13661_ gnd vdd FILL
XFILL_2__12482_ gnd vdd FILL
XSFILL89720x29050 gnd vdd FILL
XFILL_0__10873_ gnd vdd FILL
XFILL_5__14401_ gnd vdd FILL
XFILL_5__11613_ gnd vdd FILL
X_15856_ _15856_/A _15856_/B gnd _15866_/B vdd NAND2X1
XFILL_4__13042_ gnd vdd FILL
XFILL_5__12593_ gnd vdd FILL
XFILL_4__10254_ gnd vdd FILL
XFILL_5__15381_ gnd vdd FILL
XFILL_2__14221_ gnd vdd FILL
XFILL_0__15400_ gnd vdd FILL
XFILL_0__12612_ gnd vdd FILL
XFILL_3__13772_ gnd vdd FILL
XFILL_2_BUFX2_insert760 gnd vdd FILL
XFILL_2__11433_ gnd vdd FILL
XFILL_1__14951_ gnd vdd FILL
XFILL_0__13592_ gnd vdd FILL
X_14807_ _10738_/Q gnd _14809_/B vdd INVX1
XFILL_2_BUFX2_insert771 gnd vdd FILL
XFILL_0__7110_ gnd vdd FILL
XFILL_6__12903_ gnd vdd FILL
XFILL_0__16380_ gnd vdd FILL
XFILL_0__8090_ gnd vdd FILL
XSFILL59080x70050 gnd vdd FILL
XFILL_3__15511_ gnd vdd FILL
XFILL_2_BUFX2_insert782 gnd vdd FILL
XFILL_5__14332_ gnd vdd FILL
XSFILL89320x31050 gnd vdd FILL
XFILL_5__11544_ gnd vdd FILL
XFILL_3__12723_ gnd vdd FILL
X_15787_ _15787_/A gnd _15787_/Y vdd INVX1
XFILL_2_BUFX2_insert793 gnd vdd FILL
XFILL_2__14152_ gnd vdd FILL
X_12999_ _6886_/A gnd _12999_/Y vdd INVX1
XFILL_4__10185_ gnd vdd FILL
XFILL_1__13902_ gnd vdd FILL
XFILL_0__15331_ gnd vdd FILL
XSFILL109480x37050 gnd vdd FILL
XFILL_2__11364_ gnd vdd FILL
XFILL_0__7041_ gnd vdd FILL
XFILL_1__14882_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1077 gnd vdd FILL
X_14738_ _14738_/A _7364_/A _7876_/A _13865_/B gnd _14738_/Y vdd AOI22X1
XFILL_5__14263_ gnd vdd FILL
XFILL_2__13103_ gnd vdd FILL
XFILL_5__11475_ gnd vdd FILL
XFILL_3__15442_ gnd vdd FILL
XFILL_3__12654_ gnd vdd FILL
XFILL_2__10315_ gnd vdd FILL
XFILL112280x76050 gnd vdd FILL
XFILL_1__13833_ gnd vdd FILL
XFILL_4__14993_ gnd vdd FILL
XFILL_2__11295_ gnd vdd FILL
XFILL_0__15262_ gnd vdd FILL
XFILL_2__14083_ gnd vdd FILL
XSFILL54040x17050 gnd vdd FILL
XFILL_5__16002_ gnd vdd FILL
XFILL_0__12474_ gnd vdd FILL
XFILL_5__13214_ gnd vdd FILL
XFILL_5__6967_ gnd vdd FILL
XFILL_5__9755_ gnd vdd FILL
XFILL_5__10426_ gnd vdd FILL
XFILL_5__14194_ gnd vdd FILL
XFILL_3__11605_ gnd vdd FILL
X_14669_ _16076_/A _14344_/B _14290_/C _7663_/Q gnd _14680_/A vdd AOI22X1
XSFILL94440x22050 gnd vdd FILL
XFILL_0__14213_ gnd vdd FILL
XFILL_3__15373_ gnd vdd FILL
XFILL_2__13034_ gnd vdd FILL
XFILL_2__10246_ gnd vdd FILL
XFILL_4__13944_ gnd vdd FILL
XFILL_3__12585_ gnd vdd FILL
XFILL_3__8770_ gnd vdd FILL
XFILL_2__9977_ gnd vdd FILL
XFILL_0__11425_ gnd vdd FILL
XFILL_0__15193_ gnd vdd FILL
X_16408_ _16408_/A gnd _16410_/A vdd INVX1
XFILL_5__8706_ gnd vdd FILL
XFILL_1__13764_ gnd vdd FILL
XFILL_1__10976_ gnd vdd FILL
XFILL_5__13145_ gnd vdd FILL
XFILL_5__6898_ gnd vdd FILL
XFILL_3__14324_ gnd vdd FILL
XFILL_0__8992_ gnd vdd FILL
XFILL_1__15503_ gnd vdd FILL
XFILL_3__11536_ gnd vdd FILL
XFILL_3__7721_ gnd vdd FILL
XFILL_1__12715_ gnd vdd FILL
XFILL_4__13875_ gnd vdd FILL
XFILL_0__14144_ gnd vdd FILL
XFILL_2__10177_ gnd vdd FILL
XFILL_5__8637_ gnd vdd FILL
XFILL_0__11356_ gnd vdd FILL
XBUFX2_insert770 _13301_/Y gnd _7878_/B vdd BUFX2
X_16339_ _16339_/A gnd _16341_/A vdd INVX1
XFILL_1__13695_ gnd vdd FILL
XBUFX2_insert781 _10911_/Y gnd _12123_/B vdd BUFX2
X_9270_ _9228_/A _7222_/B gnd _9270_/Y vdd NAND2X1
XFILL_4__15614_ gnd vdd FILL
XBUFX2_insert792 _15052_/Y gnd _15321_/C vdd BUFX2
XFILL_0__7943_ gnd vdd FILL
XFILL_3__14255_ gnd vdd FILL
XFILL_5__10288_ gnd vdd FILL
XFILL_4__12826_ gnd vdd FILL
XFILL_2__8859_ gnd vdd FILL
XSFILL18680x36050 gnd vdd FILL
XFILL_0__10307_ gnd vdd FILL
XFILL_1__15434_ gnd vdd FILL
XFILL_3__11467_ gnd vdd FILL
XFILL_1__12646_ gnd vdd FILL
XFILL_2__14985_ gnd vdd FILL
XFILL_0__14075_ gnd vdd FILL
XFILL_5__8568_ gnd vdd FILL
XFILL_5__12027_ gnd vdd FILL
XFILL_0__11287_ gnd vdd FILL
X_8221_ _8221_/A gnd _8223_/A vdd INVX1
XFILL_4__12757_ gnd vdd FILL
XFILL_4__15545_ gnd vdd FILL
XFILL_3__10418_ gnd vdd FILL
XFILL_0__7874_ gnd vdd FILL
XFILL_6__9100_ gnd vdd FILL
XSFILL84360x74050 gnd vdd FILL
XFILL_3__14186_ gnd vdd FILL
XFILL_0__13026_ gnd vdd FILL
XFILL_2__13936_ gnd vdd FILL
XFILL_1__15365_ gnd vdd FILL
XFILL_3__7583_ gnd vdd FILL
XFILL_3__11398_ gnd vdd FILL
XFILL_0__10238_ gnd vdd FILL
XFILL_1__12577_ gnd vdd FILL
XFILL_0__9613_ gnd vdd FILL
X_8152_ _8152_/Q _8152_/CLK _8664_/R vdd _8152_/D gnd vdd DFFSR
XFILL_4__11708_ gnd vdd FILL
XFILL_5__8499_ gnd vdd FILL
XFILL_3__13137_ gnd vdd FILL
XFILL_1__14316_ gnd vdd FILL
XFILL_4__15476_ gnd vdd FILL
XFILL_2__13867_ gnd vdd FILL
XSFILL59160x50050 gnd vdd FILL
XFILL_1__11528_ gnd vdd FILL
X_7103_ _7055_/A _8255_/B gnd _7104_/C vdd NAND2X1
XFILL_0__10169_ gnd vdd FILL
XFILL_1__15296_ gnd vdd FILL
XFILL_0__9544_ gnd vdd FILL
X_8083_ _8081_/Y _8082_/A _8083_/C gnd _8159_/D vdd OAI21X1
XFILL_4__11639_ gnd vdd FILL
XFILL_2__15606_ gnd vdd FILL
XFILL_4__14427_ gnd vdd FILL
XSFILL109560x17050 gnd vdd FILL
XFILL_3__9253_ gnd vdd FILL
XFILL_5__13978_ gnd vdd FILL
XFILL_1__14247_ gnd vdd FILL
XFILL_1__11459_ gnd vdd FILL
XFILL_2__13798_ gnd vdd FILL
XSFILL38840x49050 gnd vdd FILL
XFILL_5__15717_ gnd vdd FILL
XFILL_0__14977_ gnd vdd FILL
X_7034_ _7061_/A _6906_/B gnd _7034_/Y vdd NAND2X1
XFILL_0__9475_ gnd vdd FILL
XFILL_3__8204_ gnd vdd FILL
XFILL112360x56050 gnd vdd FILL
XFILL_3__12019_ gnd vdd FILL
XFILL_4__14358_ gnd vdd FILL
XFILL_2__15537_ gnd vdd FILL
XFILL_2__12749_ gnd vdd FILL
XFILL_1__14178_ gnd vdd FILL
XFILL_0__13928_ gnd vdd FILL
XFILL_4__13309_ gnd vdd FILL
XFILL_5__15648_ gnd vdd FILL
XFILL_3__8135_ gnd vdd FILL
XFILL_4__14289_ gnd vdd FILL
XFILL_1__13129_ gnd vdd FILL
XFILL_2__15468_ gnd vdd FILL
XFILL_0__13859_ gnd vdd FILL
XSFILL79320x63050 gnd vdd FILL
XFILL_0__8357_ gnd vdd FILL
XFILL_4__16028_ gnd vdd FILL
XFILL_2__14419_ gnd vdd FILL
XFILL_5__15579_ gnd vdd FILL
XFILL_3__8066_ gnd vdd FILL
X_8985_ _8983_/Y _8969_/A _8985_/C gnd _8985_/Y vdd OAI21X1
XFILL_2__15399_ gnd vdd FILL
XFILL_0__7308_ gnd vdd FILL
XSFILL18760x16050 gnd vdd FILL
XFILL_1__7081_ gnd vdd FILL
X_7936_ _7937_/B _8576_/B gnd _7936_/Y vdd NAND2X1
XFILL_3__15709_ gnd vdd FILL
XSFILL114520x72050 gnd vdd FILL
XSFILL44040x49050 gnd vdd FILL
XFILL_0__15529_ gnd vdd FILL
XFILL_0__7239_ gnd vdd FILL
X_7867_ _7917_/Q gnd _7867_/Y vdd INVX1
XFILL_4__7830_ gnd vdd FILL
X_9606_ _9597_/A _9478_/B gnd _9607_/C vdd NAND2X1
XSFILL18600x80050 gnd vdd FILL
XFILL_3__8968_ gnd vdd FILL
X_7798_ _7894_/Q gnd _7798_/Y vdd INVX1
XFILL_4__7761_ gnd vdd FILL
XFILL_5_BUFX2_insert100 gnd vdd FILL
XFILL_4__9500_ gnd vdd FILL
X_9537_ _9583_/Q gnd _9537_/Y vdd INVX1
XFILL_1__7983_ gnd vdd FILL
XSFILL38920x29050 gnd vdd FILL
XFILL112440x36050 gnd vdd FILL
XFILL_4__7692_ gnd vdd FILL
XFILL_3__8899_ gnd vdd FILL
XFILL_1__9722_ gnd vdd FILL
XFILL_1__6934_ gnd vdd FILL
X_9468_ _9468_/A gnd _9470_/A vdd INVX1
X_10350_ _10302_/A _7781_/CLK _8670_/R vdd _10350_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert800 gnd vdd FILL
XSFILL39000x38050 gnd vdd FILL
XFILL_1__9653_ gnd vdd FILL
XFILL_4_BUFX2_insert811 gnd vdd FILL
X_8419_ _8349_/A _7651_/CLK _7011_/R vdd _8351_/Y gnd vdd DFFSR
XFILL_1__6865_ gnd vdd FILL
XSFILL49160x82050 gnd vdd FILL
X_9399_ _9399_/A _9398_/A _9399_/C gnd _9399_/Y vdd OAI21X1
XSFILL79400x43050 gnd vdd FILL
XFILL_4_BUFX2_insert822 gnd vdd FILL
XFILL_4__9362_ gnd vdd FILL
XFILL_4_BUFX2_insert833 gnd vdd FILL
XSFILL3640x69050 gnd vdd FILL
XFILL_1__8604_ gnd vdd FILL
X_10281_ _10343_/Q gnd _10281_/Y vdd INVX1
XFILL_4_BUFX2_insert844 gnd vdd FILL
XFILL_4_BUFX2_insert855 gnd vdd FILL
XFILL_4_BUFX2_insert866 gnd vdd FILL
XFILL_4__8313_ gnd vdd FILL
XFILL_4__9293_ gnd vdd FILL
X_12020_ _12084_/A _12713_/A _12084_/C gnd _12022_/B vdd NAND3X1
XFILL_4_BUFX2_insert877 gnd vdd FILL
XFILL_6__9229_ gnd vdd FILL
XSFILL114600x52050 gnd vdd FILL
XFILL_4_BUFX2_insert888 gnd vdd FILL
XFILL_4_BUFX2_insert899 gnd vdd FILL
XSFILL44120x29050 gnd vdd FILL
XFILL_4__8244_ gnd vdd FILL
XSFILL69080x33050 gnd vdd FILL
XFILL_1__8466_ gnd vdd FILL
X_13971_ _8596_/A _13864_/B _14403_/C _8544_/Q gnd _13971_/Y vdd AOI22X1
XFILL_1__7417_ gnd vdd FILL
XFILL_1__8397_ gnd vdd FILL
XFILL_2__7190_ gnd vdd FILL
X_15710_ _7782_/Q gnd _15711_/D vdd INVX1
X_12922_ _12125_/B _9050_/CLK _9050_/R vdd _12922_/D gnd vdd DFFSR
XFILL_1__7348_ gnd vdd FILL
XFILL_4__7057_ gnd vdd FILL
X_15641_ _15641_/A _15641_/B gnd _15650_/A vdd NAND2X1
XFILL_5_BUFX2_insert0 gnd vdd FILL
XSFILL23800x51050 gnd vdd FILL
X_12853_ _12929_/Q gnd _12853_/Y vdd INVX1
XFILL_1_BUFX2_insert701 gnd vdd FILL
XFILL_1_BUFX2_insert712 gnd vdd FILL
XSFILL89240x46050 gnd vdd FILL
XFILL_5__7870_ gnd vdd FILL
XFILL_1_BUFX2_insert723 gnd vdd FILL
X_11804_ _11444_/Y _11778_/B _11804_/C gnd _11805_/C vdd OAI21X1
XFILL_1_BUFX2_insert734 gnd vdd FILL
X_15572_ _15550_/Y _15571_/Y _15572_/C gnd _15572_/Y vdd NOR3X1
XFILL_1__9018_ gnd vdd FILL
X_12784_ _12782_/Y _12789_/A _12784_/C gnd _12820_/D vdd OAI21X1
XFILL_1_BUFX2_insert745 gnd vdd FILL
XFILL_2__9900_ gnd vdd FILL
XFILL_1_BUFX2_insert756 gnd vdd FILL
XSFILL3720x49050 gnd vdd FILL
XFILL_1_BUFX2_insert767 gnd vdd FILL
X_14523_ _9580_/Q gnd _14524_/A vdd INVX1
XFILL_1_BUFX2_insert778 gnd vdd FILL
XFILL_5__11260_ gnd vdd FILL
X_11735_ _11267_/Y _11682_/B _11734_/Y gnd _11735_/Y vdd OAI21X1
XFILL_1_BUFX2_insert789 gnd vdd FILL
XFILL_4__11990_ gnd vdd FILL
XFILL_2__11080_ gnd vdd FILL
XFILL_1__10830_ gnd vdd FILL
XSFILL94360x37050 gnd vdd FILL
XFILL_5__9540_ gnd vdd FILL
XFILL_4__7959_ gnd vdd FILL
X_14454_ _14454_/A gnd _14454_/Y vdd INVX1
XFILL_4__10941_ gnd vdd FILL
XFILL_4_BUFX2_insert16 gnd vdd FILL
XFILL_2__10031_ gnd vdd FILL
X_11666_ _11060_/Y _11573_/C gnd _11666_/Y vdd NAND2X1
XFILL_5__11191_ gnd vdd FILL
XFILL_2__9762_ gnd vdd FILL
XFILL_3__12370_ gnd vdd FILL
XFILL_4_BUFX2_insert27 gnd vdd FILL
XFILL_0__11210_ gnd vdd FILL
XFILL_2__6974_ gnd vdd FILL
XFILL_1__10761_ gnd vdd FILL
XFILL_4_BUFX2_insert38 gnd vdd FILL
XFILL_5__9471_ gnd vdd FILL
X_13405_ _13381_/B _13381_/A gnd _13718_/A vdd AND2X2
XSFILL69160x13050 gnd vdd FILL
XFILL_0__12190_ gnd vdd FILL
XFILL_4_BUFX2_insert49 gnd vdd FILL
XFILL_5__10142_ gnd vdd FILL
X_10617_ _13530_/A gnd _10617_/Y vdd INVX1
XFILL_4__13660_ gnd vdd FILL
XFILL_2__8713_ gnd vdd FILL
X_14385_ _8809_/Q gnd _14386_/D vdd INVX1
XFILL_3__11321_ gnd vdd FILL
XFILL_1__12500_ gnd vdd FILL
XFILL_4__10872_ gnd vdd FILL
X_11597_ _11597_/A _11596_/Y _11587_/C gnd _11597_/Y vdd AOI21X1
XFILL_0__11141_ gnd vdd FILL
XFILL_1__10692_ gnd vdd FILL
X_16124_ _16124_/A _16102_/Y _15651_/C gnd _12902_/B vdd AOI21X1
XFILL_1__13480_ gnd vdd FILL
XFILL_4__9629_ gnd vdd FILL
X_13336_ _13209_/B _13288_/B _13282_/B gnd _13337_/C vdd AOI21X1
XFILL_4__12611_ gnd vdd FILL
XFILL_3__14040_ gnd vdd FILL
XFILL_5__14950_ gnd vdd FILL
X_10548_ _10548_/A _10548_/B _10547_/Y gnd _10602_/D vdd OAI21X1
XFILL_4__13591_ gnd vdd FILL
XFILL_2__8644_ gnd vdd FILL
XFILL_3__11252_ gnd vdd FILL
XSFILL104360x22050 gnd vdd FILL
XFILL_1__12431_ gnd vdd FILL
XFILL_2__14770_ gnd vdd FILL
XFILL_5__8353_ gnd vdd FILL
XFILL_2__11982_ gnd vdd FILL
XSFILL104520x5050 gnd vdd FILL
XFILL_0__11072_ gnd vdd FILL
X_16055_ _9839_/Q gnd _16055_/Y vdd INVX1
XFILL_5__13901_ gnd vdd FILL
X_13267_ _13263_/C _13266_/Y gnd _13268_/B vdd NAND2X1
XFILL_4__15330_ gnd vdd FILL
XFILL_5__14881_ gnd vdd FILL
X_10479_ _16070_/A _8815_/CLK _8047_/R vdd _10435_/Y gnd vdd DFFSR
XFILL_2__13721_ gnd vdd FILL
XFILL_2__10933_ gnd vdd FILL
XFILL_2__8575_ gnd vdd FILL
XFILL_1__12362_ gnd vdd FILL
XFILL_5__7304_ gnd vdd FILL
XFILL_0__10023_ gnd vdd FILL
XFILL_3__11183_ gnd vdd FILL
XFILL_0__14900_ gnd vdd FILL
XFILL_1__15150_ gnd vdd FILL
XSFILL8840x82050 gnd vdd FILL
X_15006_ _15953_/A gnd _15356_/C vdd INVX4
X_12218_ _12218_/A _12214_/Y _12217_/Y gnd _12218_/Y vdd NAND3X1
XFILL_0__15880_ gnd vdd FILL
XFILL_5__13832_ gnd vdd FILL
XFILL_4__15261_ gnd vdd FILL
XFILL_0__7590_ gnd vdd FILL
XSFILL59080x65050 gnd vdd FILL
X_13198_ _12184_/A _13175_/CLK _13199_/R vdd _13150_/Y gnd vdd DFFSR
XFILL_4__12473_ gnd vdd FILL
XFILL_1__11313_ gnd vdd FILL
XFILL_3__10134_ gnd vdd FILL
XFILL_1__14101_ gnd vdd FILL
XFILL_2__13652_ gnd vdd FILL
XSFILL99480x70050 gnd vdd FILL
XFILL_3__15991_ gnd vdd FILL
XFILL_0__14831_ gnd vdd FILL
XFILL_1__15081_ gnd vdd FILL
XFILL_1__12293_ gnd vdd FILL
XFILL_5__7235_ gnd vdd FILL
XFILL_4__14212_ gnd vdd FILL
X_12149_ _12134_/A _12856_/A gnd _12150_/C vdd NAND2X1
XFILL_4__11424_ gnd vdd FILL
XFILL_2__12603_ gnd vdd FILL
XFILL_4__15192_ gnd vdd FILL
XFILL_5__13763_ gnd vdd FILL
XSFILL79080x9050 gnd vdd FILL
XFILL_5__10975_ gnd vdd FILL
XFILL_2__16371_ gnd vdd FILL
XFILL_2__7457_ gnd vdd FILL
XFILL_1__14032_ gnd vdd FILL
XFILL_3__14942_ gnd vdd FILL
XFILL_1__11244_ gnd vdd FILL
XFILL_3__10065_ gnd vdd FILL
XFILL_2__13583_ gnd vdd FILL
XFILL_0__11974_ gnd vdd FILL
XFILL_2__10795_ gnd vdd FILL
XFILL_5__7166_ gnd vdd FILL
XFILL_0__14762_ gnd vdd FILL
XFILL_5__15502_ gnd vdd FILL
XFILL_5__12714_ gnd vdd FILL
XFILL_6__10176_ gnd vdd FILL
XFILL_4__14143_ gnd vdd FILL
XFILL_0__9260_ gnd vdd FILL
XFILL_2__15322_ gnd vdd FILL
XSFILL94440x17050 gnd vdd FILL
XFILL_4__11355_ gnd vdd FILL
XFILL_3__14873_ gnd vdd FILL
XFILL_2__12534_ gnd vdd FILL
XFILL_5__13694_ gnd vdd FILL
XFILL_0__10925_ gnd vdd FILL
XFILL_0__13713_ gnd vdd FILL
XFILL_1__11175_ gnd vdd FILL
XFILL_0__8211_ gnd vdd FILL
XSFILL13800x83050 gnd vdd FILL
X_15908_ _15908_/A _15905_/Y gnd _15908_/Y vdd NOR2X1
XFILL_5__7097_ gnd vdd FILL
XFILL_0__14693_ gnd vdd FILL
XFILL_4__10306_ gnd vdd FILL
XFILL_5__15433_ gnd vdd FILL
XFILL_5__12645_ gnd vdd FILL
XFILL_3__13824_ gnd vdd FILL
XFILL_6__14984_ gnd vdd FILL
XFILL_2__9127_ gnd vdd FILL
XFILL_4__14074_ gnd vdd FILL
XFILL_0_BUFX2_insert1003 gnd vdd FILL
XFILL_1__10126_ gnd vdd FILL
XFILL_2__15253_ gnd vdd FILL
XFILL_4__11286_ gnd vdd FILL
XSFILL79240x78050 gnd vdd FILL
XFILL_0_BUFX2_insert1014 gnd vdd FILL
XFILL_2__12465_ gnd vdd FILL
XSFILL94280x3050 gnd vdd FILL
XFILL_0_BUFX2_insert1025 gnd vdd FILL
XFILL_1__15983_ gnd vdd FILL
XFILL_0__13644_ gnd vdd FILL
XFILL_0__8142_ gnd vdd FILL
XFILL_4__13025_ gnd vdd FILL
XFILL_6__13935_ gnd vdd FILL
XFILL_0_BUFX2_insert1036 gnd vdd FILL
XFILL_2__14204_ gnd vdd FILL
XFILL_5__15364_ gnd vdd FILL
X_15839_ _15839_/A _15838_/Y gnd _15840_/B vdd NOR2X1
XFILL_4__10237_ gnd vdd FILL
XFILL_5__12576_ gnd vdd FILL
XFILL_3__13755_ gnd vdd FILL
XFILL_0_BUFX2_insert1047 gnd vdd FILL
X_8770_ _8753_/B _9794_/B gnd _8771_/C vdd NAND2X1
XFILL_2__11416_ gnd vdd FILL
XFILL_3__10967_ gnd vdd FILL
XFILL_2__15184_ gnd vdd FILL
XFILL_2_BUFX2_insert590 gnd vdd FILL
XFILL_1__14934_ gnd vdd FILL
XFILL_0_BUFX2_insert1058 gnd vdd FILL
XFILL_1__10057_ gnd vdd FILL
XFILL_3__9940_ gnd vdd FILL
XFILL_0__16363_ gnd vdd FILL
XFILL_2__12396_ gnd vdd FILL
XFILL_0__13575_ gnd vdd FILL
XFILL_0_BUFX2_insert1069 gnd vdd FILL
XFILL_0__10787_ gnd vdd FILL
XFILL_5__14315_ gnd vdd FILL
XFILL_3__12706_ gnd vdd FILL
XFILL_0__8073_ gnd vdd FILL
XFILL_5__11527_ gnd vdd FILL
X_7721_ _7721_/A gnd _7723_/A vdd INVX1
XFILL_2__8009_ gnd vdd FILL
XFILL_2__14135_ gnd vdd FILL
XFILL_4__10168_ gnd vdd FILL
XFILL_5__15295_ gnd vdd FILL
XFILL_3__9871_ gnd vdd FILL
XFILL_3__13686_ gnd vdd FILL
XFILL_0__15314_ gnd vdd FILL
XFILL_0__12526_ gnd vdd FILL
XFILL_2__11347_ gnd vdd FILL
XFILL_5__9807_ gnd vdd FILL
XFILL_3__10898_ gnd vdd FILL
XFILL_1__14865_ gnd vdd FILL
XFILL_0__16294_ gnd vdd FILL
XFILL_5__7999_ gnd vdd FILL
XFILL_5__14246_ gnd vdd FILL
XFILL_3__12637_ gnd vdd FILL
XFILL_6__13797_ gnd vdd FILL
XFILL_3__8822_ gnd vdd FILL
X_7652_ _7584_/A _9188_/CLK _8801_/R vdd _7652_/D gnd vdd DFFSR
XFILL_5__11458_ gnd vdd FILL
XFILL_3__15425_ gnd vdd FILL
XFILL_1__13816_ gnd vdd FILL
XFILL_2__14066_ gnd vdd FILL
XFILL_4__14976_ gnd vdd FILL
XFILL_0__12457_ gnd vdd FILL
XFILL_0__15245_ gnd vdd FILL
XSFILL59160x45050 gnd vdd FILL
XFILL_6__8531_ gnd vdd FILL
XFILL_2__11278_ gnd vdd FILL
XFILL_5__9738_ gnd vdd FILL
XFILL_1__14796_ gnd vdd FILL
XFILL_6__15536_ gnd vdd FILL
XFILL_6__12748_ gnd vdd FILL
XFILL_5__10409_ gnd vdd FILL
XFILL_3__15356_ gnd vdd FILL
XFILL_5__14177_ gnd vdd FILL
XFILL_2__13017_ gnd vdd FILL
X_7583_ _7583_/A _7624_/A _7583_/C gnd _7583_/Y vdd OAI21X1
XFILL_5__11389_ gnd vdd FILL
XFILL_4__13927_ gnd vdd FILL
XFILL_3__12568_ gnd vdd FILL
XFILL_0__11408_ gnd vdd FILL
XFILL_3__8753_ gnd vdd FILL
XFILL_0__15176_ gnd vdd FILL
XFILL_1__13747_ gnd vdd FILL
XFILL_1__10959_ gnd vdd FILL
XFILL_0__12388_ gnd vdd FILL
XFILL111880x44050 gnd vdd FILL
XFILL_5__13128_ gnd vdd FILL
XFILL_5__9669_ gnd vdd FILL
XFILL_3__14307_ gnd vdd FILL
X_9322_ _9266_/A _9705_/CLK _7914_/R vdd _9268_/Y gnd vdd DFFSR
XFILL_0__8975_ gnd vdd FILL
XFILL_3__7704_ gnd vdd FILL
XFILL_3__11519_ gnd vdd FILL
XFILL_4__13858_ gnd vdd FILL
XFILL_3__15287_ gnd vdd FILL
XFILL_0__14127_ gnd vdd FILL
XFILL_3__12499_ gnd vdd FILL
XFILL_0__11339_ gnd vdd FILL
XFILL_1__13678_ gnd vdd FILL
XFILL_0__7926_ gnd vdd FILL
XFILL_6__15398_ gnd vdd FILL
X_9253_ _9251_/Y _9277_/B _9252_/Y gnd _9253_/Y vdd OAI21X1
XFILL_3__14238_ gnd vdd FILL
XFILL_4_BUFX2_insert107 gnd vdd FILL
XSFILL109400x76050 gnd vdd FILL
XFILL_3__7635_ gnd vdd FILL
XFILL_1__15417_ gnd vdd FILL
XFILL_1__12629_ gnd vdd FILL
XFILL_4__13789_ gnd vdd FILL
XFILL_0__14058_ gnd vdd FILL
XFILL_2__14968_ gnd vdd FILL
XFILL_1__16397_ gnd vdd FILL
XSFILL8680x4050 gnd vdd FILL
X_8204_ _8246_/A _6924_/B gnd _8204_/Y vdd NAND2X1
XFILL_6__14349_ gnd vdd FILL
XSFILL54040x6050 gnd vdd FILL
XFILL_4__15528_ gnd vdd FILL
XFILL_0__7857_ gnd vdd FILL
X_9184_ _9184_/Q _7791_/CLK _9711_/R vdd _9184_/D gnd vdd DFFSR
XFILL_3__14169_ gnd vdd FILL
XFILL_0__13009_ gnd vdd FILL
XFILL_2__13919_ gnd vdd FILL
XFILL_3__7566_ gnd vdd FILL
XFILL_1__15348_ gnd vdd FILL
XFILL_2__14899_ gnd vdd FILL
X_8135_ _8177_/Q gnd _8137_/A vdd INVX1
XFILL_3_BUFX2_insert807 gnd vdd FILL
XFILL_3_BUFX2_insert818 gnd vdd FILL
XFILL_4__15459_ gnd vdd FILL
XSFILL114520x67050 gnd vdd FILL
XFILL_3_BUFX2_insert829 gnd vdd FILL
XFILL_3__7497_ gnd vdd FILL
XFILL_1__15279_ gnd vdd FILL
XFILL_0__9527_ gnd vdd FILL
XFILL_1__8320_ gnd vdd FILL
X_8066_ _8066_/A gnd _8066_/Y vdd INVX1
XFILL_3__9236_ gnd vdd FILL
X_7017_ _6959_/A _7916_/CLK _9580_/R vdd _7017_/D gnd vdd DFFSR
XFILL_1__8251_ gnd vdd FILL
XFILL_3__9167_ gnd vdd FILL
XFILL_1__7202_ gnd vdd FILL
XFILL_3__8118_ gnd vdd FILL
XFILL_1__8182_ gnd vdd FILL
XFILL_0__9389_ gnd vdd FILL
XFILL_3__9098_ gnd vdd FILL
XFILL_6__9916_ gnd vdd FILL
XFILL_4__9980_ gnd vdd FILL
XSFILL23720x66050 gnd vdd FILL
X_8968_ _8968_/A gnd _8968_/Y vdd INVX1
XFILL112040x33050 gnd vdd FILL
XFILL_1__7064_ gnd vdd FILL
X_7919_ _7919_/Q _9568_/CLK _8431_/R vdd _7875_/Y gnd vdd DFFSR
XFILL_4__8862_ gnd vdd FILL
X_8899_ _8899_/A _8902_/B _8898_/Y gnd _8943_/D vdd OAI21X1
XSFILL113720x19050 gnd vdd FILL
XFILL_0_CLKBUF1_insert112 gnd vdd FILL
XFILL_0_CLKBUF1_insert123 gnd vdd FILL
XSFILL39400x54050 gnd vdd FILL
XFILL_0_BUFX2_insert708 gnd vdd FILL
XFILL_4__7813_ gnd vdd FILL
XFILL_0_CLKBUF1_insert134 gnd vdd FILL
XFILL_0_BUFX2_insert719 gnd vdd FILL
XFILL_0_CLKBUF1_insert145 gnd vdd FILL
X_11520_ _11569_/C _11520_/B _11518_/Y gnd _11521_/A vdd AOI21X1
XFILL_0_CLKBUF1_insert156 gnd vdd FILL
XFILL_0_CLKBUF1_insert167 gnd vdd FILL
XFILL_0_CLKBUF1_insert178 gnd vdd FILL
XFILL_4__7744_ gnd vdd FILL
XFILL_0_CLKBUF1_insert189 gnd vdd FILL
X_11451_ _11297_/Y _11451_/B gnd _11550_/A vdd NOR2X1
XSFILL69080x28050 gnd vdd FILL
XFILL_1__7966_ gnd vdd FILL
X_10402_ _10402_/A _10372_/B _10401_/Y gnd _10402_/Y vdd OAI21X1
XFILL_4__7675_ gnd vdd FILL
X_14170_ _14170_/A _14170_/B gnd _14171_/A vdd NOR2X1
XFILL_1__6917_ gnd vdd FILL
X_11382_ _12238_/Y _11031_/B _11381_/Y gnd _11382_/Y vdd OAI21X1
XFILL_4__9414_ gnd vdd FILL
X_13121_ _11929_/A gnd _13123_/A vdd INVX1
XSFILL104280x37050 gnd vdd FILL
X_10333_ _10333_/Q _7261_/CLK _8669_/R vdd _10253_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert630 gnd vdd FILL
XFILL_1__9636_ gnd vdd FILL
XFILL_4_BUFX2_insert641 gnd vdd FILL
XFILL_1__6848_ gnd vdd FILL
XFILL_4__9345_ gnd vdd FILL
XFILL_4_BUFX2_insert652 gnd vdd FILL
XFILL_4_BUFX2_insert663 gnd vdd FILL
XFILL_4_BUFX2_insert674 gnd vdd FILL
X_13052_ _6875_/A _8169_/CLK _8937_/R vdd _13052_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert685 gnd vdd FILL
X_10264_ _10264_/A _8600_/B gnd _10265_/C vdd NAND2X1
XFILL_2__8360_ gnd vdd FILL
XFILL_4_BUFX2_insert696 gnd vdd FILL
XFILL_4__9276_ gnd vdd FILL
X_12003_ _12007_/A _12355_/A _12059_/C gnd _12006_/A vdd NAND3X1
XFILL112120x13050 gnd vdd FILL
XFILL_2__7311_ gnd vdd FILL
XFILL_1__8518_ gnd vdd FILL
X_10195_ _10229_/Q gnd _10197_/A vdd INVX1
XSFILL74040x83050 gnd vdd FILL
XFILL_4__8227_ gnd vdd FILL
XFILL_1__9498_ gnd vdd FILL
XFILL_5__10760_ gnd vdd FILL
XSFILL38840x6050 gnd vdd FILL
XFILL_1__8449_ gnd vdd FILL
XFILL_2__7242_ gnd vdd FILL
XFILL_2__10580_ gnd vdd FILL
XSFILL13480x36050 gnd vdd FILL
X_13954_ _8724_/A gnd _13956_/A vdd INVX1
XFILL_4__11140_ gnd vdd FILL
XFILL_5__10691_ gnd vdd FILL
XFILL_4__7109_ gnd vdd FILL
XFILL_3__11870_ gnd vdd FILL
XFILL_2__7173_ gnd vdd FILL
XFILL_4__8089_ gnd vdd FILL
XFILL_0__11690_ gnd vdd FILL
X_12905_ vdd _16164_/Y gnd _12905_/Y vdd NAND2X1
XFILL_5__12430_ gnd vdd FILL
XFILL_5__8971_ gnd vdd FILL
X_13885_ _13883_/Y _13885_/B _13880_/Y gnd _13885_/Y vdd NAND3X1
XSFILL94760x53050 gnd vdd FILL
XFILL_3__10821_ gnd vdd FILL
XFILL_4__11071_ gnd vdd FILL
XFILL_2__12250_ gnd vdd FILL
XFILL_0__10641_ gnd vdd FILL
XFILL_6__13720_ gnd vdd FILL
XFILL_1__12980_ gnd vdd FILL
XSFILL84200x11050 gnd vdd FILL
XFILL_4__10022_ gnd vdd FILL
X_15624_ _15624_/A _16213_/B gnd _15627_/B vdd NOR2X1
XFILL_5__12361_ gnd vdd FILL
X_12836_ vdd _12836_/B gnd _12837_/C vdd NAND2X1
XFILL_1_BUFX2_insert520 gnd vdd FILL
XFILL_1_BUFX2_insert531 gnd vdd FILL
XFILL_3__13540_ gnd vdd FILL
XFILL_2__11201_ gnd vdd FILL
XFILL_3__10752_ gnd vdd FILL
XFILL_0__13360_ gnd vdd FILL
XFILL_1__11931_ gnd vdd FILL
XFILL_1_BUFX2_insert542 gnd vdd FILL
XFILL_2__12181_ gnd vdd FILL
XFILL_1_BUFX2_insert553 gnd vdd FILL
XFILL_0__10572_ gnd vdd FILL
XFILL_5__7853_ gnd vdd FILL
XFILL_5__14100_ gnd vdd FILL
X_15555_ _15555_/A _15555_/B gnd _15560_/A vdd NOR2X1
XFILL_5__11312_ gnd vdd FILL
XFILL_1_BUFX2_insert564 gnd vdd FILL
X_12767_ _12767_/A gnd _12767_/Y vdd INVX1
XFILL_1_BUFX2_insert575 gnd vdd FILL
XFILL_4__14830_ gnd vdd FILL
XFILL_5__12292_ gnd vdd FILL
XSFILL109400x50 gnd vdd FILL
XFILL_5__15080_ gnd vdd FILL
XFILL_3__13471_ gnd vdd FILL
XFILL_0__12311_ gnd vdd FILL
XFILL_2__11132_ gnd vdd FILL
XFILL_3__10683_ gnd vdd FILL
XFILL_1_BUFX2_insert586 gnd vdd FILL
XFILL_1__14650_ gnd vdd FILL
XFILL_0__13291_ gnd vdd FILL
X_14506_ _14506_/A _15948_/B _14506_/C _15937_/C gnd _14506_/Y vdd OAI22X1
XFILL_1_BUFX2_insert597 gnd vdd FILL
XFILL_1__11862_ gnd vdd FILL
XFILL_3__15210_ gnd vdd FILL
XFILL_6__16370_ gnd vdd FILL
XFILL_5__14031_ gnd vdd FILL
X_11718_ _11718_/A gnd _12473_/B vdd INVX1
XFILL_5__11243_ gnd vdd FILL
XFILL_3__12422_ gnd vdd FILL
X_15486_ _13940_/A _15581_/C _15544_/A _13937_/B gnd _15486_/Y vdd OAI22X1
XFILL_6__13582_ gnd vdd FILL
X_12698_ _12792_/Q gnd _12700_/A vdd INVX1
XFILL_1__13601_ gnd vdd FILL
XFILL_4__11973_ gnd vdd FILL
XFILL_3__16190_ gnd vdd FILL
XFILL_0__15030_ gnd vdd FILL
XFILL_2__15940_ gnd vdd FILL
XFILL_2__11063_ gnd vdd FILL
XFILL_4__14761_ gnd vdd FILL
XFILL_1__10813_ gnd vdd FILL
XFILL_0__12242_ gnd vdd FILL
XFILL_1__14581_ gnd vdd FILL
XFILL_6__15321_ gnd vdd FILL
XFILL_5__9523_ gnd vdd FILL
XSFILL64040x1050 gnd vdd FILL
XSFILL99480x65050 gnd vdd FILL
XSFILL103640x1050 gnd vdd FILL
XFILL_1__11793_ gnd vdd FILL
X_14437_ _14437_/A _14437_/B gnd _14438_/A vdd NOR2X1
XSFILL74120x63050 gnd vdd FILL
X_11649_ _11641_/C gnd _11649_/Y vdd INVX2
XFILL_4__13712_ gnd vdd FILL
XFILL_3__15141_ gnd vdd FILL
XFILL_5__11174_ gnd vdd FILL
XFILL_3__12353_ gnd vdd FILL
XFILL_4__10924_ gnd vdd FILL
XFILL_1__16320_ gnd vdd FILL
XFILL_2__10014_ gnd vdd FILL
XFILL_2__9745_ gnd vdd FILL
XFILL_2__6957_ gnd vdd FILL
XFILL_4__14692_ gnd vdd FILL
XFILL_1__13532_ gnd vdd FILL
XFILL_2__15871_ gnd vdd FILL
XFILL_1__10744_ gnd vdd FILL
XFILL_0__12173_ gnd vdd FILL
XFILL_5__10125_ gnd vdd FILL
XFILL_6__12464_ gnd vdd FILL
XFILL_0__8760_ gnd vdd FILL
X_14368_ _8495_/A gnd _14370_/D vdd INVX1
XFILL_3__11304_ gnd vdd FILL
XFILL_5__15982_ gnd vdd FILL
XFILL_4__13643_ gnd vdd FILL
XFILL_2__14822_ gnd vdd FILL
XFILL_3__15072_ gnd vdd FILL
XSFILL13560x16050 gnd vdd FILL
XFILL_2__9676_ gnd vdd FILL
XFILL_3__12284_ gnd vdd FILL
XFILL_0__11124_ gnd vdd FILL
XFILL_1__16251_ gnd vdd FILL
XFILL_1__13463_ gnd vdd FILL
X_16107_ _16107_/A gnd _16107_/Y vdd INVX1
XFILL_2__6888_ gnd vdd FILL
XFILL_5__8405_ gnd vdd FILL
XFILL_1__10675_ gnd vdd FILL
XSFILL3400x26050 gnd vdd FILL
X_13319_ _13305_/A _13244_/B _13316_/Y gnd _13320_/B vdd OAI21X1
XFILL_5__9385_ gnd vdd FILL
XFILL_0__7711_ gnd vdd FILL
XSFILL53960x21050 gnd vdd FILL
XFILL_6__11415_ gnd vdd FILL
XFILL_6__15183_ gnd vdd FILL
XFILL_3__14023_ gnd vdd FILL
XFILL_5__10056_ gnd vdd FILL
XFILL_5__14933_ gnd vdd FILL
XFILL_1__15202_ gnd vdd FILL
X_14299_ _10343_/Q gnd _14299_/Y vdd INVX1
XFILL_4__16362_ gnd vdd FILL
XFILL_4__13574_ gnd vdd FILL
XFILL_3__7420_ gnd vdd FILL
XFILL_2__8627_ gnd vdd FILL
XFILL_3__11235_ gnd vdd FILL
XFILL_1__12414_ gnd vdd FILL
XSFILL109480x50050 gnd vdd FILL
XFILL_4__10786_ gnd vdd FILL
XFILL_2__14753_ gnd vdd FILL
XFILL_5__8336_ gnd vdd FILL
XFILL_1__16182_ gnd vdd FILL
XFILL_2__11965_ gnd vdd FILL
XFILL_0__15932_ gnd vdd FILL
XFILL_0__11055_ gnd vdd FILL
X_16038_ _15384_/A _14623_/Y _16037_/Y gnd _16039_/B vdd OAI21X1
XFILL_6__14134_ gnd vdd FILL
XFILL_1__13394_ gnd vdd FILL
XSFILL13800x3050 gnd vdd FILL
XFILL_4__15313_ gnd vdd FILL
XFILL_5__14864_ gnd vdd FILL
XFILL_4__12525_ gnd vdd FILL
XFILL_2__13704_ gnd vdd FILL
XFILL_3__7351_ gnd vdd FILL
XFILL_2__10916_ gnd vdd FILL
XFILL_4__16293_ gnd vdd FILL
XSFILL54040x30050 gnd vdd FILL
XFILL_0__10006_ gnd vdd FILL
XFILL_1__15133_ gnd vdd FILL
XFILL_3__11166_ gnd vdd FILL
XFILL_1__12345_ gnd vdd FILL
XFILL_2__14684_ gnd vdd FILL
XFILL_5__8267_ gnd vdd FILL
XFILL_2__11896_ gnd vdd FILL
XFILL_0__15863_ gnd vdd FILL
XFILL_5__13815_ gnd vdd FILL
XFILL_4__15244_ gnd vdd FILL
XFILL_2__7509_ gnd vdd FILL
XFILL_4__12456_ gnd vdd FILL
XFILL_0__7573_ gnd vdd FILL
XFILL_3__10117_ gnd vdd FILL
XFILL_6__11277_ gnd vdd FILL
XFILL_2__13635_ gnd vdd FILL
XFILL_5__14795_ gnd vdd FILL
XFILL_3__15974_ gnd vdd FILL
XFILL_0__14814_ gnd vdd FILL
XFILL_1__15064_ gnd vdd FILL
XFILL_2__8489_ gnd vdd FILL
XFILL_3__11097_ gnd vdd FILL
XFILL_5__7218_ gnd vdd FILL
XFILL_1__12276_ gnd vdd FILL
XFILL_0__15794_ gnd vdd FILL
XFILL_4__11407_ gnd vdd FILL
XFILL_5__8198_ gnd vdd FILL
XFILL_3__9021_ gnd vdd FILL
XFILL_5__13746_ gnd vdd FILL
X_9940_ _9941_/B _9940_/B gnd _9940_/Y vdd NAND2X1
XFILL_5__10958_ gnd vdd FILL
XSFILL43880x73050 gnd vdd FILL
XFILL_4__15175_ gnd vdd FILL
XFILL_3__10048_ gnd vdd FILL
XFILL_4__12387_ gnd vdd FILL
XFILL_1__14015_ gnd vdd FILL
XFILL_2__16354_ gnd vdd FILL
XFILL_3__14925_ gnd vdd FILL
XFILL_2__13566_ gnd vdd FILL
XFILL_1__11227_ gnd vdd FILL
XFILL_2__10778_ gnd vdd FILL
XFILL_0_BUFX2_insert14 gnd vdd FILL
XFILL_0__14745_ gnd vdd FILL
XFILL_0__11957_ gnd vdd FILL
XFILL_0__9243_ gnd vdd FILL
XFILL_0_BUFX2_insert25 gnd vdd FILL
XFILL_2__15305_ gnd vdd FILL
XFILL_4__14126_ gnd vdd FILL
XFILL_0_BUFX2_insert36 gnd vdd FILL
XFILL_4__11338_ gnd vdd FILL
X_9871_ _9920_/B _8719_/B gnd _9872_/C vdd NAND2X1
XFILL_5__13677_ gnd vdd FILL
XFILL_2__12517_ gnd vdd FILL
XSFILL48920x10050 gnd vdd FILL
XFILL_3__14856_ gnd vdd FILL
XFILL_2__16285_ gnd vdd FILL
XFILL_5__10889_ gnd vdd FILL
XFILL_0_BUFX2_insert47 gnd vdd FILL
XFILL_1__11158_ gnd vdd FILL
XFILL_0__10908_ gnd vdd FILL
XFILL_0_BUFX2_insert58 gnd vdd FILL
XFILL_2__13497_ gnd vdd FILL
XFILL_0_BUFX2_insert69 gnd vdd FILL
XFILL_0__14676_ gnd vdd FILL
XFILL_5__15416_ gnd vdd FILL
XFILL_5__12628_ gnd vdd FILL
XFILL_0__11888_ gnd vdd FILL
X_8822_ _8918_/Q gnd _8822_/Y vdd INVX1
XFILL_4__14057_ gnd vdd FILL
XFILL_3__13807_ gnd vdd FILL
XFILL_2__15236_ gnd vdd FILL
XFILL_5__16396_ gnd vdd FILL
XFILL_1__10109_ gnd vdd FILL
XFILL_4__11269_ gnd vdd FILL
XFILL_2__12448_ gnd vdd FILL
XFILL_0__16415_ gnd vdd FILL
XFILL_0__13627_ gnd vdd FILL
XFILL_3__11999_ gnd vdd FILL
XFILL_1__15966_ gnd vdd FILL
XFILL_3__14787_ gnd vdd FILL
XFILL_1__11089_ gnd vdd FILL
XFILL_0__8125_ gnd vdd FILL
XFILL_4__13008_ gnd vdd FILL
XFILL_5__15347_ gnd vdd FILL
X_8753_ _8753_/A _8753_/B _8752_/Y gnd _8753_/Y vdd OAI21X1
XFILL_6_CLKBUF1_insert1083 gnd vdd FILL
XFILL_3__9923_ gnd vdd FILL
XFILL_2__15167_ gnd vdd FILL
XFILL_3__13738_ gnd vdd FILL
XFILL_1__14917_ gnd vdd FILL
XFILL_0__16346_ gnd vdd FILL
XFILL_2__12379_ gnd vdd FILL
XFILL_6_BUFX2_insert725 gnd vdd FILL
XFILL_1__15897_ gnd vdd FILL
XFILL_6__9632_ gnd vdd FILL
XFILL_0__13558_ gnd vdd FILL
XFILL_0__8056_ gnd vdd FILL
X_7704_ _7684_/B _9624_/B gnd _7705_/C vdd NAND2X1
XFILL_2__14118_ gnd vdd FILL
XFILL_5__15278_ gnd vdd FILL
X_8684_ _8632_/A _9453_/CLK _9453_/R vdd _8634_/Y gnd vdd DFFSR
XFILL_3__13669_ gnd vdd FILL
XFILL_1__14848_ gnd vdd FILL
XFILL_0__12509_ gnd vdd FILL
XFILL_2__15098_ gnd vdd FILL
XFILL_3__9854_ gnd vdd FILL
XFILL_0__16277_ gnd vdd FILL
XFILL_5__14229_ gnd vdd FILL
XSFILL54120x10050 gnd vdd FILL
XFILL_0__13489_ gnd vdd FILL
XFILL_3__15408_ gnd vdd FILL
X_7635_ _7669_/Q gnd _7637_/A vdd INVX1
XFILL_2__14049_ gnd vdd FILL
XFILL_4__14959_ gnd vdd FILL
XFILL_3__16388_ gnd vdd FILL
XFILL_0__15228_ gnd vdd FILL
XFILL_3__9785_ gnd vdd FILL
XFILL_3__6997_ gnd vdd FILL
XFILL_1__14779_ gnd vdd FILL
XFILL_1__7820_ gnd vdd FILL
X_7566_ _7646_/Q gnd _7566_/Y vdd INVX1
XFILL_3__15339_ gnd vdd FILL
XFILL_3__8736_ gnd vdd FILL
XFILL_1_CLKBUF1_insert207 gnd vdd FILL
XFILL_1_CLKBUF1_insert218 gnd vdd FILL
XSFILL43960x53050 gnd vdd FILL
XFILL_0__15159_ gnd vdd FILL
X_9305_ _9215_/A _8921_/CLK _9049_/R vdd _9217_/Y gnd vdd DFFSR
XFILL_0__8958_ gnd vdd FILL
XFILL_1__7751_ gnd vdd FILL
XFILL_1__16449_ gnd vdd FILL
XFILL_4__7460_ gnd vdd FILL
XSFILL84040x46050 gnd vdd FILL
X_7497_ _7495_/Y _7416_/B _7497_/C gnd _7537_/D vdd OAI21X1
XFILL_6__8376_ gnd vdd FILL
XSFILL99640x25050 gnd vdd FILL
X_9236_ _9312_/Q gnd _9238_/A vdd INVX1
XSFILL44040x62050 gnd vdd FILL
XFILL_1__7682_ gnd vdd FILL
XFILL_0__8889_ gnd vdd FILL
XFILL_3__7618_ gnd vdd FILL
XFILL_3__8598_ gnd vdd FILL
XFILL_6__7327_ gnd vdd FILL
XFILL111960x19050 gnd vdd FILL
XFILL_1__9421_ gnd vdd FILL
X_9167_ _9165_/Y _9163_/A _9167_/C gnd _9203_/D vdd OAI21X1
XFILL_4__9130_ gnd vdd FILL
XFILL_3_BUFX2_insert604 gnd vdd FILL
XFILL_3__7549_ gnd vdd FILL
XFILL_3_BUFX2_insert615 gnd vdd FILL
XFILL_3_BUFX2_insert626 gnd vdd FILL
X_8118_ _8118_/A _7094_/B gnd _8119_/C vdd NAND2X1
XFILL_1__9352_ gnd vdd FILL
XFILL_3_BUFX2_insert637 gnd vdd FILL
XSFILL23880x20050 gnd vdd FILL
XFILL112040x28050 gnd vdd FILL
X_9098_ _9098_/A _9151_/A _9097_/Y gnd _9098_/Y vdd OAI21X1
XFILL_3_BUFX2_insert648 gnd vdd FILL
XFILL_3_BUFX2_insert659 gnd vdd FILL
XSFILL59880x6050 gnd vdd FILL
XFILL_3__9219_ gnd vdd FILL
XFILL_4__8012_ gnd vdd FILL
XFILL_1__9283_ gnd vdd FILL
XSFILL38120x23050 gnd vdd FILL
X_8049_ _8049_/Q _7786_/CLK _7153_/R vdd _8049_/D gnd vdd DFFSR
XSFILL89560x77050 gnd vdd FILL
XFILL_1__8234_ gnd vdd FILL
X_10951_ _10940_/Y gnd _10955_/A vdd INVX1
XSFILL68840x78050 gnd vdd FILL
XFILL_1__7116_ gnd vdd FILL
X_13670_ _10114_/A gnd _15233_/C vdd INVX1
X_10882_ _10882_/A _10882_/B gnd _10882_/Y vdd NOR2X1
XSFILL109480x7050 gnd vdd FILL
XFILL_1__8096_ gnd vdd FILL
XFILL_4__8914_ gnd vdd FILL
X_12621_ _12621_/A gnd _12621_/Y vdd INVX1
XSFILL94280x70050 gnd vdd FILL
XFILL_4__9894_ gnd vdd FILL
XFILL_1__7047_ gnd vdd FILL
XFILL_4__8845_ gnd vdd FILL
X_15340_ _13794_/Y _16002_/A gnd _15343_/A vdd NOR2X1
XFILL_0_BUFX2_insert505 gnd vdd FILL
XFILL_0_BUFX2_insert516 gnd vdd FILL
X_12552_ _12055_/B _13180_/CLK _13180_/R vdd _12492_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert527 gnd vdd FILL
XFILL_2__7860_ gnd vdd FILL
XFILL_0_BUFX2_insert538 gnd vdd FILL
XFILL_0_BUFX2_insert549 gnd vdd FILL
X_11503_ _11503_/A _11500_/Y _11503_/C gnd _11504_/C vdd AOI21X1
XFILL_4__8776_ gnd vdd FILL
XSFILL33160x66050 gnd vdd FILL
X_15271_ _13722_/A _15025_/B _15756_/D _15270_/Y gnd _15272_/B vdd OAI22X1
X_12483_ _12483_/A vdd _12482_/Y gnd _12549_/D vdd OAI21X1
XFILL_1__8998_ gnd vdd FILL
X_14222_ _8870_/A gnd _14222_/Y vdd INVX1
XFILL_4__7727_ gnd vdd FILL
X_11434_ _11542_/A _11107_/B gnd _11435_/A vdd NAND2X1
XFILL_2__9530_ gnd vdd FILL
XFILL_1__7949_ gnd vdd FILL
X_14153_ _14152_/Y _14153_/B gnd _14154_/C vdd NOR2X1
XFILL_4__10640_ gnd vdd FILL
X_11365_ _11200_/Y _11848_/A gnd _11366_/C vdd NAND2X1
X_13104_ _13168_/B _12022_/Y gnd _13104_/Y vdd NAND2X1
XFILL_5__9170_ gnd vdd FILL
XFILL_6__11200_ gnd vdd FILL
X_10316_ _10316_/A _10318_/A _10315_/Y gnd _10316_/Y vdd OAI21X1
XFILL_4__7589_ gnd vdd FILL
XFILL_4_BUFX2_insert460 gnd vdd FILL
XCLKBUF1_insert206 CLKBUF1_insert206/A gnd _7389_/CLK vdd CLKBUF1
XFILL_5__11930_ gnd vdd FILL
X_14084_ _14084_/A _14084_/B gnd _14085_/C vdd NOR2X1
XFILL_3__11020_ gnd vdd FILL
XFILL_4_BUFX2_insert471 gnd vdd FILL
XFILL_4__10571_ gnd vdd FILL
X_11296_ _11313_/B _11295_/Y gnd _11303_/B vdd NAND2X1
XFILL_1__9619_ gnd vdd FILL
XCLKBUF1_insert217 CLKBUF1_insert218/A gnd _7661_/CLK vdd CLKBUF1
XFILL_5__8121_ gnd vdd FILL
XFILL_4_BUFX2_insert482 gnd vdd FILL
XFILL_2__9392_ gnd vdd FILL
XFILL112360x50 gnd vdd FILL
XFILL_2__11750_ gnd vdd FILL
XFILL_4_BUFX2_insert493 gnd vdd FILL
XFILL_1__10391_ gnd vdd FILL
X_13035_ _6898_/A gnd _13035_/Y vdd INVX1
XFILL_4__12310_ gnd vdd FILL
X_10247_ _10247_/A _10325_/B _10246_/Y gnd _10247_/Y vdd OAI21X1
XFILL_4__13290_ gnd vdd FILL
XFILL_2__10701_ gnd vdd FILL
XSFILL28920x74050 gnd vdd FILL
XFILL_2__8343_ gnd vdd FILL
XFILL_5__11861_ gnd vdd FILL
XSFILL94360x50050 gnd vdd FILL
XFILL_1__12130_ gnd vdd FILL
XFILL_4__9259_ gnd vdd FILL
XFILL_2__11681_ gnd vdd FILL
XFILL_5__13600_ gnd vdd FILL
XFILL_0__12860_ gnd vdd FILL
XFILL_5__10812_ gnd vdd FILL
XFILL_4__12241_ gnd vdd FILL
XFILL_6__11062_ gnd vdd FILL
XFILL_5__14580_ gnd vdd FILL
XFILL_2__13420_ gnd vdd FILL
X_10178_ _10193_/A _6978_/B gnd _10179_/C vdd NAND2X1
XFILL_2__10632_ gnd vdd FILL
XFILL_1__12061_ gnd vdd FILL
XFILL_3__12971_ gnd vdd FILL
XFILL_5__11792_ gnd vdd FILL
XFILL_2__8274_ gnd vdd FILL
XFILL_0__11811_ gnd vdd FILL
XSFILL29000x83050 gnd vdd FILL
XFILL_5__13531_ gnd vdd FILL
XFILL_5__10743_ gnd vdd FILL
XFILL_3__11922_ gnd vdd FILL
XFILL_4__12172_ gnd vdd FILL
XFILL_2__7225_ gnd vdd FILL
XFILL_3__14710_ gnd vdd FILL
XFILL_1__11012_ gnd vdd FILL
XFILL_2__13351_ gnd vdd FILL
XFILL_3__15690_ gnd vdd FILL
X_14986_ _14986_/A _14981_/Y _16035_/B gnd _14986_/Y vdd NAND3X1
XSFILL85000x9050 gnd vdd FILL
XFILL_0__14530_ gnd vdd FILL
XFILL_2__10563_ gnd vdd FILL
XFILL_0__11742_ gnd vdd FILL
XFILL_3_CLKBUF1_insert140 gnd vdd FILL
XFILL_4__11123_ gnd vdd FILL
XFILL_5__16250_ gnd vdd FILL
XFILL_5__13462_ gnd vdd FILL
XFILL_2__12302_ gnd vdd FILL
X_13937_ _14410_/A _13937_/B _14718_/B _15464_/B gnd _13941_/B vdd OAI22X1
XFILL_3_CLKBUF1_insert151 gnd vdd FILL
XFILL_3__14641_ gnd vdd FILL
XFILL_3_CLKBUF1_insert162 gnd vdd FILL
XFILL_1__15820_ gnd vdd FILL
XFILL_2__16070_ gnd vdd FILL
XFILL_5__10674_ gnd vdd FILL
XFILL_3__11853_ gnd vdd FILL
XFILL_2__13282_ gnd vdd FILL
XFILL_0__14461_ gnd vdd FILL
XFILL_5__15201_ gnd vdd FILL
XFILL_3_CLKBUF1_insert173 gnd vdd FILL
XFILL_0__11673_ gnd vdd FILL
XFILL_2__10494_ gnd vdd FILL
XFILL_5__12413_ gnd vdd FILL
XFILL_3_CLKBUF1_insert184 gnd vdd FILL
XFILL_5__8954_ gnd vdd FILL
XFILL_3_CLKBUF1_insert195 gnd vdd FILL
X_13868_ _13867_/Y _13868_/B _14593_/C _13866_/Y gnd _13868_/Y vdd OAI22X1
XFILL_5__16181_ gnd vdd FILL
XFILL_2__15021_ gnd vdd FILL
XFILL_4__15931_ gnd vdd FILL
XFILL_4__11054_ gnd vdd FILL
XFILL_3__10804_ gnd vdd FILL
XFILL_3__14572_ gnd vdd FILL
XFILL_0__16200_ gnd vdd FILL
XFILL_5__13393_ gnd vdd FILL
XFILL_2__12233_ gnd vdd FILL
XFILL_0__10624_ gnd vdd FILL
XFILL_0__13412_ gnd vdd FILL
XFILL_2__7087_ gnd vdd FILL
XFILL_1__15751_ gnd vdd FILL
XFILL_3__11784_ gnd vdd FILL
XFILL_1__12963_ gnd vdd FILL
XFILL_0__14392_ gnd vdd FILL
X_12819_ _12779_/A _12692_/CLK _12692_/R vdd _12819_/D gnd vdd DFFSR
XFILL_6__10915_ gnd vdd FILL
XFILL_1_BUFX2_insert350 gnd vdd FILL
XFILL_4__10005_ gnd vdd FILL
X_15607_ _15603_/Y _15606_/Y gnd _15607_/Y vdd NOR2X1
XFILL_5__15132_ gnd vdd FILL
XSFILL53960x16050 gnd vdd FILL
XFILL_5__8885_ gnd vdd FILL
XFILL_5__12344_ gnd vdd FILL
XFILL_3__16311_ gnd vdd FILL
XFILL_3__13523_ gnd vdd FILL
X_13799_ _8413_/Q gnd _13799_/Y vdd INVX1
XFILL_3__6920_ gnd vdd FILL
XFILL_1__14702_ gnd vdd FILL
XFILL_1_BUFX2_insert361 gnd vdd FILL
XFILL_4__15862_ gnd vdd FILL
XFILL_1_BUFX2_insert372 gnd vdd FILL
XSFILL109480x45050 gnd vdd FILL
XFILL_1__11914_ gnd vdd FILL
XFILL_2__12164_ gnd vdd FILL
XFILL_0__16131_ gnd vdd FILL
XFILL_0__13343_ gnd vdd FILL
XFILL_1__15682_ gnd vdd FILL
XFILL_0__10555_ gnd vdd FILL
XFILL_1_BUFX2_insert383 gnd vdd FILL
XFILL_1__12894_ gnd vdd FILL
XFILL_0__9930_ gnd vdd FILL
XFILL_5__7836_ gnd vdd FILL
XFILL_1_BUFX2_insert394 gnd vdd FILL
XFILL_4__14813_ gnd vdd FILL
XFILL_5__15063_ gnd vdd FILL
X_15538_ _15978_/C _8474_/A _7578_/A _15662_/A gnd _15542_/B vdd AOI22X1
XFILL_3__16242_ gnd vdd FILL
XFILL_3__13454_ gnd vdd FILL
XFILL_5__12275_ gnd vdd FILL
XFILL_2__11115_ gnd vdd FILL
XFILL_1__14633_ gnd vdd FILL
XFILL_3__6851_ gnd vdd FILL
XFILL_4__15793_ gnd vdd FILL
XFILL_3__10666_ gnd vdd FILL
XSFILL54040x25050 gnd vdd FILL
XFILL_0__13274_ gnd vdd FILL
XFILL_2__12095_ gnd vdd FILL
XFILL_0__16062_ gnd vdd FILL
XFILL_1__11845_ gnd vdd FILL
XFILL_5__14014_ gnd vdd FILL
XFILL_0__10486_ gnd vdd FILL
XFILL_3__12405_ gnd vdd FILL
X_15469_ _15841_/C _13956_/D _13959_/D _15813_/C gnd _15469_/Y vdd OAI22X1
XFILL_0__9861_ gnd vdd FILL
X_7420_ _7420_/A gnd _7422_/A vdd INVX1
XFILL_5__11226_ gnd vdd FILL
XFILL_3__16173_ gnd vdd FILL
XFILL_4__14744_ gnd vdd FILL
XFILL_2__15923_ gnd vdd FILL
XFILL_4__11956_ gnd vdd FILL
XFILL_0__15013_ gnd vdd FILL
XFILL_3__13385_ gnd vdd FILL
XFILL_0__12225_ gnd vdd FILL
XFILL_2__11046_ gnd vdd FILL
XFILL_2__7989_ gnd vdd FILL
XFILL_1__14564_ gnd vdd FILL
XFILL_5__9506_ gnd vdd FILL
XFILL_1__11776_ gnd vdd FILL
XFILL_5__11157_ gnd vdd FILL
XFILL_3__15124_ gnd vdd FILL
XFILL_5__7698_ gnd vdd FILL
XFILL_0__9792_ gnd vdd FILL
XFILL_4__10907_ gnd vdd FILL
X_7351_ _7351_/A _7308_/A _7350_/Y gnd _7351_/Y vdd OAI21X1
XFILL_1__16303_ gnd vdd FILL
XFILL_3__8521_ gnd vdd FILL
XFILL_3__12336_ gnd vdd FILL
XFILL_2__9728_ gnd vdd FILL
XSFILL43880x68050 gnd vdd FILL
XFILL_4__14675_ gnd vdd FILL
XFILL_1__13515_ gnd vdd FILL
XFILL_4__11887_ gnd vdd FILL
XFILL_2__15854_ gnd vdd FILL
XFILL_0__12156_ gnd vdd FILL
XFILL_1__14495_ gnd vdd FILL
XFILL_5__10108_ gnd vdd FILL
XFILL_0__8743_ gnd vdd FILL
XSFILL83480x54050 gnd vdd FILL
XFILL_4__16414_ gnd vdd FILL
X_7282_ _7282_/Q _7282_/CLK _9054_/R vdd _7244_/Y gnd vdd DFFSR
XFILL_4__13626_ gnd vdd FILL
XFILL_3__15055_ gnd vdd FILL
XFILL_5__15965_ gnd vdd FILL
XFILL_5__11088_ gnd vdd FILL
XFILL_2__14805_ gnd vdd FILL
XFILL_1__16234_ gnd vdd FILL
XFILL_3__8452_ gnd vdd FILL
XFILL_3__12267_ gnd vdd FILL
XFILL_0__11107_ gnd vdd FILL
XFILL_2__9659_ gnd vdd FILL
XFILL_1__13446_ gnd vdd FILL
XSFILL18680x44050 gnd vdd FILL
XFILL_2__15785_ gnd vdd FILL
XFILL_2__12997_ gnd vdd FILL
XFILL_1__10658_ gnd vdd FILL
XFILL_0__12087_ gnd vdd FILL
XSFILL74200x38050 gnd vdd FILL
X_9021_ _9019_/Y _8961_/B _9021_/C gnd _9069_/D vdd OAI21X1
XFILL_5__10039_ gnd vdd FILL
XFILL_5__9368_ gnd vdd FILL
XFILL_3__14006_ gnd vdd FILL
XSFILL23960x4050 gnd vdd FILL
XFILL_5__14916_ gnd vdd FILL
XFILL_4__16345_ gnd vdd FILL
XFILL_3__11218_ gnd vdd FILL
XFILL_5__15896_ gnd vdd FILL
XFILL_2__14736_ gnd vdd FILL
XFILL_4__10769_ gnd vdd FILL
XFILL_4__13557_ gnd vdd FILL
XSFILL84360x82050 gnd vdd FILL
XFILL_0__15915_ gnd vdd FILL
XFILL_3__8383_ gnd vdd FILL
XFILL_1__16165_ gnd vdd FILL
XFILL_2__11948_ gnd vdd FILL
XFILL_3__12198_ gnd vdd FILL
XFILL_0__11038_ gnd vdd FILL
XFILL_5__8319_ gnd vdd FILL
XFILL_1__13377_ gnd vdd FILL
XFILL_6__8092_ gnd vdd FILL
XFILL_5__9299_ gnd vdd FILL
XFILL_0__7625_ gnd vdd FILL
XSFILL49000x14050 gnd vdd FILL
XFILL_5__14847_ gnd vdd FILL
XFILL_4__12508_ gnd vdd FILL
XFILL_3__7334_ gnd vdd FILL
XFILL_3__11149_ gnd vdd FILL
XFILL_1__15116_ gnd vdd FILL
XFILL_4__16276_ gnd vdd FILL
XFILL_1__12328_ gnd vdd FILL
XFILL_2__14667_ gnd vdd FILL
XFILL_4__13488_ gnd vdd FILL
XFILL_2__11879_ gnd vdd FILL
XFILL_6__7043_ gnd vdd FILL
XFILL_1__16096_ gnd vdd FILL
XFILL_0__15846_ gnd vdd FILL
XFILL112440x8050 gnd vdd FILL
XFILL_4__15227_ gnd vdd FILL
XFILL_0__7556_ gnd vdd FILL
XFILL_2__13618_ gnd vdd FILL
XFILL_4__12439_ gnd vdd FILL
XFILL_2__16406_ gnd vdd FILL
XFILL_5__14778_ gnd vdd FILL
XFILL_3__15957_ gnd vdd FILL
XFILL_1__15047_ gnd vdd FILL
XFILL_2__14598_ gnd vdd FILL
XFILL_1__12259_ gnd vdd FILL
XFILL_0__15777_ gnd vdd FILL
XFILL112360x64050 gnd vdd FILL
XFILL_0__12989_ gnd vdd FILL
XFILL_3__9004_ gnd vdd FILL
X_9923_ _9921_/Y _9937_/A _9923_/C gnd _9967_/D vdd OAI21X1
XFILL_5__13729_ gnd vdd FILL
XFILL_0__7487_ gnd vdd FILL
XFILL_2__16337_ gnd vdd FILL
XFILL_4__15158_ gnd vdd FILL
XFILL_3__14908_ gnd vdd FILL
XFILL_2__13549_ gnd vdd FILL
XFILL_3__7196_ gnd vdd FILL
XFILL_0__14728_ gnd vdd FILL
XFILL_3__15888_ gnd vdd FILL
XFILL_0__9226_ gnd vdd FILL
XFILL_4__14109_ gnd vdd FILL
X_9854_ _9852_/Y _9902_/B _9854_/C gnd _9944_/D vdd OAI21X1
XFILL_3__14839_ gnd vdd FILL
XFILL_4__15089_ gnd vdd FILL
XFILL_2__16268_ gnd vdd FILL
XSFILL79320x71050 gnd vdd FILL
XFILL_0__14659_ gnd vdd FILL
X_8805_ _8805_/Q _7781_/CLK _9566_/R vdd _8741_/Y gnd vdd DFFSR
XSFILL114120x59050 gnd vdd FILL
XSFILL43960x48050 gnd vdd FILL
XFILL_0__9157_ gnd vdd FILL
XFILL_2__15219_ gnd vdd FILL
XFILL_5__16379_ gnd vdd FILL
XFILL_6_BUFX2_insert500 gnd vdd FILL
X_9785_ _9785_/A _9785_/B gnd _9786_/C vdd NAND2X1
XFILL_2__16199_ gnd vdd FILL
XFILL_1__15949_ gnd vdd FILL
XFILL_4__6960_ gnd vdd FILL
X_6997_ _6997_/A _6937_/B _6996_/Y gnd _6997_/Y vdd OAI21X1
XFILL_0__8108_ gnd vdd FILL
XSFILL18760x24050 gnd vdd FILL
XFILL_0__9088_ gnd vdd FILL
X_8736_ _8736_/A gnd _8736_/Y vdd INVX1
XSFILL114520x80050 gnd vdd FILL
XFILL_3__9906_ gnd vdd FILL
XFILL_0__16329_ gnd vdd FILL
XFILL_4__6891_ gnd vdd FILL
XFILL_6_BUFX2_insert577 gnd vdd FILL
XFILL_4__8630_ gnd vdd FILL
X_8667_ _8667_/Q _8679_/CLK _9959_/R vdd _8583_/Y gnd vdd DFFSR
XFILL_1__8852_ gnd vdd FILL
X_7618_ _7570_/A _7490_/B gnd _7619_/C vdd NAND2X1
XSFILL23880x15050 gnd vdd FILL
X_8598_ _8596_/Y _8657_/A _8598_/C gnd _8598_/Y vdd OAI21X1
XFILL_3__9768_ gnd vdd FILL
XFILL_1__7803_ gnd vdd FILL
XSFILL108600x41050 gnd vdd FILL
XFILL_1__8783_ gnd vdd FILL
XSFILL38920x37050 gnd vdd FILL
X_7549_ _7624_/A _7037_/B gnd _7549_/Y vdd NAND2X1
XFILL_3__8719_ gnd vdd FILL
XFILL112440x44050 gnd vdd FILL
XFILL_4__8492_ gnd vdd FILL
XFILL_1__7734_ gnd vdd FILL
XSFILL79800x49050 gnd vdd FILL
XFILL_4__7443_ gnd vdd FILL
X_11150_ _11147_/Y _11150_/B _11150_/C gnd _11150_/Y vdd OAI21X1
X_9219_ _9228_/A _9859_/B gnd _9219_/Y vdd NAND2X1
XFILL_4__7374_ gnd vdd FILL
XFILL_3_BUFX2_insert401 gnd vdd FILL
X_10101_ _10067_/A _9589_/CLK _7413_/R vdd _10101_/D gnd vdd DFFSR
XSFILL3640x77050 gnd vdd FILL
XFILL_1__9404_ gnd vdd FILL
XFILL_3_BUFX2_insert412 gnd vdd FILL
X_11081_ _11081_/A _11081_/B _11081_/C gnd _11086_/A vdd AOI21X1
XFILL_4__9113_ gnd vdd FILL
XFILL_3_BUFX2_insert423 gnd vdd FILL
XFILL_3_BUFX2_insert434 gnd vdd FILL
XFILL_1__7596_ gnd vdd FILL
XFILL_3_BUFX2_insert445 gnd vdd FILL
XFILL_3_BUFX2_insert456 gnd vdd FILL
X_10032_ _10024_/B _6960_/B gnd _10033_/C vdd NAND2X1
XSFILL114600x60050 gnd vdd FILL
XFILL_1__9335_ gnd vdd FILL
XFILL_3_BUFX2_insert467 gnd vdd FILL
XSFILL44120x37050 gnd vdd FILL
XFILL_3_BUFX2_insert478 gnd vdd FILL
XFILL_4__9044_ gnd vdd FILL
XFILL_3_BUFX2_insert489 gnd vdd FILL
X_14840_ _9587_/Q gnd _14840_/Y vdd INVX1
XSFILL69080x41050 gnd vdd FILL
XFILL_1__9266_ gnd vdd FILL
XFILL_1__8217_ gnd vdd FILL
X_14771_ _16127_/B _14506_/A _14718_/C _14771_/D gnd _14771_/Y vdd OAI22X1
X_11983_ _12084_/A gnd _11983_/Y vdd INVX8
X_13722_ _13722_/A _14865_/B _13467_/A _13722_/D gnd _13722_/Y vdd OAI22X1
X_10934_ _12779_/A _10934_/B _10933_/Y gnd _10934_/Y vdd NAND3X1
XFILL_0_BUFX2_insert6 gnd vdd FILL
XFILL_1__8148_ gnd vdd FILL
XFILL_4_CLKBUF1_insert202 gnd vdd FILL
X_13653_ _9090_/A gnd _13653_/Y vdd INVX1
XSFILL49640x68050 gnd vdd FILL
X_16441_ _16393_/A _7269_/CLK _8165_/R vdd _16441_/D gnd vdd DFFSR
XFILL_4_CLKBUF1_insert213 gnd vdd FILL
XFILL_4_CLKBUF1_insert224 gnd vdd FILL
XFILL_5__10390_ gnd vdd FILL
X_10865_ _14774_/D _8433_/CLK _8433_/R vdd _10865_/D gnd vdd DFFSR
XFILL_2__8961_ gnd vdd FILL
XFILL_1__8079_ gnd vdd FILL
XSFILL18760x5050 gnd vdd FILL
XSFILL89240x54050 gnd vdd FILL
X_12604_ vdd memoryOutData[12] gnd _12604_/Y vdd NAND2X1
XFILL_0_BUFX2_insert302 gnd vdd FILL
X_16372_ _15747_/A gnd _16374_/A vdd INVX1
XFILL_4__9877_ gnd vdd FILL
XFILL_3__10520_ gnd vdd FILL
X_13584_ _13584_/A _13583_/Y _14791_/C gnd _13584_/Y vdd AOI21X1
XFILL_0_BUFX2_insert313 gnd vdd FILL
X_10796_ _10796_/A gnd _10798_/A vdd INVX1
XFILL_2__8892_ gnd vdd FILL
XFILL_0_BUFX2_insert324 gnd vdd FILL
X_15323_ _15321_/Y _15322_/Y gnd _15323_/Y vdd NOR2X1
XFILL_5__7621_ gnd vdd FILL
XFILL_4__8828_ gnd vdd FILL
XFILL_0_BUFX2_insert335 gnd vdd FILL
X_12535_ _12343_/A _13175_/CLK _13199_/R vdd _12535_/D gnd vdd DFFSR
XFILL_5__12060_ gnd vdd FILL
XFILL_6__10631_ gnd vdd FILL
XFILL_0_BUFX2_insert346 gnd vdd FILL
XFILL_4__11810_ gnd vdd FILL
XFILL_2__7843_ gnd vdd FILL
XFILL_0_BUFX2_insert357 gnd vdd FILL
XFILL_3__10451_ gnd vdd FILL
XFILL_4__12790_ gnd vdd FILL
XFILL_0_BUFX2_insert368 gnd vdd FILL
XSFILL28920x69050 gnd vdd FILL
XFILL_1__11630_ gnd vdd FILL
XFILL_5__7552_ gnd vdd FILL
XFILL_0_BUFX2_insert379 gnd vdd FILL
XFILL_0__10271_ gnd vdd FILL
XFILL_5__11011_ gnd vdd FILL
XFILL_4__8759_ gnd vdd FILL
X_15254_ _8666_/Q gnd _15255_/C vdd INVX1
X_12466_ _12023_/B gnd _12468_/A vdd INVX1
XFILL_3__13170_ gnd vdd FILL
XFILL_0__12010_ gnd vdd FILL
XFILL_4__11741_ gnd vdd FILL
XFILL_3__10382_ gnd vdd FILL
X_14205_ _14196_/Y _14197_/Y _14205_/C gnd _14216_/A vdd NAND3X1
XFILL_1__11561_ gnd vdd FILL
XFILL_5__7483_ gnd vdd FILL
X_11417_ _11414_/Y _11417_/B _11417_/C gnd _11417_/Y vdd AOI21X1
X_15185_ _15185_/A _15185_/B gnd _15208_/A vdd NOR2X1
XFILL_3__12121_ gnd vdd FILL
XFILL_1__13300_ gnd vdd FILL
XFILL_4__14460_ gnd vdd FILL
X_12397_ _12553_/Q gnd _12397_/Y vdd INVX1
XFILL_4__11672_ gnd vdd FILL
XFILL_2__9513_ gnd vdd FILL
XFILL_1__10512_ gnd vdd FILL
XFILL_2__12851_ gnd vdd FILL
XFILL_6__15020_ gnd vdd FILL
XFILL_5__9222_ gnd vdd FILL
XFILL_1__14280_ gnd vdd FILL
X_14136_ _7840_/A gnd _14138_/A vdd INVX1
XFILL_1__11492_ gnd vdd FILL
XFILL_4__10623_ gnd vdd FILL
XFILL_4__13411_ gnd vdd FILL
XFILL_5__15750_ gnd vdd FILL
X_11348_ _11348_/A _11226_/B _11347_/Y gnd _11348_/Y vdd OAI21X1
XFILL_5__12962_ gnd vdd FILL
XFILL_3__12052_ gnd vdd FILL
XSFILL104360x30050 gnd vdd FILL
XFILL_2__11802_ gnd vdd FILL
XFILL_1__13231_ gnd vdd FILL
XFILL_2__15570_ gnd vdd FILL
XFILL_4__14391_ gnd vdd FILL
XFILL_2__12782_ gnd vdd FILL
XFILL_1__10443_ gnd vdd FILL
XFILL_5__9153_ gnd vdd FILL
XFILL_5__14701_ gnd vdd FILL
XFILL_0__13961_ gnd vdd FILL
XFILL_5_BUFX2_insert1003 gnd vdd FILL
XFILL_5__11913_ gnd vdd FILL
X_14067_ _8802_/Q gnd _14067_/Y vdd INVX1
XFILL_4_BUFX2_insert290 gnd vdd FILL
XFILL_4__16130_ gnd vdd FILL
XSFILL74280x12050 gnd vdd FILL
XFILL_3__11003_ gnd vdd FILL
XFILL_4__13342_ gnd vdd FILL
XFILL_5__15681_ gnd vdd FILL
XFILL_5_BUFX2_insert1014 gnd vdd FILL
XFILL_2__14521_ gnd vdd FILL
XFILL_4__10554_ gnd vdd FILL
X_11279_ _12270_/Y _12156_/Y gnd _11279_/Y vdd NOR2X1
XFILL_5_BUFX2_insert1025 gnd vdd FILL
XFILL_0__15700_ gnd vdd FILL
XFILL_5__8104_ gnd vdd FILL
XFILL_5__12893_ gnd vdd FILL
XFILL_2__9375_ gnd vdd FILL
XFILL_2__11733_ gnd vdd FILL
XFILL_0__12912_ gnd vdd FILL
XFILL_1__13162_ gnd vdd FILL
XFILL_1__10374_ gnd vdd FILL
XFILL_5_BUFX2_insert1036 gnd vdd FILL
X_13018_ vdd _13018_/B gnd _13019_/C vdd NAND2X1
XFILL_5__9084_ gnd vdd FILL
XFILL_5__14632_ gnd vdd FILL
XFILL_5_BUFX2_insert1047 gnd vdd FILL
XSFILL89320x34050 gnd vdd FILL
XFILL_0__13892_ gnd vdd FILL
XFILL_4__13273_ gnd vdd FILL
XSFILL59080x73050 gnd vdd FILL
XFILL_0__8390_ gnd vdd FILL
XFILL_3__15811_ gnd vdd FILL
XFILL_5_BUFX2_insert1058 gnd vdd FILL
XFILL_2__8326_ gnd vdd FILL
XFILL_4__16061_ gnd vdd FILL
XFILL_5__11844_ gnd vdd FILL
XFILL_2__14452_ gnd vdd FILL
XFILL_1__12113_ gnd vdd FILL
XFILL_5_BUFX2_insert1069 gnd vdd FILL
XFILL_0__15631_ gnd vdd FILL
XFILL_2__11664_ gnd vdd FILL
XFILL_0__12843_ gnd vdd FILL
XFILL_1__13093_ gnd vdd FILL
XFILL_4__15012_ gnd vdd FILL
XFILL_3_BUFX2_insert990 gnd vdd FILL
XFILL_0__7341_ gnd vdd FILL
XFILL_4__12224_ gnd vdd FILL
XFILL_5__14563_ gnd vdd FILL
XFILL_2__13403_ gnd vdd FILL
XFILL_3__7050_ gnd vdd FILL
XFILL_2__10615_ gnd vdd FILL
XFILL_2__8257_ gnd vdd FILL
XFILL_3__15742_ gnd vdd FILL
XFILL_5__11775_ gnd vdd FILL
XFILL_1__12044_ gnd vdd FILL
XFILL_2__14383_ gnd vdd FILL
XFILL_3__12954_ gnd vdd FILL
XFILL_0__15562_ gnd vdd FILL
XFILL_5__16302_ gnd vdd FILL
XFILL_2__11595_ gnd vdd FILL
XFILL_0__12774_ gnd vdd FILL
XFILL_5__13514_ gnd vdd FILL
X_6920_ _7004_/Q gnd _6920_/Y vdd INVX1
XFILL_2__7208_ gnd vdd FILL
XFILL_2__16122_ gnd vdd FILL
XFILL_6__15853_ gnd vdd FILL
XFILL_4__12155_ gnd vdd FILL
XFILL_2__13334_ gnd vdd FILL
XFILL_5__14494_ gnd vdd FILL
XFILL_3__11905_ gnd vdd FILL
X_14969_ _10067_/A gnd _14969_/Y vdd INVX1
XSFILL94440x25050 gnd vdd FILL
XFILL_3__15673_ gnd vdd FILL
XFILL_0__14513_ gnd vdd FILL
XFILL_2__8188_ gnd vdd FILL
XFILL_3__12885_ gnd vdd FILL
XFILL_2__10546_ gnd vdd FILL
XFILL_0__11725_ gnd vdd FILL
XFILL_0__9011_ gnd vdd FILL
XFILL_5__16233_ gnd vdd FILL
XFILL_4__11106_ gnd vdd FILL
XFILL_0__15493_ gnd vdd FILL
XFILL_5__9986_ gnd vdd FILL
XFILL_5__13445_ gnd vdd FILL
XFILL_3__14624_ gnd vdd FILL
XFILL_6__12996_ gnd vdd FILL
XFILL_4__12086_ gnd vdd FILL
XFILL_5__10657_ gnd vdd FILL
X_6851_ _6851_/A gnd memoryAddress[13] vdd BUFX2
XFILL_1__15803_ gnd vdd FILL
XFILL_2__16053_ gnd vdd FILL
XFILL_3_BUFX2_insert1040 gnd vdd FILL
XFILL_3__11836_ gnd vdd FILL
XFILL_2__13265_ gnd vdd FILL
XFILL_3_BUFX2_insert1051 gnd vdd FILL
XFILL_0__14444_ gnd vdd FILL
XFILL_3_BUFX2_insert1062 gnd vdd FILL
XFILL_1__13995_ gnd vdd FILL
XFILL_6__7730_ gnd vdd FILL
XFILL_0__11656_ gnd vdd FILL
XFILL_4__15914_ gnd vdd FILL
XFILL_3_BUFX2_insert1073 gnd vdd FILL
XFILL_6__11947_ gnd vdd FILL
XFILL_4__11037_ gnd vdd FILL
XFILL_2__15004_ gnd vdd FILL
XFILL_5__16164_ gnd vdd FILL
XFILL_3_BUFX2_insert1084 gnd vdd FILL
XFILL_5__13376_ gnd vdd FILL
X_9570_ _9570_/Q _7010_/CLK _7413_/R vdd _9570_/D gnd vdd DFFSR
XFILL_2__12216_ gnd vdd FILL
XFILL_3__14555_ gnd vdd FILL
XFILL_3__11767_ gnd vdd FILL
XFILL_1__15734_ gnd vdd FILL
XFILL_3__7952_ gnd vdd FILL
XSFILL18680x39050 gnd vdd FILL
XFILL_0__14375_ gnd vdd FILL
XFILL_0__11587_ gnd vdd FILL
XSFILL104440x10050 gnd vdd FILL
XFILL_5__15115_ gnd vdd FILL
XFILL_5__8868_ gnd vdd FILL
X_8521_ _8519_/Y _8440_/B _8521_/C gnd _8561_/D vdd OAI21X1
XFILL_5__12327_ gnd vdd FILL
XFILL_5__16095_ gnd vdd FILL
XFILL_4__15845_ gnd vdd FILL
XFILL_3__13506_ gnd vdd FILL
XFILL_3__14486_ gnd vdd FILL
XFILL_3__6903_ gnd vdd FILL
XSFILL33720x42050 gnd vdd FILL
XFILL_0__16114_ gnd vdd FILL
XFILL_2__12147_ gnd vdd FILL
XFILL_0__13326_ gnd vdd FILL
XFILL_1__15665_ gnd vdd FILL
XFILL_5_BUFX2_insert507 gnd vdd FILL
XFILL_3__7883_ gnd vdd FILL
XFILL_6__9400_ gnd vdd FILL
XFILL_3__11698_ gnd vdd FILL
XFILL_0__10538_ gnd vdd FILL
XFILL_5_BUFX2_insert518 gnd vdd FILL
XFILL_5__7819_ gnd vdd FILL
XFILL_1__12877_ gnd vdd FILL
XFILL_5__15046_ gnd vdd FILL
XFILL_0__9913_ gnd vdd FILL
XFILL_5_BUFX2_insert529 gnd vdd FILL
XFILL_3__16225_ gnd vdd FILL
X_8452_ _8452_/A _8460_/A _8451_/Y gnd _8452_/Y vdd OAI21X1
XFILL_3__13437_ gnd vdd FILL
XFILL_5__12258_ gnd vdd FILL
XFILL_1__14616_ gnd vdd FILL
XFILL_3__10649_ gnd vdd FILL
XFILL_4__15776_ gnd vdd FILL
XFILL_3__9622_ gnd vdd FILL
XFILL_0__16045_ gnd vdd FILL
XFILL_2__12078_ gnd vdd FILL
XFILL_4__12988_ gnd vdd FILL
XSFILL89400x14050 gnd vdd FILL
XFILL_1__11828_ gnd vdd FILL
XFILL_0__13257_ gnd vdd FILL
XSFILL59160x53050 gnd vdd FILL
XFILL_1__15596_ gnd vdd FILL
X_7403_ _7403_/Q _7147_/CLK _7531_/R vdd _7351_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert880 gnd vdd FILL
XFILL_5__11209_ gnd vdd FILL
XFILL_0_BUFX2_insert891 gnd vdd FILL
XFILL_4__14727_ gnd vdd FILL
XFILL_2__15906_ gnd vdd FILL
X_8383_ _8321_/B _7359_/B gnd _8384_/C vdd NAND2X1
XFILL_5__12189_ gnd vdd FILL
XFILL_3__13368_ gnd vdd FILL
XFILL_4__11939_ gnd vdd FILL
XFILL_2__11029_ gnd vdd FILL
XFILL_3__16156_ gnd vdd FILL
XFILL_1__14547_ gnd vdd FILL
XFILL_0__12208_ gnd vdd FILL
XFILL_3__9553_ gnd vdd FILL
XFILL_1__11759_ gnd vdd FILL
XFILL_3_BUFX2_insert40 gnd vdd FILL
X_7334_ _7398_/Q gnd _7334_/Y vdd INVX1
XFILL112360x59050 gnd vdd FILL
XFILL_0__9775_ gnd vdd FILL
XFILL_3__12319_ gnd vdd FILL
XFILL_3__15107_ gnd vdd FILL
XFILL_3_BUFX2_insert51 gnd vdd FILL
XFILL_0__6987_ gnd vdd FILL
XFILL_3__8504_ gnd vdd FILL
XFILL_4__14658_ gnd vdd FILL
XFILL_3__16087_ gnd vdd FILL
XFILL_3__13299_ gnd vdd FILL
XFILL_3__9484_ gnd vdd FILL
XFILL_0__12139_ gnd vdd FILL
XFILL_2__15837_ gnd vdd FILL
XFILL_1__14478_ gnd vdd FILL
XFILL_3_BUFX2_insert62 gnd vdd FILL
XFILL_3_BUFX2_insert73 gnd vdd FILL
XFILL_0__8726_ gnd vdd FILL
XFILL_4__13609_ gnd vdd FILL
XFILL_3_BUFX2_insert84 gnd vdd FILL
XFILL_5__15948_ gnd vdd FILL
XFILL_1__16217_ gnd vdd FILL
XFILL_3_BUFX2_insert95 gnd vdd FILL
XFILL_3__15038_ gnd vdd FILL
X_7265_ _7191_/A _9953_/CLK _7276_/R vdd _7265_/D gnd vdd DFFSR
XFILL_4__14589_ gnd vdd FILL
XFILL_1__13429_ gnd vdd FILL
XSFILL24280x60050 gnd vdd FILL
XFILL_2__15768_ gnd vdd FILL
X_9004_ _9004_/A gnd _9004_/Y vdd INVX1
XSFILL79320x66050 gnd vdd FILL
XFILL_1__7450_ gnd vdd FILL
XFILL_4__16328_ gnd vdd FILL
XFILL_0__8657_ gnd vdd FILL
X_7196_ _7196_/A _7207_/A _7196_/C gnd _7266_/D vdd OAI21X1
XFILL_5__15879_ gnd vdd FILL
XFILL_2__14719_ gnd vdd FILL
XFILL_3__8366_ gnd vdd FILL
XFILL_1__16148_ gnd vdd FILL
XFILL_2__15699_ gnd vdd FILL
XFILL_0__7608_ gnd vdd FILL
XFILL_0__8588_ gnd vdd FILL
XFILL_1__7381_ gnd vdd FILL
XFILL_3__7317_ gnd vdd FILL
XSFILL18760x19050 gnd vdd FILL
XFILL_4__16259_ gnd vdd FILL
XSFILL114520x75050 gnd vdd FILL
XSFILL8600x29050 gnd vdd FILL
XFILL_0__15829_ gnd vdd FILL
XFILL_4__7090_ gnd vdd FILL
XFILL_1__16079_ gnd vdd FILL
XFILL_2_BUFX2_insert408 gnd vdd FILL
XFILL_1__9120_ gnd vdd FILL
XFILL_2_BUFX2_insert419 gnd vdd FILL
XFILL_3__7248_ gnd vdd FILL
XSFILL79480x4050 gnd vdd FILL
X_9906_ _9906_/A gnd _9908_/A vdd INVX1
XFILL_3__7179_ gnd vdd FILL
XFILL_1__8002_ gnd vdd FILL
XFILL_0__9209_ gnd vdd FILL
X_9837_ _9837_/Q _8038_/CLK _8038_/R vdd _9789_/Y gnd vdd DFFSR
XFILL_4__9800_ gnd vdd FILL
XFILL112440x39050 gnd vdd FILL
XFILL_4__7992_ gnd vdd FILL
X_9768_ _9768_/A _9789_/B _9767_/Y gnd _9768_/Y vdd OAI21X1
XSFILL23720x74050 gnd vdd FILL
XFILL_6_BUFX2_insert341 gnd vdd FILL
XFILL_4__9731_ gnd vdd FILL
XFILL_4__6943_ gnd vdd FILL
XBUFX2_insert407 _10920_/Y gnd _12368_/A vdd BUFX2
X_10650_ _15566_/A gnd _10650_/Y vdd INVX1
XFILL_6_BUFX2_insert352 gnd vdd FILL
X_8719_ _8740_/A _8719_/B gnd _8720_/C vdd NAND2X1
XFILL_6__7859_ gnd vdd FILL
XBUFX2_insert418 _15050_/Y gnd _15801_/A vdd BUFX2
XBUFX2_insert429 _15047_/Y gnd _15351_/D vdd BUFX2
XSFILL24360x40050 gnd vdd FILL
X_9699_ _9699_/Q _7651_/CLK _7011_/R vdd _9699_/D gnd vdd DFFSR
XFILL_4__9662_ gnd vdd FILL
XFILL_4__6874_ gnd vdd FILL
XFILL_1__8904_ gnd vdd FILL
X_10581_ _10579_/Y _10581_/B _10580_/Y gnd _10581_/Y vdd OAI21X1
XFILL_4__8613_ gnd vdd FILL
XFILL_1__9884_ gnd vdd FILL
X_12320_ _12312_/A _12340_/B _12312_/C gnd _12320_/Y vdd NAND3X1
XFILL_6__9529_ gnd vdd FILL
XFILL_4__9593_ gnd vdd FILL
XFILL_1__8835_ gnd vdd FILL
X_12251_ _12255_/A gnd _12255_/C gnd _12254_/A vdd NAND3X1
XSFILL115240x21050 gnd vdd FILL
XFILL_1__8766_ gnd vdd FILL
XSFILL69080x36050 gnd vdd FILL
XFILL_4__8475_ gnd vdd FILL
X_11202_ _12201_/Y _12330_/Y gnd _11202_/Y vdd AND2X2
XFILL_1__7717_ gnd vdd FILL
X_12182_ _12201_/B _12889_/A gnd _12183_/C vdd NAND2X1
XFILL_4__7426_ gnd vdd FILL
XFILL_2__7490_ gnd vdd FILL
XFILL_1__8697_ gnd vdd FILL
XSFILL104280x45050 gnd vdd FILL
X_11133_ _12168_/Y _11150_/B gnd _11133_/Y vdd NOR2X1
XFILL_4__7357_ gnd vdd FILL
XFILL_3_BUFX2_insert231 gnd vdd FILL
XSFILL73960x82050 gnd vdd FILL
XFILL_3_BUFX2_insert242 gnd vdd FILL
X_15941_ _9836_/Q _15390_/B _15940_/Y gnd _15941_/Y vdd AOI21X1
X_11064_ _12153_/Y gnd _11064_/Y vdd INVX2
XFILL_3_BUFX2_insert253 gnd vdd FILL
XFILL_2__9160_ gnd vdd FILL
XFILL_1__7579_ gnd vdd FILL
XFILL_3_BUFX2_insert264 gnd vdd FILL
XSFILL89240x49050 gnd vdd FILL
XFILL_3_BUFX2_insert275 gnd vdd FILL
XFILL112120x21050 gnd vdd FILL
XFILL_3_BUFX2_insert286 gnd vdd FILL
XFILL_4__7288_ gnd vdd FILL
X_10015_ _10015_/A _10066_/B _10014_/Y gnd _10015_/Y vdd OAI21X1
XFILL_2__8111_ gnd vdd FILL
X_15872_ _9394_/A _15945_/C _16148_/C gnd _15873_/C vdd NAND3X1
XFILL_4__10270_ gnd vdd FILL
XFILL_3_BUFX2_insert297 gnd vdd FILL
XFILL_2__9091_ gnd vdd FILL
XFILL_4__9027_ gnd vdd FILL
XFILL_2_BUFX2_insert920 gnd vdd FILL
XFILL_2_BUFX2_insert931 gnd vdd FILL
X_14823_ _10442_/A _14389_/B _13853_/C _6986_/A gnd _14832_/A vdd AOI22X1
XFILL_2_BUFX2_insert942 gnd vdd FILL
XFILL_1__9249_ gnd vdd FILL
XFILL_2__10400_ gnd vdd FILL
XFILL_2_BUFX2_insert953 gnd vdd FILL
XFILL_5__11560_ gnd vdd FILL
XFILL_2_BUFX2_insert964 gnd vdd FILL
XFILL_2__11380_ gnd vdd FILL
XFILL_2_BUFX2_insert975 gnd vdd FILL
XFILL_5__10511_ gnd vdd FILL
XFILL_2_BUFX2_insert986 gnd vdd FILL
X_11966_ _11955_/B _12091_/B gnd _11967_/C vdd NAND2X1
XFILL_2_BUFX2_insert997 gnd vdd FILL
X_14754_ _14746_/Y _14754_/B _14754_/C gnd _14765_/A vdd NAND3X1
XSFILL8520x1050 gnd vdd FILL
XFILL_5__11491_ gnd vdd FILL
XFILL_0__11510_ gnd vdd FILL
XFILL_0__12490_ gnd vdd FILL
XFILL_5__13230_ gnd vdd FILL
X_10917_ _10920_/B _10944_/B gnd _16450_/C vdd NOR2X1
XFILL_5__9771_ gnd vdd FILL
X_13705_ _13705_/A _13705_/B gnd _13705_/Y vdd NOR2X1
XSFILL69160x16050 gnd vdd FILL
XFILL_5__10442_ gnd vdd FILL
X_14685_ _8001_/A gnd _14686_/D vdd INVX1
XFILL_3__11621_ gnd vdd FILL
XFILL_5__6983_ gnd vdd FILL
X_11897_ _11975_/A _12352_/A gnd _11897_/Y vdd NAND2X1
XFILL_4__13960_ gnd vdd FILL
XFILL_2__10262_ gnd vdd FILL
XFILL_0__11441_ gnd vdd FILL
XFILL_1__13780_ gnd vdd FILL
XFILL_2__9993_ gnd vdd FILL
XFILL_5__8722_ gnd vdd FILL
XFILL_4__9929_ gnd vdd FILL
X_16424_ _16342_/A _7147_/CLK _7133_/R vdd _16424_/D gnd vdd DFFSR
X_13636_ _13636_/A _13636_/B gnd _13637_/B vdd NOR2X1
XFILL_1__10992_ gnd vdd FILL
XFILL_6__11732_ gnd vdd FILL
XFILL_4__12911_ gnd vdd FILL
XFILL_2__12001_ gnd vdd FILL
XFILL_5__13161_ gnd vdd FILL
XFILL_3__14340_ gnd vdd FILL
XFILL_5__10373_ gnd vdd FILL
X_10848_ _10848_/Q _8433_/CLK _7921_/R vdd _10774_/Y gnd vdd DFFSR
XFILL_3__11552_ gnd vdd FILL
XFILL_1__12731_ gnd vdd FILL
XFILL_0_BUFX2_insert110 gnd vdd FILL
XFILL_4__13891_ gnd vdd FILL
XFILL_0__14160_ gnd vdd FILL
XSFILL104520x8050 gnd vdd FILL
XFILL_2__10193_ gnd vdd FILL
XBUFX2_insert930 _12435_/Y gnd _8273_/B vdd BUFX2
XFILL_0__11372_ gnd vdd FILL
XFILL_5__8653_ gnd vdd FILL
XFILL_5__12112_ gnd vdd FILL
XBUFX2_insert941 _12426_/Y gnd _7752_/B vdd BUFX2
XFILL_4__15630_ gnd vdd FILL
X_16355_ gnd gnd gnd _16356_/C vdd NAND2X1
XFILL_3__10503_ gnd vdd FILL
X_13567_ _13567_/A _13567_/B gnd _13571_/C vdd NOR2X1
XFILL_4__12842_ gnd vdd FILL
X_10779_ _10762_/B _8987_/B gnd _10780_/C vdd NAND2X1
XFILL_5__13092_ gnd vdd FILL
XBUFX2_insert952 _13365_/Y gnd _10773_/A vdd BUFX2
XFILL_3__14271_ gnd vdd FILL
XBUFX2_insert963 _13361_/Y gnd _10405_/B vdd BUFX2
XFILL_0__13111_ gnd vdd FILL
XFILL_1__15450_ gnd vdd FILL
XFILL_3__11483_ gnd vdd FILL
XFILL_0__10323_ gnd vdd FILL
XFILL_1__12662_ gnd vdd FILL
XSFILL8040x66050 gnd vdd FILL
XBUFX2_insert974 _16451_/Y gnd _13153_/B vdd BUFX2
XFILL_2__8875_ gnd vdd FILL
XFILL_5__7604_ gnd vdd FILL
XFILL_0__14091_ gnd vdd FILL
X_15306_ _15384_/A _13774_/Y _13777_/Y _15384_/D gnd _15308_/B vdd OAI22X1
X_12518_ vdd _12093_/A gnd _12518_/Y vdd NAND2X1
XFILL_0__6910_ gnd vdd FILL
XBUFX2_insert985 _13351_/Y gnd _10054_/B vdd BUFX2
XFILL_3__13222_ gnd vdd FILL
XFILL_5__8584_ gnd vdd FILL
XFILL_3__16010_ gnd vdd FILL
XFILL_5__12043_ gnd vdd FILL
X_16286_ _16285_/Y _16286_/B gnd _16296_/B vdd NAND2X1
XBUFX2_insert996 _14998_/Y gnd _14999_/A vdd BUFX2
XSFILL59080x68050 gnd vdd FILL
XFILL_4__15561_ gnd vdd FILL
XFILL_1__14401_ gnd vdd FILL
XFILL_3__10434_ gnd vdd FILL
XFILL_6__11594_ gnd vdd FILL
X_13498_ _13496_/Y _14778_/B _14887_/B _13497_/Y gnd _13498_/Y vdd OAI22X1
XFILL_0__7890_ gnd vdd FILL
XFILL_4__12773_ gnd vdd FILL
XFILL_1__11613_ gnd vdd FILL
XFILL_2__13952_ gnd vdd FILL
XFILL_2__7826_ gnd vdd FILL
XFILL_0__13042_ gnd vdd FILL
XFILL_0__10254_ gnd vdd FILL
XFILL_1__15381_ gnd vdd FILL
XFILL_1__12593_ gnd vdd FILL
XSFILL99480x73050 gnd vdd FILL
XFILL_0__6841_ gnd vdd FILL
X_12449_ vdd _12449_/B gnd _12449_/Y vdd NAND2X1
X_15237_ _15237_/A gnd _15239_/A vdd INVX1
XSFILL49320x45050 gnd vdd FILL
XFILL_4__14512_ gnd vdd FILL
XFILL_3__13153_ gnd vdd FILL
XFILL_2__12903_ gnd vdd FILL
XFILL_4__11724_ gnd vdd FILL
XFILL_2__7757_ gnd vdd FILL
XFILL_1__14332_ gnd vdd FILL
XFILL_3__10365_ gnd vdd FILL
XFILL_4__15492_ gnd vdd FILL
XFILL_2__13883_ gnd vdd FILL
XFILL_1__11544_ gnd vdd FILL
XFILL_5__15802_ gnd vdd FILL
XFILL_0__10185_ gnd vdd FILL
XFILL_5__7466_ gnd vdd FILL
X_15168_ _9177_/Q gnd _15169_/C vdd INVX1
XFILL_3__12104_ gnd vdd FILL
XFILL_4__14443_ gnd vdd FILL
XFILL_2__12834_ gnd vdd FILL
XFILL_2__15622_ gnd vdd FILL
XFILL_5__13994_ gnd vdd FILL
XFILL_3__13084_ gnd vdd FILL
XFILL_4__11655_ gnd vdd FILL
XFILL_2__7688_ gnd vdd FILL
XFILL_1__14263_ gnd vdd FILL
XFILL_3__10296_ gnd vdd FILL
XFILL_0__8511_ gnd vdd FILL
XFILL_1__11475_ gnd vdd FILL
X_14119_ _14115_/Y _14119_/B gnd _14120_/C vdd NOR2X1
X_7050_ _7048_/Y _7068_/B _7050_/C gnd _7050_/Y vdd OAI21X1
XFILL_0__14993_ gnd vdd FILL
XFILL_5__15733_ gnd vdd FILL
XFILL_1__16002_ gnd vdd FILL
XFILL_3__12035_ gnd vdd FILL
XFILL_3__8220_ gnd vdd FILL
XFILL_0__9491_ gnd vdd FILL
X_15099_ _8407_/Q _15978_/B _15978_/C _8441_/A gnd _15099_/Y vdd AOI22X1
XFILL_1__13214_ gnd vdd FILL
XFILL_2__15553_ gnd vdd FILL
XFILL_2__9427_ gnd vdd FILL
XFILL_4__14374_ gnd vdd FILL
XFILL_4__11586_ gnd vdd FILL
XFILL_2__12765_ gnd vdd FILL
XFILL_1__10426_ gnd vdd FILL
XFILL_1__14194_ gnd vdd FILL
XFILL_5__9136_ gnd vdd FILL
XSFILL94280x6050 gnd vdd FILL
XFILL_0__13944_ gnd vdd FILL
XFILL_4__16113_ gnd vdd FILL
XFILL_0__8442_ gnd vdd FILL
XFILL_4__13325_ gnd vdd FILL
XFILL_5__15664_ gnd vdd FILL
XFILL_2__9358_ gnd vdd FILL
XFILL_2__14504_ gnd vdd FILL
XFILL_5__12876_ gnd vdd FILL
XFILL_2__11716_ gnd vdd FILL
XFILL_4__10537_ gnd vdd FILL
XFILL_1__13145_ gnd vdd FILL
XFILL_2__15484_ gnd vdd FILL
XFILL_2__12696_ gnd vdd FILL
XFILL_0__13875_ gnd vdd FILL
XFILL_5__14615_ gnd vdd FILL
XFILL_0__8373_ gnd vdd FILL
XFILL_3__7102_ gnd vdd FILL
XFILL_4__16044_ gnd vdd FILL
XFILL_5__11827_ gnd vdd FILL
XFILL_4__13256_ gnd vdd FILL
XFILL_2__14435_ gnd vdd FILL
XFILL_5__15595_ gnd vdd FILL
XFILL_0__15614_ gnd vdd FILL
XFILL_2__9289_ gnd vdd FILL
XFILL_2__11647_ gnd vdd FILL
XFILL_3__8082_ gnd vdd FILL
XFILL_3__13986_ gnd vdd FILL
XFILL_1__10288_ gnd vdd FILL
XFILL_0__12826_ gnd vdd FILL
XFILL_5__8018_ gnd vdd FILL
XFILL_6__15905_ gnd vdd FILL
XFILL_0__7324_ gnd vdd FILL
XFILL_5__14546_ gnd vdd FILL
XFILL_4__12207_ gnd vdd FILL
XSFILL43880x81050 gnd vdd FILL
X_7952_ _7950_/Y _7937_/B _7952_/C gnd _7952_/Y vdd OAI21X1
XFILL_3__15725_ gnd vdd FILL
XFILL_3__7033_ gnd vdd FILL
XFILL_5__11758_ gnd vdd FILL
XFILL_1__12027_ gnd vdd FILL
XFILL_2__14366_ gnd vdd FILL
XFILL_4__10399_ gnd vdd FILL
XFILL_0__15545_ gnd vdd FILL
XFILL_2__11578_ gnd vdd FILL
XFILL_0__12757_ gnd vdd FILL
XSFILL59160x48050 gnd vdd FILL
X_6903_ _6903_/A _6948_/A gnd _6904_/C vdd NAND2X1
XFILL_5__10709_ gnd vdd FILL
XFILL_2__13317_ gnd vdd FILL
XFILL_5__14477_ gnd vdd FILL
XFILL_4__12138_ gnd vdd FILL
XFILL_2__16105_ gnd vdd FILL
XFILL_3__15656_ gnd vdd FILL
X_7883_ _7824_/B _7883_/B gnd _7884_/C vdd NAND2X1
XFILL_2__10529_ gnd vdd FILL
XFILL_5__11689_ gnd vdd FILL
XFILL_3__12868_ gnd vdd FILL
XSFILL74200x51050 gnd vdd FILL
XFILL_0__11708_ gnd vdd FILL
XFILL_2__14297_ gnd vdd FILL
XFILL_5__16216_ gnd vdd FILL
XFILL_0__15476_ gnd vdd FILL
XFILL_5__13428_ gnd vdd FILL
X_9622_ _9622_/A _9652_/B _9621_/Y gnd _9622_/Y vdd OAI21X1
XFILL_3__14607_ gnd vdd FILL
XFILL_2__16036_ gnd vdd FILL
XFILL_4__12069_ gnd vdd FILL
XFILL_0__7186_ gnd vdd FILL
XFILL_2__13248_ gnd vdd FILL
XFILL_3__11819_ gnd vdd FILL
XFILL_3__15587_ gnd vdd FILL
XFILL_0__14427_ gnd vdd FILL
XFILL_3__8984_ gnd vdd FILL
XFILL_1__13978_ gnd vdd FILL
XFILL_0__11639_ gnd vdd FILL
XSFILL64280x39050 gnd vdd FILL
XFILL_6__14718_ gnd vdd FILL
XFILL_5__16147_ gnd vdd FILL
XFILL_5__13359_ gnd vdd FILL
X_9553_ _9554_/B _8401_/B gnd _9553_/Y vdd NAND2X1
XSFILL109400x79050 gnd vdd FILL
XFILL_3__14538_ gnd vdd FILL
XFILL_3__7935_ gnd vdd FILL
XFILL_1__15717_ gnd vdd FILL
XFILL_0__14358_ gnd vdd FILL
XSFILL8680x7050 gnd vdd FILL
X_8504_ _8556_/Q gnd _8504_/Y vdd INVX1
XFILL_5_BUFX2_insert304 gnd vdd FILL
XFILL_1__6950_ gnd vdd FILL
XFILL_4__15828_ gnd vdd FILL
XSFILL54040x9050 gnd vdd FILL
XFILL_5__16078_ gnd vdd FILL
XFILL_5_BUFX2_insert315 gnd vdd FILL
X_9484_ _9551_/B _9100_/B gnd _9484_/Y vdd NAND2X1
XFILL_5_BUFX2_insert326 gnd vdd FILL
XSFILL64680x60050 gnd vdd FILL
XSFILL89400x7050 gnd vdd FILL
XFILL_0__13309_ gnd vdd FILL
XFILL_3__14469_ gnd vdd FILL
XBUFX2_insert16 _14989_/Y gnd _16208_/B vdd BUFX2
XFILL_1__15648_ gnd vdd FILL
XFILL_5_BUFX2_insert337 gnd vdd FILL
XSFILL38840x70050 gnd vdd FILL
XFILL_3__7866_ gnd vdd FILL
XBUFX2_insert27 _13320_/Y gnd _8469_/A vdd BUFX2
XFILL_5__15029_ gnd vdd FILL
XFILL_5_BUFX2_insert348 gnd vdd FILL
XFILL_0__14289_ gnd vdd FILL
X_8435_ _8435_/Q _8429_/CLK _9203_/R vdd _8399_/Y gnd vdd DFFSR
XFILL_3__16208_ gnd vdd FILL
XFILL_6__7575_ gnd vdd FILL
XFILL_5_BUFX2_insert359 gnd vdd FILL
XBUFX2_insert38 _13265_/Y gnd _6955_/B vdd BUFX2
XBUFX2_insert49 _13381_/Y gnd _13680_/B vdd BUFX2
XFILL_1__6881_ gnd vdd FILL
XFILL_4__15759_ gnd vdd FILL
XFILL_3__9605_ gnd vdd FILL
XSFILL2680x82050 gnd vdd FILL
XFILL_0__16028_ gnd vdd FILL
XSFILL95000x30050 gnd vdd FILL
XFILL_1__15579_ gnd vdd FILL
XFILL_1__8620_ gnd vdd FILL
XFILL_6__16319_ gnd vdd FILL
X_8366_ _8364_/Y _8365_/A _8366_/C gnd _8366_/Y vdd OAI21X1
XSFILL33800x17050 gnd vdd FILL
XFILL_3__16139_ gnd vdd FILL
XFILL_3__9536_ gnd vdd FILL
XSFILL43960x61050 gnd vdd FILL
XFILL_6__9245_ gnd vdd FILL
X_7317_ _7354_/B _7317_/B gnd _7317_/Y vdd NAND2X1
XFILL_0__9758_ gnd vdd FILL
XFILL_4__8260_ gnd vdd FILL
XSFILL59240x28050 gnd vdd FILL
X_8297_ _8297_/Q _8297_/CLK _7796_/R vdd _8297_/D gnd vdd DFFSR
XFILL_3__9467_ gnd vdd FILL
XFILL_1__7502_ gnd vdd FILL
XFILL_0__8709_ gnd vdd FILL
XFILL_1__8482_ gnd vdd FILL
X_7248_ _7248_/A gnd _7250_/A vdd INVX1
XFILL_4__7211_ gnd vdd FILL
XSFILL44040x70050 gnd vdd FILL
XFILL_4__8191_ gnd vdd FILL
XFILL_3__9398_ gnd vdd FILL
XFILL111960x27050 gnd vdd FILL
XFILL_1__7433_ gnd vdd FILL
X_7179_ _7261_/Q gnd _7181_/A vdd INVX1
XSFILL23720x69050 gnd vdd FILL
XFILL_3__8349_ gnd vdd FILL
XFILL112040x36050 gnd vdd FILL
XFILL_1__7364_ gnd vdd FILL
XFILL_2_BUFX2_insert227 gnd vdd FILL
XFILL_4__7073_ gnd vdd FILL
XFILL_1__9103_ gnd vdd FILL
XFILL_2_BUFX2_insert238 gnd vdd FILL
XSFILL38920x50050 gnd vdd FILL
XFILL_2_BUFX2_insert249 gnd vdd FILL
XFILL_1__7295_ gnd vdd FILL
X_11820_ _11812_/Y _11811_/Y _11820_/C gnd _12449_/B vdd OAI21X1
XFILL_1__9034_ gnd vdd FILL
XFILL_1_BUFX2_insert905 gnd vdd FILL
XFILL_1_BUFX2_insert916 gnd vdd FILL
XFILL_1_BUFX2_insert927 gnd vdd FILL
XFILL_1_BUFX2_insert938 gnd vdd FILL
X_11751_ _11257_/Y _11386_/Y _11751_/C gnd _11752_/B vdd OAI21X1
XFILL_1_BUFX2_insert949 gnd vdd FILL
X_10702_ _10678_/A _8526_/B gnd _10703_/C vdd NAND2X1
XFILL_4__7975_ gnd vdd FILL
X_14470_ _9835_/Q _14470_/B _14469_/Y gnd _14472_/A vdd AOI21X1
X_11682_ _11279_/Y _11682_/B _11681_/Y gnd _11683_/B vdd OAI21X1
XSFILL84120x34050 gnd vdd FILL
XFILL_2__6990_ gnd vdd FILL
XBUFX2_insert226 _12432_/Y gnd _7502_/B vdd BUFX2
XFILL_4__6926_ gnd vdd FILL
X_13421_ _8918_/Q gnd _13421_/Y vdd INVX1
X_10633_ _10700_/B _9353_/B gnd _10634_/C vdd NAND2X1
XBUFX2_insert237 _12348_/Y gnd _6906_/B vdd BUFX2
XBUFX2_insert248 _10922_/Y gnd _14265_/C vdd BUFX2
XSFILL44120x50050 gnd vdd FILL
XBUFX2_insert259 _12423_/Y gnd _7877_/B vdd BUFX2
XFILL_1__9936_ gnd vdd FILL
XFILL_4__9645_ gnd vdd FILL
X_16140_ _16140_/A _16139_/Y gnd _16140_/Y vdd NOR2X1
X_13352_ _13259_/C _13352_/B gnd _13352_/Y vdd NOR2X1
XFILL_4__6857_ gnd vdd FILL
X_10564_ _10608_/Q gnd _10566_/A vdd INVX1
XFILL_5_CLKBUF1_insert116 gnd vdd FILL
XSFILL23800x49050 gnd vdd FILL
XFILL_5_CLKBUF1_insert127 gnd vdd FILL
XFILL_2__8660_ gnd vdd FILL
XFILL_5_BUFX2_insert860 gnd vdd FILL
XFILL_1__9867_ gnd vdd FILL
XFILL_5_CLKBUF1_insert138 gnd vdd FILL
XFILL_5_CLKBUF1_insert149 gnd vdd FILL
XFILL_5_BUFX2_insert871 gnd vdd FILL
X_12303_ _12327_/A gnd _12319_/C gnd _12306_/A vdd NAND3X1
XFILL_5_BUFX2_insert882 gnd vdd FILL
X_16071_ _16071_/A gnd _16071_/Y vdd INVX1
X_13283_ _13283_/A _13230_/Y gnd _13295_/A vdd NOR2X1
XFILL_2__7611_ gnd vdd FILL
X_10495_ _10495_/A gnd _10495_/Y vdd INVX1
XFILL_5_BUFX2_insert893 gnd vdd FILL
XFILL_2__8591_ gnd vdd FILL
XFILL_5__7320_ gnd vdd FILL
XFILL_4__8527_ gnd vdd FILL
X_15022_ _15022_/A _15197_/B _15633_/D _13445_/Y gnd _15026_/B vdd OAI22X1
XFILL_1__9798_ gnd vdd FILL
X_12234_ _12231_/Y _12234_/B _12234_/C gnd _11025_/A vdd NAND3X1
XBUFX2_insert1090 rst gnd BUFX2_insert524/A vdd BUFX2
XFILL_3__10150_ gnd vdd FILL
XFILL_2__7542_ gnd vdd FILL
XSFILL38840x9050 gnd vdd FILL
XFILL_1__8749_ gnd vdd FILL
XFILL_2__10880_ gnd vdd FILL
XFILL_5__7251_ gnd vdd FILL
XFILL_4__8458_ gnd vdd FILL
X_12165_ _12165_/A _12150_/B _12165_/C gnd _12165_/Y vdd OAI21X1
XFILL_4__11440_ gnd vdd FILL
XFILL_2__7473_ gnd vdd FILL
XFILL_5__10991_ gnd vdd FILL
XFILL_1__11260_ gnd vdd FILL
XFILL_5__7182_ gnd vdd FILL
X_11116_ _12177_/Y _12298_/Y gnd _11116_/Y vdd NOR2X1
XFILL_5__12730_ gnd vdd FILL
XFILL_0__11990_ gnd vdd FILL
XFILL_4__8389_ gnd vdd FILL
XFILL_2__9212_ gnd vdd FILL
X_12096_ _11988_/B _12770_/A _12096_/C gnd _12098_/B vdd NAND3X1
XFILL_4__11371_ gnd vdd FILL
XSFILL3720x70050 gnd vdd FILL
XFILL_1__11191_ gnd vdd FILL
XFILL_0__10941_ gnd vdd FILL
XSFILL84200x14050 gnd vdd FILL
X_15924_ _14465_/Y _15924_/B _16000_/A _14463_/B gnd _15926_/A vdd OAI22X1
XFILL_4__13110_ gnd vdd FILL
X_11047_ _11045_/Y _11046_/Y gnd _11640_/C vdd NOR2X1
XFILL_4__10322_ gnd vdd FILL
XFILL_2__9143_ gnd vdd FILL
XFILL_5__12661_ gnd vdd FILL
XFILL_4__14090_ gnd vdd FILL
XSFILL103880x13050 gnd vdd FILL
XFILL_2__11501_ gnd vdd FILL
XSFILL28920x82050 gnd vdd FILL
XFILL_3__13840_ gnd vdd FILL
XFILL_1__10142_ gnd vdd FILL
XFILL_2__12481_ gnd vdd FILL
XFILL_0__13660_ gnd vdd FILL
XFILL_5__14400_ gnd vdd FILL
XFILL_0__10872_ gnd vdd FILL
XFILL_5__11612_ gnd vdd FILL
XFILL_4__10253_ gnd vdd FILL
XFILL_5__15380_ gnd vdd FILL
XFILL_2__14220_ gnd vdd FILL
X_15855_ _15969_/C _7786_/Q _8170_/Q _16011_/D gnd _15856_/A vdd AOI22X1
XFILL_4__13041_ gnd vdd FILL
XFILL_5__12592_ gnd vdd FILL
XFILL_2__11432_ gnd vdd FILL
XFILL_3__10983_ gnd vdd FILL
XFILL_0__12611_ gnd vdd FILL
XFILL_3__13771_ gnd vdd FILL
XFILL_2_BUFX2_insert750 gnd vdd FILL
XFILL_1__14950_ gnd vdd FILL
XFILL_2_BUFX2_insert761 gnd vdd FILL
XFILL_0__13591_ gnd vdd FILL
X_14806_ _14805_/Y _13868_/B _14593_/C _14804_/Y gnd _14810_/A vdd OAI22X1
XFILL_5__14331_ gnd vdd FILL
XFILL_2_BUFX2_insert772 gnd vdd FILL
XFILL_3__15510_ gnd vdd FILL
XFILL_5__11543_ gnd vdd FILL
XFILL_3__12722_ gnd vdd FILL
XFILL_2__14151_ gnd vdd FILL
X_15786_ _15786_/A _15786_/B gnd _15812_/A vdd NOR2X1
XFILL_2_BUFX2_insert783 gnd vdd FILL
XFILL_4__10184_ gnd vdd FILL
XFILL_1__13901_ gnd vdd FILL
X_12998_ _12996_/Y vdd _12998_/C gnd _13062_/D vdd OAI21X1
XFILL_0__15330_ gnd vdd FILL
XFILL_2_BUFX2_insert794 gnd vdd FILL
XFILL_2__11363_ gnd vdd FILL
XFILL_1__14881_ gnd vdd FILL
XFILL_0__7040_ gnd vdd FILL
XSFILL99480x68050 gnd vdd FILL
XFILL_0_CLKBUF1_insert1078 gnd vdd FILL
XFILL_5__14262_ gnd vdd FILL
XFILL_2__13102_ gnd vdd FILL
X_14737_ _14737_/A _14737_/B gnd _14740_/C vdd NOR2X1
XFILL_2__10314_ gnd vdd FILL
XSFILL74120x66050 gnd vdd FILL
X_11949_ _11949_/A _11955_/B _11949_/C gnd _6858_/A vdd OAI21X1
XFILL_5__11474_ gnd vdd FILL
XFILL_3__15441_ gnd vdd FILL
XFILL_3__12653_ gnd vdd FILL
XFILL_1__13832_ gnd vdd FILL
XFILL_4__14992_ gnd vdd FILL
XFILL_2__14082_ gnd vdd FILL
XFILL_5__16001_ gnd vdd FILL
XFILL_2__11294_ gnd vdd FILL
XFILL_0__15261_ gnd vdd FILL
XFILL_5__13213_ gnd vdd FILL
XFILL_5__9754_ gnd vdd FILL
XFILL_0__12473_ gnd vdd FILL
XFILL_5__6966_ gnd vdd FILL
XFILL_6__15552_ gnd vdd FILL
XFILL_5__10425_ gnd vdd FILL
XFILL_5__14193_ gnd vdd FILL
XFILL_3__11604_ gnd vdd FILL
X_14668_ _14668_/A _14668_/B gnd _14692_/A vdd NOR2X1
XFILL_4__13943_ gnd vdd FILL
XFILL_2__13033_ gnd vdd FILL
XFILL_3__15372_ gnd vdd FILL
XFILL_0__14212_ gnd vdd FILL
XFILL_3__12584_ gnd vdd FILL
XFILL_2__10245_ gnd vdd FILL
XSFILL13560x19050 gnd vdd FILL
XFILL_5__8705_ gnd vdd FILL
XFILL_2__9976_ gnd vdd FILL
XFILL_1__13763_ gnd vdd FILL
XFILL_0__11424_ gnd vdd FILL
XFILL_1__10975_ gnd vdd FILL
XFILL_0__15192_ gnd vdd FILL
X_16407_ _16407_/A gnd _16406_/Y gnd _16407_/Y vdd OAI21X1
XFILL_6__14503_ gnd vdd FILL
X_13619_ _7167_/A _13619_/B _13864_/C _8447_/A gnd _13622_/A vdd AOI22X1
XFILL_5__13144_ gnd vdd FILL
XFILL_5__9685_ gnd vdd FILL
XSFILL53960x24050 gnd vdd FILL
XFILL_3__14323_ gnd vdd FILL
XFILL_5__6897_ gnd vdd FILL
XFILL_3__11535_ gnd vdd FILL
XFILL_0__8991_ gnd vdd FILL
XFILL_1__15502_ gnd vdd FILL
XFILL_3__7720_ gnd vdd FILL
XFILL_1__12714_ gnd vdd FILL
XFILL_4__13874_ gnd vdd FILL
X_14599_ _10606_/Q gnd _14599_/Y vdd INVX1
XFILL_2__10176_ gnd vdd FILL
XFILL_0__14143_ gnd vdd FILL
XBUFX2_insert760 _13412_/Y gnd _13633_/C vdd BUFX2
XFILL_5__8636_ gnd vdd FILL
XFILL_1__13694_ gnd vdd FILL
XFILL_0__11355_ gnd vdd FILL
XFILL_4__15613_ gnd vdd FILL
XSFILL3800x50050 gnd vdd FILL
XBUFX2_insert771 _13301_/Y gnd _7800_/B vdd BUFX2
XSFILL13800x6050 gnd vdd FILL
XFILL_0__7942_ gnd vdd FILL
X_16338_ _16336_/Y gnd _16338_/C gnd _16338_/Y vdd OAI21X1
XFILL_4__12825_ gnd vdd FILL
XBUFX2_insert782 _10911_/Y gnd _12150_/B vdd BUFX2
XFILL_3__14254_ gnd vdd FILL
XFILL_5__10287_ gnd vdd FILL
XBUFX2_insert793 _13334_/Y gnd _9401_/A vdd BUFX2
XFILL_1__15433_ gnd vdd FILL
XFILL_3__11466_ gnd vdd FILL
XFILL_1__12645_ gnd vdd FILL
XFILL_2__8858_ gnd vdd FILL
XSFILL54040x33050 gnd vdd FILL
XFILL_0__10306_ gnd vdd FILL
XFILL_2__14984_ gnd vdd FILL
XFILL_0__14074_ gnd vdd FILL
XFILL_0__11286_ gnd vdd FILL
XFILL_5__8567_ gnd vdd FILL
XFILL_5__12026_ gnd vdd FILL
X_8220_ _8218_/Y _8232_/B _8220_/C gnd _8290_/D vdd OAI21X1
XFILL_6__14365_ gnd vdd FILL
XFILL_4__15544_ gnd vdd FILL
XFILL_3__10417_ gnd vdd FILL
XFILL_0__7873_ gnd vdd FILL
X_16269_ _7156_/Q gnd _16269_/Y vdd INVX1
XFILL_2__7809_ gnd vdd FILL
XFILL_4__12756_ gnd vdd FILL
XFILL_3__14185_ gnd vdd FILL
XFILL_1__15364_ gnd vdd FILL
XFILL_0__13025_ gnd vdd FILL
XFILL_3__7582_ gnd vdd FILL
XFILL_2__13935_ gnd vdd FILL
XFILL_3__11397_ gnd vdd FILL
XFILL_0__10237_ gnd vdd FILL
XFILL_6__13316_ gnd vdd FILL
XFILL_1__12576_ gnd vdd FILL
XFILL_6__16104_ gnd vdd FILL
XFILL_2__8789_ gnd vdd FILL
XFILL_0__9612_ gnd vdd FILL
XFILL_6__7291_ gnd vdd FILL
XFILL_3__13136_ gnd vdd FILL
XFILL_4__11707_ gnd vdd FILL
X_8151_ _8057_/A _8151_/CLK _8664_/R vdd _8151_/D gnd vdd DFFSR
XFILL_5__8498_ gnd vdd FILL
XFILL_1__14315_ gnd vdd FILL
XFILL_4__15475_ gnd vdd FILL
XFILL_1__11527_ gnd vdd FILL
XFILL_2__13866_ gnd vdd FILL
XFILL_0__10168_ gnd vdd FILL
XSFILL109320x4050 gnd vdd FILL
XFILL_1__15295_ gnd vdd FILL
X_7102_ _7150_/Q gnd _7102_/Y vdd INVX1
XFILL_5__7449_ gnd vdd FILL
XFILL_0__9543_ gnd vdd FILL
XFILL_4__14426_ gnd vdd FILL
XFILL_3__9252_ gnd vdd FILL
XFILL_5__13977_ gnd vdd FILL
X_8082_ _8082_/A _9362_/B gnd _8083_/C vdd NAND2X1
XFILL_4__11638_ gnd vdd FILL
XFILL_2__15605_ gnd vdd FILL
XSFILL48920x13050 gnd vdd FILL
XFILL_1__14246_ gnd vdd FILL
XSFILL18680x52050 gnd vdd FILL
XFILL_3__10279_ gnd vdd FILL
XFILL_2__13797_ gnd vdd FILL
XFILL_1__11458_ gnd vdd FILL
XSFILL74200x46050 gnd vdd FILL
XFILL_0__14976_ gnd vdd FILL
XFILL_0__9474_ gnd vdd FILL
XFILL_5__15716_ gnd vdd FILL
XFILL_3__12018_ gnd vdd FILL
X_7033_ _7127_/Q gnd _7035_/A vdd INVX1
XFILL_3__8203_ gnd vdd FILL
XFILL_4__14357_ gnd vdd FILL
XFILL_2__12748_ gnd vdd FILL
XFILL_2__15536_ gnd vdd FILL
XFILL_1__10409_ gnd vdd FILL
XFILL_4__11569_ gnd vdd FILL
XFILL_1__14177_ gnd vdd FILL
XFILL_5__9119_ gnd vdd FILL
XFILL_0__13927_ gnd vdd FILL
XFILL_1__11389_ gnd vdd FILL
XSFILL49000x22050 gnd vdd FILL
XFILL_4__13308_ gnd vdd FILL
XFILL_5__15647_ gnd vdd FILL
XFILL_5__12859_ gnd vdd FILL
XFILL_3__8134_ gnd vdd FILL
XFILL_1__13128_ gnd vdd FILL
XFILL_4__14288_ gnd vdd FILL
XFILL_2__15467_ gnd vdd FILL
XFILL_0__13858_ gnd vdd FILL
XFILL_6__9932_ gnd vdd FILL
XFILL_0__8356_ gnd vdd FILL
XFILL_4__16027_ gnd vdd FILL
XFILL_4__13239_ gnd vdd FILL
XFILL_5__15578_ gnd vdd FILL
XFILL_3__8065_ gnd vdd FILL
X_8984_ _8969_/A _8472_/B gnd _8985_/C vdd NAND2X1
XFILL_2__14418_ gnd vdd FILL
XFILL_2__15398_ gnd vdd FILL
XFILL_3__13969_ gnd vdd FILL
XFILL_0__7307_ gnd vdd FILL
XSFILL38840x65050 gnd vdd FILL
XFILL112360x72050 gnd vdd FILL
XFILL_0__13789_ gnd vdd FILL
XFILL_5__14529_ gnd vdd FILL
X_7935_ _8025_/Q gnd _7935_/Y vdd INVX1
XFILL_1__7080_ gnd vdd FILL
XFILL_3__15708_ gnd vdd FILL
XSFILL54120x13050 gnd vdd FILL
XFILL_2__14349_ gnd vdd FILL
XFILL_0__15528_ gnd vdd FILL
XFILL_0__7238_ gnd vdd FILL
XFILL_3__15639_ gnd vdd FILL
X_7866_ _7866_/A _7821_/B _7865_/Y gnd _7866_/Y vdd OAI21X1
XFILL_0__15459_ gnd vdd FILL
X_9605_ _9691_/Q gnd _9605_/Y vdd INVX1
XFILL_0__7169_ gnd vdd FILL
XFILL_2__16019_ gnd vdd FILL
X_7797_ _7763_/A _7010_/CLK _7413_/R vdd _7797_/D gnd vdd DFFSR
XFILL_3__8967_ gnd vdd FILL
XFILL_4__7760_ gnd vdd FILL
XSFILL38840x50 gnd vdd FILL
X_9536_ _9534_/Y _9535_/A _9536_/C gnd _9582_/D vdd OAI21X1
XFILL_5_BUFX2_insert101 gnd vdd FILL
XSFILL18760x32050 gnd vdd FILL
XFILL_1__7982_ gnd vdd FILL
XSFILL44040x65050 gnd vdd FILL
XFILL_4__7691_ gnd vdd FILL
XFILL_6__7627_ gnd vdd FILL
XFILL_3__8898_ gnd vdd FILL
XFILL_1__6933_ gnd vdd FILL
XFILL_1__9721_ gnd vdd FILL
XSFILL58600x80050 gnd vdd FILL
X_9467_ _9467_/A _9466_/A _9467_/C gnd _9559_/D vdd OAI21X1
XFILL_3__7849_ gnd vdd FILL
X_8418_ _8418_/Q _7778_/CLK _8418_/R vdd _8418_/D gnd vdd DFFSR
XFILL_1__6864_ gnd vdd FILL
XFILL_4_BUFX2_insert801 gnd vdd FILL
XFILL_1__9652_ gnd vdd FILL
X_9398_ _9398_/A _7222_/B gnd _9399_/C vdd NAND2X1
XFILL_4_BUFX2_insert812 gnd vdd FILL
XFILL_4_BUFX2_insert823 gnd vdd FILL
XFILL_4__9361_ gnd vdd FILL
XFILL_4_BUFX2_insert834 gnd vdd FILL
X_10280_ _10280_/A _10280_/B _10279_/Y gnd _10342_/D vdd OAI21X1
XFILL_1__8603_ gnd vdd FILL
X_8349_ _8349_/A gnd _8349_/Y vdd INVX1
XFILL_4_BUFX2_insert845 gnd vdd FILL
XFILL_4_BUFX2_insert856 gnd vdd FILL
XFILL_4__8312_ gnd vdd FILL
XFILL_3__9519_ gnd vdd FILL
XFILL112440x52050 gnd vdd FILL
XFILL_4__9292_ gnd vdd FILL
XFILL_4_BUFX2_insert867 gnd vdd FILL
XSFILL64200x78050 gnd vdd FILL
XFILL_4_BUFX2_insert878 gnd vdd FILL
XFILL_4_BUFX2_insert889 gnd vdd FILL
XFILL_4__8243_ gnd vdd FILL
XFILL_1__8465_ gnd vdd FILL
XSFILL113720x40050 gnd vdd FILL
XFILL_1__7416_ gnd vdd FILL
X_13970_ _13970_/A _13966_/Y gnd _13973_/C vdd NOR2X1
XFILL_1__8396_ gnd vdd FILL
XFILL_4__7125_ gnd vdd FILL
XSFILL18840x12050 gnd vdd FILL
XSFILL94280x73050 gnd vdd FILL
X_12921_ _12829_/A _8180_/CLK _7391_/R vdd _12831_/Y gnd vdd DFFSR
XSFILL44120x45050 gnd vdd FILL
XFILL_1__7347_ gnd vdd FILL
XFILL_4__7056_ gnd vdd FILL
XSFILL84520x50050 gnd vdd FILL
X_15640_ _15637_/Y _15640_/B gnd _15641_/B vdd NOR2X1
XSFILL99320x10050 gnd vdd FILL
XFILL_5_BUFX2_insert1 gnd vdd FILL
X_12852_ _12850_/Y vdd _12851_/Y gnd _12852_/Y vdd OAI21X1
XFILL_1_BUFX2_insert702 gnd vdd FILL
XFILL_1_BUFX2_insert713 gnd vdd FILL
XFILL_1_BUFX2_insert724 gnd vdd FILL
XFILL_1__9017_ gnd vdd FILL
X_11803_ _11026_/C _11732_/B _11764_/D _11025_/Y gnd _11804_/C vdd AOI22X1
X_12783_ _12789_/A memoryOutData[29] gnd _12784_/C vdd NAND2X1
X_15571_ _15571_/A _15564_/Y gnd _15571_/Y vdd NAND2X1
XFILL_1_BUFX2_insert735 gnd vdd FILL
XSFILL73560x74050 gnd vdd FILL
XFILL_1_BUFX2_insert746 gnd vdd FILL
XFILL_1_BUFX2_insert757 gnd vdd FILL
XSFILL23800x1050 gnd vdd FILL
XFILL_1_BUFX2_insert768 gnd vdd FILL
X_14522_ _14522_/A _14572_/C _14522_/C gnd _14526_/A vdd AOI21X1
X_11734_ _11731_/B _11764_/A _11733_/Y gnd _11734_/Y vdd AOI21X1
XFILL_1_BUFX2_insert779 gnd vdd FILL
XFILL_4__7958_ gnd vdd FILL
X_14453_ _14451_/Y _13614_/C _13467_/A _14452_/Y gnd _14453_/Y vdd OAI22X1
X_11665_ _11762_/B _11641_/Y _11664_/Y gnd _11674_/B vdd NOR3X1
XFILL_4__10940_ gnd vdd FILL
XFILL_2__10030_ gnd vdd FILL
XFILL_5__11190_ gnd vdd FILL
XFILL_2__6973_ gnd vdd FILL
XSFILL89240x62050 gnd vdd FILL
XFILL_2__9761_ gnd vdd FILL
XSFILL53880x39050 gnd vdd FILL
XFILL_4_BUFX2_insert17 gnd vdd FILL
XFILL_1__10760_ gnd vdd FILL
XFILL_4_BUFX2_insert28 gnd vdd FILL
XFILL_4__6909_ gnd vdd FILL
X_13404_ _13372_/A _13404_/B _13718_/B gnd _13879_/B vdd NAND3X1
X_10616_ _10616_/A _10700_/B _10615_/Y gnd _10616_/Y vdd OAI21X1
XFILL_5__9470_ gnd vdd FILL
XFILL_4_BUFX2_insert39 gnd vdd FILL
X_14384_ _8879_/A gnd _15820_/A vdd INVX1
XFILL_5__10141_ gnd vdd FILL
XFILL_3__11320_ gnd vdd FILL
XFILL_4__7889_ gnd vdd FILL
XFILL_1__9919_ gnd vdd FILL
XFILL_2__8712_ gnd vdd FILL
X_11596_ _11431_/Y _11616_/B _11301_/Y gnd _11596_/Y vdd OAI21X1
XSFILL3720x65050 gnd vdd FILL
XFILL_4__10871_ gnd vdd FILL
XFILL_0__11140_ gnd vdd FILL
XFILL_4__9628_ gnd vdd FILL
X_13335_ _13335_/A gnd _13335_/Y vdd INVX1
X_16123_ _16123_/A _16123_/B gnd _16124_/A vdd NOR2X1
XFILL_6__11431_ gnd vdd FILL
XFILL_1__10691_ gnd vdd FILL
XFILL_4__12610_ gnd vdd FILL
X_10547_ _10548_/B _9011_/B gnd _10547_/Y vdd NAND2X1
XFILL_3__11251_ gnd vdd FILL
XSFILL28920x77050 gnd vdd FILL
XFILL_1__12430_ gnd vdd FILL
XFILL_4__13590_ gnd vdd FILL
XSFILL28120x58050 gnd vdd FILL
XFILL_2__8643_ gnd vdd FILL
XFILL_5_BUFX2_insert690 gnd vdd FILL
XFILL_2__11981_ gnd vdd FILL
XFILL_0__11071_ gnd vdd FILL
XFILL_5__8352_ gnd vdd FILL
XFILL_6__14150_ gnd vdd FILL
XFILL_5__13900_ gnd vdd FILL
X_13266_ _13266_/A _13262_/B _13260_/B _13295_/C gnd _13266_/Y vdd AOI22X1
X_16054_ _9967_/Q gnd _16056_/D vdd INVX1
XFILL_5__14880_ gnd vdd FILL
X_10478_ _10430_/A _8165_/CLK _8165_/R vdd _10432_/Y gnd vdd DFFSR
XFILL_2__10932_ gnd vdd FILL
XFILL_0__10022_ gnd vdd FILL
XFILL_2__13720_ gnd vdd FILL
XFILL_2__8574_ gnd vdd FILL
XFILL_3__11182_ gnd vdd FILL
XFILL_1__12361_ gnd vdd FILL
XFILL_5__7303_ gnd vdd FILL
X_15005_ _15000_/A _14982_/Y _14981_/Y gnd _15005_/Y vdd NAND3X1
X_12217_ _6870_/A _12289_/B _12289_/C gnd gnd _12217_/Y vdd AOI22X1
XFILL_5__13831_ gnd vdd FILL
X_13197_ _13145_/A _13201_/CLK _13201_/R vdd _13197_/D gnd vdd DFFSR
XFILL_3__10133_ gnd vdd FILL
XFILL_1__14100_ gnd vdd FILL
XFILL_4__15260_ gnd vdd FILL
XFILL_2__13651_ gnd vdd FILL
XFILL_4__12472_ gnd vdd FILL
XFILL_1__11312_ gnd vdd FILL
XFILL_3__15990_ gnd vdd FILL
XFILL_0__14830_ gnd vdd FILL
XFILL_1__15080_ gnd vdd FILL
XFILL_6__13032_ gnd vdd FILL
XFILL_1__12292_ gnd vdd FILL
XFILL_5__7234_ gnd vdd FILL
XSFILL7960x70050 gnd vdd FILL
XFILL_4__14211_ gnd vdd FILL
X_12148_ _13186_/Q gnd _12150_/A vdd INVX1
XFILL_2__12602_ gnd vdd FILL
XFILL_5__13762_ gnd vdd FILL
XFILL_4__11423_ gnd vdd FILL
XFILL_5__10974_ gnd vdd FILL
XFILL_4__15191_ gnd vdd FILL
XFILL_2__7456_ gnd vdd FILL
XFILL_1__14031_ gnd vdd FILL
XFILL_3__14941_ gnd vdd FILL
XFILL_3__10064_ gnd vdd FILL
XFILL_2__16370_ gnd vdd FILL
XFILL_2__13582_ gnd vdd FILL
XFILL_1__11243_ gnd vdd FILL
XFILL_5__15501_ gnd vdd FILL
XFILL_5__7165_ gnd vdd FILL
XFILL_0__14761_ gnd vdd FILL
XFILL_2__10794_ gnd vdd FILL
XFILL_5__12713_ gnd vdd FILL
XFILL_0__11973_ gnd vdd FILL
XSFILL74280x20050 gnd vdd FILL
X_12079_ _12047_/A _12508_/A _12011_/C gnd _12082_/A vdd NAND3X1
XFILL_4__14142_ gnd vdd FILL
XFILL_2__15321_ gnd vdd FILL
XFILL_2__12533_ gnd vdd FILL
XFILL_5__13693_ gnd vdd FILL
XFILL_4__11354_ gnd vdd FILL
XFILL_3__14872_ gnd vdd FILL
XFILL_0__13712_ gnd vdd FILL
XFILL_0__10924_ gnd vdd FILL
XFILL_0__8210_ gnd vdd FILL
XFILL_1__11174_ gnd vdd FILL
X_15907_ _15906_/Y _16213_/B _16208_/B _14484_/Y gnd _15908_/A vdd OAI22X1
XFILL_5__7096_ gnd vdd FILL
XFILL_0__14692_ gnd vdd FILL
XFILL_5__15432_ gnd vdd FILL
XSFILL59080x81050 gnd vdd FILL
XFILL_5__12644_ gnd vdd FILL
XSFILL89320x42050 gnd vdd FILL
XFILL_4__10305_ gnd vdd FILL
XSFILL53960x19050 gnd vdd FILL
XFILL_3__13823_ gnd vdd FILL
XFILL_2__15252_ gnd vdd FILL
XFILL_2__9126_ gnd vdd FILL
XFILL_4__14073_ gnd vdd FILL
XFILL_4__11285_ gnd vdd FILL
XFILL_1__10125_ gnd vdd FILL
XFILL_2__12464_ gnd vdd FILL
XSFILL109480x48050 gnd vdd FILL
XFILL_0__13643_ gnd vdd FILL
XFILL_0_BUFX2_insert1004 gnd vdd FILL
XFILL_0__8141_ gnd vdd FILL
XFILL_1__15982_ gnd vdd FILL
XFILL_0_BUFX2_insert1015 gnd vdd FILL
XFILL_2__14203_ gnd vdd FILL
XFILL_5__15363_ gnd vdd FILL
XFILL_4__13024_ gnd vdd FILL
XFILL_0_BUFX2_insert1026 gnd vdd FILL
X_15838_ _15953_/A _15837_/Y _15521_/C _14376_/Y gnd _15838_/Y vdd OAI22X1
XFILL_4__10236_ gnd vdd FILL
XFILL_5__12575_ gnd vdd FILL
XFILL_0_BUFX2_insert1037 gnd vdd FILL
XFILL_2__11415_ gnd vdd FILL
XFILL_2__15183_ gnd vdd FILL
XFILL_3__13754_ gnd vdd FILL
XFILL_0_BUFX2_insert1048 gnd vdd FILL
XFILL_2_BUFX2_insert580 gnd vdd FILL
XFILL_3__10966_ gnd vdd FILL
XFILL_2_BUFX2_insert591 gnd vdd FILL
XFILL_2__12395_ gnd vdd FILL
XFILL_0__16362_ gnd vdd FILL
XFILL_1__10056_ gnd vdd FILL
XFILL_1__14933_ gnd vdd FILL
XFILL_0_BUFX2_insert1059 gnd vdd FILL
XFILL_5__14314_ gnd vdd FILL
XFILL_0__13574_ gnd vdd FILL
X_7720_ _7718_/Y _7744_/B _7719_/Y gnd _7720_/Y vdd OAI21X1
XFILL_0__8072_ gnd vdd FILL
XFILL_0__10786_ gnd vdd FILL
XFILL_5__11526_ gnd vdd FILL
XFILL_2__8008_ gnd vdd FILL
XFILL_3__12705_ gnd vdd FILL
XFILL_4__10167_ gnd vdd FILL
XFILL_2__14134_ gnd vdd FILL
XSFILL94440x33050 gnd vdd FILL
X_15769_ _15769_/A _15769_/B _15758_/Y gnd _15769_/Y vdd NOR3X1
XFILL_5__15294_ gnd vdd FILL
XFILL_0__15313_ gnd vdd FILL
XFILL_2__11346_ gnd vdd FILL
XFILL_5__9806_ gnd vdd FILL
XFILL_1__14864_ gnd vdd FILL
XFILL_3__9870_ gnd vdd FILL
XFILL_3__10897_ gnd vdd FILL
XFILL_3__13685_ gnd vdd FILL
XFILL_0__12525_ gnd vdd FILL
XFILL_0__16293_ gnd vdd FILL
XFILL_5__14245_ gnd vdd FILL
XFILL_5__7998_ gnd vdd FILL
X_7651_ _7581_/A _7651_/CLK _7665_/R vdd _7583_/Y gnd vdd DFFSR
XFILL_3__15424_ gnd vdd FILL
XFILL_5__11457_ gnd vdd FILL
XFILL_3__12636_ gnd vdd FILL
XFILL_1__13815_ gnd vdd FILL
XFILL_2__14065_ gnd vdd FILL
XFILL_4__14975_ gnd vdd FILL
XFILL_0__15244_ gnd vdd FILL
XFILL_2__11277_ gnd vdd FILL
XFILL_5__9737_ gnd vdd FILL
XFILL_1__14795_ gnd vdd FILL
XFILL_0__12456_ gnd vdd FILL
XFILL_5__10408_ gnd vdd FILL
XFILL_5__6949_ gnd vdd FILL
XFILL_2__13016_ gnd vdd FILL
XFILL_5__14176_ gnd vdd FILL
XFILL_4__13926_ gnd vdd FILL
XFILL_3__15355_ gnd vdd FILL
X_7582_ _7624_/A _9374_/B gnd _7583_/C vdd NAND2X1
XFILL_5__11388_ gnd vdd FILL
XFILL_3__12567_ gnd vdd FILL
XFILL_1__13746_ gnd vdd FILL
XSFILL18680x47050 gnd vdd FILL
XFILL_0__11407_ gnd vdd FILL
XFILL_3__8752_ gnd vdd FILL
XFILL_1__10958_ gnd vdd FILL
XFILL_0__15175_ gnd vdd FILL
XFILL_0__12387_ gnd vdd FILL
XFILL_5__13127_ gnd vdd FILL
X_9321_ _9321_/Q _7916_/CLK _7276_/R vdd _9265_/Y gnd vdd DFFSR
XFILL_5__9668_ gnd vdd FILL
XFILL_3__14306_ gnd vdd FILL
XFILL_0__8974_ gnd vdd FILL
XFILL_4__13857_ gnd vdd FILL
XFILL_3__7703_ gnd vdd FILL
XFILL_3__11518_ gnd vdd FILL
XFILL_0__14126_ gnd vdd FILL
XFILL_3__12498_ gnd vdd FILL
XFILL_2__10159_ gnd vdd FILL
XFILL_3__15286_ gnd vdd FILL
XSFILL34200x57050 gnd vdd FILL
XFILL_1__13677_ gnd vdd FILL
XBUFX2_insert590 BUFX2_insert556/A gnd _9580_/R vdd BUFX2
XFILL_5__8619_ gnd vdd FILL
XFILL_0__11338_ gnd vdd FILL
XFILL_1__10889_ gnd vdd FILL
XFILL_5__9599_ gnd vdd FILL
X_9252_ _9277_/B _9380_/B gnd _9252_/Y vdd NAND2X1
XSFILL49000x17050 gnd vdd FILL
XFILL_4_BUFX2_insert108 gnd vdd FILL
XFILL_3__14237_ gnd vdd FILL
XFILL_3__11449_ gnd vdd FILL
XFILL_1__15416_ gnd vdd FILL
XFILL_1__12628_ gnd vdd FILL
XFILL_4__13788_ gnd vdd FILL
XSFILL89400x22050 gnd vdd FILL
XFILL_3__7634_ gnd vdd FILL
XFILL_0__14057_ gnd vdd FILL
XFILL_2__14967_ gnd vdd FILL
XFILL_1__16396_ gnd vdd FILL
X_8203_ _8203_/A gnd _8205_/A vdd INVX1
XFILL_5__12009_ gnd vdd FILL
XFILL_6__7343_ gnd vdd FILL
XFILL_0__11269_ gnd vdd FILL
XFILL_4__15527_ gnd vdd FILL
XFILL_4__12739_ gnd vdd FILL
XFILL_0__7856_ gnd vdd FILL
X_9183_ _9105_/A _7274_/CLK _7274_/R vdd _9107_/Y gnd vdd DFFSR
XFILL_1__15347_ gnd vdd FILL
XFILL_3__14168_ gnd vdd FILL
XFILL_0__13008_ gnd vdd FILL
XFILL_2__13918_ gnd vdd FILL
XFILL_3__7565_ gnd vdd FILL
XFILL_2__14898_ gnd vdd FILL
XFILL112360x67050 gnd vdd FILL
X_8134_ _8134_/A _8133_/A _8134_/C gnd _8176_/D vdd OAI21X1
XFILL_3__13119_ gnd vdd FILL
XFILL_4__15458_ gnd vdd FILL
XFILL_3_BUFX2_insert808 gnd vdd FILL
XFILL_3__14099_ gnd vdd FILL
XFILL_2__13849_ gnd vdd FILL
XFILL_3__7496_ gnd vdd FILL
XFILL_3_BUFX2_insert819 gnd vdd FILL
XFILL_1__15278_ gnd vdd FILL
XFILL_0__9526_ gnd vdd FILL
XFILL_4__14409_ gnd vdd FILL
X_8065_ _8065_/A _8079_/A _8064_/Y gnd _8065_/Y vdd OAI21X1
XFILL_1__14229_ gnd vdd FILL
XFILL_4__15389_ gnd vdd FILL
XFILL_3__9235_ gnd vdd FILL
XFILL_0__14959_ gnd vdd FILL
XSFILL79320x74050 gnd vdd FILL
XFILL_1__8250_ gnd vdd FILL
X_7016_ _6956_/A _7016_/CLK _8424_/R vdd _7016_/D gnd vdd DFFSR
XFILL_2__15519_ gnd vdd FILL
XFILL_3__9166_ gnd vdd FILL
XFILL_1__7201_ gnd vdd FILL
XFILL_0__9388_ gnd vdd FILL
XSFILL18760x27050 gnd vdd FILL
XSFILL114520x83050 gnd vdd FILL
XFILL_3__8117_ gnd vdd FILL
XFILL_3__9097_ gnd vdd FILL
XSFILL33800x30050 gnd vdd FILL
XFILL_0__8339_ gnd vdd FILL
X_8967_ _8965_/Y _9005_/A _8967_/C gnd _9051_/D vdd OAI21X1
X_7918_ _7918_/Q _8942_/CLK _9561_/R vdd _7872_/Y gnd vdd DFFSR
XFILL_1__7063_ gnd vdd FILL
XSFILL23880x18050 gnd vdd FILL
X_8898_ _8902_/B _9794_/B gnd _8898_/Y vdd NAND2X1
XFILL_4__8861_ gnd vdd FILL
XFILL_6__9777_ gnd vdd FILL
X_7849_ _7911_/Q gnd _7851_/A vdd INVX1
XFILL_0_CLKBUF1_insert113 gnd vdd FILL
XFILL_4__7812_ gnd vdd FILL
XFILL_0_CLKBUF1_insert124 gnd vdd FILL
XFILL112440x47050 gnd vdd FILL
XFILL_0_BUFX2_insert709 gnd vdd FILL
XFILL_0_CLKBUF1_insert135 gnd vdd FILL
XFILL_6__8728_ gnd vdd FILL
XFILL_0_CLKBUF1_insert146 gnd vdd FILL
XFILL_3__9999_ gnd vdd FILL
XFILL_0_CLKBUF1_insert157 gnd vdd FILL
XFILL_0_CLKBUF1_insert168 gnd vdd FILL
XFILL_4__7743_ gnd vdd FILL
XFILL_0_CLKBUF1_insert179 gnd vdd FILL
X_11450_ _11301_/Y gnd _11451_/B vdd INVX1
XSFILL39000x49050 gnd vdd FILL
X_9519_ _9577_/Q gnd _9519_/Y vdd INVX1
XFILL_1__7965_ gnd vdd FILL
X_10401_ _10372_/B _7329_/B gnd _10401_/Y vdd NAND2X1
XFILL_4__7674_ gnd vdd FILL
X_11381_ _11026_/A _11026_/B _11785_/A gnd _11381_/Y vdd OAI21X1
XFILL_1__6916_ gnd vdd FILL
XFILL_4__9413_ gnd vdd FILL
X_13120_ _13118_/Y _13155_/A _13120_/C gnd _13188_/D vdd OAI21X1
X_10332_ _10332_/Q _7781_/CLK _8670_/R vdd _10332_/D gnd vdd DFFSR
XSFILL114600x63050 gnd vdd FILL
XFILL_4_BUFX2_insert620 gnd vdd FILL
XFILL_1__9635_ gnd vdd FILL
XFILL_4_BUFX2_insert631 gnd vdd FILL
XFILL_1__6847_ gnd vdd FILL
XFILL_4_BUFX2_insert642 gnd vdd FILL
XFILL_4__9344_ gnd vdd FILL
XFILL_4_BUFX2_insert653 gnd vdd FILL
X_13051_ _6874_/A _13184_/CLK _8033_/R vdd _13051_/D gnd vdd DFFSR
X_10263_ _15509_/D gnd _10265_/A vdd INVX1
XFILL_4_BUFX2_insert664 gnd vdd FILL
XFILL_4_BUFX2_insert675 gnd vdd FILL
XFILL_4_BUFX2_insert686 gnd vdd FILL
X_12002_ _12002_/A _12000_/Y _12001_/Y gnd _13089_/B vdd NAND3X1
XFILL_4_BUFX2_insert697 gnd vdd FILL
XFILL_4__9275_ gnd vdd FILL
XFILL_2__7310_ gnd vdd FILL
XFILL_1__8517_ gnd vdd FILL
X_10194_ _10194_/A _10193_/A _10194_/C gnd _10194_/Y vdd OAI21X1
XFILL_1__9497_ gnd vdd FILL
XFILL_4__8226_ gnd vdd FILL
XFILL_2__7241_ gnd vdd FILL
XFILL_1__8448_ gnd vdd FILL
X_13953_ _13942_/Y _13953_/B gnd _13975_/B vdd NOR2X1
XFILL_1__8379_ gnd vdd FILL
XFILL_2__7172_ gnd vdd FILL
XFILL_5__10690_ gnd vdd FILL
XSFILL89240x57050 gnd vdd FILL
XFILL_4__7108_ gnd vdd FILL
XSFILL18760x8050 gnd vdd FILL
XFILL_4__8088_ gnd vdd FILL
XFILL_5__8970_ gnd vdd FILL
X_12904_ _12946_/Q gnd _12904_/Y vdd INVX1
XFILL_4__11070_ gnd vdd FILL
X_13884_ _16425_/Q _14344_/B _13884_/C _10846_/Q gnd _13885_/B vdd AOI22X1
XFILL_3__10820_ gnd vdd FILL
XFILL_4__7039_ gnd vdd FILL
XFILL_0__10640_ gnd vdd FILL
XFILL_4__10021_ gnd vdd FILL
X_15623_ _8864_/A gnd _15624_/A vdd INVX1
XFILL_1_BUFX2_insert510 gnd vdd FILL
X_12835_ _12923_/Q gnd _12837_/A vdd INVX1
XFILL_5__12360_ gnd vdd FILL
XFILL_2__11200_ gnd vdd FILL
XFILL_3__10751_ gnd vdd FILL
XFILL_1_BUFX2_insert521 gnd vdd FILL
XFILL_1_BUFX2_insert532 gnd vdd FILL
XFILL_2__12180_ gnd vdd FILL
XFILL_1__11930_ gnd vdd FILL
XSFILL94360x48050 gnd vdd FILL
XFILL_1_BUFX2_insert543 gnd vdd FILL
XFILL_0__10571_ gnd vdd FILL
XFILL_5__7852_ gnd vdd FILL
XSFILL33960x2050 gnd vdd FILL
XFILL_5__11311_ gnd vdd FILL
XFILL_1_BUFX2_insert554 gnd vdd FILL
X_15554_ _15633_/D _15553_/Y _15321_/C _15554_/D gnd _15555_/B vdd OAI22X1
X_12766_ _12764_/Y _12777_/A _12766_/C gnd _12814_/D vdd OAI21X1
XFILL_1_BUFX2_insert565 gnd vdd FILL
XFILL_5__12291_ gnd vdd FILL
XFILL_2__11131_ gnd vdd FILL
XFILL_3__13470_ gnd vdd FILL
XFILL_3__10682_ gnd vdd FILL
XFILL_0__12310_ gnd vdd FILL
XFILL_1_BUFX2_insert576 gnd vdd FILL
XFILL_1__11861_ gnd vdd FILL
XFILL_1_BUFX2_insert587 gnd vdd FILL
XFILL_0__13290_ gnd vdd FILL
XFILL_1_BUFX2_insert598 gnd vdd FILL
XFILL_5__14030_ gnd vdd FILL
X_14505_ _9708_/Q gnd _15937_/C vdd INVX1
XSFILL69160x24050 gnd vdd FILL
X_11717_ _11716_/Y _11717_/B gnd _11718_/A vdd NOR2X1
XFILL_5__11242_ gnd vdd FILL
XFILL_1__13600_ gnd vdd FILL
X_12697_ _12695_/Y _10944_/C _12697_/C gnd _12791_/D vdd OAI21X1
XFILL_3__12421_ gnd vdd FILL
XFILL_2__9813_ gnd vdd FILL
X_15485_ _15484_/Y _16311_/A _14999_/A _15485_/D gnd _15487_/B vdd OAI22X1
XFILL_4__14760_ gnd vdd FILL
XFILL_1__10812_ gnd vdd FILL
XFILL_4__11972_ gnd vdd FILL
XFILL_2__11062_ gnd vdd FILL
XFILL_1__14580_ gnd vdd FILL
XFILL_0__12241_ gnd vdd FILL
XFILL_5__9522_ gnd vdd FILL
XFILL_1__11792_ gnd vdd FILL
XSFILL7960x65050 gnd vdd FILL
X_11648_ _11646_/A _11647_/Y _11648_/C gnd _11661_/B vdd AOI21X1
XFILL_4__13711_ gnd vdd FILL
X_14436_ _14200_/C _14436_/B _14377_/B _14436_/D gnd _14437_/A vdd OAI22X1
XFILL_3__12352_ gnd vdd FILL
XFILL_4__10923_ gnd vdd FILL
XSFILL104360x33050 gnd vdd FILL
XFILL_2__10013_ gnd vdd FILL
XFILL_3__15140_ gnd vdd FILL
XFILL_5__11173_ gnd vdd FILL
XFILL_2__9744_ gnd vdd FILL
XFILL_4__14691_ gnd vdd FILL
XFILL_1__13531_ gnd vdd FILL
XFILL_1__10743_ gnd vdd FILL
XFILL_2__6956_ gnd vdd FILL
XFILL_2__15870_ gnd vdd FILL
XFILL_0__12172_ gnd vdd FILL
XFILL_5__10124_ gnd vdd FILL
XFILL_3__11303_ gnd vdd FILL
XSFILL74280x15050 gnd vdd FILL
XFILL_4__13642_ gnd vdd FILL
X_14367_ _14358_/Y _14367_/B _14366_/Y gnd _14380_/A vdd NAND3X1
X_11579_ _11578_/Y _11579_/B gnd _11580_/A vdd NOR2X1
XFILL_5__15981_ gnd vdd FILL
XFILL_2__14821_ gnd vdd FILL
XFILL_3__15071_ gnd vdd FILL
XSFILL79320x1050 gnd vdd FILL
XFILL_1__16250_ gnd vdd FILL
XFILL_3__12283_ gnd vdd FILL
XFILL_1__13462_ gnd vdd FILL
XFILL_2__9675_ gnd vdd FILL
XFILL_5__8404_ gnd vdd FILL
XFILL_0__11123_ gnd vdd FILL
X_16106_ _16106_/A _16106_/B _14705_/C _16225_/C gnd _16110_/B vdd OAI22X1
XFILL_2__6887_ gnd vdd FILL
XFILL_1__10674_ gnd vdd FILL
X_13318_ _13297_/C _13317_/Y gnd _13318_/Y vdd NOR2X1
XFILL_5__9384_ gnd vdd FILL
XFILL_0__7710_ gnd vdd FILL
XFILL_1__15201_ gnd vdd FILL
XFILL_3__14022_ gnd vdd FILL
XSFILL89320x37050 gnd vdd FILL
XFILL_5__14932_ gnd vdd FILL
X_14298_ _14298_/A _14290_/Y _14297_/Y gnd _14311_/A vdd NAND3X1
XFILL_4__16361_ gnd vdd FILL
XFILL_3__11234_ gnd vdd FILL
XFILL_5__10055_ gnd vdd FILL
XFILL_1__12413_ gnd vdd FILL
XFILL_4__13573_ gnd vdd FILL
XFILL_2__8626_ gnd vdd FILL
XFILL_1__16181_ gnd vdd FILL
XFILL_0__15931_ gnd vdd FILL
XFILL_4__10785_ gnd vdd FILL
XFILL_2__11964_ gnd vdd FILL
XFILL_2__14752_ gnd vdd FILL
XFILL_0__11054_ gnd vdd FILL
XSFILL99480x81050 gnd vdd FILL
XFILL_5__8335_ gnd vdd FILL
XFILL_1__13393_ gnd vdd FILL
X_16037_ _8894_/A _16037_/B _16037_/C gnd _16037_/Y vdd NAND3X1
XFILL_4__15312_ gnd vdd FILL
X_13249_ _13244_/A _13305_/B gnd _13249_/Y vdd NOR2X1
XFILL_5__14863_ gnd vdd FILL
XFILL_4__12524_ gnd vdd FILL
XFILL_3__7350_ gnd vdd FILL
XFILL_2__10915_ gnd vdd FILL
XFILL_4__16292_ gnd vdd FILL
XFILL_3__11165_ gnd vdd FILL
XFILL_2__13703_ gnd vdd FILL
XFILL_0__10005_ gnd vdd FILL
XFILL_1__15132_ gnd vdd FILL
XFILL_1__12344_ gnd vdd FILL
XFILL_2__11895_ gnd vdd FILL
XFILL_2__14683_ gnd vdd FILL
XFILL_0__15862_ gnd vdd FILL
XFILL_5__8266_ gnd vdd FILL
XFILL_5__13814_ gnd vdd FILL
XFILL_3__10116_ gnd vdd FILL
XFILL_4__15243_ gnd vdd FILL
XFILL_0__7572_ gnd vdd FILL
XFILL_5__14794_ gnd vdd FILL
XFILL_2__7508_ gnd vdd FILL
XFILL_4__12455_ gnd vdd FILL
XSFILL94440x28050 gnd vdd FILL
XFILL_2__13634_ gnd vdd FILL
XFILL_3__15973_ gnd vdd FILL
XFILL_0__14813_ gnd vdd FILL
XFILL_1__15063_ gnd vdd FILL
XFILL_3__11096_ gnd vdd FILL
XFILL_2__8488_ gnd vdd FILL
XFILL_5__7217_ gnd vdd FILL
XFILL_1__12275_ gnd vdd FILL
XFILL_0__15793_ gnd vdd FILL
XFILL_5__13745_ gnd vdd FILL
XFILL_4__11406_ gnd vdd FILL
XFILL_5__8197_ gnd vdd FILL
XFILL_3__9020_ gnd vdd FILL
XFILL_5__10957_ gnd vdd FILL
XFILL_4__15174_ gnd vdd FILL
XFILL_3__10047_ gnd vdd FILL
XFILL_1__14014_ gnd vdd FILL
XFILL_3__14924_ gnd vdd FILL
XFILL_2__7439_ gnd vdd FILL
XFILL_4__12386_ gnd vdd FILL
XFILL_2__16353_ gnd vdd FILL
XFILL_2__13565_ gnd vdd FILL
XFILL_1__11226_ gnd vdd FILL
XFILL_2__10777_ gnd vdd FILL
XFILL_0__14744_ gnd vdd FILL
XFILL_0__11956_ gnd vdd FILL
XFILL_0_BUFX2_insert15 gnd vdd FILL
XFILL_0__9242_ gnd vdd FILL
XFILL_4__14125_ gnd vdd FILL
X_9870_ _9870_/A gnd _9870_/Y vdd INVX1
XFILL_0_BUFX2_insert26 gnd vdd FILL
XFILL_2__15304_ gnd vdd FILL
XFILL_5__13676_ gnd vdd FILL
XFILL_2__12516_ gnd vdd FILL
XFILL_4__11337_ gnd vdd FILL
XFILL_3__14855_ gnd vdd FILL
XFILL_5__10888_ gnd vdd FILL
XFILL_0_BUFX2_insert37 gnd vdd FILL
XFILL_0__10907_ gnd vdd FILL
XFILL_0_BUFX2_insert48 gnd vdd FILL
XFILL_2__16284_ gnd vdd FILL
XFILL_2__13496_ gnd vdd FILL
XFILL_1__11157_ gnd vdd FILL
XFILL_5__7079_ gnd vdd FILL
XFILL_0_BUFX2_insert59 gnd vdd FILL
XFILL_0__14675_ gnd vdd FILL
XFILL_5__12627_ gnd vdd FILL
XFILL_0__11887_ gnd vdd FILL
XFILL_5__15415_ gnd vdd FILL
X_8821_ _8821_/Q _9834_/CLK _7793_/R vdd _8821_/D gnd vdd DFFSR
XFILL_0__9173_ gnd vdd FILL
XFILL_5__16395_ gnd vdd FILL
XFILL_3__13806_ gnd vdd FILL
XFILL_4__14056_ gnd vdd FILL
XFILL_2__9109_ gnd vdd FILL
XFILL_2__15235_ gnd vdd FILL
XFILL_2__12447_ gnd vdd FILL
XFILL_0__16414_ gnd vdd FILL
XFILL_1__10108_ gnd vdd FILL
XFILL_4__11268_ gnd vdd FILL
XFILL_0__13626_ gnd vdd FILL
XFILL_3__14786_ gnd vdd FILL
XFILL_0__8124_ gnd vdd FILL
XFILL_3__11998_ gnd vdd FILL
XFILL_1__15965_ gnd vdd FILL
XFILL_1__11088_ gnd vdd FILL
XFILL_5__15346_ gnd vdd FILL
XFILL_4__13007_ gnd vdd FILL
X_8752_ _8753_/B _8624_/B gnd _8752_/Y vdd NAND2X1
XFILL_3__9922_ gnd vdd FILL
XFILL_2__15166_ gnd vdd FILL
XFILL_3__13737_ gnd vdd FILL
XFILL_6__14897_ gnd vdd FILL
XFILL_4__11199_ gnd vdd FILL
XFILL_3__10949_ gnd vdd FILL
XFILL_1__10039_ gnd vdd FILL
XFILL_0__16345_ gnd vdd FILL
XFILL_6_BUFX2_insert715 gnd vdd FILL
XFILL_2__12378_ gnd vdd FILL
XFILL_1__14916_ gnd vdd FILL
XSFILL59160x56050 gnd vdd FILL
XFILL_0__13557_ gnd vdd FILL
XSFILL89400x17050 gnd vdd FILL
XFILL_1__15896_ gnd vdd FILL
XFILL_0__8055_ gnd vdd FILL
X_7703_ _7703_/A gnd _7705_/A vdd INVX1
XFILL_0__10769_ gnd vdd FILL
XFILL_5__11509_ gnd vdd FILL
XFILL_6__13848_ gnd vdd FILL
XFILL_5__15277_ gnd vdd FILL
X_8683_ _8683_/Q _9963_/CLK _9963_/R vdd _8631_/Y gnd vdd DFFSR
XFILL_5__12489_ gnd vdd FILL
XFILL_2__14117_ gnd vdd FILL
XFILL_2__11329_ gnd vdd FILL
XFILL_3__13668_ gnd vdd FILL
XFILL_0__12508_ gnd vdd FILL
XFILL_2__15097_ gnd vdd FILL
XFILL_3__9853_ gnd vdd FILL
XFILL_1__14847_ gnd vdd FILL
XFILL_0__16276_ gnd vdd FILL
XFILL_5__14228_ gnd vdd FILL
XFILL_0__13488_ gnd vdd FILL
XFILL_3__15407_ gnd vdd FILL
X_7634_ _7632_/Y _7577_/B _7634_/C gnd _7668_/D vdd OAI21X1
XFILL_3__12619_ gnd vdd FILL
XFILL_2__14048_ gnd vdd FILL
XFILL_4__14958_ gnd vdd FILL
XFILL_3__16387_ gnd vdd FILL
XFILL_0__15227_ gnd vdd FILL
XFILL_3__13599_ gnd vdd FILL
XFILL_0__12439_ gnd vdd FILL
XFILL_3__9784_ gnd vdd FILL
XFILL_1__14778_ gnd vdd FILL
XFILL_3__6996_ gnd vdd FILL
XSFILL13640x12050 gnd vdd FILL
XFILL_5__14159_ gnd vdd FILL
XFILL_6__9493_ gnd vdd FILL
XFILL_4__13909_ gnd vdd FILL
X_7565_ _7563_/Y _7606_/A _7565_/C gnd _7645_/D vdd OAI21X1
XFILL_3__15338_ gnd vdd FILL
XFILL_3__8735_ gnd vdd FILL
XFILL_4__14889_ gnd vdd FILL
XFILL_1_CLKBUF1_insert208 gnd vdd FILL
XFILL_0__15158_ gnd vdd FILL
XFILL_1__13729_ gnd vdd FILL
XFILL_6__8444_ gnd vdd FILL
X_9304_ _9304_/Q _7143_/CLK _7015_/R vdd _9214_/Y gnd vdd DFFSR
XSFILL79320x69050 gnd vdd FILL
XFILL_1_CLKBUF1_insert219 gnd vdd FILL
XFILL_6__15449_ gnd vdd FILL
XFILL_0__8957_ gnd vdd FILL
XFILL_1__7750_ gnd vdd FILL
X_7496_ _7416_/B _7496_/B gnd _7497_/C vdd NAND2X1
XFILL_0__14109_ gnd vdd FILL
XFILL_3__15269_ gnd vdd FILL
XFILL_2__15999_ gnd vdd FILL
XFILL_0__15089_ gnd vdd FILL
X_9235_ _9233_/Y _9282_/A _9235_/C gnd _9311_/D vdd OAI21X1
XFILL_1__7681_ gnd vdd FILL
XSFILL114520x78050 gnd vdd FILL
XFILL_0__8888_ gnd vdd FILL
XFILL_3__7617_ gnd vdd FILL
XFILL_1__16379_ gnd vdd FILL
XFILL_3__8597_ gnd vdd FILL
XFILL_1__9420_ gnd vdd FILL
X_9166_ _9163_/A _8654_/B gnd _9167_/C vdd NAND2X1
XFILL_0__7839_ gnd vdd FILL
XSFILL33800x25050 gnd vdd FILL
XFILL_3_BUFX2_insert605 gnd vdd FILL
XFILL_3__7548_ gnd vdd FILL
X_8117_ _8171_/Q gnd _8117_/Y vdd INVX1
XFILL_3_BUFX2_insert616 gnd vdd FILL
XFILL_3_BUFX2_insert627 gnd vdd FILL
XSFILL28760x3050 gnd vdd FILL
XFILL_1__9351_ gnd vdd FILL
X_9097_ _9151_/A _9737_/B gnd _9097_/Y vdd NAND2X1
XFILL_3_BUFX2_insert638 gnd vdd FILL
XFILL_3_BUFX2_insert649 gnd vdd FILL
XFILL_3__7479_ gnd vdd FILL
XFILL_0__9509_ gnd vdd FILL
X_8048_ _8048_/Q _8289_/CLK _7152_/R vdd _8006_/Y gnd vdd DFFSR
XFILL_1__9282_ gnd vdd FILL
XFILL_6__7188_ gnd vdd FILL
XFILL_3__9218_ gnd vdd FILL
XFILL_4__8011_ gnd vdd FILL
XFILL_1__8233_ gnd vdd FILL
XFILL_3__9149_ gnd vdd FILL
XSFILL23720x77050 gnd vdd FILL
X_10950_ _10957_/B _10936_/B _10950_/C gnd _10956_/C vdd NAND3X1
XFILL112040x44050 gnd vdd FILL
X_9999_ _9975_/B _9615_/B gnd _9999_/Y vdd NAND2X1
XFILL_1__7115_ gnd vdd FILL
X_10881_ _10881_/A _10881_/B gnd _10882_/B vdd NAND2X1
XFILL_1__8095_ gnd vdd FILL
XFILL_4__8913_ gnd vdd FILL
X_12620_ _12618_/Y vdd _12620_/C gnd _12680_/D vdd OAI21X1
XFILL_4__9893_ gnd vdd FILL
XFILL_1__7046_ gnd vdd FILL
XFILL_4__8844_ gnd vdd FILL
X_12551_ _11936_/B _12537_/CLK _12536_/R vdd _12551_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert506 gnd vdd FILL
XSFILL69080x39050 gnd vdd FILL
XFILL_0_BUFX2_insert517 gnd vdd FILL
XFILL_0_BUFX2_insert528 gnd vdd FILL
XFILL_0_BUFX2_insert539 gnd vdd FILL
X_11502_ _11502_/A _11502_/B gnd _11503_/A vdd NOR2X1
XFILL_4__8775_ gnd vdd FILL
X_12482_ vdd _12482_/B gnd _12482_/Y vdd NAND2X1
X_15270_ _8667_/Q gnd _15270_/Y vdd INVX1
XFILL_1__8997_ gnd vdd FILL
XFILL_4__7726_ gnd vdd FILL
X_14221_ _14221_/A gnd _14223_/D vdd INVX1
X_11433_ _11431_/Y _11616_/B _11433_/C gnd _11433_/Y vdd OAI21X1
XFILL_1__7948_ gnd vdd FILL
X_14152_ _14152_/A _13843_/C _14200_/C _14151_/Y gnd _14152_/Y vdd OAI22X1
X_11364_ _11484_/B gnd _11364_/Y vdd INVX8
XSFILL23800x57050 gnd vdd FILL
XFILL_1__7879_ gnd vdd FILL
X_10315_ _10318_/A _7499_/B gnd _10315_/Y vdd NAND2X1
X_13103_ _13103_/A gnd _13105_/A vdd INVX1
XFILL_4__7588_ gnd vdd FILL
XFILL_4_BUFX2_insert450 gnd vdd FILL
X_14083_ _14083_/A _13843_/C _13574_/C _14083_/D gnd _14084_/A vdd OAI22X1
XFILL_4_BUFX2_insert461 gnd vdd FILL
X_11295_ _11294_/Y gnd _11295_/Y vdd INVX1
XFILL_1__9618_ gnd vdd FILL
XCLKBUF1_insert207 CLKBUF1_insert192/A gnd _8429_/CLK vdd CLKBUF1
XFILL_4__10570_ gnd vdd FILL
XFILL_4_BUFX2_insert472 gnd vdd FILL
XCLKBUF1_insert218 CLKBUF1_insert218/A gnd _8038_/CLK vdd CLKBUF1
XFILL_5__8120_ gnd vdd FILL
XFILL_4_BUFX2_insert483 gnd vdd FILL
XFILL_2__9391_ gnd vdd FILL
X_13034_ _13032_/Y vdd _13034_/C gnd _13074_/D vdd OAI21X1
XFILL_1__10390_ gnd vdd FILL
XFILL_4_BUFX2_insert494 gnd vdd FILL
X_10246_ _10325_/B _6918_/B gnd _10246_/Y vdd NAND2X1
XFILL_2__10700_ gnd vdd FILL
XFILL_5__11860_ gnd vdd FILL
XFILL_1__9549_ gnd vdd FILL
XFILL_2__8342_ gnd vdd FILL
XFILL_2__11680_ gnd vdd FILL
XFILL_4__9258_ gnd vdd FILL
XFILL_5__10811_ gnd vdd FILL
XFILL_4__12240_ gnd vdd FILL
X_10177_ _10177_/A gnd _10179_/A vdd INVX1
XFILL_2__10631_ gnd vdd FILL
XFILL_5__11791_ gnd vdd FILL
XFILL_2__8273_ gnd vdd FILL
XFILL_1__12060_ gnd vdd FILL
XFILL_3__12970_ gnd vdd FILL
XFILL_4__8209_ gnd vdd FILL
XFILL_0__11810_ gnd vdd FILL
XFILL_0__12790_ gnd vdd FILL
XFILL_5__13530_ gnd vdd FILL
XSFILL69160x19050 gnd vdd FILL
XFILL_5__10742_ gnd vdd FILL
XFILL_2__7224_ gnd vdd FILL
XFILL_2__13350_ gnd vdd FILL
X_14985_ _12764_/A _14984_/Y gnd _16035_/B vdd NOR2X1
XFILL_3__11921_ gnd vdd FILL
XFILL_4__12171_ gnd vdd FILL
XFILL_1__11011_ gnd vdd FILL
XFILL_2__10562_ gnd vdd FILL
XFILL_0__11741_ gnd vdd FILL
XFILL_6__14820_ gnd vdd FILL
XFILL_3_CLKBUF1_insert130 gnd vdd FILL
XFILL_5__13461_ gnd vdd FILL
XFILL_2__12301_ gnd vdd FILL
XFILL_4__11122_ gnd vdd FILL
X_13936_ _7700_/A gnd _13937_/B vdd INVX1
XFILL_3__14640_ gnd vdd FILL
XFILL_3_CLKBUF1_insert141 gnd vdd FILL
XFILL_5__10673_ gnd vdd FILL
XSFILL104360x28050 gnd vdd FILL
XFILL_2__13281_ gnd vdd FILL
XFILL_3_CLKBUF1_insert152 gnd vdd FILL
XFILL_3__11852_ gnd vdd FILL
XFILL_0__14460_ gnd vdd FILL
XFILL_5__15200_ gnd vdd FILL
XFILL_3_CLKBUF1_insert163 gnd vdd FILL
XFILL_2__10493_ gnd vdd FILL
XFILL_5__12412_ gnd vdd FILL
XFILL_0__11672_ gnd vdd FILL
XFILL_5__8953_ gnd vdd FILL
XFILL_3_CLKBUF1_insert174 gnd vdd FILL
XFILL_3_CLKBUF1_insert185 gnd vdd FILL
XFILL_5__16180_ gnd vdd FILL
XFILL_4__15930_ gnd vdd FILL
XFILL_2__15020_ gnd vdd FILL
XFILL_6__11963_ gnd vdd FILL
XFILL_4__11053_ gnd vdd FILL
X_13867_ _8206_/A gnd _13867_/Y vdd INVX1
XFILL_5__13392_ gnd vdd FILL
XFILL_2__12232_ gnd vdd FILL
XFILL_3__10803_ gnd vdd FILL
XFILL_3_CLKBUF1_insert196 gnd vdd FILL
XFILL_3__14571_ gnd vdd FILL
XFILL_0__13411_ gnd vdd FILL
XFILL_2__7086_ gnd vdd FILL
XFILL_0__10623_ gnd vdd FILL
XFILL_1__12962_ gnd vdd FILL
XFILL_3__11783_ gnd vdd FILL
XFILL_1__15750_ gnd vdd FILL
XFILL_0__14391_ gnd vdd FILL
X_15606_ _16314_/D _15606_/B _16309_/A _15604_/Y gnd _15606_/Y vdd OAI22X1
XFILL_5__15131_ gnd vdd FILL
X_12818_ _12818_/Q _12692_/CLK _12692_/R vdd _12818_/D gnd vdd DFFSR
XFILL_5__12343_ gnd vdd FILL
XFILL_1_BUFX2_insert340 gnd vdd FILL
XFILL_3__16310_ gnd vdd FILL
XFILL_5__8884_ gnd vdd FILL
XFILL_4__10004_ gnd vdd FILL
XFILL_1_BUFX2_insert351 gnd vdd FILL
XFILL_6__14682_ gnd vdd FILL
XFILL_3__13522_ gnd vdd FILL
XFILL_4__15861_ gnd vdd FILL
X_13798_ _13798_/A _13868_/B gnd _13804_/A vdd NOR2X1
XFILL_1__11913_ gnd vdd FILL
XFILL_2__12163_ gnd vdd FILL
XFILL_1__14701_ gnd vdd FILL
XFILL_0__16130_ gnd vdd FILL
XFILL_1_BUFX2_insert362 gnd vdd FILL
XFILL_0__13342_ gnd vdd FILL
XFILL_1_BUFX2_insert373 gnd vdd FILL
XFILL_1__15681_ gnd vdd FILL
XFILL_1__12893_ gnd vdd FILL
XFILL_0__10554_ gnd vdd FILL
XFILL_5__7835_ gnd vdd FILL
XFILL_6__13633_ gnd vdd FILL
XFILL_4__14812_ gnd vdd FILL
XFILL_5__15062_ gnd vdd FILL
X_15537_ _16166_/A _15537_/B _8034_/Q _15081_/Y gnd _15537_/Y vdd AOI22X1
XFILL_1_BUFX2_insert384 gnd vdd FILL
X_12749_ _12809_/Q gnd _12751_/A vdd INVX1
XFILL_3__16241_ gnd vdd FILL
XFILL_5__12274_ gnd vdd FILL
XFILL_2__11114_ gnd vdd FILL
XFILL_1_BUFX2_insert395 gnd vdd FILL
XFILL_1__14632_ gnd vdd FILL
XFILL_3__13453_ gnd vdd FILL
XFILL_4__15792_ gnd vdd FILL
XFILL_3__10665_ gnd vdd FILL
XSFILL89720x53050 gnd vdd FILL
XFILL_2__12094_ gnd vdd FILL
XFILL_3__6850_ gnd vdd FILL
XFILL_0__16061_ gnd vdd FILL
XFILL_1__11844_ gnd vdd FILL
XFILL_0__13273_ gnd vdd FILL
XFILL_5__14013_ gnd vdd FILL
XFILL_5__11225_ gnd vdd FILL
XFILL_0__9860_ gnd vdd FILL
XFILL_3__12404_ gnd vdd FILL
XFILL_6__10776_ gnd vdd FILL
XFILL_4__14743_ gnd vdd FILL
X_15468_ _15225_/A _7572_/A _7520_/Q _15383_/D gnd _15468_/Y vdd AOI22X1
XFILL_2__15922_ gnd vdd FILL
XFILL_3__16172_ gnd vdd FILL
XFILL_4__11955_ gnd vdd FILL
XFILL_0__15012_ gnd vdd FILL
XSFILL13560x27050 gnd vdd FILL
XFILL_2__11045_ gnd vdd FILL
XFILL_1__14563_ gnd vdd FILL
XFILL_5__9505_ gnd vdd FILL
XFILL_3__13384_ gnd vdd FILL
XFILL_0__12224_ gnd vdd FILL
XFILL_2__7988_ gnd vdd FILL
XFILL_1__11775_ gnd vdd FILL
XFILL_6__12515_ gnd vdd FILL
XSFILL53960x32050 gnd vdd FILL
X_14419_ _9906_/A gnd _14419_/Y vdd INVX1
XFILL_4__10906_ gnd vdd FILL
X_7350_ _7308_/A _7222_/B gnd _7350_/Y vdd NAND2X1
XFILL_5__11156_ gnd vdd FILL
XFILL_3__15123_ gnd vdd FILL
XFILL_6__13495_ gnd vdd FILL
XFILL_5__7697_ gnd vdd FILL
XFILL_6__16283_ gnd vdd FILL
XFILL_0__9791_ gnd vdd FILL
XFILL_2__9727_ gnd vdd FILL
XSFILL78760x77050 gnd vdd FILL
X_15399_ _16425_/Q _15680_/B _15680_/C gnd _15399_/Y vdd NAND3X1
XSFILL109480x61050 gnd vdd FILL
XFILL_3__8520_ gnd vdd FILL
XFILL_1__16302_ gnd vdd FILL
XFILL_3__12335_ gnd vdd FILL
XFILL_4__14674_ gnd vdd FILL
XFILL_1__13514_ gnd vdd FILL
XFILL_4__11886_ gnd vdd FILL
XFILL_2__6939_ gnd vdd FILL
XFILL_2__15853_ gnd vdd FILL
XFILL_1__14494_ gnd vdd FILL
XSFILL94280x9050 gnd vdd FILL
XFILL_0__12155_ gnd vdd FILL
XFILL_6__15234_ gnd vdd FILL
XFILL_5__10107_ gnd vdd FILL
XFILL_4__16413_ gnd vdd FILL
XFILL_4__13625_ gnd vdd FILL
XFILL_0__8742_ gnd vdd FILL
XFILL_2__14804_ gnd vdd FILL
XFILL_3__15054_ gnd vdd FILL
XFILL_5__15964_ gnd vdd FILL
XFILL_5__11087_ gnd vdd FILL
X_7281_ _7281_/Q _9205_/CLK _8433_/R vdd _7281_/D gnd vdd DFFSR
XFILL_4__10837_ gnd vdd FILL
XFILL_1__16233_ gnd vdd FILL
XFILL_3__8451_ gnd vdd FILL
XFILL_1__13445_ gnd vdd FILL
XSFILL54040x41050 gnd vdd FILL
XFILL_2__9658_ gnd vdd FILL
XFILL_3__12266_ gnd vdd FILL
XFILL_0__11106_ gnd vdd FILL
XFILL_1__10657_ gnd vdd FILL
XFILL_2__15784_ gnd vdd FILL
X_9020_ _8961_/B _7868_/B gnd _9021_/C vdd NAND2X1
XFILL_2__12996_ gnd vdd FILL
XFILL_0__12086_ gnd vdd FILL
XFILL_5__9367_ gnd vdd FILL
XSFILL69640x20050 gnd vdd FILL
XFILL_5__10038_ gnd vdd FILL
XFILL_4__16344_ gnd vdd FILL
XFILL_6__12377_ gnd vdd FILL
XFILL_3__14005_ gnd vdd FILL
XFILL_5__14915_ gnd vdd FILL
XFILL_2__8609_ gnd vdd FILL
XFILL_4__13556_ gnd vdd FILL
XFILL_3__11217_ gnd vdd FILL
XFILL_4__10768_ gnd vdd FILL
XFILL_5__15895_ gnd vdd FILL
XFILL_2__14735_ gnd vdd FILL
XFILL_3__12197_ gnd vdd FILL
XFILL_1__16164_ gnd vdd FILL
XFILL_0__15914_ gnd vdd FILL
XFILL_3__8382_ gnd vdd FILL
XFILL_1__13376_ gnd vdd FILL
XFILL_2__11947_ gnd vdd FILL
XFILL_0__11037_ gnd vdd FILL
XFILL_5__8318_ gnd vdd FILL
XFILL_6__11328_ gnd vdd FILL
XFILL_4__12507_ gnd vdd FILL
XFILL_5__9298_ gnd vdd FILL
XFILL_0__7624_ gnd vdd FILL
XFILL_6__15096_ gnd vdd FILL
XFILL_5__14846_ gnd vdd FILL
XFILL_3__11148_ gnd vdd FILL
XFILL_1__15115_ gnd vdd FILL
XFILL_4__16275_ gnd vdd FILL
XFILL_3__7333_ gnd vdd FILL
XFILL_4__13487_ gnd vdd FILL
XFILL_1__12327_ gnd vdd FILL
XFILL_4__10699_ gnd vdd FILL
XFILL_1__16095_ gnd vdd FILL
XFILL_0__15845_ gnd vdd FILL
XFILL_2__14666_ gnd vdd FILL
XFILL_2__11878_ gnd vdd FILL
XFILL_5__8249_ gnd vdd FILL
XFILL_6__14047_ gnd vdd FILL
XFILL_4__15226_ gnd vdd FILL
XFILL_0__7555_ gnd vdd FILL
XFILL_2__16405_ gnd vdd FILL
XFILL_4__12438_ gnd vdd FILL
XFILL_2__13617_ gnd vdd FILL
XFILL_5__11989_ gnd vdd FILL
XFILL_3__15956_ gnd vdd FILL
XFILL_1__15046_ gnd vdd FILL
XFILL_3__11079_ gnd vdd FILL
XSFILL48920x21050 gnd vdd FILL
XFILL_5__14777_ gnd vdd FILL
XFILL_2__10829_ gnd vdd FILL
XFILL_1__12258_ gnd vdd FILL
XSFILL49400x28050 gnd vdd FILL
XFILL_2__14597_ gnd vdd FILL
XFILL_0__15776_ gnd vdd FILL
XFILL_0__12988_ gnd vdd FILL
XFILL_0__7486_ gnd vdd FILL
X_9922_ _9937_/A _9282_/B gnd _9923_/C vdd NAND2X1
XFILL_4__15157_ gnd vdd FILL
XFILL_5__13728_ gnd vdd FILL
XFILL_3__14907_ gnd vdd FILL
XFILL_3__9003_ gnd vdd FILL
XFILL_4__12369_ gnd vdd FILL
XFILL_2__16336_ gnd vdd FILL
XFILL_1__11209_ gnd vdd FILL
XFILL_3__7195_ gnd vdd FILL
XFILL_0__14727_ gnd vdd FILL
XFILL_2__13548_ gnd vdd FILL
XFILL_3__15887_ gnd vdd FILL
XFILL_1__12189_ gnd vdd FILL
XFILL_0__11939_ gnd vdd FILL
XFILL_0__9225_ gnd vdd FILL
XSFILL49000x30050 gnd vdd FILL
XFILL_4__14108_ gnd vdd FILL
XFILL_5__13659_ gnd vdd FILL
XSFILL37960x45050 gnd vdd FILL
X_9853_ _9902_/B _9981_/B gnd _9854_/C vdd NAND2X1
XFILL_3__14838_ gnd vdd FILL
XFILL_4__15088_ gnd vdd FILL
XFILL_2__16267_ gnd vdd FILL
XFILL_0__14658_ gnd vdd FILL
XFILL_2__13479_ gnd vdd FILL
XFILL_0__9156_ gnd vdd FILL
X_8804_ _8736_/A _8161_/CLK _7140_/R vdd _8804_/D gnd vdd DFFSR
XFILL_4__14039_ gnd vdd FILL
XFILL_2__15218_ gnd vdd FILL
X_9784_ _9836_/Q gnd _9786_/A vdd INVX1
XFILL_5__16378_ gnd vdd FILL
XFILL_0__13609_ gnd vdd FILL
X_6996_ _6937_/B _7508_/B gnd _6996_/Y vdd NAND2X1
XFILL_3__14769_ gnd vdd FILL
XSFILL38840x73050 gnd vdd FILL
XFILL_2__16198_ gnd vdd FILL
XFILL_1__15948_ gnd vdd FILL
XFILL_0__8107_ gnd vdd FILL
XFILL112360x80050 gnd vdd FILL
XFILL_0__14589_ gnd vdd FILL
XFILL_0__9087_ gnd vdd FILL
XFILL_5__15329_ gnd vdd FILL
XFILL_6__7875_ gnd vdd FILL
X_8735_ _8735_/A _8698_/A _8735_/C gnd _8803_/D vdd OAI21X1
XSFILL54120x21050 gnd vdd FILL
XFILL_3__9905_ gnd vdd FILL
XFILL_0__16328_ gnd vdd FILL
XFILL_2__15149_ gnd vdd FILL
XFILL_6_BUFX2_insert556 gnd vdd FILL
XFILL_4__6890_ gnd vdd FILL
XFILL_1__15879_ gnd vdd FILL
XFILL_6_BUFX2_insert567 gnd vdd FILL
X_8666_ _8666_/Q _9306_/CLK _9306_/R vdd _8666_/D gnd vdd DFFSR
XFILL_0__16259_ gnd vdd FILL
XSFILL43960x64050 gnd vdd FILL
X_7617_ _7663_/Q gnd _7619_/A vdd INVX1
XFILL_1__8851_ gnd vdd FILL
X_8597_ _8657_/A _7317_/B gnd _8598_/C vdd NAND2X1
XFILL_3__9767_ gnd vdd FILL
XFILL_3__6979_ gnd vdd FILL
XSFILL18760x40050 gnd vdd FILL
XSFILL99640x36050 gnd vdd FILL
XFILL_1__7802_ gnd vdd FILL
X_7548_ _7548_/A gnd _7550_/A vdd INVX1
XFILL_3__8718_ gnd vdd FILL
XSFILL44040x73050 gnd vdd FILL
XFILL_1__8782_ gnd vdd FILL
XFILL_0__9989_ gnd vdd FILL
XFILL_4__8491_ gnd vdd FILL
XFILL_1__7733_ gnd vdd FILL
X_7479_ _7479_/A _7503_/B _7478_/Y gnd _7479_/Y vdd OAI21X1
XFILL_4__7442_ gnd vdd FILL
XFILL_3__8649_ gnd vdd FILL
X_9218_ _9306_/Q gnd _9220_/A vdd INVX1
X_10100_ _10100_/Q _9834_/CLK _7793_/R vdd _10066_/Y gnd vdd DFFSR
XSFILL109640x21050 gnd vdd FILL
XFILL_4__7373_ gnd vdd FILL
XFILL_3_BUFX2_insert402 gnd vdd FILL
XFILL_1__9403_ gnd vdd FILL
X_11080_ _11079_/Y gnd _11081_/B vdd INVX1
X_9149_ _9147_/Y _9101_/B _9148_/Y gnd _9149_/Y vdd OAI21X1
XFILL_3_BUFX2_insert413 gnd vdd FILL
XFILL_3_BUFX2_insert424 gnd vdd FILL
XFILL_4__9112_ gnd vdd FILL
XFILL_1__7595_ gnd vdd FILL
XFILL112440x60050 gnd vdd FILL
X_10031_ _15846_/A gnd _10031_/Y vdd INVX1
XFILL_3_BUFX2_insert435 gnd vdd FILL
XFILL_3_BUFX2_insert446 gnd vdd FILL
XFILL_1__9334_ gnd vdd FILL
XFILL_3_BUFX2_insert457 gnd vdd FILL
XFILL_3_BUFX2_insert468 gnd vdd FILL
XFILL_3_BUFX2_insert479 gnd vdd FILL
XSFILL114520x6050 gnd vdd FILL
XFILL_4__9043_ gnd vdd FILL
XFILL_1__9265_ gnd vdd FILL
XSFILL114200x55050 gnd vdd FILL
XFILL_1__8216_ gnd vdd FILL
X_14770_ _9457_/Q gnd _14771_/D vdd INVX1
X_11982_ _11980_/Y _11895_/B _11982_/C gnd _6869_/A vdd OAI21X1
XSFILL18840x20050 gnd vdd FILL
XSFILL94280x81050 gnd vdd FILL
X_13721_ _8453_/A gnd _13722_/D vdd INVX1
X_10933_ _12782_/A gnd _10933_/Y vdd INVX1
XFILL_1__8147_ gnd vdd FILL
XFILL_0_BUFX2_insert7 gnd vdd FILL
X_16440_ _16390_/A _7269_/CLK _9061_/R vdd _16392_/Y gnd vdd DFFSR
XFILL_4_CLKBUF1_insert203 gnd vdd FILL
X_13652_ _9434_/Q gnd _15213_/A vdd INVX1
X_10864_ _16107_/A _7664_/CLK _7920_/R vdd _10864_/D gnd vdd DFFSR
XFILL_1__8078_ gnd vdd FILL
XFILL_4_CLKBUF1_insert214 gnd vdd FILL
XFILL_2__8960_ gnd vdd FILL
X_12603_ _12675_/Q gnd _12605_/A vdd INVX1
XFILL_4__9876_ gnd vdd FILL
XFILL112120x19050 gnd vdd FILL
X_16371_ _16369_/Y gnd _16371_/C gnd _16433_/D vdd OAI21X1
XFILL_0_BUFX2_insert303 gnd vdd FILL
X_10795_ _10795_/A _10797_/A _10795_/C gnd _10855_/D vdd OAI21X1
X_13583_ _13571_/Y _13582_/Y gnd _13583_/Y vdd NOR2X1
XFILL_0_BUFX2_insert314 gnd vdd FILL
XFILL_2__8891_ gnd vdd FILL
XFILL_5__7620_ gnd vdd FILL
XFILL_4__8827_ gnd vdd FILL
XFILL_0_BUFX2_insert325 gnd vdd FILL
X_15322_ _15322_/A _13781_/Y _13780_/Y _15322_/D gnd _15322_/Y vdd OAI22X1
X_12534_ _12534_/A vdd _12533_/Y gnd _12566_/D vdd OAI21X1
XFILL_0_BUFX2_insert336 gnd vdd FILL
XFILL_0_BUFX2_insert347 gnd vdd FILL
XFILL_3__10450_ gnd vdd FILL
XFILL_2__7842_ gnd vdd FILL
XFILL_0_BUFX2_insert358 gnd vdd FILL
XFILL_0_BUFX2_insert369 gnd vdd FILL
XFILL_0__10270_ gnd vdd FILL
XFILL_5__7551_ gnd vdd FILL
XFILL_4__8758_ gnd vdd FILL
XFILL_5__11010_ gnd vdd FILL
X_15253_ _15251_/Y _15924_/B _16000_/A _15252_/Y gnd _15253_/Y vdd OAI22X1
X_12465_ _12465_/A vdd _12464_/Y gnd _12465_/Y vdd OAI21X1
XFILL_4__11740_ gnd vdd FILL
XFILL_3__10381_ gnd vdd FILL
XSFILL89240x70050 gnd vdd FILL
XSFILL53880x47050 gnd vdd FILL
XFILL_6__12300_ gnd vdd FILL
XFILL_4__7709_ gnd vdd FILL
XFILL_1__11560_ gnd vdd FILL
X_14204_ _14204_/A _14203_/Y gnd _14205_/C vdd NOR2X1
XFILL_6__13280_ gnd vdd FILL
XFILL_5__7482_ gnd vdd FILL
X_11416_ _11416_/A _11212_/A gnd _11417_/B vdd NOR2X1
X_15184_ _15184_/A _15178_/Y _15184_/C gnd _15185_/A vdd NAND3X1
XFILL_2__9512_ gnd vdd FILL
X_12396_ _12394_/Y _12395_/A _12396_/C gnd _12396_/Y vdd OAI21X1
XFILL_6__10492_ gnd vdd FILL
XFILL_3__12120_ gnd vdd FILL
XFILL_1__10511_ gnd vdd FILL
XSFILL3720x73050 gnd vdd FILL
XFILL_4__11671_ gnd vdd FILL
XSFILL68920x69050 gnd vdd FILL
XFILL_2__12850_ gnd vdd FILL
XFILL_5__9221_ gnd vdd FILL
XFILL_1__11491_ gnd vdd FILL
X_14135_ _14470_/B _9760_/A _14135_/C _13621_/B gnd _14143_/B vdd AOI22X1
XFILL_4__13410_ gnd vdd FILL
X_11347_ _10996_/Y _11223_/B gnd _11347_/Y vdd NAND2X1
XFILL_5__12961_ gnd vdd FILL
XFILL_3__12051_ gnd vdd FILL
XFILL_4__10622_ gnd vdd FILL
XFILL_1__13230_ gnd vdd FILL
XFILL_4__14390_ gnd vdd FILL
XFILL_2__11801_ gnd vdd FILL
XFILL_2__12781_ gnd vdd FILL
XFILL_1__10442_ gnd vdd FILL
XSFILL94360x61050 gnd vdd FILL
XFILL_5__9152_ gnd vdd FILL
XFILL_0__13960_ gnd vdd FILL
XFILL_4_BUFX2_insert280 gnd vdd FILL
XFILL_5__11912_ gnd vdd FILL
XFILL_6__12162_ gnd vdd FILL
XFILL_5__14700_ gnd vdd FILL
XFILL_3__11002_ gnd vdd FILL
XSFILL69000x78050 gnd vdd FILL
XFILL_4__13341_ gnd vdd FILL
XFILL_5__15680_ gnd vdd FILL
X_14066_ _8930_/Q gnd _14068_/A vdd INVX1
X_11278_ _11278_/A _11278_/B gnd _11278_/Y vdd NOR2X1
XFILL_4_BUFX2_insert291 gnd vdd FILL
XFILL_5__12892_ gnd vdd FILL
XFILL_2__14520_ gnd vdd FILL
XFILL_4__10553_ gnd vdd FILL
XFILL_5_BUFX2_insert1004 gnd vdd FILL
XFILL_5__8103_ gnd vdd FILL
XFILL_0__12911_ gnd vdd FILL
XFILL_1__13161_ gnd vdd FILL
XFILL_5_BUFX2_insert1015 gnd vdd FILL
XFILL_2__9374_ gnd vdd FILL
XFILL_2__11732_ gnd vdd FILL
XFILL_5_BUFX2_insert1026 gnd vdd FILL
XFILL_1__10373_ gnd vdd FILL
XFILL_6__11113_ gnd vdd FILL
XFILL_5_BUFX2_insert1037 gnd vdd FILL
X_13017_ _6892_/A gnd _13017_/Y vdd INVX1
X_10229_ _10229_/Q _7537_/CLK _7537_/R vdd _10197_/Y gnd vdd DFFSR
XFILL_0__13891_ gnd vdd FILL
XFILL_5__9083_ gnd vdd FILL
XFILL_5__14631_ gnd vdd FILL
XFILL_5_BUFX2_insert1048 gnd vdd FILL
XFILL_3__15810_ gnd vdd FILL
XFILL_4__16060_ gnd vdd FILL
XFILL_5__11843_ gnd vdd FILL
XSFILL103720x80050 gnd vdd FILL
XFILL_4__13272_ gnd vdd FILL
XFILL_1__12112_ gnd vdd FILL
XFILL_2__8325_ gnd vdd FILL
XFILL_2__14451_ gnd vdd FILL
XFILL_5_BUFX2_insert1059 gnd vdd FILL
XFILL_0__15630_ gnd vdd FILL
XFILL_2__11663_ gnd vdd FILL
XFILL_0__12842_ gnd vdd FILL
XFILL_1__13092_ gnd vdd FILL
XFILL_4__15011_ gnd vdd FILL
XFILL_0__7340_ gnd vdd FILL
XSFILL64040x7050 gnd vdd FILL
XFILL_5__14562_ gnd vdd FILL
XFILL_3_BUFX2_insert980 gnd vdd FILL
XFILL_4__12223_ gnd vdd FILL
XFILL_3_BUFX2_insert991 gnd vdd FILL
XSFILL74120x69050 gnd vdd FILL
XFILL_2__13402_ gnd vdd FILL
XFILL_2__10614_ gnd vdd FILL
XFILL_5__11774_ gnd vdd FILL
XFILL_3__15741_ gnd vdd FILL
XFILL_2__8256_ gnd vdd FILL
XFILL_1__12043_ gnd vdd FILL
XFILL_3__12953_ gnd vdd FILL
XFILL_2__14382_ gnd vdd FILL
XFILL_0__15561_ gnd vdd FILL
XFILL_2__11594_ gnd vdd FILL
XFILL_0__12773_ gnd vdd FILL
XFILL_5__16301_ gnd vdd FILL
XFILL_5__13513_ gnd vdd FILL
XFILL_5__14493_ gnd vdd FILL
XFILL_2__7207_ gnd vdd FILL
XFILL_2__16121_ gnd vdd FILL
XFILL_3__11904_ gnd vdd FILL
X_14968_ _9973_/Q _13751_/C _14968_/C gnd _14976_/B vdd AOI21X1
XFILL_4__12154_ gnd vdd FILL
XFILL_2__13333_ gnd vdd FILL
XFILL_3__15672_ gnd vdd FILL
XSFILL49720x64050 gnd vdd FILL
XFILL_0__14512_ gnd vdd FILL
XFILL_2__10545_ gnd vdd FILL
XFILL_2__8187_ gnd vdd FILL
XFILL_0__11724_ gnd vdd FILL
XFILL_0__9010_ gnd vdd FILL
XFILL_3__12884_ gnd vdd FILL
XFILL_0__15492_ gnd vdd FILL
XFILL_5__9985_ gnd vdd FILL
XFILL_5__16232_ gnd vdd FILL
XSFILL89320x50050 gnd vdd FILL
XFILL_5__13444_ gnd vdd FILL
XSFILL53960x27050 gnd vdd FILL
XFILL_4__11105_ gnd vdd FILL
X_13919_ _13919_/A gnd _13919_/Y vdd INVX1
XFILL_3__14623_ gnd vdd FILL
XFILL_5__10656_ gnd vdd FILL
X_6850_ _6850_/A gnd memoryAddress[12] vdd BUFX2
XFILL_2__13264_ gnd vdd FILL
XFILL_4__12085_ gnd vdd FILL
XFILL_1__15802_ gnd vdd FILL
XFILL_2__16052_ gnd vdd FILL
XFILL_3_BUFX2_insert1030 gnd vdd FILL
X_14899_ _7888_/A gnd _16272_/A vdd INVX1
XFILL_3__11835_ gnd vdd FILL
XSFILL109480x56050 gnd vdd FILL
XFILL_3_BUFX2_insert1041 gnd vdd FILL
XSFILL59000x50 gnd vdd FILL
XFILL_0__14443_ gnd vdd FILL
XFILL_1__13994_ gnd vdd FILL
XFILL_3_BUFX2_insert1052 gnd vdd FILL
XFILL_0__11655_ gnd vdd FILL
XSFILL13800x9050 gnd vdd FILL
XFILL_5__16163_ gnd vdd FILL
XFILL_4__15913_ gnd vdd FILL
XFILL_5__13375_ gnd vdd FILL
XFILL_2__15003_ gnd vdd FILL
XFILL_2__12215_ gnd vdd FILL
XFILL_4__11036_ gnd vdd FILL
XFILL_3_BUFX2_insert1063 gnd vdd FILL
XFILL_3__14554_ gnd vdd FILL
XFILL_2__7069_ gnd vdd FILL
XFILL_3__7951_ gnd vdd FILL
XFILL_3_BUFX2_insert1085 gnd vdd FILL
XSFILL54040x36050 gnd vdd FILL
XFILL_1__15733_ gnd vdd FILL
XFILL_3__11766_ gnd vdd FILL
XFILL_0__14374_ gnd vdd FILL
XFILL_5__15114_ gnd vdd FILL
X_8520_ _8440_/B _7496_/B gnd _8521_/C vdd NAND2X1
XFILL_0__11586_ gnd vdd FILL
XFILL_5__8867_ gnd vdd FILL
XFILL_5__12326_ gnd vdd FILL
XFILL_5__16094_ gnd vdd FILL
XFILL_3__13505_ gnd vdd FILL
XFILL_3__6902_ gnd vdd FILL
XFILL_0__16113_ gnd vdd FILL
XFILL_4__15844_ gnd vdd FILL
XFILL_2__12146_ gnd vdd FILL
XFILL_3__14485_ gnd vdd FILL
XFILL_0__13325_ gnd vdd FILL
XFILL_1__15664_ gnd vdd FILL
XFILL_3__7882_ gnd vdd FILL
XFILL_5__7818_ gnd vdd FILL
XFILL_1__12876_ gnd vdd FILL
XFILL_3__11697_ gnd vdd FILL
XFILL_0__10537_ gnd vdd FILL
XFILL_5_BUFX2_insert508 gnd vdd FILL
XFILL_5__15045_ gnd vdd FILL
XFILL_0__9912_ gnd vdd FILL
XFILL_6__7591_ gnd vdd FILL
XFILL_3__16224_ gnd vdd FILL
X_8451_ _8460_/A _9347_/B gnd _8451_/Y vdd NAND2X1
XFILL_5_BUFX2_insert519 gnd vdd FILL
XFILL_5__12257_ gnd vdd FILL
XFILL_4__15775_ gnd vdd FILL
XFILL_3__9621_ gnd vdd FILL
XFILL_3__13436_ gnd vdd FILL
XSFILL43880x79050 gnd vdd FILL
XFILL_0__16044_ gnd vdd FILL
XFILL_1__14615_ gnd vdd FILL
XFILL_2__12077_ gnd vdd FILL
XFILL_3__10648_ gnd vdd FILL
XFILL_4__12987_ gnd vdd FILL
XFILL_1__11827_ gnd vdd FILL
XFILL_0__13256_ gnd vdd FILL
XFILL_0_BUFX2_insert870 gnd vdd FILL
X_7402_ _7402_/Q _9705_/CLK _7914_/R vdd _7402_/D gnd vdd DFFSR
XFILL_1__15595_ gnd vdd FILL
XFILL_5__11208_ gnd vdd FILL
XFILL_5__7749_ gnd vdd FILL
XFILL_4__14726_ gnd vdd FILL
X_8382_ _8430_/Q gnd _8384_/A vdd INVX1
XFILL_2__15905_ gnd vdd FILL
XFILL_5__12188_ gnd vdd FILL
XFILL_4__11938_ gnd vdd FILL
XFILL_0_BUFX2_insert881 gnd vdd FILL
XFILL_2__11028_ gnd vdd FILL
XFILL_3__16155_ gnd vdd FILL
XFILL_0_BUFX2_insert892 gnd vdd FILL
XSFILL18680x55050 gnd vdd FILL
XFILL_3__13367_ gnd vdd FILL
XFILL_0__12207_ gnd vdd FILL
XSFILL48920x16050 gnd vdd FILL
XFILL_3__9552_ gnd vdd FILL
XFILL_1__14546_ gnd vdd FILL
XFILL_3__10579_ gnd vdd FILL
XFILL_1__11758_ gnd vdd FILL
XSFILL74200x49050 gnd vdd FILL
X_7333_ _7331_/Y _7359_/A _7333_/C gnd _7397_/D vdd OAI21X1
XFILL_3_BUFX2_insert30 gnd vdd FILL
XFILL_0__10399_ gnd vdd FILL
XFILL_5__11139_ gnd vdd FILL
XFILL_3__15106_ gnd vdd FILL
XFILL_3__8503_ gnd vdd FILL
XFILL_0__9774_ gnd vdd FILL
XFILL_4__14657_ gnd vdd FILL
XFILL_3__12318_ gnd vdd FILL
XFILL_0__6986_ gnd vdd FILL
XFILL_3_BUFX2_insert41 gnd vdd FILL
XFILL_4__11869_ gnd vdd FILL
XFILL_2__15836_ gnd vdd FILL
XFILL_1__10709_ gnd vdd FILL
XFILL_3__16086_ gnd vdd FILL
XFILL_3__9483_ gnd vdd FILL
XFILL_3__13298_ gnd vdd FILL
XFILL_1__14477_ gnd vdd FILL
XFILL_0__12138_ gnd vdd FILL
XFILL_5__9419_ gnd vdd FILL
XFILL_3_BUFX2_insert52 gnd vdd FILL
XFILL_3_BUFX2_insert63 gnd vdd FILL
XFILL_1__11689_ gnd vdd FILL
XFILL_3_BUFX2_insert74 gnd vdd FILL
XFILL_4__13608_ gnd vdd FILL
XFILL_0__8725_ gnd vdd FILL
XSFILL49000x25050 gnd vdd FILL
XFILL_3__15037_ gnd vdd FILL
XFILL_5__15947_ gnd vdd FILL
X_7264_ _7188_/A _7535_/CLK _8682_/R vdd _7264_/D gnd vdd DFFSR
XFILL_4__14588_ gnd vdd FILL
XFILL_1__16216_ gnd vdd FILL
XFILL_1__13428_ gnd vdd FILL
XFILL_3_BUFX2_insert85 gnd vdd FILL
XFILL_3__12249_ gnd vdd FILL
XFILL_3_BUFX2_insert96 gnd vdd FILL
XFILL_2__15767_ gnd vdd FILL
XFILL_6__8143_ gnd vdd FILL
XFILL_0__12069_ gnd vdd FILL
XFILL_2__12979_ gnd vdd FILL
X_9003_ _9001_/Y _9005_/A _9002_/Y gnd _9063_/D vdd OAI21X1
XFILL_4__16327_ gnd vdd FILL
XFILL_4__13539_ gnd vdd FILL
XFILL_0__8656_ gnd vdd FILL
X_7195_ _7207_/A _7579_/B gnd _7196_/C vdd NAND2X1
XFILL_2__14718_ gnd vdd FILL
XFILL_5__15878_ gnd vdd FILL
XFILL_1__13359_ gnd vdd FILL
XFILL_3__8365_ gnd vdd FILL
XFILL_1__16147_ gnd vdd FILL
XSFILL38840x68050 gnd vdd FILL
XFILL_2__15698_ gnd vdd FILL
XFILL112360x75050 gnd vdd FILL
XFILL_0__7607_ gnd vdd FILL
XFILL_5__14829_ gnd vdd FILL
XFILL_1__7380_ gnd vdd FILL
XSFILL54120x16050 gnd vdd FILL
XFILL_4__16258_ gnd vdd FILL
XFILL_0__8587_ gnd vdd FILL
XFILL_3__7316_ gnd vdd FILL
XFILL_2__14649_ gnd vdd FILL
XFILL_1__16078_ gnd vdd FILL
XFILL_0__15828_ gnd vdd FILL
XFILL_4__15209_ gnd vdd FILL
XFILL_2_BUFX2_insert409 gnd vdd FILL
XFILL_4__16189_ gnd vdd FILL
XFILL_1__15029_ gnd vdd FILL
XFILL_3__15939_ gnd vdd FILL
XFILL_3__7247_ gnd vdd FILL
XSFILL79320x82050 gnd vdd FILL
XSFILL43960x59050 gnd vdd FILL
XFILL_0__15759_ gnd vdd FILL
X_9905_ _9903_/Y _9896_/B _9905_/C gnd _9961_/D vdd OAI21X1
XFILL_2__16319_ gnd vdd FILL
XFILL_0__7469_ gnd vdd FILL
XFILL_3__7178_ gnd vdd FILL
XFILL_1__8001_ gnd vdd FILL
XFILL_0__9208_ gnd vdd FILL
XFILL_6__8976_ gnd vdd FILL
XSFILL18760x35050 gnd vdd FILL
XSFILL8600x45050 gnd vdd FILL
X_9836_ _9836_/Q _7020_/CLK _8053_/R vdd _9836_/D gnd vdd DFFSR
XSFILL44040x68050 gnd vdd FILL
XFILL_4__7991_ gnd vdd FILL
XFILL_6__7927_ gnd vdd FILL
XFILL_0__9139_ gnd vdd FILL
X_9767_ _9789_/B _7975_/B gnd _9767_/Y vdd NAND2X1
XFILL_4__9730_ gnd vdd FILL
X_6979_ _6979_/A _6982_/B _6979_/C gnd _7023_/D vdd OAI21X1
XFILL_4__6942_ gnd vdd FILL
XFILL_6_BUFX2_insert331 gnd vdd FILL
XBUFX2_insert408 _10920_/Y gnd _12380_/A vdd BUFX2
X_8718_ _8718_/A gnd _8718_/Y vdd INVX1
XBUFX2_insert419 _14991_/Y gnd _15044_/C vdd BUFX2
X_9698_ _9698_/Q _8680_/CLK _8418_/R vdd _9628_/Y gnd vdd DFFSR
XFILL_4__9661_ gnd vdd FILL
XSFILL109640x16050 gnd vdd FILL
XFILL_4__6873_ gnd vdd FILL
XFILL_1__8903_ gnd vdd FILL
X_10580_ _10581_/B _9172_/B gnd _10580_/Y vdd NAND2X1
X_8649_ _8647_/Y _8607_/B _8649_/C gnd _8689_/D vdd OAI21X1
XFILL_4__8612_ gnd vdd FILL
XSFILL38920x48050 gnd vdd FILL
XFILL_1__9883_ gnd vdd FILL
XFILL112440x55050 gnd vdd FILL
XFILL_4__9592_ gnd vdd FILL
XFILL_1__8834_ gnd vdd FILL
X_12250_ _12247_/Y _12250_/B _12250_/C gnd _12250_/Y vdd NAND3X1
XSFILL39000x57050 gnd vdd FILL
XFILL_1__8765_ gnd vdd FILL
X_11201_ _12204_/Y _12334_/Y gnd _11201_/Y vdd NOR2X1
XFILL_4__8474_ gnd vdd FILL
X_12181_ _13145_/A gnd _12183_/A vdd INVX1
XFILL_1__7716_ gnd vdd FILL
XFILL_4__7425_ gnd vdd FILL
XFILL_1__8696_ gnd vdd FILL
X_11132_ _11300_/A gnd _11149_/A vdd INVX1
XSFILL18840x15050 gnd vdd FILL
XSFILL94280x76050 gnd vdd FILL
XSFILL44120x48050 gnd vdd FILL
XFILL_4__7356_ gnd vdd FILL
X_15940_ _14515_/A _15940_/B gnd _15940_/Y vdd NOR2X1
XFILL_3_BUFX2_insert232 gnd vdd FILL
X_11063_ _12266_/Y gnd _11063_/Y vdd INVX1
XSFILL69080x52050 gnd vdd FILL
XFILL_3_BUFX2_insert243 gnd vdd FILL
XSFILL99320x13050 gnd vdd FILL
XFILL_3_BUFX2_insert254 gnd vdd FILL
XFILL_1__7578_ gnd vdd FILL
XSFILL85080x7050 gnd vdd FILL
XFILL_3_BUFX2_insert265 gnd vdd FILL
X_10014_ _10066_/B _7326_/B gnd _10014_/Y vdd NAND2X1
XFILL_4__7287_ gnd vdd FILL
XFILL_3_BUFX2_insert276 gnd vdd FILL
XFILL_3_BUFX2_insert287 gnd vdd FILL
XFILL_2__8110_ gnd vdd FILL
X_15871_ _15871_/A _15870_/Y gnd _15877_/A vdd NOR2X1
XFILL_2__9090_ gnd vdd FILL
XFILL_3_BUFX2_insert298 gnd vdd FILL
XSFILL73560x77050 gnd vdd FILL
XFILL_2_BUFX2_insert910 gnd vdd FILL
XFILL_4__9026_ gnd vdd FILL
XSFILL104280x61050 gnd vdd FILL
XFILL_2_BUFX2_insert921 gnd vdd FILL
XSFILL23800x4050 gnd vdd FILL
X_14822_ _14820_/Y _14821_/Y _14819_/Y gnd _14833_/B vdd NAND3X1
XFILL_2_BUFX2_insert932 gnd vdd FILL
XFILL_1__9248_ gnd vdd FILL
XFILL_2_BUFX2_insert943 gnd vdd FILL
XFILL_2_BUFX2_insert954 gnd vdd FILL
XFILL_2_BUFX2_insert965 gnd vdd FILL
XFILL_5__10510_ gnd vdd FILL
XFILL_2_BUFX2_insert976 gnd vdd FILL
XSFILL23800x70050 gnd vdd FILL
X_14753_ _14753_/A _14753_/B gnd _14754_/C vdd NOR2X1
X_11965_ _13157_/A gnd _11967_/A vdd INVX1
XFILL_5__11490_ gnd vdd FILL
XFILL_2_BUFX2_insert987 gnd vdd FILL
XSFILL89240x65050 gnd vdd FILL
XFILL_2_BUFX2_insert998 gnd vdd FILL
XFILL_5__9770_ gnd vdd FILL
X_13704_ _14946_/A _13704_/B _14768_/D _13704_/D gnd _13705_/B vdd OAI22X1
X_10916_ _10898_/Y _10906_/Y gnd _10944_/B vdd NAND2X1
XFILL_5__6982_ gnd vdd FILL
XFILL_5__10441_ gnd vdd FILL
X_14684_ _8687_/Q gnd _16083_/C vdd INVX1
XFILL_3__11620_ gnd vdd FILL
X_11896_ _11896_/A gnd _11896_/Y vdd INVX1
XFILL_2__10261_ gnd vdd FILL
XSFILL3720x68050 gnd vdd FILL
XFILL_2__9992_ gnd vdd FILL
XFILL_5__8721_ gnd vdd FILL
XFILL_0__11440_ gnd vdd FILL
XFILL_4__9928_ gnd vdd FILL
X_16423_ _16339_/A _8165_/CLK _8165_/R vdd _16423_/D gnd vdd DFFSR
XFILL_1__10991_ gnd vdd FILL
X_13635_ _13635_/A _13635_/B _13634_/Y gnd _13636_/B vdd NAND3X1
XFILL_4__12910_ gnd vdd FILL
XFILL_2__12000_ gnd vdd FILL
XFILL_5__13160_ gnd vdd FILL
XFILL_5__10372_ gnd vdd FILL
X_10847_ _13922_/A _7007_/CLK _9332_/R vdd _10847_/D gnd vdd DFFSR
XFILL_1__12730_ gnd vdd FILL
XFILL_3__11551_ gnd vdd FILL
XFILL_4__13890_ gnd vdd FILL
XSFILL94360x56050 gnd vdd FILL
XFILL_0_BUFX2_insert100 gnd vdd FILL
XFILL_2__10192_ gnd vdd FILL
XFILL_5__8652_ gnd vdd FILL
XFILL_4__9859_ gnd vdd FILL
XFILL_5__12111_ gnd vdd FILL
XBUFX2_insert920 _15069_/Y gnd _15848_/A vdd BUFX2
XFILL_0__11371_ gnd vdd FILL
X_16354_ _13980_/A gnd _16356_/A vdd INVX1
XBUFX2_insert931 _12435_/Y gnd _8401_/B vdd BUFX2
XFILL_4__12841_ gnd vdd FILL
XFILL_5__13091_ gnd vdd FILL
XBUFX2_insert942 _12426_/Y gnd _8136_/B vdd BUFX2
XFILL_3__10502_ gnd vdd FILL
X_13566_ _13564_/Y _14317_/C _13587_/C _13565_/Y gnd _13567_/B vdd OAI22X1
X_10778_ _10778_/A gnd _10778_/Y vdd INVX1
XFILL_0__13110_ gnd vdd FILL
XBUFX2_insert953 _13365_/Y gnd _10822_/B vdd BUFX2
XFILL_3__14270_ gnd vdd FILL
XFILL_1__12661_ gnd vdd FILL
XBUFX2_insert964 _13361_/Y gnd _10372_/B vdd BUFX2
XFILL_0__10322_ gnd vdd FILL
XFILL_2__8874_ gnd vdd FILL
XFILL_5__7603_ gnd vdd FILL
XFILL_3__11482_ gnd vdd FILL
X_15305_ _15662_/A _7560_/A _7432_/A _15383_/D gnd _15305_/Y vdd AOI22X1
XSFILL69160x32050 gnd vdd FILL
XFILL_0__14090_ gnd vdd FILL
X_12517_ _12091_/B gnd _12519_/A vdd INVX1
XBUFX2_insert975 _16451_/Y gnd _13155_/A vdd BUFX2
XFILL_5__12042_ gnd vdd FILL
XFILL_5__8583_ gnd vdd FILL
XFILL_3__13221_ gnd vdd FILL
XBUFX2_insert986 _13351_/Y gnd _9975_/B vdd BUFX2
XFILL_4__15560_ gnd vdd FILL
X_16285_ _15969_/C _7763_/A _8147_/A _16011_/D gnd _16285_/Y vdd AOI22X1
XFILL_4__12772_ gnd vdd FILL
XBUFX2_insert997 _14998_/Y gnd _15563_/A vdd BUFX2
XFILL_1__14400_ gnd vdd FILL
XFILL_1__11612_ gnd vdd FILL
XFILL_3__10433_ gnd vdd FILL
X_13497_ _13497_/A gnd _13497_/Y vdd INVX1
XFILL_2__7825_ gnd vdd FILL
XFILL_1__15380_ gnd vdd FILL
XFILL_2__13951_ gnd vdd FILL
XFILL_0__13041_ gnd vdd FILL
XFILL_1__12592_ gnd vdd FILL
XFILL_0__10253_ gnd vdd FILL
X_15236_ _16235_/A _15235_/Y _13679_/Y _16225_/C gnd _15236_/Y vdd OAI22X1
XFILL_4__14511_ gnd vdd FILL
X_12448_ _12352_/A gnd _12448_/Y vdd INVX1
XFILL_0__6840_ gnd vdd FILL
XSFILL104360x41050 gnd vdd FILL
XFILL_4__11723_ gnd vdd FILL
XFILL_3__13152_ gnd vdd FILL
XFILL_2__12902_ gnd vdd FILL
XFILL_1__14331_ gnd vdd FILL
XFILL_3__10364_ gnd vdd FILL
XFILL_4__15491_ gnd vdd FILL
XFILL_2__7756_ gnd vdd FILL
XFILL_1__11543_ gnd vdd FILL
XFILL_2__13882_ gnd vdd FILL
XFILL_0__10184_ gnd vdd FILL
XFILL_5__15801_ gnd vdd FILL
XFILL_5__7465_ gnd vdd FILL
XSFILL74280x23050 gnd vdd FILL
XFILL_3__12103_ gnd vdd FILL
XFILL_4__14442_ gnd vdd FILL
X_15167_ _15167_/A _15167_/B _14791_/C gnd _15167_/Y vdd AOI21X1
XFILL_2__15621_ gnd vdd FILL
X_12379_ _12035_/B gnd _12381_/A vdd INVX1
XFILL_4__11654_ gnd vdd FILL
XFILL_3__10295_ gnd vdd FILL
XFILL_1__14262_ gnd vdd FILL
XFILL_2__12833_ gnd vdd FILL
XFILL_5__13993_ gnd vdd FILL
XFILL_3__13083_ gnd vdd FILL
XFILL_1__11474_ gnd vdd FILL
XFILL_2__7687_ gnd vdd FILL
XFILL_0__8510_ gnd vdd FILL
XFILL_0__14992_ gnd vdd FILL
X_14118_ _14118_/A _13630_/B _13479_/C _14118_/D gnd _14119_/B vdd OAI22X1
XFILL_5__15732_ gnd vdd FILL
XSFILL89320x45050 gnd vdd FILL
XFILL_1__13213_ gnd vdd FILL
XFILL_1__16001_ gnd vdd FILL
XFILL_3__12034_ gnd vdd FILL
X_15098_ _15025_/B gnd _15978_/B vdd INVX4
XFILL_4__14373_ gnd vdd FILL
XFILL_0__9490_ gnd vdd FILL
XFILL_2__9426_ gnd vdd FILL
XFILL_2__15552_ gnd vdd FILL
XFILL_1__10425_ gnd vdd FILL
XFILL_4__11585_ gnd vdd FILL
XFILL_2__12764_ gnd vdd FILL
XFILL_1__14193_ gnd vdd FILL
XFILL_5__9135_ gnd vdd FILL
XFILL_0__13943_ gnd vdd FILL
XFILL_4__16112_ gnd vdd FILL
XFILL_4__13324_ gnd vdd FILL
X_14049_ _9442_/Q gnd _14049_/Y vdd INVX1
XFILL_0__8441_ gnd vdd FILL
XFILL_4__10536_ gnd vdd FILL
XFILL_5__15663_ gnd vdd FILL
XFILL_2__14503_ gnd vdd FILL
XFILL_5__12875_ gnd vdd FILL
XFILL_2__9357_ gnd vdd FILL
XFILL_1__13144_ gnd vdd FILL
XFILL_2__11715_ gnd vdd FILL
XFILL_2__15483_ gnd vdd FILL
XFILL_2__12695_ gnd vdd FILL
XFILL_0__13874_ gnd vdd FILL
XFILL_5__14614_ gnd vdd FILL
XFILL_4__16043_ gnd vdd FILL
XFILL_5__11826_ gnd vdd FILL
XFILL_0__8372_ gnd vdd FILL
XFILL_3__7101_ gnd vdd FILL
XFILL_4__13255_ gnd vdd FILL
XSFILL94440x36050 gnd vdd FILL
XFILL_5__15594_ gnd vdd FILL
XFILL_2__14434_ gnd vdd FILL
XFILL_0__15613_ gnd vdd FILL
XFILL_3__13985_ gnd vdd FILL
XFILL_0__12825_ gnd vdd FILL
XFILL_2__9288_ gnd vdd FILL
XFILL_2__11646_ gnd vdd FILL
XFILL_3__8081_ gnd vdd FILL
XFILL_5__8017_ gnd vdd FILL
XFILL_1__10287_ gnd vdd FILL
XFILL_0__7323_ gnd vdd FILL
XFILL_4__12206_ gnd vdd FILL
X_7951_ _7937_/B _9615_/B gnd _7952_/C vdd NAND2X1
XFILL_3__15724_ gnd vdd FILL
XFILL_5__14545_ gnd vdd FILL
XFILL_5__11757_ gnd vdd FILL
XFILL_3__7032_ gnd vdd FILL
XFILL_1__12026_ gnd vdd FILL
XSFILL69240x12050 gnd vdd FILL
XFILL_2__8239_ gnd vdd FILL
XFILL_0__15544_ gnd vdd FILL
XFILL_2__14365_ gnd vdd FILL
XFILL_4__10398_ gnd vdd FILL
XFILL_2__11577_ gnd vdd FILL
XFILL_0__12756_ gnd vdd FILL
X_6902_ _6998_/Q gnd _6902_/Y vdd INVX1
XFILL_5__10708_ gnd vdd FILL
XFILL_5__14476_ gnd vdd FILL
XFILL_4__12137_ gnd vdd FILL
XFILL_2__16104_ gnd vdd FILL
XFILL_2__13316_ gnd vdd FILL
XFILL_3__15655_ gnd vdd FILL
X_7882_ _7922_/Q gnd _7882_/Y vdd INVX1
XFILL_2__10528_ gnd vdd FILL
XFILL_5__11688_ gnd vdd FILL
XFILL_3__12867_ gnd vdd FILL
XFILL_0__11707_ gnd vdd FILL
XFILL_0__15475_ gnd vdd FILL
XSFILL104440x21050 gnd vdd FILL
XFILL_2__14296_ gnd vdd FILL
XFILL_5__16215_ gnd vdd FILL
XFILL_5__13427_ gnd vdd FILL
XFILL_5__10639_ gnd vdd FILL
XFILL_3__14606_ gnd vdd FILL
XFILL_6__15766_ gnd vdd FILL
XFILL_0__7185_ gnd vdd FILL
X_9621_ _9652_/B _7061_/B gnd _9621_/Y vdd NAND2X1
XFILL_2__16035_ gnd vdd FILL
XFILL_4__12068_ gnd vdd FILL
XFILL_3__11818_ gnd vdd FILL
XFILL_2__13247_ gnd vdd FILL
XFILL_3__15586_ gnd vdd FILL
XFILL_0__14426_ gnd vdd FILL
XFILL_3__8983_ gnd vdd FILL
XFILL_0__11638_ gnd vdd FILL
XFILL_1__13977_ gnd vdd FILL
XFILL_5__13358_ gnd vdd FILL
X_9552_ _9552_/A gnd _9554_/A vdd INVX1
XFILL_5__9899_ gnd vdd FILL
XFILL_4__11019_ gnd vdd FILL
XFILL_5__16146_ gnd vdd FILL
XFILL_3__14537_ gnd vdd FILL
XFILL_1__15716_ gnd vdd FILL
XFILL_3__7934_ gnd vdd FILL
XFILL_3__11749_ gnd vdd FILL
XSFILL59160x64050 gnd vdd FILL
XFILL_0__14357_ gnd vdd FILL
XSFILL89400x25050 gnd vdd FILL
X_8503_ _8503_/A _8503_/B _8502_/Y gnd _8503_/Y vdd OAI21X1
XFILL_5__12309_ gnd vdd FILL
XFILL_0__11569_ gnd vdd FILL
XFILL_5_BUFX2_insert305 gnd vdd FILL
XFILL_5__16077_ gnd vdd FILL
XFILL_5__13289_ gnd vdd FILL
X_9483_ _9565_/Q gnd _9485_/A vdd INVX1
XFILL_4__15827_ gnd vdd FILL
XFILL_0__13308_ gnd vdd FILL
XFILL_3__14468_ gnd vdd FILL
XFILL_5_BUFX2_insert316 gnd vdd FILL
XFILL_2__12129_ gnd vdd FILL
XFILL_1__15647_ gnd vdd FILL
XFILL_3__7865_ gnd vdd FILL
XFILL_5_BUFX2_insert327 gnd vdd FILL
XFILL_5_BUFX2_insert338 gnd vdd FILL
XFILL_1__12859_ gnd vdd FILL
XBUFX2_insert17 _13443_/Y gnd _14506_/C vdd BUFX2
XFILL_0__14288_ gnd vdd FILL
XFILL_3__16207_ gnd vdd FILL
X_8434_ _8394_/A _7662_/CLK _8166_/R vdd _8434_/D gnd vdd DFFSR
XBUFX2_insert28 _13320_/Y gnd _8460_/A vdd BUFX2
XFILL_5__15028_ gnd vdd FILL
XFILL_5_BUFX2_insert349 gnd vdd FILL
XFILL_3__9604_ gnd vdd FILL
XFILL_3__13419_ gnd vdd FILL
XBUFX2_insert39 _13265_/Y gnd _6985_/B vdd BUFX2
XFILL_0__16027_ gnd vdd FILL
XFILL_1__6880_ gnd vdd FILL
XFILL_4__15758_ gnd vdd FILL
XFILL_0__13239_ gnd vdd FILL
XFILL_3__14399_ gnd vdd FILL
XFILL_1__15578_ gnd vdd FILL
XSFILL94520x16050 gnd vdd FILL
XSFILL13640x20050 gnd vdd FILL
XFILL_4__14709_ gnd vdd FILL
X_8365_ _8365_/A _9005_/B gnd _8366_/C vdd NAND2X1
XSFILL79080x15050 gnd vdd FILL
XFILL_3__16138_ gnd vdd FILL
XFILL_4__15689_ gnd vdd FILL
XFILL_3__9535_ gnd vdd FILL
XSFILL24280x71050 gnd vdd FILL
XFILL_1__14529_ gnd vdd FILL
XSFILL39080x31050 gnd vdd FILL
X_7316_ _7316_/A gnd _7318_/A vdd INVX1
XFILL_0__9757_ gnd vdd FILL
XFILL_0__6969_ gnd vdd FILL
XFILL_2__15819_ gnd vdd FILL
X_8296_ _8236_/A _7912_/CLK _7911_/R vdd _8238_/Y gnd vdd DFFSR
XFILL_3__16069_ gnd vdd FILL
XFILL_3__9466_ gnd vdd FILL
XFILL_1__7501_ gnd vdd FILL
XFILL_0__8708_ gnd vdd FILL
X_7247_ _7245_/Y _7168_/A _7247_/C gnd _7283_/D vdd OAI21X1
XFILL_1__8481_ gnd vdd FILL
XFILL_4__7210_ gnd vdd FILL
XFILL_3__9397_ gnd vdd FILL
XFILL_4__8190_ gnd vdd FILL
XFILL_0__8639_ gnd vdd FILL
XFILL_1__7432_ gnd vdd FILL
XSFILL33800x33050 gnd vdd FILL
X_7178_ _7178_/A _7184_/B _7177_/Y gnd _7260_/D vdd OAI21X1
XFILL_3__8348_ gnd vdd FILL
XFILL_1__7363_ gnd vdd FILL
XFILL_4__7072_ gnd vdd FILL
XFILL_2_BUFX2_insert228 gnd vdd FILL
XFILL_1__9102_ gnd vdd FILL
XSFILL19240x60050 gnd vdd FILL
XFILL_2_BUFX2_insert239 gnd vdd FILL
XFILL_1__7294_ gnd vdd FILL
XFILL_1__9033_ gnd vdd FILL
XFILL_1_BUFX2_insert906 gnd vdd FILL
XFILL_1_BUFX2_insert917 gnd vdd FILL
XFILL_1_BUFX2_insert928 gnd vdd FILL
XFILL112040x52050 gnd vdd FILL
X_11750_ _11257_/Y _11386_/Y gnd _11750_/Y vdd AND2X2
XFILL_1_BUFX2_insert939 gnd vdd FILL
X_9819_ _9733_/A _8679_/CLK _7131_/R vdd _9819_/D gnd vdd DFFSR
XFILL_4__7974_ gnd vdd FILL
X_10701_ _10739_/Q gnd _10701_/Y vdd INVX1
X_11681_ _11278_/Y _11681_/B gnd _11681_/Y vdd NAND2X1
XFILL_4__6925_ gnd vdd FILL
XBUFX2_insert227 _12432_/Y gnd _8654_/B vdd BUFX2
X_13420_ _13416_/Y _13420_/B _13420_/C _13417_/Y gnd _13420_/Y vdd OAI22X1
X_10632_ _10716_/Q gnd _10632_/Y vdd INVX1
XBUFX2_insert238 _12348_/Y gnd _9466_/B vdd BUFX2
XFILL_1__9935_ gnd vdd FILL
XSFILL114600x66050 gnd vdd FILL
XBUFX2_insert249 _10922_/Y gnd _14402_/C vdd BUFX2
XFILL_4__9644_ gnd vdd FILL
XFILL_4__6856_ gnd vdd FILL
X_13351_ _13351_/A _13348_/Y gnd _13351_/Y vdd NOR2X1
X_10563_ _10563_/A _10548_/B _10562_/Y gnd _10607_/D vdd OAI21X1
XSFILL69080x47050 gnd vdd FILL
XFILL_5_CLKBUF1_insert117 gnd vdd FILL
XFILL_1__9866_ gnd vdd FILL
XFILL_5_BUFX2_insert850 gnd vdd FILL
XFILL_5_CLKBUF1_insert128 gnd vdd FILL
X_12302_ _12302_/A _12300_/Y _12302_/C gnd _12302_/Y vdd NAND3X1
XFILL_5_BUFX2_insert861 gnd vdd FILL
XFILL_5_CLKBUF1_insert139 gnd vdd FILL
XFILL_5_BUFX2_insert872 gnd vdd FILL
X_16070_ _16070_/A _15175_/B _16069_/Y gnd _16070_/Y vdd AOI21X1
X_13282_ _13295_/C _13282_/B gnd _13291_/A vdd NAND2X1
XFILL_2__7610_ gnd vdd FILL
XFILL_5_BUFX2_insert883 gnd vdd FILL
X_10494_ _10494_/A _10539_/B _10494_/C gnd _10584_/D vdd OAI21X1
XFILL_5_BUFX2_insert894 gnd vdd FILL
XFILL_2__8590_ gnd vdd FILL
XFILL_4__8526_ gnd vdd FILL
XFILL_1__9797_ gnd vdd FILL
X_15021_ _16232_/B _15636_/B gnd _15197_/B vdd NAND2X1
X_12233_ _6874_/A _12277_/B _12309_/C _12701_/A gnd _12234_/C vdd AOI22X1
XBUFX2_insert1091 rst gnd BUFX2_insert494/A vdd BUFX2
XFILL_1__8748_ gnd vdd FILL
XFILL_4__8457_ gnd vdd FILL
XFILL_5__7250_ gnd vdd FILL
X_12164_ _12134_/A _12871_/A gnd _12165_/C vdd NAND2X1
XFILL_5__10990_ gnd vdd FILL
XFILL_2__7472_ gnd vdd FILL
X_11115_ _11113_/Y _11115_/B gnd _11115_/Y vdd NOR2X1
XFILL_5__7181_ gnd vdd FILL
XFILL_4__8388_ gnd vdd FILL
XFILL_6__10191_ gnd vdd FILL
X_12095_ _12111_/A _11969_/B _12111_/C gnd _12098_/A vdd NAND3X1
XSFILL113800x18050 gnd vdd FILL
XFILL_2__9211_ gnd vdd FILL
XFILL_4__11370_ gnd vdd FILL
XFILL_0__10940_ gnd vdd FILL
XFILL_4__7339_ gnd vdd FILL
XFILL_1__11190_ gnd vdd FILL
X_15923_ _15923_/A _15923_/B gnd _15923_/Y vdd NOR2X1
X_11046_ _12266_/Y _12153_/Y gnd _11046_/Y vdd XOR2X1
XFILL_5__12660_ gnd vdd FILL
XFILL_4__10321_ gnd vdd FILL
XFILL_2__9142_ gnd vdd FILL
XFILL_2__11500_ gnd vdd FILL
XFILL_2__12480_ gnd vdd FILL
XFILL_1__10141_ gnd vdd FILL
XFILL_0__10871_ gnd vdd FILL
XFILL_5__11611_ gnd vdd FILL
X_15854_ _15972_/C gnd _16011_/D vdd INVX2
XFILL_4__13040_ gnd vdd FILL
XFILL_6__13950_ gnd vdd FILL
XFILL_5__12591_ gnd vdd FILL
XFILL_4__10252_ gnd vdd FILL
XFILL_2__11431_ gnd vdd FILL
XFILL_0__12610_ gnd vdd FILL
XFILL_3__13770_ gnd vdd FILL
XFILL_4__9009_ gnd vdd FILL
XFILL_2_BUFX2_insert740 gnd vdd FILL
XFILL_2_BUFX2_insert751 gnd vdd FILL
XFILL_3__10982_ gnd vdd FILL
X_14805_ _8266_/A gnd _14805_/Y vdd INVX1
XFILL_0__13590_ gnd vdd FILL
XFILL_5__14330_ gnd vdd FILL
XSFILL69160x27050 gnd vdd FILL
XFILL_2_BUFX2_insert762 gnd vdd FILL
XFILL_5__11542_ gnd vdd FILL
XFILL_2_BUFX2_insert773 gnd vdd FILL
XFILL_3__12721_ gnd vdd FILL
X_15785_ _15778_/Y _15779_/Y _15785_/C gnd _15786_/A vdd NAND3X1
XSFILL68920x82050 gnd vdd FILL
X_12997_ vdd _12997_/B gnd _12998_/C vdd NAND2X1
XFILL_2__14150_ gnd vdd FILL
XFILL_4__10183_ gnd vdd FILL
XFILL_1__13900_ gnd vdd FILL
XFILL_2_BUFX2_insert784 gnd vdd FILL
XFILL_2__11362_ gnd vdd FILL
XFILL_2_BUFX2_insert795 gnd vdd FILL
XFILL_1__14880_ gnd vdd FILL
XSFILL84200x30050 gnd vdd FILL
XFILL_5__14261_ gnd vdd FILL
X_14736_ _14735_/Y _14045_/A _14872_/C _16104_/B gnd _14737_/B vdd OAI22X1
XFILL_2__13101_ gnd vdd FILL
X_11948_ _11955_/B _12403_/A gnd _11949_/C vdd NAND2X1
XFILL_2__10313_ gnd vdd FILL
XFILL_3__15440_ gnd vdd FILL
XFILL_5__11473_ gnd vdd FILL
XFILL_3__12652_ gnd vdd FILL
XFILL_4__14991_ gnd vdd FILL
XSFILL104360x36050 gnd vdd FILL
XFILL_2__14081_ gnd vdd FILL
XFILL_0_CLKBUF1_insert1079 gnd vdd FILL
XFILL_1__13831_ gnd vdd FILL
XFILL_2__11293_ gnd vdd FILL
XFILL_0__15260_ gnd vdd FILL
XFILL_5__13212_ gnd vdd FILL
XFILL_5__16000_ gnd vdd FILL
XFILL_5__9753_ gnd vdd FILL
XFILL_0__12472_ gnd vdd FILL
XFILL_5__6965_ gnd vdd FILL
XFILL_5__10424_ gnd vdd FILL
XFILL_6__12763_ gnd vdd FILL
XFILL_5__14192_ gnd vdd FILL
XFILL_2__13032_ gnd vdd FILL
XFILL_3__11603_ gnd vdd FILL
X_14667_ _14667_/A _14667_/B _14666_/Y gnd _14668_/B vdd NAND3X1
XFILL_4__13942_ gnd vdd FILL
X_11879_ _11874_/B _11879_/B gnd _11879_/Y vdd NAND2X1
XFILL_3__15371_ gnd vdd FILL
XFILL_0__14211_ gnd vdd FILL
XFILL_2__10244_ gnd vdd FILL
XSFILL79320x4050 gnd vdd FILL
XFILL_5__8704_ gnd vdd FILL
XFILL_3__12583_ gnd vdd FILL
XFILL_2__9975_ gnd vdd FILL
XFILL_0__11423_ gnd vdd FILL
XFILL_1__10974_ gnd vdd FILL
XFILL_0__15191_ gnd vdd FILL
XFILL_1__13762_ gnd vdd FILL
X_16406_ gnd gnd gnd _16406_/Y vdd NAND2X1
X_13618_ _13618_/A _13618_/B gnd _13622_/C vdd NOR2X1
XFILL_5__13143_ gnd vdd FILL
XFILL_5__9684_ gnd vdd FILL
XFILL_3__14322_ gnd vdd FILL
XFILL_5__6896_ gnd vdd FILL
X_14598_ _14598_/A gnd _14598_/Y vdd INVX1
XFILL_4__13873_ gnd vdd FILL
XFILL_1__15501_ gnd vdd FILL
XFILL_3__11534_ gnd vdd FILL
XFILL_0__8990_ gnd vdd FILL
XFILL112200x12050 gnd vdd FILL
XFILL_1__12713_ gnd vdd FILL
XFILL_2__10175_ gnd vdd FILL
XFILL_0__14142_ gnd vdd FILL
XFILL_5__8635_ gnd vdd FILL
XBUFX2_insert750 _13344_/Y gnd _9737_/A vdd BUFX2
XFILL_1__13693_ gnd vdd FILL
XFILL_0__11354_ gnd vdd FILL
XBUFX2_insert761 _13412_/Y gnd _14718_/C vdd BUFX2
X_16337_ gnd gnd gnd _16338_/C vdd NAND2X1
XSFILL74120x82050 gnd vdd FILL
XFILL_4__15612_ gnd vdd FILL
XFILL_4__12824_ gnd vdd FILL
XFILL_0__7941_ gnd vdd FILL
XBUFX2_insert772 _13301_/Y gnd _7814_/A vdd BUFX2
X_13549_ _9468_/A gnd _15157_/B vdd INVX1
XFILL_6__11645_ gnd vdd FILL
XFILL_3__14253_ gnd vdd FILL
XFILL_5__10286_ gnd vdd FILL
XBUFX2_insert783 _10911_/Y gnd _12117_/B vdd BUFX2
XFILL_1__12644_ gnd vdd FILL
XFILL_2__8857_ gnd vdd FILL
XFILL_0__10305_ gnd vdd FILL
XFILL_1__15432_ gnd vdd FILL
XFILL_3__11465_ gnd vdd FILL
XBUFX2_insert794 _13334_/Y gnd _9420_/B vdd BUFX2
XFILL_2__14983_ gnd vdd FILL
XFILL_0__14073_ gnd vdd FILL
XFILL_5__8566_ gnd vdd FILL
XFILL_5__12025_ gnd vdd FILL
XFILL_0__11285_ gnd vdd FILL
XFILL_4__15543_ gnd vdd FILL
X_16268_ _16268_/A _15680_/B _15680_/C gnd _16268_/Y vdd NAND3X1
XFILL_0__7872_ gnd vdd FILL
XFILL_2__7808_ gnd vdd FILL
XFILL_4__12755_ gnd vdd FILL
XFILL_3__10416_ gnd vdd FILL
XFILL_3__14184_ gnd vdd FILL
XFILL_0__13024_ gnd vdd FILL
XFILL_2__13934_ gnd vdd FILL
XFILL_1__12575_ gnd vdd FILL
XFILL_1__15363_ gnd vdd FILL
XFILL_3__11396_ gnd vdd FILL
XFILL_3__7581_ gnd vdd FILL
XFILL_0__10236_ gnd vdd FILL
XFILL_2__8788_ gnd vdd FILL
XFILL_0__9611_ gnd vdd FILL
X_15219_ _15219_/A _15218_/Y _15219_/C gnd _15230_/B vdd NAND3X1
XSFILL53960x40050 gnd vdd FILL
X_8150_ _8150_/Q _8022_/CLK _9046_/R vdd _8150_/D gnd vdd DFFSR
XFILL_5__8497_ gnd vdd FILL
XFILL_4__11706_ gnd vdd FILL
XFILL_6__10527_ gnd vdd FILL
X_16199_ _15169_/D _16198_/Y _16199_/C _16199_/D gnd _16200_/B vdd OAI22X1
XFILL_3__13135_ gnd vdd FILL
XFILL_4__15474_ gnd vdd FILL
XFILL_2__7739_ gnd vdd FILL
XFILL_1__14314_ gnd vdd FILL
XFILL_1__11526_ gnd vdd FILL
XFILL_2__13865_ gnd vdd FILL
XFILL_1__15294_ gnd vdd FILL
X_7101_ _7099_/Y _7100_/A _7101_/C gnd _7101_/Y vdd OAI21X1
XFILL_0__10167_ gnd vdd FILL
XFILL_5__7448_ gnd vdd FILL
XFILL_0__9542_ gnd vdd FILL
XFILL_4__14425_ gnd vdd FILL
XFILL_4__11637_ gnd vdd FILL
X_8081_ _8159_/Q gnd _8081_/Y vdd INVX1
XFILL_2__15604_ gnd vdd FILL
XFILL_3__9251_ gnd vdd FILL
XFILL_1__14245_ gnd vdd FILL
XFILL_5__13976_ gnd vdd FILL
XFILL_3__10278_ gnd vdd FILL
XFILL_1__11457_ gnd vdd FILL
XFILL_2__13796_ gnd vdd FILL
XFILL_5__15715_ gnd vdd FILL
X_7032_ _7030_/Y _7068_/B _7032_/C gnd _7126_/D vdd OAI21X1
XFILL_5__7379_ gnd vdd FILL
XFILL_0__14975_ gnd vdd FILL
XSFILL104440x16050 gnd vdd FILL
XFILL_0__9473_ gnd vdd FILL
XFILL_3__12017_ gnd vdd FILL
XFILL_3__8202_ gnd vdd FILL
XFILL_4__14356_ gnd vdd FILL
XFILL_2__9409_ gnd vdd FILL
XFILL_1__10408_ gnd vdd FILL
XFILL_2__15535_ gnd vdd FILL
XFILL_4__11568_ gnd vdd FILL
XFILL_2__12747_ gnd vdd FILL
XFILL_1__14176_ gnd vdd FILL
XSFILL33720x48050 gnd vdd FILL
XFILL_5__9118_ gnd vdd FILL
XFILL_1__11388_ gnd vdd FILL
XFILL_0__13926_ gnd vdd FILL
XFILL_4__13307_ gnd vdd FILL
XFILL_5__15646_ gnd vdd FILL
XFILL_4__10519_ gnd vdd FILL
XFILL_1__13127_ gnd vdd FILL
XFILL_5__12858_ gnd vdd FILL
XFILL_3__8133_ gnd vdd FILL
XFILL_4__14287_ gnd vdd FILL
XFILL_4__11499_ gnd vdd FILL
XFILL_2__15466_ gnd vdd FILL
XFILL_0__13857_ gnd vdd FILL
XFILL_4__16026_ gnd vdd FILL
XSFILL59160x59050 gnd vdd FILL
XFILL_4__13238_ gnd vdd FILL
XFILL_0__8355_ gnd vdd FILL
XFILL_5__11809_ gnd vdd FILL
XFILL_5__15577_ gnd vdd FILL
XFILL_2__14417_ gnd vdd FILL
XFILL_5__12789_ gnd vdd FILL
XFILL_3__8064_ gnd vdd FILL
X_8983_ _9057_/Q gnd _8983_/Y vdd INVX1
XFILL_2__11629_ gnd vdd FILL
XFILL_3__13968_ gnd vdd FILL
XFILL_2__15397_ gnd vdd FILL
XFILL_0__7306_ gnd vdd FILL
XFILL_0__13788_ gnd vdd FILL
XFILL_5__14528_ gnd vdd FILL
XFILL_3__15707_ gnd vdd FILL
XFILL_4__13169_ gnd vdd FILL
XFILL_1__12009_ gnd vdd FILL
X_7934_ _7934_/A _7931_/B _7933_/Y gnd _8024_/D vdd OAI21X1
XFILL_2__14348_ gnd vdd FILL
XFILL_0__12739_ gnd vdd FILL
XFILL_0__15527_ gnd vdd FILL
XFILL_3__13899_ gnd vdd FILL
XFILL_6__15818_ gnd vdd FILL
XSFILL13640x15050 gnd vdd FILL
XFILL_0__7237_ gnd vdd FILL
XFILL_5__14459_ gnd vdd FILL
XFILL_3__15638_ gnd vdd FILL
X_7865_ _7821_/B _9017_/B gnd _7865_/Y vdd NAND2X1
XFILL_2__14279_ gnd vdd FILL
XFILL_0__15458_ gnd vdd FILL
XFILL_0__7168_ gnd vdd FILL
X_9604_ _9602_/Y _9613_/B _9603_/Y gnd _9690_/D vdd OAI21X1
XFILL_2__16018_ gnd vdd FILL
XFILL_3__15569_ gnd vdd FILL
X_7796_ _7796_/Q _8297_/CLK _7796_/R vdd _7796_/D gnd vdd DFFSR
XSFILL38840x81050 gnd vdd FILL
XSFILL38040x62050 gnd vdd FILL
XFILL_0__14409_ gnd vdd FILL
XFILL_3__8966_ gnd vdd FILL
XFILL_0__15389_ gnd vdd FILL
XFILL_5__16129_ gnd vdd FILL
XFILL_0__7099_ gnd vdd FILL
X_9535_ _9535_/A _8511_/B gnd _9536_/C vdd NAND2X1
XFILL_1__7981_ gnd vdd FILL
XFILL_5_BUFX2_insert102 gnd vdd FILL
XFILL_4__7690_ gnd vdd FILL
XFILL_3__8897_ gnd vdd FILL
XFILL_1__9720_ gnd vdd FILL
XFILL_1__6932_ gnd vdd FILL
X_9466_ _9466_/A _9466_/B gnd _9467_/C vdd NAND2X1
XFILL_3__7848_ gnd vdd FILL
XSFILL43960x72050 gnd vdd FILL
X_8417_ _8343_/A _7268_/CLK _8688_/R vdd _8417_/D gnd vdd DFFSR
XSFILL28760x6050 gnd vdd FILL
XFILL_1__9651_ gnd vdd FILL
X_9397_ _9451_/Q gnd _9399_/A vdd INVX1
XFILL_1__6863_ gnd vdd FILL
XFILL_4_BUFX2_insert802 gnd vdd FILL
XFILL_4__9360_ gnd vdd FILL
XFILL_4_BUFX2_insert813 gnd vdd FILL
XFILL_1__8602_ gnd vdd FILL
XFILL_4_BUFX2_insert824 gnd vdd FILL
XFILL_0__9809_ gnd vdd FILL
XFILL_4_BUFX2_insert835 gnd vdd FILL
X_8348_ _8346_/Y _8356_/A _8348_/C gnd _8418_/D vdd OAI21X1
XSFILL44040x81050 gnd vdd FILL
XFILL_4__8311_ gnd vdd FILL
XFILL_3__9518_ gnd vdd FILL
XFILL_4_BUFX2_insert846 gnd vdd FILL
XFILL_4_BUFX2_insert857 gnd vdd FILL
XFILL_4__9291_ gnd vdd FILL
XFILL111960x38050 gnd vdd FILL
XFILL_4_BUFX2_insert868 gnd vdd FILL
XFILL_1__8533_ gnd vdd FILL
XFILL_4_BUFX2_insert879 gnd vdd FILL
X_8279_ _8185_/A _9447_/CLK _9447_/R vdd _8279_/D gnd vdd DFFSR
XFILL_4__8242_ gnd vdd FILL
XFILL_1__8464_ gnd vdd FILL
XFILL_1__7415_ gnd vdd FILL
XSFILL38920x61050 gnd vdd FILL
XSFILL38120x42050 gnd vdd FILL
XFILL_1__8395_ gnd vdd FILL
XFILL_4__7124_ gnd vdd FILL
X_12920_ _12119_/B _8180_/CLK _7391_/R vdd _12920_/D gnd vdd DFFSR
XFILL_1__7346_ gnd vdd FILL
XFILL_4__7055_ gnd vdd FILL
XSFILL39000x70050 gnd vdd FILL
X_12851_ vdd _12851_/B gnd _12851_/Y vdd NAND2X1
XFILL_5_BUFX2_insert2 gnd vdd FILL
XFILL_1_BUFX2_insert703 gnd vdd FILL
X_11802_ _11802_/A _11786_/Y _11802_/C gnd _11808_/C vdd NAND3X1
XFILL_1_BUFX2_insert714 gnd vdd FILL
XFILL_1__9016_ gnd vdd FILL
X_15570_ _15569_/Y _15565_/Y _15570_/C gnd _15571_/A vdd NOR3X1
X_12782_ _12782_/A gnd _12782_/Y vdd INVX1
XFILL_1_BUFX2_insert725 gnd vdd FILL
XFILL_1_BUFX2_insert736 gnd vdd FILL
XFILL_1_BUFX2_insert747 gnd vdd FILL
X_14521_ _14520_/Y _13978_/B gnd _14522_/C vdd NOR2X1
XFILL_1_BUFX2_insert758 gnd vdd FILL
X_11733_ _11268_/Y _11366_/B _11733_/C gnd _11733_/Y vdd OAI21X1
XFILL_1_BUFX2_insert769 gnd vdd FILL
XFILL_4__7957_ gnd vdd FILL
X_14452_ _8555_/Q gnd _14452_/Y vdd INVX1
XSFILL89800x5050 gnd vdd FILL
X_11664_ _11649_/Y _11664_/B gnd _11664_/Y vdd NOR2X1
XSFILL105160x79050 gnd vdd FILL
XFILL_2__9760_ gnd vdd FILL
XFILL_2__6972_ gnd vdd FILL
XFILL_4_BUFX2_insert18 gnd vdd FILL
XFILL_4__6908_ gnd vdd FILL
XFILL_4_BUFX2_insert29 gnd vdd FILL
X_13403_ _9718_/A gnd _13403_/Y vdd INVX1
XFILL112120x27050 gnd vdd FILL
XFILL_5__10140_ gnd vdd FILL
X_10615_ _8183_/A _10615_/B gnd _10615_/Y vdd NAND2X1
XFILL_4__7888_ gnd vdd FILL
XFILL_1__9918_ gnd vdd FILL
X_14383_ _14383_/A _13978_/B _14545_/B _15841_/D gnd _14387_/B vdd OAI22X1
XFILL_2__8711_ gnd vdd FILL
XFILL_4__10870_ gnd vdd FILL
X_11595_ _11121_/Y _11129_/Y _11595_/C gnd _11599_/C vdd NAND3X1
XSFILL23400x62050 gnd vdd FILL
XFILL_4__9627_ gnd vdd FILL
XSFILL64040x12050 gnd vdd FILL
X_16122_ _16122_/A _16122_/B _16112_/Y gnd _16123_/B vdd NAND3X1
XFILL_4__6839_ gnd vdd FILL
XFILL_1__10690_ gnd vdd FILL
X_13334_ _13259_/C _13270_/A gnd _13334_/Y vdd NOR2X1
X_10546_ _15878_/A gnd _10548_/A vdd INVX1
XFILL_5_BUFX2_insert680 gnd vdd FILL
XFILL_1__9849_ gnd vdd FILL
XFILL_2__8642_ gnd vdd FILL
XFILL_3__11250_ gnd vdd FILL
XFILL_2__11980_ gnd vdd FILL
XFILL_5__8351_ gnd vdd FILL
XFILL_0__11070_ gnd vdd FILL
XFILL_5_BUFX2_insert691 gnd vdd FILL
X_16053_ _16048_/Y _16053_/B _16052_/Y gnd _16059_/C vdd NOR3X1
X_13265_ _13297_/C _13265_/B gnd _13265_/Y vdd NOR2X1
X_10477_ _10427_/A _8038_/CLK _7789_/R vdd _10477_/D gnd vdd DFFSR
XFILL_3__11181_ gnd vdd FILL
XFILL_2__10931_ gnd vdd FILL
XFILL_0__10021_ gnd vdd FILL
XFILL_4__8509_ gnd vdd FILL
XFILL_1__12360_ gnd vdd FILL
XFILL_2__8573_ gnd vdd FILL
XFILL_5__7302_ gnd vdd FILL
XFILL_6__13100_ gnd vdd FILL
X_15004_ _16306_/C gnd _15695_/D vdd INVX2
X_12216_ _12216_/A _12216_/B gnd _12216_/Y vdd AND2X2
XFILL_4__9489_ gnd vdd FILL
XFILL_5__13830_ gnd vdd FILL
XFILL_6__11292_ gnd vdd FILL
X_13196_ _13196_/Q _13175_/CLK _13199_/R vdd _13196_/D gnd vdd DFFSR
XFILL_4__12471_ gnd vdd FILL
XFILL_3__10132_ gnd vdd FILL
XFILL_1__11311_ gnd vdd FILL
XSFILL3720x81050 gnd vdd FILL
XSFILL14360x78050 gnd vdd FILL
XFILL_2__13650_ gnd vdd FILL
XFILL_1__12291_ gnd vdd FILL
XFILL_5__7233_ gnd vdd FILL
XFILL_4__14210_ gnd vdd FILL
XFILL_6__10243_ gnd vdd FILL
XSFILL29160x38050 gnd vdd FILL
XSFILL84200x25050 gnd vdd FILL
X_12147_ _12147_/A _12122_/A _12146_/Y gnd _12147_/Y vdd OAI21X1
XFILL_4__11422_ gnd vdd FILL
XFILL_2__12601_ gnd vdd FILL
XFILL_5__10973_ gnd vdd FILL
XFILL_3__10063_ gnd vdd FILL
XFILL_4__15190_ gnd vdd FILL
XFILL_5__13761_ gnd vdd FILL
XFILL_1__14030_ gnd vdd FILL
XFILL_3__14940_ gnd vdd FILL
XFILL_2__7455_ gnd vdd FILL
XFILL_1__11242_ gnd vdd FILL
XFILL_2__10793_ gnd vdd FILL
XFILL_2__13581_ gnd vdd FILL
XFILL_0__14760_ gnd vdd FILL
XFILL_0__11972_ gnd vdd FILL
XFILL_5__15500_ gnd vdd FILL
XFILL_5__7164_ gnd vdd FILL
XFILL_5__12712_ gnd vdd FILL
XFILL_4__14141_ gnd vdd FILL
XFILL_2__15320_ gnd vdd FILL
X_12078_ _12078_/A _12078_/B _12077_/Y gnd _13146_/B vdd NAND3X1
XFILL_5__13692_ gnd vdd FILL
XFILL_4__11353_ gnd vdd FILL
XFILL_3__14871_ gnd vdd FILL
XFILL_2__12532_ gnd vdd FILL
XFILL_0__13711_ gnd vdd FILL
XFILL_0__10923_ gnd vdd FILL
XFILL_1__11173_ gnd vdd FILL
XFILL_0__14691_ gnd vdd FILL
XFILL_4__10304_ gnd vdd FILL
XFILL_5__7095_ gnd vdd FILL
X_15906_ _8939_/Q gnd _15906_/Y vdd INVX1
XFILL_5__15431_ gnd vdd FILL
X_11029_ _12238_/Y _11030_/A gnd _11034_/B vdd XNOR2X1
XFILL_3__13822_ gnd vdd FILL
XFILL_2__9125_ gnd vdd FILL
XFILL_5__12643_ gnd vdd FILL
XFILL_4__14072_ gnd vdd FILL
XFILL_1__10124_ gnd vdd FILL
XFILL_2__15251_ gnd vdd FILL
XFILL_4__11284_ gnd vdd FILL
XFILL_0__13642_ gnd vdd FILL
XFILL_2__12463_ gnd vdd FILL
XFILL_1__15981_ gnd vdd FILL
XFILL_0_BUFX2_insert1005 gnd vdd FILL
XSFILL99480x79050 gnd vdd FILL
XFILL_0_BUFX2_insert1016 gnd vdd FILL
XFILL_4__13023_ gnd vdd FILL
XFILL_0__8140_ gnd vdd FILL
X_15837_ _15837_/A gnd _15837_/Y vdd INVX1
XFILL_2__14202_ gnd vdd FILL
XFILL_5__12574_ gnd vdd FILL
XFILL_5__15362_ gnd vdd FILL
XFILL_4__10235_ gnd vdd FILL
XFILL_2_BUFX2_insert570 gnd vdd FILL
XFILL_3__13753_ gnd vdd FILL
XFILL_0_BUFX2_insert1027 gnd vdd FILL
XFILL_2__11414_ gnd vdd FILL
XFILL_0_BUFX2_insert1038 gnd vdd FILL
XFILL_3__10965_ gnd vdd FILL
XFILL_2__15182_ gnd vdd FILL
XFILL_2__12394_ gnd vdd FILL
XFILL_1__14932_ gnd vdd FILL
XFILL_0__16361_ gnd vdd FILL
XFILL_1__10055_ gnd vdd FILL
XFILL_2_BUFX2_insert581 gnd vdd FILL
XFILL_0_BUFX2_insert1049 gnd vdd FILL
XFILL_0__13573_ gnd vdd FILL
XFILL_2_BUFX2_insert592 gnd vdd FILL
XFILL_0__10785_ gnd vdd FILL
XFILL_5__14313_ gnd vdd FILL
XFILL_5__11525_ gnd vdd FILL
XFILL_0__8071_ gnd vdd FILL
XFILL_3__12704_ gnd vdd FILL
X_15768_ _15762_/Y _15767_/Y gnd _15769_/A vdd NAND2X1
XFILL_2__8007_ gnd vdd FILL
XFILL_4__10166_ gnd vdd FILL
XFILL_2__14133_ gnd vdd FILL
XFILL_5__15293_ gnd vdd FILL
XFILL_0__15312_ gnd vdd FILL
XFILL_3__13684_ gnd vdd FILL
XFILL_0__12524_ gnd vdd FILL
XFILL_2__11345_ gnd vdd FILL
XFILL_5__9805_ gnd vdd FILL
XFILL_1__14863_ gnd vdd FILL
XFILL_3__10896_ gnd vdd FILL
XFILL_0__16292_ gnd vdd FILL
XFILL_6__15603_ gnd vdd FILL
X_14719_ _9028_/A gnd _14719_/Y vdd INVX1
XSFILL53960x35050 gnd vdd FILL
XFILL_5__7997_ gnd vdd FILL
XFILL_5__14244_ gnd vdd FILL
X_7650_ _7578_/A _7778_/CLK _8418_/R vdd _7650_/D gnd vdd DFFSR
XFILL_5__11456_ gnd vdd FILL
XFILL_3__15423_ gnd vdd FILL
XFILL_3__12635_ gnd vdd FILL
X_15699_ _15698_/Y _16228_/B gnd _15699_/Y vdd NOR2X1
XFILL_1__13814_ gnd vdd FILL
XSFILL109480x64050 gnd vdd FILL
XFILL_0__15243_ gnd vdd FILL
XFILL_2__14064_ gnd vdd FILL
XFILL_4__14974_ gnd vdd FILL
XFILL_2__11276_ gnd vdd FILL
XFILL_0__12455_ gnd vdd FILL
XFILL_5__10407_ gnd vdd FILL
XFILL_5__6948_ gnd vdd FILL
XFILL_5__9736_ gnd vdd FILL
XFILL_1__14794_ gnd vdd FILL
XSFILL38760x1050 gnd vdd FILL
XFILL_5__14175_ gnd vdd FILL
XSFILL28760x11050 gnd vdd FILL
XFILL_3__15354_ gnd vdd FILL
XFILL_2__13015_ gnd vdd FILL
X_7581_ _7581_/A gnd _7583_/A vdd INVX1
XFILL_5__11387_ gnd vdd FILL
XFILL_4__13925_ gnd vdd FILL
XSFILL54040x44050 gnd vdd FILL
XFILL_0__11406_ gnd vdd FILL
XFILL_3__8751_ gnd vdd FILL
XFILL_0__15174_ gnd vdd FILL
XFILL_1__13745_ gnd vdd FILL
XFILL_1__10957_ gnd vdd FILL
XFILL_5__13126_ gnd vdd FILL
XFILL_0__12386_ gnd vdd FILL
X_9320_ _9320_/Q _7912_/CLK _7911_/R vdd _9262_/Y gnd vdd DFFSR
XFILL_5__9667_ gnd vdd FILL
XFILL_3__14305_ gnd vdd FILL
XFILL_5__6879_ gnd vdd FILL
XFILL_6__15465_ gnd vdd FILL
XFILL_2__8909_ gnd vdd FILL
XFILL_0__8973_ gnd vdd FILL
XFILL_3__7702_ gnd vdd FILL
XFILL_3__11517_ gnd vdd FILL
XFILL_4__13856_ gnd vdd FILL
XFILL_0__14125_ gnd vdd FILL
XFILL_2__10158_ gnd vdd FILL
XFILL_3__15285_ gnd vdd FILL
XFILL_2__9889_ gnd vdd FILL
XFILL_3__12497_ gnd vdd FILL
XFILL_5__8618_ gnd vdd FILL
XFILL_0__11337_ gnd vdd FILL
XBUFX2_insert580 BUFX2_insert524/A gnd _9447_/R vdd BUFX2
XFILL_1__13676_ gnd vdd FILL
XBUFX2_insert591 BUFX2_insert607/A gnd _8278_/R vdd BUFX2
XFILL_1__10888_ gnd vdd FILL
XFILL_6__14416_ gnd vdd FILL
X_9251_ _9317_/Q gnd _9251_/Y vdd INVX1
XFILL_5__9598_ gnd vdd FILL
XFILL_6__8391_ gnd vdd FILL
XFILL_3__14236_ gnd vdd FILL
XFILL_5__10269_ gnd vdd FILL
XSFILL104040x13050 gnd vdd FILL
XFILL_4__13787_ gnd vdd FILL
XFILL_3__11448_ gnd vdd FILL
XFILL_1__15415_ gnd vdd FILL
XFILL_3__7633_ gnd vdd FILL
XFILL_1__12627_ gnd vdd FILL
XFILL_0__14056_ gnd vdd FILL
XFILL_4_BUFX2_insert109 gnd vdd FILL
XFILL_2__14966_ gnd vdd FILL
XFILL_4__10999_ gnd vdd FILL
XFILL_1__16395_ gnd vdd FILL
X_8202_ _8202_/A _8232_/B _8202_/C gnd _8202_/Y vdd OAI21X1
XFILL_5__12008_ gnd vdd FILL
XFILL_0__11268_ gnd vdd FILL
XFILL_4__12738_ gnd vdd FILL
X_9182_ _9102_/A _8537_/CLK _9054_/R vdd _9182_/D gnd vdd DFFSR
XFILL_4__15526_ gnd vdd FILL
XFILL_0__7855_ gnd vdd FILL
XFILL_3__14167_ gnd vdd FILL
XFILL_0__13007_ gnd vdd FILL
XFILL_2__13917_ gnd vdd FILL
XSFILL48920x24050 gnd vdd FILL
XFILL_3__7564_ gnd vdd FILL
XFILL_1__15346_ gnd vdd FILL
XFILL_3__11379_ gnd vdd FILL
XSFILL74200x57050 gnd vdd FILL
XFILL_2__14897_ gnd vdd FILL
X_8133_ _8133_/A _9797_/B gnd _8134_/C vdd NAND2X1
XFILL_0__11199_ gnd vdd FILL
XFILL_3__13118_ gnd vdd FILL
XFILL_6__14278_ gnd vdd FILL
XFILL_4__15457_ gnd vdd FILL
XFILL_2__13848_ gnd vdd FILL
XFILL_3_BUFX2_insert809 gnd vdd FILL
XFILL_1__11509_ gnd vdd FILL
XFILL_3__14098_ gnd vdd FILL
XFILL_6__9012_ gnd vdd FILL
XFILL_6__16017_ gnd vdd FILL
XSFILL99160x61050 gnd vdd FILL
XFILL_1__12489_ gnd vdd FILL
XFILL_3__7495_ gnd vdd FILL
XFILL_1__15277_ gnd vdd FILL
XFILL_0__9525_ gnd vdd FILL
XFILL_6__13229_ gnd vdd FILL
XSFILL49000x33050 gnd vdd FILL
X_8064_ _8079_/A _7424_/B gnd _8064_/Y vdd NAND2X1
XFILL_4__14408_ gnd vdd FILL
XFILL_4__15388_ gnd vdd FILL
XFILL_3__9234_ gnd vdd FILL
XFILL_5__13959_ gnd vdd FILL
XFILL_1__14228_ gnd vdd FILL
XFILL_2__13779_ gnd vdd FILL
XFILL_0__14958_ gnd vdd FILL
X_7015_ _7015_/Q _8551_/CLK _7015_/R vdd _7015_/D gnd vdd DFFSR
XFILL_4__14339_ gnd vdd FILL
XFILL_2__15518_ gnd vdd FILL
XFILL_3__9165_ gnd vdd FILL
XFILL_1__14159_ gnd vdd FILL
XFILL_0__13909_ gnd vdd FILL
XFILL_1__7200_ gnd vdd FILL
XFILL112360x83050 gnd vdd FILL
XFILL_5__15629_ gnd vdd FILL
XFILL_0__14889_ gnd vdd FILL
XFILL_3__8116_ gnd vdd FILL
XFILL_0__9387_ gnd vdd FILL
XFILL_2__15449_ gnd vdd FILL
XFILL_3__9096_ gnd vdd FILL
XFILL_4__16009_ gnd vdd FILL
XFILL_0__8338_ gnd vdd FILL
X_8966_ _9005_/A _9094_/B gnd _8967_/C vdd NAND2X1
XSFILL43960x67050 gnd vdd FILL
XFILL_1__7062_ gnd vdd FILL
X_7917_ _7917_/Q _8947_/CLK _9069_/R vdd _7917_/D gnd vdd DFFSR
XFILL_0__8269_ gnd vdd FILL
XFILL_4__8860_ gnd vdd FILL
X_8897_ _8943_/Q gnd _8899_/A vdd INVX1
XSFILL18760x43050 gnd vdd FILL
XSFILL8600x53050 gnd vdd FILL
X_7848_ _7848_/A _7872_/B _7847_/Y gnd _7848_/Y vdd OAI21X1
XFILL_4__7811_ gnd vdd FILL
XFILL_0_CLKBUF1_insert114 gnd vdd FILL
XFILL_3__9998_ gnd vdd FILL
XFILL_0_CLKBUF1_insert125 gnd vdd FILL
XFILL_0_CLKBUF1_insert136 gnd vdd FILL
XFILL_0_CLKBUF1_insert147 gnd vdd FILL
XFILL_0_CLKBUF1_insert158 gnd vdd FILL
XFILL_4__7742_ gnd vdd FILL
XFILL_0_CLKBUF1_insert169 gnd vdd FILL
XSFILL18680x50 gnd vdd FILL
X_7779_ _7709_/A _7530_/CLK _7665_/R vdd _7711_/Y gnd vdd DFFSR
X_9518_ _9516_/Y _9535_/A _9518_/C gnd _9576_/D vdd OAI21X1
XFILL_1__7964_ gnd vdd FILL
X_10400_ _14146_/B gnd _10402_/A vdd INVX1
XSFILL110120x12050 gnd vdd FILL
XFILL_4__7673_ gnd vdd FILL
X_11380_ _11021_/Y gnd _11380_/Y vdd INVX1
XFILL_6__8589_ gnd vdd FILL
XFILL_1__6915_ gnd vdd FILL
XSFILL38920x56050 gnd vdd FILL
XFILL_4__9412_ gnd vdd FILL
X_9449_ _9449_/Q _7786_/CLK _9964_/R vdd _9449_/D gnd vdd DFFSR
XFILL112440x63050 gnd vdd FILL
XFILL_4_BUFX2_insert610 gnd vdd FILL
X_10331_ _13700_/A _7640_/CLK _7896_/R vdd _10247_/Y gnd vdd DFFSR
XFILL_1__9634_ gnd vdd FILL
XFILL_4_BUFX2_insert621 gnd vdd FILL
XFILL_4_BUFX2_insert632 gnd vdd FILL
XFILL_1__6846_ gnd vdd FILL
XFILL_4__9343_ gnd vdd FILL
XSFILL114520x9050 gnd vdd FILL
XFILL_4_BUFX2_insert643 gnd vdd FILL
X_13050_ _6873_/A _7005_/CLK _7133_/R vdd _12962_/Y gnd vdd DFFSR
XSFILL39000x65050 gnd vdd FILL
XFILL_4_BUFX2_insert654 gnd vdd FILL
X_10262_ _10262_/A _10271_/B _10261_/Y gnd _10336_/D vdd OAI21X1
XFILL_4_BUFX2_insert665 gnd vdd FILL
XFILL_4_BUFX2_insert676 gnd vdd FILL
XSFILL114200x58050 gnd vdd FILL
X_12001_ _12449_/B _12105_/B _12001_/C gnd gnd _12001_/Y vdd AOI22X1
XFILL_4_BUFX2_insert687 gnd vdd FILL
XFILL_4__9274_ gnd vdd FILL
XFILL_4_BUFX2_insert698 gnd vdd FILL
XFILL_1__8516_ gnd vdd FILL
X_10193_ _10193_/A _8273_/B gnd _10194_/C vdd NAND2X1
XFILL_1__9496_ gnd vdd FILL
XFILL_4__8225_ gnd vdd FILL
XSFILL44120x56050 gnd vdd FILL
XFILL_1__8447_ gnd vdd FILL
XFILL_2__7240_ gnd vdd FILL
XSFILL59720x35050 gnd vdd FILL
XSFILL84520x61050 gnd vdd FILL
XSFILL69080x60050 gnd vdd FILL
X_13952_ _13952_/A _13952_/B _13952_/C gnd _13953_/B vdd NAND3X1
XSFILL99320x21050 gnd vdd FILL
XFILL_1__8378_ gnd vdd FILL
XFILL_2__7171_ gnd vdd FILL
XFILL_4__7107_ gnd vdd FILL
XFILL_4__8087_ gnd vdd FILL
X_12903_ _12901_/Y vdd _12903_/C gnd _12945_/D vdd OAI21X1
X_13883_ _9438_/Q _13883_/B _13883_/C gnd _13883_/Y vdd AOI21X1
XFILL_1__7329_ gnd vdd FILL
XFILL_4__7038_ gnd vdd FILL
X_15622_ _15622_/A _15621_/Y _15239_/B _14157_/C gnd _15622_/Y vdd OAI22X1
XFILL_6__10930_ gnd vdd FILL
XFILL_4__10020_ gnd vdd FILL
X_12834_ _12832_/Y vdd _12834_/C gnd _12922_/D vdd OAI21X1
XFILL_1_BUFX2_insert500 gnd vdd FILL
XSFILL38200x17050 gnd vdd FILL
XFILL_1_BUFX2_insert511 gnd vdd FILL
XFILL_1_BUFX2_insert522 gnd vdd FILL
XFILL_3__10750_ gnd vdd FILL
XSFILL84840x50 gnd vdd FILL
XFILL_0__10570_ gnd vdd FILL
XFILL_1_BUFX2_insert533 gnd vdd FILL
XFILL_5__7851_ gnd vdd FILL
XFILL_5__11310_ gnd vdd FILL
XFILL_1_BUFX2_insert544 gnd vdd FILL
X_15553_ _6938_/A gnd _15553_/Y vdd INVX1
X_12765_ _12777_/A memoryOutData[23] gnd _12766_/C vdd NAND2X1
XFILL_5__12290_ gnd vdd FILL
XFILL_1_BUFX2_insert555 gnd vdd FILL
XFILL_2__11130_ gnd vdd FILL
XSFILL89240x73050 gnd vdd FILL
XFILL_1_BUFX2_insert566 gnd vdd FILL
XFILL_3__10681_ gnd vdd FILL
XFILL_1__11860_ gnd vdd FILL
XFILL_1_BUFX2_insert577 gnd vdd FILL
X_14504_ _14504_/A gnd _15948_/B vdd INVX1
XSFILL3480x14050 gnd vdd FILL
XFILL_1_BUFX2_insert588 gnd vdd FILL
X_11716_ _11716_/A _11716_/B _11710_/Y gnd _11716_/Y vdd OAI21X1
XFILL_4__8989_ gnd vdd FILL
XFILL_5__11241_ gnd vdd FILL
XFILL_3__12420_ gnd vdd FILL
XFILL_2__9812_ gnd vdd FILL
XFILL_1_BUFX2_insert599 gnd vdd FILL
X_15484_ _7188_/A gnd _15484_/Y vdd INVX1
X_12696_ memoryOutData[0] _10944_/C gnd _12697_/C vdd NAND2X1
XFILL_4__11971_ gnd vdd FILL
XFILL_2__11061_ gnd vdd FILL
XSFILL3720x76050 gnd vdd FILL
XFILL_1__10811_ gnd vdd FILL
XFILL_0__12240_ gnd vdd FILL
XFILL_5__9521_ gnd vdd FILL
XSFILL100040x5050 gnd vdd FILL
XFILL_1__11791_ gnd vdd FILL
X_14435_ _7090_/A gnd _14436_/B vdd INVX1
XSFILL54760x78050 gnd vdd FILL
XFILL_4__10922_ gnd vdd FILL
XFILL_2__10012_ gnd vdd FILL
X_11647_ _11748_/A _11658_/A _11621_/C gnd _11647_/Y vdd OAI21X1
XFILL_4__13710_ gnd vdd FILL
XFILL_5__11172_ gnd vdd FILL
XFILL_2__9743_ gnd vdd FILL
XFILL_3__12351_ gnd vdd FILL
XFILL_4__14690_ gnd vdd FILL
XFILL_1__10742_ gnd vdd FILL
XFILL_1__13530_ gnd vdd FILL
XFILL_2__6955_ gnd vdd FILL
XSFILL94360x64050 gnd vdd FILL
XFILL_0__12171_ gnd vdd FILL
XFILL_5__10123_ gnd vdd FILL
XFILL_6__15250_ gnd vdd FILL
XFILL_4__13641_ gnd vdd FILL
X_14366_ _14366_/A _14366_/B gnd _14366_/Y vdd NOR2X1
XFILL_3__11302_ gnd vdd FILL
XFILL_5__15980_ gnd vdd FILL
XFILL_2__14820_ gnd vdd FILL
XFILL_3__15070_ gnd vdd FILL
X_11578_ _11576_/Y _11578_/B _11575_/Y gnd _11578_/Y vdd OAI21X1
XFILL_2__9674_ gnd vdd FILL
XFILL_3__12282_ gnd vdd FILL
XFILL_5__8403_ gnd vdd FILL
XFILL_0__11122_ gnd vdd FILL
XFILL_6__14201_ gnd vdd FILL
XFILL_1__13461_ gnd vdd FILL
X_16105_ _16105_/A _15175_/B _16104_/Y gnd _16111_/C vdd AOI21X1
XSFILL69160x40050 gnd vdd FILL
XFILL_2__6886_ gnd vdd FILL
XFILL_1__10673_ gnd vdd FILL
X_13317_ _13289_/B _13303_/B _13316_/Y gnd _13317_/Y vdd OAI21X1
XFILL_5__9383_ gnd vdd FILL
X_10529_ _10557_/B _9633_/B gnd _10529_/Y vdd NAND2X1
XFILL_3__14021_ gnd vdd FILL
XFILL_5__10054_ gnd vdd FILL
XFILL_5__14931_ gnd vdd FILL
XFILL_1__15200_ gnd vdd FILL
XFILL_2__8625_ gnd vdd FILL
XFILL_4__16360_ gnd vdd FILL
XFILL_4__13572_ gnd vdd FILL
XFILL_3__11233_ gnd vdd FILL
X_14297_ _14293_/Y _14296_/Y gnd _14297_/Y vdd NOR2X1
XFILL_1__12412_ gnd vdd FILL
XFILL_4__10784_ gnd vdd FILL
XFILL_2__14751_ gnd vdd FILL
XFILL_5__8334_ gnd vdd FILL
XFILL_1__13392_ gnd vdd FILL
XFILL_1__16180_ gnd vdd FILL
XFILL_0__15930_ gnd vdd FILL
XFILL_2__11963_ gnd vdd FILL
XFILL_0__11053_ gnd vdd FILL
X_16036_ _16036_/A _16036_/B _16036_/C gnd _16036_/Y vdd OAI21X1
XSFILL48840x39050 gnd vdd FILL
X_13248_ _13248_/A gnd _13305_/B vdd INVX1
XFILL_4__15311_ gnd vdd FILL
XFILL_4__12523_ gnd vdd FILL
XFILL_6__11344_ gnd vdd FILL
XFILL_5__14862_ gnd vdd FILL
XFILL_4__16291_ gnd vdd FILL
XFILL_2__13702_ gnd vdd FILL
XFILL_2__10914_ gnd vdd FILL
XFILL_1__12343_ gnd vdd FILL
XFILL_3__11164_ gnd vdd FILL
XFILL_0__10004_ gnd vdd FILL
XFILL_1__15131_ gnd vdd FILL
XFILL_2__14682_ gnd vdd FILL
XFILL_2__11894_ gnd vdd FILL
XFILL_5__8265_ gnd vdd FILL
XFILL_0__15861_ gnd vdd FILL
XFILL_5__13813_ gnd vdd FILL
XFILL_4__15242_ gnd vdd FILL
XFILL_6__14063_ gnd vdd FILL
XFILL_3__10115_ gnd vdd FILL
X_13179_ _12127_/A _12537_/CLK _12536_/R vdd _13179_/D gnd vdd DFFSR
XFILL_2__7507_ gnd vdd FILL
XFILL_4__12454_ gnd vdd FILL
XSFILL89880x10050 gnd vdd FILL
XFILL_0__7571_ gnd vdd FILL
XFILL_2__13633_ gnd vdd FILL
XFILL_5__14793_ gnd vdd FILL
XFILL_3__15972_ gnd vdd FILL
XFILL_2__8487_ gnd vdd FILL
XFILL_0__14812_ gnd vdd FILL
XFILL_1__15062_ gnd vdd FILL
XFILL_5__7216_ gnd vdd FILL
XFILL_1__12274_ gnd vdd FILL
XFILL_3__11095_ gnd vdd FILL
XFILL_5__8196_ gnd vdd FILL
XFILL_0__15792_ gnd vdd FILL
XFILL_4__11405_ gnd vdd FILL
XFILL_5__13744_ gnd vdd FILL
XFILL_4__15173_ gnd vdd FILL
XFILL_5__10956_ gnd vdd FILL
XFILL_2__7438_ gnd vdd FILL
XFILL_3__10046_ gnd vdd FILL
XFILL_4__12385_ gnd vdd FILL
XFILL_1__14013_ gnd vdd FILL
XFILL_2__16352_ gnd vdd FILL
XFILL_1__11225_ gnd vdd FILL
XFILL_3__14923_ gnd vdd FILL
XSFILL109480x59050 gnd vdd FILL
XFILL_2__13564_ gnd vdd FILL
XFILL_0__11955_ gnd vdd FILL
XFILL_2__10776_ gnd vdd FILL
XFILL_0__14743_ gnd vdd FILL
XFILL_4__14124_ gnd vdd FILL
XFILL_0__9241_ gnd vdd FILL
XFILL_2__15303_ gnd vdd FILL
XFILL_0_BUFX2_insert16 gnd vdd FILL
XFILL_4__11336_ gnd vdd FILL
XFILL_5__13675_ gnd vdd FILL
XFILL_3__14854_ gnd vdd FILL
XFILL_2__12515_ gnd vdd FILL
XFILL_5__10887_ gnd vdd FILL
XFILL_0_BUFX2_insert27 gnd vdd FILL
XFILL_0__10906_ gnd vdd FILL
XFILL_2__7369_ gnd vdd FILL
XFILL_1__11156_ gnd vdd FILL
XFILL_2__16283_ gnd vdd FILL
XFILL_2__13495_ gnd vdd FILL
XFILL_0_BUFX2_insert38 gnd vdd FILL
XFILL_5__15414_ gnd vdd FILL
XFILL_0__11886_ gnd vdd FILL
XFILL_5__7078_ gnd vdd FILL
XFILL_0_BUFX2_insert49 gnd vdd FILL
XFILL_0__14674_ gnd vdd FILL
XFILL_3__13805_ gnd vdd FILL
XFILL_5__12626_ gnd vdd FILL
XSFILL94440x44050 gnd vdd FILL
XFILL_4__14055_ gnd vdd FILL
XFILL_2__9108_ gnd vdd FILL
X_8820_ _8820_/Q _7647_/CLK _9823_/R vdd _8820_/D gnd vdd DFFSR
XFILL_0__9172_ gnd vdd FILL
XFILL_2__15234_ gnd vdd FILL
XFILL_1__10107_ gnd vdd FILL
XFILL_4__11267_ gnd vdd FILL
XFILL_5__16394_ gnd vdd FILL
XFILL_2__12446_ gnd vdd FILL
XFILL_0__16413_ gnd vdd FILL
XFILL_3__14785_ gnd vdd FILL
XFILL_0__13625_ gnd vdd FILL
XFILL_3__11997_ gnd vdd FILL
XFILL_1__15964_ gnd vdd FILL
XFILL_1__11087_ gnd vdd FILL
XFILL_0__10837_ gnd vdd FILL
XFILL_0__8123_ gnd vdd FILL
XFILL_4__13006_ gnd vdd FILL
XFILL_5__15345_ gnd vdd FILL
XFILL_2__9039_ gnd vdd FILL
XFILL_3__9921_ gnd vdd FILL
XFILL_3__13736_ gnd vdd FILL
X_8751_ _8809_/Q gnd _8753_/A vdd INVX1
XFILL_3__10948_ gnd vdd FILL
XFILL_1__10038_ gnd vdd FILL
XFILL_2__15165_ gnd vdd FILL
XFILL_1__14915_ gnd vdd FILL
XFILL_4__11198_ gnd vdd FILL
XFILL_0__16344_ gnd vdd FILL
XFILL_2__12377_ gnd vdd FILL
XFILL_6_BUFX2_insert705 gnd vdd FILL
XFILL_0__13556_ gnd vdd FILL
XFILL_0__10768_ gnd vdd FILL
XFILL_1__15895_ gnd vdd FILL
XFILL_6__6842_ gnd vdd FILL
X_7702_ _7700_/Y _7753_/B _7702_/C gnd _7702_/Y vdd OAI21X1
XFILL_5__11508_ gnd vdd FILL
XFILL_0__8054_ gnd vdd FILL
XFILL_4__10149_ gnd vdd FILL
XFILL_5__12488_ gnd vdd FILL
XFILL_2__14116_ gnd vdd FILL
XFILL_5__15276_ gnd vdd FILL
XFILL_3__13667_ gnd vdd FILL
XFILL_0__12507_ gnd vdd FILL
XFILL_3__9852_ gnd vdd FILL
XFILL_2__11328_ gnd vdd FILL
X_8682_ _8626_/A _9716_/CLK _8682_/R vdd _8682_/D gnd vdd DFFSR
XFILL_1__14846_ gnd vdd FILL
XSFILL18680x58050 gnd vdd FILL
XFILL_3__10879_ gnd vdd FILL
XFILL_2__15096_ gnd vdd FILL
XFILL_0__13487_ gnd vdd FILL
XFILL_0__16275_ gnd vdd FILL
XFILL_3__15406_ gnd vdd FILL
XFILL_5__14227_ gnd vdd FILL
XFILL_0__10699_ gnd vdd FILL
XSFILL58280x44050 gnd vdd FILL
XFILL_5__11439_ gnd vdd FILL
XFILL_3__12618_ gnd vdd FILL
X_7633_ _7577_/B _8401_/B gnd _7634_/C vdd NAND2X1
XFILL_3__16386_ gnd vdd FILL
XFILL_2__14047_ gnd vdd FILL
XFILL_4__14957_ gnd vdd FILL
XFILL_3__9783_ gnd vdd FILL
XFILL_3__13598_ gnd vdd FILL
XFILL_0__15226_ gnd vdd FILL
XFILL_0__12438_ gnd vdd FILL
XFILL_2__11259_ gnd vdd FILL
XFILL_5__9719_ gnd vdd FILL
XFILL_3__6995_ gnd vdd FILL
XFILL_1__14777_ gnd vdd FILL
XFILL_1__11989_ gnd vdd FILL
X_7564_ _7606_/A _7564_/B gnd _7565_/C vdd NAND2X1
XFILL_3__15337_ gnd vdd FILL
XFILL_5__14158_ gnd vdd FILL
XFILL_4__13908_ gnd vdd FILL
XFILL_3__8734_ gnd vdd FILL
XFILL_0__15157_ gnd vdd FILL
XFILL_1__13728_ gnd vdd FILL
XFILL_4__14888_ gnd vdd FILL
XFILL_0__12369_ gnd vdd FILL
XFILL_5__13109_ gnd vdd FILL
X_9303_ _9303_/Q _9447_/CLK _9447_/R vdd _9211_/Y gnd vdd DFFSR
XFILL_1_CLKBUF1_insert209 gnd vdd FILL
XSFILL109560x39050 gnd vdd FILL
XFILL_0__8956_ gnd vdd FILL
XFILL_5__14089_ gnd vdd FILL
XFILL_4__13839_ gnd vdd FILL
X_7495_ _7495_/A gnd _7495_/Y vdd INVX1
XFILL_0__14108_ gnd vdd FILL
XFILL_3__15268_ gnd vdd FILL
XFILL_2__15998_ gnd vdd FILL
XFILL_1__13659_ gnd vdd FILL
XFILL_0__15088_ gnd vdd FILL
XFILL111880x71050 gnd vdd FILL
XFILL112360x78050 gnd vdd FILL
XFILL_3__14219_ gnd vdd FILL
X_9234_ _9282_/A _9362_/B gnd _9235_/C vdd NAND2X1
XFILL_1__7680_ gnd vdd FILL
XFILL_0__8887_ gnd vdd FILL
XFILL_3__7616_ gnd vdd FILL
XFILL_3__15199_ gnd vdd FILL
XFILL_0__14039_ gnd vdd FILL
XFILL_2__14949_ gnd vdd FILL
XFILL_1__16378_ gnd vdd FILL
XFILL_3__8596_ gnd vdd FILL
XSFILL64280x63050 gnd vdd FILL
XSFILL99080x8050 gnd vdd FILL
X_9165_ _9203_/Q gnd _9165_/Y vdd INVX1
XFILL_4__15509_ gnd vdd FILL
XFILL_0__7838_ gnd vdd FILL
XFILL_1__15329_ gnd vdd FILL
XFILL_3__7547_ gnd vdd FILL
XFILL_3_BUFX2_insert606 gnd vdd FILL
X_8116_ _8116_/A _8133_/A _8116_/C gnd _8116_/Y vdd OAI21X1
XFILL_3_BUFX2_insert617 gnd vdd FILL
XFILL_1__9350_ gnd vdd FILL
X_9096_ _9180_/Q gnd _9098_/A vdd INVX1
XFILL_3_BUFX2_insert628 gnd vdd FILL
XFILL_3__7478_ gnd vdd FILL
XFILL_3_BUFX2_insert639 gnd vdd FILL
XFILL_0__9508_ gnd vdd FILL
X_8047_ _8001_/A _8815_/CLK _8047_/R vdd _8003_/Y gnd vdd DFFSR
XFILL_3__9217_ gnd vdd FILL
XFILL_4__8010_ gnd vdd FILL
XSFILL18760x38050 gnd vdd FILL
XFILL_1__9281_ gnd vdd FILL
XSFILL73800x25050 gnd vdd FILL
XSFILL8600x48050 gnd vdd FILL
XFILL_1__8232_ gnd vdd FILL
XSFILL33800x41050 gnd vdd FILL
XFILL_3__9148_ gnd vdd FILL
XSFILL85080x42050 gnd vdd FILL
XSFILL59240x52050 gnd vdd FILL
XFILL_3__9079_ gnd vdd FILL
X_9998_ _9998_/A gnd _9998_/Y vdd INVX1
XSFILL22840x65050 gnd vdd FILL
XFILL_1__7114_ gnd vdd FILL
X_10880_ _10879_/Y _10878_/Y gnd _10881_/B vdd NOR2X1
XFILL111960x51050 gnd vdd FILL
XFILL_1__8094_ gnd vdd FILL
X_8949_ _8915_/A _9205_/CLK _8433_/R vdd _8949_/D gnd vdd DFFSR
XFILL_4__8912_ gnd vdd FILL
XFILL_4__9892_ gnd vdd FILL
XFILL112440x58050 gnd vdd FILL
XFILL_1__7045_ gnd vdd FILL
XFILL_4__8843_ gnd vdd FILL
XFILL112360x3050 gnd vdd FILL
X_12550_ _12388_/A _12669_/CLK _9050_/R vdd _12486_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert507 gnd vdd FILL
XFILL_0_BUFX2_insert518 gnd vdd FILL
XFILL_0_BUFX2_insert529 gnd vdd FILL
XFILL_4__8774_ gnd vdd FILL
X_11501_ _11494_/A _11186_/Y _11415_/C gnd _11502_/A vdd OAI21X1
X_12481_ _12385_/A gnd _12483_/A vdd INVX1
XSFILL114360x12050 gnd vdd FILL
XFILL_1__8996_ gnd vdd FILL
XFILL_4__7725_ gnd vdd FILL
X_14220_ _14218_/Y _14865_/B _14567_/D _14219_/Y gnd _14224_/B vdd OAI22X1
XSFILL18840x18050 gnd vdd FILL
X_11432_ _11289_/C gnd _11616_/B vdd INVX2
XSFILL94280x79050 gnd vdd FILL
XFILL_1__7947_ gnd vdd FILL
X_14151_ _7072_/A gnd _14151_/Y vdd INVX1
XSFILL99320x16050 gnd vdd FILL
X_11363_ _11227_/A _11218_/B gnd _11366_/B vdd NAND2X1
XFILL_1__7878_ gnd vdd FILL
X_13102_ _13100_/Y _13153_/B _13101_/Y gnd _13182_/D vdd OAI21X1
X_10314_ _10354_/Q gnd _10316_/A vdd INVX1
XFILL_4__7587_ gnd vdd FILL
XFILL_4_BUFX2_insert440 gnd vdd FILL
XFILL_4_BUFX2_insert451 gnd vdd FILL
X_14082_ _7325_/A gnd _14083_/A vdd INVX1
XFILL_1__9617_ gnd vdd FILL
X_11294_ _11553_/B _11117_/Y gnd _11294_/Y vdd NAND2X1
XFILL_4_BUFX2_insert462 gnd vdd FILL
XFILL_2__9390_ gnd vdd FILL
XCLKBUF1_insert208 CLKBUF1_insert192/A gnd _8942_/CLK vdd CLKBUF1
XFILL_4_BUFX2_insert473 gnd vdd FILL
XCLKBUF1_insert219 CLKBUF1_insert220/A gnd _7912_/CLK vdd CLKBUF1
XFILL_4_BUFX2_insert484 gnd vdd FILL
XSFILL23800x7050 gnd vdd FILL
X_13033_ vdd _13033_/B gnd _13034_/C vdd NAND2X1
X_10245_ _13700_/A gnd _10247_/A vdd INVX1
XFILL_4_BUFX2_insert495 gnd vdd FILL
XFILL_1__9548_ gnd vdd FILL
XFILL_2__8341_ gnd vdd FILL
XFILL_4__9257_ gnd vdd FILL
XSFILL23800x73050 gnd vdd FILL
X_10176_ _10174_/Y _10127_/A _10176_/C gnd _10222_/D vdd OAI21X1
XFILL_5__10810_ gnd vdd FILL
XFILL_5__11790_ gnd vdd FILL
XFILL_4__8208_ gnd vdd FILL
XFILL_2__10630_ gnd vdd FILL
XFILL_1__9479_ gnd vdd FILL
XFILL_2__8272_ gnd vdd FILL
XSFILL89240x68050 gnd vdd FILL
XFILL_6__10011_ gnd vdd FILL
XFILL_2__7223_ gnd vdd FILL
X_14984_ _12767_/A gnd _14984_/Y vdd INVX1
XFILL_3__11920_ gnd vdd FILL
XFILL_4__12170_ gnd vdd FILL
XFILL_1__11010_ gnd vdd FILL
XFILL_4__8139_ gnd vdd FILL
XFILL_0__11740_ gnd vdd FILL
XFILL_2__10561_ gnd vdd FILL
XFILL_3_CLKBUF1_insert120 gnd vdd FILL
XFILL_4__11121_ gnd vdd FILL
X_13935_ _9492_/A gnd _15464_/B vdd INVX1
XFILL_3_CLKBUF1_insert131 gnd vdd FILL
XFILL_5__13460_ gnd vdd FILL
XFILL_5__10672_ gnd vdd FILL
XFILL_2__12300_ gnd vdd FILL
XFILL_3_CLKBUF1_insert142 gnd vdd FILL
XFILL_3__11851_ gnd vdd FILL
XFILL_5_CLKBUF1_insert1080 gnd vdd FILL
XFILL_2__13280_ gnd vdd FILL
XFILL_3_CLKBUF1_insert153 gnd vdd FILL
XFILL_2__10492_ gnd vdd FILL
XFILL_0__11671_ gnd vdd FILL
XFILL_5__12411_ gnd vdd FILL
XFILL_3_CLKBUF1_insert164 gnd vdd FILL
XFILL_5__8952_ gnd vdd FILL
X_13866_ _8974_/A gnd _13866_/Y vdd INVX1
XFILL_5__13391_ gnd vdd FILL
XFILL_4__11052_ gnd vdd FILL
XFILL_3_CLKBUF1_insert175 gnd vdd FILL
XFILL_3__10802_ gnd vdd FILL
XFILL_3__14570_ gnd vdd FILL
XFILL_3_CLKBUF1_insert186 gnd vdd FILL
XFILL_0__13410_ gnd vdd FILL
XSFILL84600x36050 gnd vdd FILL
XFILL_2__12231_ gnd vdd FILL
XFILL_2__7085_ gnd vdd FILL
XFILL_0__10622_ gnd vdd FILL
XFILL_3__11782_ gnd vdd FILL
XFILL_3_CLKBUF1_insert197 gnd vdd FILL
XFILL_1__12961_ gnd vdd FILL
XFILL_0__14390_ gnd vdd FILL
X_15605_ _9117_/A gnd _15606_/B vdd INVX1
X_12817_ _12773_/A _12692_/CLK _12692_/R vdd _12817_/D gnd vdd DFFSR
XSFILL69160x35050 gnd vdd FILL
XFILL_1_BUFX2_insert330 gnd vdd FILL
XFILL_5__12342_ gnd vdd FILL
XFILL_5__8883_ gnd vdd FILL
XFILL_4__10003_ gnd vdd FILL
XFILL_5__15130_ gnd vdd FILL
XFILL_1_BUFX2_insert341 gnd vdd FILL
XFILL_3__13521_ gnd vdd FILL
X_13797_ _8203_/A gnd _13798_/A vdd INVX1
XFILL_1__14700_ gnd vdd FILL
XFILL_4__15860_ gnd vdd FILL
XFILL_0__13341_ gnd vdd FILL
XFILL_1__11912_ gnd vdd FILL
XFILL_2__12162_ gnd vdd FILL
XFILL_1_BUFX2_insert352 gnd vdd FILL
XFILL_1__15680_ gnd vdd FILL
XFILL_0__10553_ gnd vdd FILL
XFILL_5__7834_ gnd vdd FILL
XFILL_1_BUFX2_insert363 gnd vdd FILL
XFILL_1__12892_ gnd vdd FILL
X_15536_ _15536_/A _15535_/Y _15651_/C gnd _12857_/B vdd AOI21X1
XFILL_1_BUFX2_insert374 gnd vdd FILL
X_12748_ _12748_/A _12762_/A _12748_/C gnd _12808_/D vdd OAI21X1
XFILL_1_BUFX2_insert385 gnd vdd FILL
XFILL_3__16240_ gnd vdd FILL
XFILL_4__14811_ gnd vdd FILL
XFILL_5__15061_ gnd vdd FILL
XFILL_5__12273_ gnd vdd FILL
XFILL_1_BUFX2_insert396 gnd vdd FILL
XFILL_3__13452_ gnd vdd FILL
XSFILL104360x44050 gnd vdd FILL
XFILL_2__11113_ gnd vdd FILL
XFILL_1__14631_ gnd vdd FILL
XFILL_3__10664_ gnd vdd FILL
XFILL_2__12093_ gnd vdd FILL
XFILL_4__15791_ gnd vdd FILL
XFILL_0__16060_ gnd vdd FILL
XFILL_0__13272_ gnd vdd FILL
XFILL_1__11843_ gnd vdd FILL
XFILL_5__14012_ gnd vdd FILL
XFILL_5__7765_ gnd vdd FILL
XFILL_5__11224_ gnd vdd FILL
XFILL_3__12403_ gnd vdd FILL
X_15467_ _7008_/Q _15382_/B _16096_/C _7316_/A gnd _15472_/A vdd AOI22X1
XSFILL74280x26050 gnd vdd FILL
X_12679_ _12615_/A _12809_/CLK _12685_/R vdd _12679_/D gnd vdd DFFSR
XFILL_2__15921_ gnd vdd FILL
XFILL_3__16171_ gnd vdd FILL
XFILL_4__11954_ gnd vdd FILL
XFILL_0__15011_ gnd vdd FILL
XFILL_4__14742_ gnd vdd FILL
XFILL_2__11044_ gnd vdd FILL
XFILL_3__13383_ gnd vdd FILL
XFILL_0__12223_ gnd vdd FILL
XFILL_1__14562_ gnd vdd FILL
XFILL_5__9504_ gnd vdd FILL
XFILL_2__7987_ gnd vdd FILL
XFILL_1__11774_ gnd vdd FILL
X_14418_ _14418_/A gnd _14418_/Y vdd INVX1
XFILL_5__7696_ gnd vdd FILL
XFILL_4__10905_ gnd vdd FILL
XFILL_5__11155_ gnd vdd FILL
XFILL_3__15122_ gnd vdd FILL
XFILL_0__9790_ gnd vdd FILL
X_15398_ _15398_/A _15395_/Y _15398_/C gnd _15413_/A vdd NAND3X1
XSFILL89320x48050 gnd vdd FILL
XFILL_1__16301_ gnd vdd FILL
XFILL_3__12334_ gnd vdd FILL
XFILL_2__9726_ gnd vdd FILL
XFILL112200x20050 gnd vdd FILL
XFILL_4__11885_ gnd vdd FILL
XFILL_2__6938_ gnd vdd FILL
XFILL_2__15852_ gnd vdd FILL
XFILL_4__14673_ gnd vdd FILL
XFILL_1__13513_ gnd vdd FILL
XFILL_0__12154_ gnd vdd FILL
XFILL_1__14493_ gnd vdd FILL
XFILL_5__10106_ gnd vdd FILL
XFILL_0__8741_ gnd vdd FILL
X_14349_ _10284_/A gnd _14349_/Y vdd INVX1
XFILL_4__16412_ gnd vdd FILL
XFILL_4__13624_ gnd vdd FILL
XFILL_2__14803_ gnd vdd FILL
X_7280_ _7236_/A _7642_/CLK _8676_/R vdd _7280_/D gnd vdd DFFSR
XFILL_3__15053_ gnd vdd FILL
XFILL_5__15963_ gnd vdd FILL
XFILL_5__11086_ gnd vdd FILL
XFILL_4__10836_ gnd vdd FILL
XFILL_1__16232_ gnd vdd FILL
XFILL_3__8450_ gnd vdd FILL
XFILL_2__9657_ gnd vdd FILL
XFILL_3__12265_ gnd vdd FILL
XFILL_0__11105_ gnd vdd FILL
XFILL_1__10656_ gnd vdd FILL
XFILL_1__13444_ gnd vdd FILL
XFILL_2__6869_ gnd vdd FILL
XFILL_2__15783_ gnd vdd FILL
XFILL_0__12085_ gnd vdd FILL
XFILL_2__12995_ gnd vdd FILL
XFILL_5__9366_ gnd vdd FILL
XFILL_5__10037_ gnd vdd FILL
XFILL_3__14004_ gnd vdd FILL
XFILL_5__14914_ gnd vdd FILL
XFILL_4__16343_ gnd vdd FILL
XFILL_2__8608_ gnd vdd FILL
XFILL_4__13555_ gnd vdd FILL
XFILL_3__11216_ gnd vdd FILL
XFILL_4__10767_ gnd vdd FILL
XFILL_5__15894_ gnd vdd FILL
XSFILL13560x43050 gnd vdd FILL
XFILL_2__14734_ gnd vdd FILL
XFILL_3__8381_ gnd vdd FILL
XFILL_0__15913_ gnd vdd FILL
XFILL_2__11946_ gnd vdd FILL
XFILL_6__7110_ gnd vdd FILL
XFILL_3__12196_ gnd vdd FILL
XFILL_0__11036_ gnd vdd FILL
XFILL_5__8317_ gnd vdd FILL
XFILL_1__16163_ gnd vdd FILL
X_16019_ _16019_/A _16018_/Y gnd _16020_/C vdd NOR2X1
XFILL_1__13375_ gnd vdd FILL
XFILL_5__9297_ gnd vdd FILL
XFILL_0__7623_ gnd vdd FILL
XFILL_5__14845_ gnd vdd FILL
XFILL_4__12506_ gnd vdd FILL
XFILL_3__7332_ gnd vdd FILL
XFILL_4__13486_ gnd vdd FILL
XFILL_3__11147_ gnd vdd FILL
XSFILL69240x15050 gnd vdd FILL
XFILL_1__15114_ gnd vdd FILL
XFILL_4__16274_ gnd vdd FILL
XFILL_4__10698_ gnd vdd FILL
XFILL_2__14665_ gnd vdd FILL
XFILL_1__12326_ gnd vdd FILL
XFILL_2__11877_ gnd vdd FILL
XFILL_5__8248_ gnd vdd FILL
XFILL_1__16094_ gnd vdd FILL
XFILL_0__15844_ gnd vdd FILL
XFILL_4__12437_ gnd vdd FILL
XFILL_0__7554_ gnd vdd FILL
XFILL_4__15225_ gnd vdd FILL
XFILL_2__16404_ gnd vdd FILL
XFILL_2__13616_ gnd vdd FILL
XFILL_5__14776_ gnd vdd FILL
XFILL_2__10828_ gnd vdd FILL
XFILL_1__15045_ gnd vdd FILL
XFILL_5__11988_ gnd vdd FILL
XFILL_3__15955_ gnd vdd FILL
XFILL_1__12257_ gnd vdd FILL
XFILL_3__11078_ gnd vdd FILL
XFILL_2__14596_ gnd vdd FILL
XFILL_0__15775_ gnd vdd FILL
XSFILL104440x24050 gnd vdd FILL
XFILL_0__12987_ gnd vdd FILL
X_9921_ _9967_/Q gnd _9921_/Y vdd INVX1
XFILL_4__15156_ gnd vdd FILL
XFILL_5__13727_ gnd vdd FILL
XFILL_3__9002_ gnd vdd FILL
XFILL_5__10939_ gnd vdd FILL
XFILL_4__12368_ gnd vdd FILL
XFILL_0__7485_ gnd vdd FILL
XFILL_2__16335_ gnd vdd FILL
XFILL_3__10029_ gnd vdd FILL
XFILL_3__14906_ gnd vdd FILL
XFILL_2__13547_ gnd vdd FILL
XSFILL8680x22050 gnd vdd FILL
XFILL_1__11208_ gnd vdd FILL
XFILL_1__12188_ gnd vdd FILL
XFILL_3__7194_ gnd vdd FILL
XFILL_0__14726_ gnd vdd FILL
XFILL_2__10759_ gnd vdd FILL
XFILL_3__15886_ gnd vdd FILL
XFILL_0__9224_ gnd vdd FILL
XFILL_0__11938_ gnd vdd FILL
XFILL_4__14107_ gnd vdd FILL
XFILL_4__11319_ gnd vdd FILL
XFILL_6__15997_ gnd vdd FILL
XSFILL8120x65050 gnd vdd FILL
XFILL_5__13658_ gnd vdd FILL
X_9852_ _9852_/A gnd _9852_/Y vdd INVX1
XFILL_4__15087_ gnd vdd FILL
XFILL_3__14837_ gnd vdd FILL
XFILL_4__12299_ gnd vdd FILL
XFILL_1__11139_ gnd vdd FILL
XFILL_2__16266_ gnd vdd FILL
XFILL_2__13478_ gnd vdd FILL
XSFILL59160x67050 gnd vdd FILL
XFILL_0__11869_ gnd vdd FILL
XFILL_0__14657_ gnd vdd FILL
XFILL_5__12609_ gnd vdd FILL
XFILL_4__14038_ gnd vdd FILL
XFILL_6__14948_ gnd vdd FILL
XFILL_0__9155_ gnd vdd FILL
X_8803_ _8733_/A _7515_/CLK _7515_/R vdd _8803_/D gnd vdd DFFSR
XFILL_2__15217_ gnd vdd FILL
XFILL_5__16377_ gnd vdd FILL
X_9783_ _9781_/Y _9789_/B _9783_/C gnd _9835_/D vdd OAI21X1
XFILL_5__13589_ gnd vdd FILL
XFILL_2__12429_ gnd vdd FILL
XFILL_3__14768_ gnd vdd FILL
XSFILL74200x70050 gnd vdd FILL
XFILL_0__13608_ gnd vdd FILL
XFILL_2__16197_ gnd vdd FILL
X_6995_ _7029_/Q gnd _6997_/A vdd INVX1
XFILL_1__15947_ gnd vdd FILL
XFILL_0__8106_ gnd vdd FILL
XFILL_0__14588_ gnd vdd FILL
XFILL111880x66050 gnd vdd FILL
XFILL_5__15328_ gnd vdd FILL
X_8734_ _8698_/A _7326_/B gnd _8735_/C vdd NAND2X1
XFILL_0__9086_ gnd vdd FILL
XFILL_3__9904_ gnd vdd FILL
XFILL_2__15148_ gnd vdd FILL
XFILL_3__13719_ gnd vdd FILL
XSFILL109160x36050 gnd vdd FILL
XFILL_3__14699_ gnd vdd FILL
XFILL_0__16327_ gnd vdd FILL
XFILL_6_BUFX2_insert546 gnd vdd FILL
XFILL_0__13539_ gnd vdd FILL
XSFILL13640x23050 gnd vdd FILL
XFILL_1__15878_ gnd vdd FILL
XFILL_5__15259_ gnd vdd FILL
X_8665_ _8665_/Q _8926_/CLK _8025_/R vdd _8577_/Y gnd vdd DFFSR
XSFILL79080x18050 gnd vdd FILL
XFILL_4__15989_ gnd vdd FILL
XFILL_1__14829_ gnd vdd FILL
XFILL_2__15079_ gnd vdd FILL
XFILL_0__16258_ gnd vdd FILL
XFILL_6__9544_ gnd vdd FILL
X_7616_ _7614_/Y _7568_/B _7615_/Y gnd _7662_/D vdd OAI21X1
XFILL_1__8850_ gnd vdd FILL
XFILL_3__9766_ gnd vdd FILL
XFILL_3__16369_ gnd vdd FILL
XFILL_0__15209_ gnd vdd FILL
X_8596_ _8596_/A gnd _8596_/Y vdd INVX1
XFILL_3__6978_ gnd vdd FILL
XFILL_0__16189_ gnd vdd FILL
XFILL_1__7801_ gnd vdd FILL
XFILL_1__8781_ gnd vdd FILL
XFILL_3__8717_ gnd vdd FILL
XFILL_0__9988_ gnd vdd FILL
X_7547_ _7547_/A _7624_/A _7547_/C gnd _7639_/D vdd OAI21X1
XSFILL33800x2050 gnd vdd FILL
XFILL_4__8490_ gnd vdd FILL
XSFILL33800x36050 gnd vdd FILL
XFILL_1__7732_ gnd vdd FILL
X_7478_ _7503_/B _7222_/B gnd _7478_/Y vdd NAND2X1
XFILL_4__7441_ gnd vdd FILL
XFILL_3__8648_ gnd vdd FILL
X_9217_ _9217_/A _9232_/B _9217_/C gnd _9217_/Y vdd OAI21X1
XFILL_4__7372_ gnd vdd FILL
XFILL_3__8579_ gnd vdd FILL
XFILL_1__9402_ gnd vdd FILL
XFILL_3_BUFX2_insert403 gnd vdd FILL
X_9148_ _9101_/B _9788_/B gnd _9148_/Y vdd NAND2X1
XFILL_4__9111_ gnd vdd FILL
XFILL_1__7594_ gnd vdd FILL
XFILL_3_BUFX2_insert414 gnd vdd FILL
XFILL111960x46050 gnd vdd FILL
XFILL_3_BUFX2_insert425 gnd vdd FILL
X_10030_ _10028_/Y _9993_/A _10030_/C gnd _10088_/D vdd OAI21X1
XFILL_3_BUFX2_insert436 gnd vdd FILL
XFILL_6__7239_ gnd vdd FILL
XFILL_3_BUFX2_insert447 gnd vdd FILL
X_9079_ _8567_/A _9151_/A gnd _9080_/C vdd NAND2X1
XFILL_3_BUFX2_insert458 gnd vdd FILL
XFILL_4__9042_ gnd vdd FILL
XFILL_3_BUFX2_insert469 gnd vdd FILL
XFILL_1__9264_ gnd vdd FILL
XFILL_1__8215_ gnd vdd FILL
X_11981_ _11895_/B _12436_/A gnd _11982_/C vdd NAND2X1
X_13720_ _8411_/Q gnd _13722_/A vdd INVX1
X_10932_ _12818_/Q gnd _10934_/B vdd INVX1
XFILL_1__8146_ gnd vdd FILL
XFILL_0_BUFX2_insert8 gnd vdd FILL
X_13651_ _13879_/B _13649_/Y _14849_/B _15226_/B gnd _13651_/Y vdd OAI22X1
X_10863_ _16071_/A _7007_/CLK _9332_/R vdd _10819_/Y gnd vdd DFFSR
XFILL_4_CLKBUF1_insert204 gnd vdd FILL
XFILL_4_CLKBUF1_insert215 gnd vdd FILL
XFILL_1__8077_ gnd vdd FILL
X_12602_ _12602_/A vdd _12602_/C gnd _12674_/D vdd OAI21X1
X_16370_ gnd gnd gnd _16371_/C vdd NAND2X1
XFILL_4__9875_ gnd vdd FILL
X_13582_ _13582_/A _13582_/B _13582_/C gnd _13582_/Y vdd NAND3X1
X_10794_ _10797_/A _9258_/B gnd _10795_/C vdd NAND2X1
XFILL_0_BUFX2_insert304 gnd vdd FILL
XFILL_2__8890_ gnd vdd FILL
XFILL111960x5050 gnd vdd FILL
X_15321_ _16036_/A _15321_/B _15321_/C _15321_/D gnd _15321_/Y vdd OAI22X1
XFILL_4__8826_ gnd vdd FILL
XFILL_0_BUFX2_insert315 gnd vdd FILL
XFILL_0_BUFX2_insert326 gnd vdd FILL
X_12533_ vdd _12113_/A gnd _12533_/Y vdd NAND2X1
XFILL_0_BUFX2_insert337 gnd vdd FILL
XFILL_2__7841_ gnd vdd FILL
XFILL_0_BUFX2_insert348 gnd vdd FILL
XFILL_4__8757_ gnd vdd FILL
XFILL_5__7550_ gnd vdd FILL
XFILL_0_BUFX2_insert359 gnd vdd FILL
X_15252_ _8282_/Q gnd _15252_/Y vdd INVX1
X_12464_ vdd _12021_/A gnd _12464_/Y vdd NAND2X1
XSFILL23800x68050 gnd vdd FILL
XFILL_3__10380_ gnd vdd FILL
XFILL_1__8979_ gnd vdd FILL
X_14203_ _14203_/A _14203_/B _14203_/C _14203_/D gnd _14203_/Y vdd OAI22X1
XFILL_4__7708_ gnd vdd FILL
XFILL_5__7481_ gnd vdd FILL
X_11415_ _11414_/A _11369_/Y _11415_/C gnd _11416_/A vdd OAI21X1
X_15183_ _15183_/A _15183_/B gnd _15184_/C vdd NOR2X1
XFILL_2__9511_ gnd vdd FILL
XFILL_1__10510_ gnd vdd FILL
X_12395_ _12395_/A _12618_/A gnd _12396_/C vdd NAND2X1
XFILL_4__11670_ gnd vdd FILL
XFILL_5__9220_ gnd vdd FILL
XSFILL64040x20050 gnd vdd FILL
XFILL_1__11490_ gnd vdd FILL
X_14134_ _9376_/A _13883_/B _14878_/C _10596_/Q gnd _14143_/A vdd AOI22X1
XFILL_4__10621_ gnd vdd FILL
X_11346_ _10997_/Y _11343_/Y _11346_/C gnd _11346_/Y vdd AOI21X1
XFILL_5__12960_ gnd vdd FILL
XFILL_3__12050_ gnd vdd FILL
XFILL_2__11800_ gnd vdd FILL
XFILL_1__10441_ gnd vdd FILL
XFILL_2__12780_ gnd vdd FILL
XFILL_5__9151_ gnd vdd FILL
XFILL_4_BUFX2_insert270 gnd vdd FILL
XFILL_4__13340_ gnd vdd FILL
XFILL_5__11911_ gnd vdd FILL
X_14065_ _8290_/Q _13592_/A _14065_/C _15545_/A gnd _14065_/Y vdd AOI22X1
XFILL_3__11001_ gnd vdd FILL
XFILL_4_BUFX2_insert281 gnd vdd FILL
XFILL_4__10552_ gnd vdd FILL
X_11277_ _12270_/Y gnd _11278_/A vdd INVX1
XFILL_4_BUFX2_insert292 gnd vdd FILL
XFILL_5__8102_ gnd vdd FILL
XSFILL53880x63050 gnd vdd FILL
XFILL_5__12891_ gnd vdd FILL
XFILL_1__13160_ gnd vdd FILL
XFILL_5_BUFX2_insert1005 gnd vdd FILL
XFILL_2__9373_ gnd vdd FILL
XFILL_2__11731_ gnd vdd FILL
XFILL_5_BUFX2_insert1016 gnd vdd FILL
XFILL_0__12910_ gnd vdd FILL
XFILL_1__10372_ gnd vdd FILL
XSFILL68680x23050 gnd vdd FILL
X_13016_ _13014_/Y vdd _13016_/C gnd _13068_/D vdd OAI21X1
XFILL_5__9082_ gnd vdd FILL
XFILL_5__14630_ gnd vdd FILL
XFILL_0__13890_ gnd vdd FILL
X_10228_ _10192_/A _7156_/CLK _7775_/R vdd _10194_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert1027 gnd vdd FILL
XFILL_4__13271_ gnd vdd FILL
XFILL_5_BUFX2_insert1038 gnd vdd FILL
XFILL_2__8324_ gnd vdd FILL
XFILL_1__12111_ gnd vdd FILL
XFILL_5__11842_ gnd vdd FILL
XFILL_5_BUFX2_insert1049 gnd vdd FILL
XFILL_2__14450_ gnd vdd FILL
XFILL_1__13091_ gnd vdd FILL
XFILL_2__11662_ gnd vdd FILL
XFILL_6__15920_ gnd vdd FILL
XFILL_0__12841_ gnd vdd FILL
XFILL_4__15010_ gnd vdd FILL
XSFILL84200x33050 gnd vdd FILL
XFILL_3_BUFX2_insert970 gnd vdd FILL
XFILL_4__12222_ gnd vdd FILL
XFILL_5__14561_ gnd vdd FILL
XFILL_2__13401_ gnd vdd FILL
X_10159_ _10159_/A gnd _10161_/A vdd INVX1
XFILL_3_BUFX2_insert981 gnd vdd FILL
XFILL_2__8255_ gnd vdd FILL
XFILL_3_BUFX2_insert992 gnd vdd FILL
XSFILL104360x39050 gnd vdd FILL
XFILL_3__12952_ gnd vdd FILL
XFILL_1__12042_ gnd vdd FILL
XFILL_3__15740_ gnd vdd FILL
XFILL_5__11773_ gnd vdd FILL
XFILL_2__14381_ gnd vdd FILL
XFILL_0__12772_ gnd vdd FILL
XFILL_0__15560_ gnd vdd FILL
XFILL_5__16300_ gnd vdd FILL
XFILL_2__11593_ gnd vdd FILL
XFILL_5__13512_ gnd vdd FILL
XFILL_2__7206_ gnd vdd FILL
XFILL_2__16120_ gnd vdd FILL
XFILL_3__11903_ gnd vdd FILL
XFILL_4__12153_ gnd vdd FILL
X_14967_ _14967_/A _14320_/C gnd _14968_/C vdd NOR2X1
XFILL_5__14492_ gnd vdd FILL
XFILL_2__13332_ gnd vdd FILL
XFILL_3__15671_ gnd vdd FILL
XFILL_0__14511_ gnd vdd FILL
XFILL_2__10544_ gnd vdd FILL
XFILL_0__11723_ gnd vdd FILL
XSFILL79320x7050 gnd vdd FILL
XFILL_2__8186_ gnd vdd FILL
XFILL_3__12883_ gnd vdd FILL
XFILL_5__16231_ gnd vdd FILL
XSFILL88840x36050 gnd vdd FILL
XFILL_4__11104_ gnd vdd FILL
XFILL_0__15491_ gnd vdd FILL
XFILL_5__9984_ gnd vdd FILL
XFILL_3__14622_ gnd vdd FILL
XFILL_5__13443_ gnd vdd FILL
XFILL_6__15782_ gnd vdd FILL
X_13918_ _13909_/Y _13918_/B _13918_/C gnd _13929_/A vdd NAND3X1
XFILL_3_BUFX2_insert1020 gnd vdd FILL
XFILL_4__12084_ gnd vdd FILL
XFILL_1__15801_ gnd vdd FILL
XFILL_5__10655_ gnd vdd FILL
XFILL_2__16051_ gnd vdd FILL
XFILL_3__11834_ gnd vdd FILL
X_14898_ _14897_/Y _14898_/B gnd _14906_/A vdd NOR2X1
XFILL_2__13263_ gnd vdd FILL
XFILL_3_BUFX2_insert1031 gnd vdd FILL
XFILL_0__11654_ gnd vdd FILL
XFILL_0__14442_ gnd vdd FILL
XFILL_3_BUFX2_insert1042 gnd vdd FILL
XFILL_1__13993_ gnd vdd FILL
XFILL_6__14733_ gnd vdd FILL
X_13849_ _7518_/Q gnd _13850_/A vdd INVX1
XFILL_4__15912_ gnd vdd FILL
XFILL_3_BUFX2_insert1053 gnd vdd FILL
XSFILL49320x59050 gnd vdd FILL
XFILL_2__15002_ gnd vdd FILL
XFILL_5__16162_ gnd vdd FILL
XFILL_4__11035_ gnd vdd FILL
XFILL_3__14553_ gnd vdd FILL
XFILL_3_BUFX2_insert1064 gnd vdd FILL
XFILL_5__13374_ gnd vdd FILL
XFILL_2__12214_ gnd vdd FILL
XFILL_3__7950_ gnd vdd FILL
XFILL_1__15732_ gnd vdd FILL
XFILL_2__7068_ gnd vdd FILL
XFILL_3__11765_ gnd vdd FILL
XFILL_0__14373_ gnd vdd FILL
XFILL_3_BUFX2_insert1086 gnd vdd FILL
XFILL_0__11585_ gnd vdd FILL
XFILL_5__15113_ gnd vdd FILL
XFILL_5__8866_ gnd vdd FILL
XFILL_3__13504_ gnd vdd FILL
XFILL_5__12325_ gnd vdd FILL
XFILL_6__11876_ gnd vdd FILL
XFILL_5__16093_ gnd vdd FILL
XFILL_3__6901_ gnd vdd FILL
XFILL_4__15843_ gnd vdd FILL
XFILL_0__13324_ gnd vdd FILL
XFILL_3__14484_ gnd vdd FILL
XFILL_0__16112_ gnd vdd FILL
XFILL_2__12145_ gnd vdd FILL
XFILL_0__10536_ gnd vdd FILL
XFILL_1__15663_ gnd vdd FILL
XFILL_3__11696_ gnd vdd FILL
XFILL_3__7881_ gnd vdd FILL
XFILL_0__9911_ gnd vdd FILL
XFILL_5__7817_ gnd vdd FILL
XFILL_1__12875_ gnd vdd FILL
XFILL_6__10827_ gnd vdd FILL
X_15519_ _9367_/A _15636_/B _15995_/C gnd _15520_/C vdd NAND3X1
XFILL_5__15044_ gnd vdd FILL
XSFILL53960x43050 gnd vdd FILL
XFILL_5_BUFX2_insert509 gnd vdd FILL
XFILL_6__14595_ gnd vdd FILL
XFILL_3__16223_ gnd vdd FILL
X_8450_ _8450_/A gnd _8452_/A vdd INVX1
XFILL_3__13435_ gnd vdd FILL
XFILL_5__12256_ gnd vdd FILL
XFILL_3__9620_ gnd vdd FILL
XFILL_1__14614_ gnd vdd FILL
XFILL_3__10647_ gnd vdd FILL
XFILL_4__15774_ gnd vdd FILL
XFILL_0__13255_ gnd vdd FILL
XFILL_0__16043_ gnd vdd FILL
XFILL_2__12076_ gnd vdd FILL
XFILL_4__12986_ gnd vdd FILL
XFILL_1__11826_ gnd vdd FILL
XFILL_6__16334_ gnd vdd FILL
XFILL_1__15594_ gnd vdd FILL
XFILL_0_BUFX2_insert860 gnd vdd FILL
X_7401_ _7401_/Q _9328_/CLK _7408_/R vdd _7345_/Y gnd vdd DFFSR
XFILL_6__13546_ gnd vdd FILL
XFILL_5__11207_ gnd vdd FILL
XFILL_5__7748_ gnd vdd FILL
X_8381_ _8381_/A _8360_/B _8380_/Y gnd _8429_/D vdd OAI21X1
XFILL_5__12187_ gnd vdd FILL
XFILL_0_BUFX2_insert871 gnd vdd FILL
XFILL_4__14725_ gnd vdd FILL
XFILL_3__16154_ gnd vdd FILL
XFILL_3__9551_ gnd vdd FILL
XFILL_2__15904_ gnd vdd FILL
XFILL_3__13366_ gnd vdd FILL
XFILL_4__11937_ gnd vdd FILL
XFILL_0__12206_ gnd vdd FILL
XFILL_0_BUFX2_insert882 gnd vdd FILL
XFILL_2__11027_ gnd vdd FILL
XSFILL54040x52050 gnd vdd FILL
XFILL_1__14545_ gnd vdd FILL
XFILL_3__10578_ gnd vdd FILL
XFILL_0_BUFX2_insert893 gnd vdd FILL
XFILL_6__9260_ gnd vdd FILL
XFILL_1__11757_ gnd vdd FILL
XFILL_5__7679_ gnd vdd FILL
X_7332_ _7359_/A _8356_/B gnd _7333_/C vdd NAND2X1
XFILL_0__10398_ gnd vdd FILL
XFILL_5__11138_ gnd vdd FILL
XFILL_3__15105_ gnd vdd FILL
XFILL_3__8502_ gnd vdd FILL
XFILL_3_BUFX2_insert20 gnd vdd FILL
XFILL_0__9773_ gnd vdd FILL
XFILL_3__12317_ gnd vdd FILL
XFILL_3_BUFX2_insert31 gnd vdd FILL
XFILL_1_BUFX2_insert1090 gnd vdd FILL
XFILL_4__14656_ gnd vdd FILL
XFILL_3__16085_ gnd vdd FILL
XFILL_0__6985_ gnd vdd FILL
XFILL_3__13297_ gnd vdd FILL
XFILL_0__12137_ gnd vdd FILL
XFILL_3__9482_ gnd vdd FILL
XFILL_3_BUFX2_insert42 gnd vdd FILL
XFILL_2__15835_ gnd vdd FILL
XFILL_4__11868_ gnd vdd FILL
XFILL_1__10708_ gnd vdd FILL
XFILL_6__8211_ gnd vdd FILL
XSFILL8680x17050 gnd vdd FILL
XFILL_1__14476_ gnd vdd FILL
XFILL_5__9418_ gnd vdd FILL
XFILL_6__12428_ gnd vdd FILL
XFILL_3_BUFX2_insert53 gnd vdd FILL
XFILL_0__8724_ gnd vdd FILL
XFILL_1__11688_ gnd vdd FILL
XFILL_4__13607_ gnd vdd FILL
XFILL_6__16196_ gnd vdd FILL
XFILL_3__15036_ gnd vdd FILL
XFILL_5__15946_ gnd vdd FILL
XFILL_3_BUFX2_insert64 gnd vdd FILL
XFILL_5__11069_ gnd vdd FILL
X_7263_ _7185_/A _7274_/CLK _7274_/R vdd _7187_/Y gnd vdd DFFSR
XSFILL33880x10050 gnd vdd FILL
XFILL_3_BUFX2_insert75 gnd vdd FILL
XFILL_1__16215_ gnd vdd FILL
XFILL_3__12248_ gnd vdd FILL
XFILL_4__10819_ gnd vdd FILL
XFILL_4__14587_ gnd vdd FILL
XFILL_1__13427_ gnd vdd FILL
XFILL_3_BUFX2_insert86 gnd vdd FILL
XFILL_2__15766_ gnd vdd FILL
XFILL_4__11799_ gnd vdd FILL
XFILL_1__10639_ gnd vdd FILL
XFILL_0__12068_ gnd vdd FILL
XFILL_2__12978_ gnd vdd FILL
XFILL_3_BUFX2_insert97 gnd vdd FILL
XFILL_6__15147_ gnd vdd FILL
XFILL_5__9349_ gnd vdd FILL
X_9002_ _9005_/A _7594_/B gnd _9002_/Y vdd NAND2X1
XFILL_0__8655_ gnd vdd FILL
XFILL_4__16326_ gnd vdd FILL
X_7194_ _7194_/A gnd _7196_/A vdd INVX1
XFILL_2__14717_ gnd vdd FILL
XSFILL48920x32050 gnd vdd FILL
XFILL_4__13538_ gnd vdd FILL
XFILL_5__15877_ gnd vdd FILL
XSFILL18680x71050 gnd vdd FILL
XFILL_3__12179_ gnd vdd FILL
XFILL_2__11929_ gnd vdd FILL
XFILL_3__8364_ gnd vdd FILL
XFILL_0__11019_ gnd vdd FILL
XFILL_1__16146_ gnd vdd FILL
XSFILL19160x78050 gnd vdd FILL
XFILL_1__13358_ gnd vdd FILL
XFILL_2__15697_ gnd vdd FILL
XSFILL69160x50 gnd vdd FILL
XFILL_0__7606_ gnd vdd FILL
XSFILL74200x65050 gnd vdd FILL
XFILL_5__14828_ gnd vdd FILL
XFILL_0__8586_ gnd vdd FILL
XFILL_3__7315_ gnd vdd FILL
XFILL_4__16257_ gnd vdd FILL
XFILL_4__13469_ gnd vdd FILL
XFILL_1__12309_ gnd vdd FILL
XFILL_2__14648_ gnd vdd FILL
XFILL_0__15827_ gnd vdd FILL
XFILL_1__16077_ gnd vdd FILL
XFILL_1__13289_ gnd vdd FILL
XSFILL49000x41050 gnd vdd FILL
XFILL_4__15208_ gnd vdd FILL
XSFILL13640x18050 gnd vdd FILL
XFILL_5__14759_ gnd vdd FILL
XFILL_3__7246_ gnd vdd FILL
XFILL_4__16188_ gnd vdd FILL
XFILL_1__15028_ gnd vdd FILL
XFILL_3__15938_ gnd vdd FILL
XFILL_2__14579_ gnd vdd FILL
XFILL_0__15758_ gnd vdd FILL
X_9904_ _9896_/B _6960_/B gnd _9905_/C vdd NAND2X1
XFILL_2__16318_ gnd vdd FILL
XFILL_0__7468_ gnd vdd FILL
XFILL_4__15139_ gnd vdd FILL
XFILL_3__7177_ gnd vdd FILL
XFILL_0__14709_ gnd vdd FILL
XFILL_3__15869_ gnd vdd FILL
XFILL_1__8000_ gnd vdd FILL
XFILL_0__9207_ gnd vdd FILL
XFILL_0__15689_ gnd vdd FILL
XSFILL54120x32050 gnd vdd FILL
X_9835_ _9835_/Q _9195_/CLK _8051_/R vdd _9835_/D gnd vdd DFFSR
XFILL_2__16249_ gnd vdd FILL
XFILL_4__7990_ gnd vdd FILL
XFILL_0__9138_ gnd vdd FILL
XSFILL114680x43050 gnd vdd FILL
X_9766_ _9766_/A gnd _9768_/A vdd INVX1
XFILL_6_BUFX2_insert321 gnd vdd FILL
X_6978_ _6982_/B _6978_/B gnd _6979_/C vdd NAND2X1
XFILL_4__6941_ gnd vdd FILL
XSFILL43960x75050 gnd vdd FILL
X_8717_ _8717_/A _8759_/B _8716_/Y gnd _8717_/Y vdd OAI21X1
XBUFX2_insert409 _10920_/Y gnd _12419_/A vdd BUFX2
XSFILL28760x9050 gnd vdd FILL
XFILL_4__9660_ gnd vdd FILL
X_9697_ _9623_/A _9188_/CLK _8929_/R vdd _9697_/D gnd vdd DFFSR
XSFILL84040x68050 gnd vdd FILL
XFILL_4__6872_ gnd vdd FILL
XFILL_1__8902_ gnd vdd FILL
XSFILL18760x51050 gnd vdd FILL
XSFILL8600x61050 gnd vdd FILL
XFILL_1__9882_ gnd vdd FILL
XFILL_6_BUFX2_insert398 gnd vdd FILL
XFILL_4__8611_ gnd vdd FILL
X_8648_ _8607_/B _7240_/B gnd _8649_/C vdd NAND2X1
XFILL_4__9591_ gnd vdd FILL
XFILL_1__8833_ gnd vdd FILL
XSFILL94680x7050 gnd vdd FILL
X_8579_ _8589_/B _9475_/B gnd _8579_/Y vdd NAND2X1
XFILL_3__9749_ gnd vdd FILL
XFILL_1__8764_ gnd vdd FILL
XSFILL23880x42050 gnd vdd FILL
XFILL_4__8473_ gnd vdd FILL
X_11200_ _11198_/Y _11199_/Y gnd _11200_/Y vdd NOR2X1
XFILL_1__7715_ gnd vdd FILL
X_12180_ _12178_/Y _12179_/A _12180_/C gnd _12180_/Y vdd OAI21X1
XSFILL38120x45050 gnd vdd FILL
XFILL_6__9389_ gnd vdd FILL
XFILL_4__7424_ gnd vdd FILL
XSFILL38920x64050 gnd vdd FILL
XFILL_1__8695_ gnd vdd FILL
XFILL112440x71050 gnd vdd FILL
X_11131_ _12168_/Y _11150_/B gnd _11300_/A vdd NAND2X1
XFILL_4__7355_ gnd vdd FILL
XSFILL39000x73050 gnd vdd FILL
X_11062_ _12270_/Y _12156_/Y gnd _11062_/Y vdd XNOR2X1
XSFILL89320x2050 gnd vdd FILL
XFILL_3_BUFX2_insert233 gnd vdd FILL
XFILL_3_BUFX2_insert244 gnd vdd FILL
XFILL_1__7577_ gnd vdd FILL
XFILL_3_BUFX2_insert255 gnd vdd FILL
XFILL_4__7286_ gnd vdd FILL
X_10013_ _14098_/C gnd _10015_/A vdd INVX1
XFILL_3_BUFX2_insert266 gnd vdd FILL
X_15870_ _15870_/A _15622_/A _15948_/D _15870_/D gnd _15870_/Y vdd OAI22X1
XFILL_3_BUFX2_insert277 gnd vdd FILL
XFILL_2_BUFX2_insert900 gnd vdd FILL
XFILL_3_BUFX2_insert288 gnd vdd FILL
XFILL_4__9025_ gnd vdd FILL
XFILL_3_BUFX2_insert299 gnd vdd FILL
XSFILL18840x31050 gnd vdd FILL
X_14821_ _14180_/C _16187_/A _8522_/A _13771_/D gnd _14821_/Y vdd AOI22X1
XFILL_2_BUFX2_insert911 gnd vdd FILL
XFILL_2_BUFX2_insert922 gnd vdd FILL
XFILL_1__9247_ gnd vdd FILL
XFILL_2_BUFX2_insert933 gnd vdd FILL
XFILL_2_BUFX2_insert944 gnd vdd FILL
XFILL_2_BUFX2_insert955 gnd vdd FILL
XFILL_2_BUFX2_insert966 gnd vdd FILL
X_14752_ _13456_/A _14750_/Y _14752_/C _14751_/Y gnd _14753_/B vdd OAI22X1
XSFILL89800x8050 gnd vdd FILL
XFILL_2_BUFX2_insert977 gnd vdd FILL
X_11964_ _11962_/Y _11895_/B _11964_/C gnd _6863_/A vdd OAI21X1
XFILL_2_BUFX2_insert988 gnd vdd FILL
XFILL_2_BUFX2_insert999 gnd vdd FILL
X_13703_ _9691_/Q gnd _13704_/D vdd INVX1
X_10915_ _10915_/A _10920_/B gnd _10915_/Y vdd NOR2X1
XFILL_5__6981_ gnd vdd FILL
XFILL_5__10440_ gnd vdd FILL
XFILL_1__8129_ gnd vdd FILL
X_14683_ _14683_/A _13868_/B _13467_/A _16083_/B gnd _14687_/A vdd OAI22X1
X_11895_ _11895_/A _11895_/B _11895_/C gnd _6840_/A vdd OAI21X1
XFILL_2__10260_ gnd vdd FILL
XFILL_2__9991_ gnd vdd FILL
XFILL_5__8720_ gnd vdd FILL
XSFILL64040x15050 gnd vdd FILL
XFILL_4__9927_ gnd vdd FILL
X_13634_ _13634_/A _13633_/Y gnd _13634_/Y vdd NOR2X1
XFILL_1__10990_ gnd vdd FILL
X_16422_ _15275_/A _8792_/CLK _7896_/R vdd _16338_/Y gnd vdd DFFSR
XSFILL89640x79050 gnd vdd FILL
X_10846_ _10846_/Q _7781_/CLK _9566_/R vdd _10846_/D gnd vdd DFFSR
XFILL_5__10371_ gnd vdd FILL
XFILL_3__11550_ gnd vdd FILL
XFILL_2__10191_ gnd vdd FILL
XSFILL24040x31050 gnd vdd FILL
XBUFX2_insert910 _10913_/Y gnd _12718_/B vdd BUFX2
XFILL_5__8651_ gnd vdd FILL
XFILL_0_BUFX2_insert101 gnd vdd FILL
XSFILL39640x10050 gnd vdd FILL
XFILL_0__11370_ gnd vdd FILL
XFILL_4__9858_ gnd vdd FILL
XBUFX2_insert921 _13370_/Y gnd _14180_/C vdd BUFX2
XFILL_5__12110_ gnd vdd FILL
X_16353_ _16353_/A gnd _16352_/Y gnd _16353_/Y vdd OAI21X1
XFILL_5__13090_ gnd vdd FILL
XFILL_3__10501_ gnd vdd FILL
XFILL_6__11661_ gnd vdd FILL
XSFILL13800x50 gnd vdd FILL
X_13565_ _7548_/A gnd _13565_/Y vdd INVX1
XBUFX2_insert932 _12435_/Y gnd _8529_/B vdd BUFX2
X_10777_ _10777_/A _10792_/B _10777_/C gnd _10777_/Y vdd OAI21X1
XFILL_4__12840_ gnd vdd FILL
XSFILL89240x81050 gnd vdd FILL
XFILL_2__8873_ gnd vdd FILL
XFILL_0__10321_ gnd vdd FILL
XFILL_3__11481_ gnd vdd FILL
XBUFX2_insert943 _12426_/Y gnd _7240_/B vdd BUFX2
XBUFX2_insert954 _13365_/Y gnd _10789_/B vdd BUFX2
XFILL_1__12660_ gnd vdd FILL
X_15304_ _7004_/Q _15382_/B _16096_/C _7388_/Q gnd _15309_/A vdd AOI22X1
XFILL_5__7602_ gnd vdd FILL
XBUFX2_insert965 _13361_/Y gnd _10443_/A vdd BUFX2
X_12516_ _12516_/A vdd _12515_/Y gnd _12516_/Y vdd OAI21X1
XFILL_5__12041_ gnd vdd FILL
XFILL_5__8582_ gnd vdd FILL
XFILL_4__9789_ gnd vdd FILL
XFILL_3__13220_ gnd vdd FILL
XBUFX2_insert976 _16451_/Y gnd _13108_/B vdd BUFX2
X_16284_ _15652_/A _9555_/A _9683_/A _15652_/D gnd _16286_/B vdd AOI22X1
XFILL_6__14380_ gnd vdd FILL
XFILL_2__7824_ gnd vdd FILL
XFILL_4__12771_ gnd vdd FILL
XFILL_3__10432_ gnd vdd FILL
X_13496_ _16324_/A gnd _13496_/Y vdd INVX1
XBUFX2_insert987 _13351_/Y gnd _9979_/B vdd BUFX2
XFILL_0__13040_ gnd vdd FILL
XFILL_1__11611_ gnd vdd FILL
XFILL_2__13950_ gnd vdd FILL
XFILL_0__10252_ gnd vdd FILL
XBUFX2_insert998 _14998_/Y gnd _15920_/C vdd BUFX2
XFILL_6__13331_ gnd vdd FILL
XFILL_1__12591_ gnd vdd FILL
X_15235_ _15235_/A gnd _15235_/Y vdd INVX1
X_12447_ _12447_/A vdd _12446_/Y gnd _12447_/Y vdd OAI21X1
XFILL_4__14510_ gnd vdd FILL
XFILL_6__10543_ gnd vdd FILL
XSFILL84200x28050 gnd vdd FILL
XFILL_3__13151_ gnd vdd FILL
XFILL_2__12901_ gnd vdd FILL
XFILL_4__11722_ gnd vdd FILL
XFILL_2__7755_ gnd vdd FILL
XFILL_1__14330_ gnd vdd FILL
XFILL_3__10363_ gnd vdd FILL
XFILL_4__15490_ gnd vdd FILL
XFILL_2__13881_ gnd vdd FILL
XSFILL94360x72050 gnd vdd FILL
XFILL_1__11542_ gnd vdd FILL
XFILL_5__7464_ gnd vdd FILL
XFILL_5__15800_ gnd vdd FILL
XFILL_0__10183_ gnd vdd FILL
XFILL_3__12102_ gnd vdd FILL
X_15166_ _15166_/A _15166_/B _15165_/Y gnd _15167_/B vdd NOR3X1
XFILL_2__15620_ gnd vdd FILL
X_12378_ _12376_/Y _12419_/A _12378_/C gnd _12378_/Y vdd OAI21X1
XFILL_4__11653_ gnd vdd FILL
XFILL_4__14441_ gnd vdd FILL
XFILL_2__12832_ gnd vdd FILL
XFILL_5__13992_ gnd vdd FILL
XFILL_3__13082_ gnd vdd FILL
XFILL_3__10294_ gnd vdd FILL
XFILL_1__14261_ gnd vdd FILL
XFILL_2__7686_ gnd vdd FILL
XFILL_1__11473_ gnd vdd FILL
XFILL_6__12213_ gnd vdd FILL
X_14117_ _9059_/Q gnd _14118_/D vdd INVX1
XFILL_5__15731_ gnd vdd FILL
XFILL_0__14991_ gnd vdd FILL
X_11329_ _11173_/Y _11167_/Y _11171_/Y gnd _11330_/C vdd OAI21X1
XFILL_1__16000_ gnd vdd FILL
X_15097_ _15687_/A gnd _15978_/C vdd INVX8
XFILL_3__12033_ gnd vdd FILL
XFILL_2__9425_ gnd vdd FILL
XFILL_1__13212_ gnd vdd FILL
XFILL_2__15551_ gnd vdd FILL
XFILL_4__14372_ gnd vdd FILL
XFILL_4__11584_ gnd vdd FILL
XFILL_2__12763_ gnd vdd FILL
XFILL_1__10424_ gnd vdd FILL
XFILL_5__9134_ gnd vdd FILL
XFILL_1__14192_ gnd vdd FILL
XFILL_0__13942_ gnd vdd FILL
XFILL_0__8440_ gnd vdd FILL
X_14048_ _14047_/Y _14048_/B gnd _14075_/B vdd NOR2X1
XFILL_4__16111_ gnd vdd FILL
XFILL_4__10535_ gnd vdd FILL
XFILL_4__13323_ gnd vdd FILL
XFILL_5__15662_ gnd vdd FILL
XFILL_2__14502_ gnd vdd FILL
XFILL_2__9356_ gnd vdd FILL
XFILL_5__12874_ gnd vdd FILL
XFILL_2__11714_ gnd vdd FILL
XFILL_1__13143_ gnd vdd FILL
XFILL_2__15482_ gnd vdd FILL
XFILL_0__13873_ gnd vdd FILL
XFILL_5__14613_ gnd vdd FILL
XFILL_3__7100_ gnd vdd FILL
XFILL_4__13254_ gnd vdd FILL
XFILL_4__16042_ gnd vdd FILL
XFILL_6__12075_ gnd vdd FILL
XFILL_0__8371_ gnd vdd FILL
XFILL_5__11825_ gnd vdd FILL
XFILL_5__15593_ gnd vdd FILL
XFILL_2__14433_ gnd vdd FILL
XFILL_3__8080_ gnd vdd FILL
XFILL_0__15612_ gnd vdd FILL
XFILL_2__9287_ gnd vdd FILL
XFILL_2__11645_ gnd vdd FILL
XFILL_5__8016_ gnd vdd FILL
XFILL_3__13984_ gnd vdd FILL
XFILL_0__12824_ gnd vdd FILL
XFILL_1__10286_ gnd vdd FILL
XSFILL89320x61050 gnd vdd FILL
XFILL_0__7322_ gnd vdd FILL
XFILL_4__12205_ gnd vdd FILL
XFILL_6__11026_ gnd vdd FILL
XFILL_5__14544_ gnd vdd FILL
X_7950_ _8030_/Q gnd _7950_/Y vdd INVX1
XFILL_3__15723_ gnd vdd FILL
XFILL_3__7031_ gnd vdd FILL
XFILL_2__8238_ gnd vdd FILL
XFILL_5__11756_ gnd vdd FILL
X_15999_ _8301_/Q gnd _16000_/B vdd INVX1
XFILL_1__12025_ gnd vdd FILL
XFILL_2__14364_ gnd vdd FILL
XFILL_4__10397_ gnd vdd FILL
XFILL_0__15543_ gnd vdd FILL
XFILL_2__11576_ gnd vdd FILL
XSFILL93560x24050 gnd vdd FILL
XFILL_0__12755_ gnd vdd FILL
XFILL_4__12136_ gnd vdd FILL
XFILL_2__16103_ gnd vdd FILL
XFILL_5__10707_ gnd vdd FILL
X_6901_ _6901_/A gnd memoryWriteData[31] vdd BUFX2
XFILL_0__7253_ gnd vdd FILL
XFILL_2__13315_ gnd vdd FILL
XFILL_5__14475_ gnd vdd FILL
XSFILL28760x14050 gnd vdd FILL
XFILL_3__15654_ gnd vdd FILL
XFILL_3__12866_ gnd vdd FILL
XFILL_5__11687_ gnd vdd FILL
XFILL_2__10527_ gnd vdd FILL
X_7881_ _7881_/A _7892_/A _7880_/Y gnd _7881_/Y vdd OAI21X1
XFILL_0__11706_ gnd vdd FILL
XFILL_2__14295_ gnd vdd FILL
XFILL_5__16214_ gnd vdd FILL
XFILL_0__15474_ gnd vdd FILL
XFILL_5__13426_ gnd vdd FILL
X_9620_ _9696_/Q gnd _9622_/A vdd INVX1
XFILL_5__10638_ gnd vdd FILL
XFILL_0__7184_ gnd vdd FILL
XFILL_3__14605_ gnd vdd FILL
XFILL_2__16034_ gnd vdd FILL
XSFILL94440x52050 gnd vdd FILL
XFILL_4__12067_ gnd vdd FILL
XFILL_3__11817_ gnd vdd FILL
XFILL_2__13246_ gnd vdd FILL
XFILL_3__8982_ gnd vdd FILL
XFILL_3__15585_ gnd vdd FILL
XFILL_0__14425_ gnd vdd FILL
XFILL_1__13976_ gnd vdd FILL
XFILL_0__11637_ gnd vdd FILL
XFILL_4__11018_ gnd vdd FILL
XFILL_5__16145_ gnd vdd FILL
X_9551_ _9551_/A _9551_/B _9550_/Y gnd _9587_/D vdd OAI21X1
XFILL_5__13357_ gnd vdd FILL
XFILL_5__9898_ gnd vdd FILL
XFILL_1__15715_ gnd vdd FILL
XFILL_3__14536_ gnd vdd FILL
XFILL_3__7933_ gnd vdd FILL
XFILL_3__11748_ gnd vdd FILL
XFILL_5__10569_ gnd vdd FILL
XFILL_0__14356_ gnd vdd FILL
XFILL_2__10389_ gnd vdd FILL
XFILL_0__11568_ gnd vdd FILL
X_8502_ _8503_/B _8630_/B gnd _8502_/Y vdd NAND2X1
XFILL_5__12308_ gnd vdd FILL
XFILL_5__8849_ gnd vdd FILL
XFILL_4__15826_ gnd vdd FILL
XFILL_5__16076_ gnd vdd FILL
XFILL_5__13288_ gnd vdd FILL
XFILL_3__14467_ gnd vdd FILL
X_9482_ _9482_/A _9535_/A _9482_/C gnd _9564_/D vdd OAI21X1
XFILL_5_BUFX2_insert306 gnd vdd FILL
XFILL_2__12128_ gnd vdd FILL
XFILL_0__13307_ gnd vdd FILL
XFILL_1__15646_ gnd vdd FILL
XFILL_5_BUFX2_insert317 gnd vdd FILL
XFILL_0__10519_ gnd vdd FILL
XFILL_3__7864_ gnd vdd FILL
XFILL_3__11679_ gnd vdd FILL
XSFILL8520x76050 gnd vdd FILL
XFILL_5_BUFX2_insert328 gnd vdd FILL
XFILL_1__12858_ gnd vdd FILL
XBUFX2_insert18 _13443_/Y gnd _14203_/B vdd BUFX2
XFILL_5__15027_ gnd vdd FILL
XFILL_0__11499_ gnd vdd FILL
XFILL_0__14287_ gnd vdd FILL
XFILL_3__16206_ gnd vdd FILL
XFILL_3__13418_ gnd vdd FILL
XFILL_5_BUFX2_insert339 gnd vdd FILL
XFILL_5__12239_ gnd vdd FILL
X_8433_ _8433_/Q _8433_/CLK _8433_/R vdd _8433_/D gnd vdd DFFSR
XBUFX2_insert29 _13320_/Y gnd _8503_/B vdd BUFX2
XFILL_3__9603_ gnd vdd FILL
XFILL_4__15757_ gnd vdd FILL
XFILL_0__16026_ gnd vdd FILL
XFILL_2__12059_ gnd vdd FILL
XFILL_4__12969_ gnd vdd FILL
XFILL_3__14398_ gnd vdd FILL
XFILL_1__11809_ gnd vdd FILL
XFILL_0__13238_ gnd vdd FILL
XFILL_1__15577_ gnd vdd FILL
XFILL_1__12789_ gnd vdd FILL
XFILL_0_BUFX2_insert690 gnd vdd FILL
XFILL_4__14708_ gnd vdd FILL
XSFILL49000x36050 gnd vdd FILL
XFILL_3__13349_ gnd vdd FILL
X_8364_ _8424_/Q gnd _8364_/Y vdd INVX1
XFILL_3__16137_ gnd vdd FILL
XFILL_4__15688_ gnd vdd FILL
XFILL_3__9534_ gnd vdd FILL
XFILL_1__14528_ gnd vdd FILL
XFILL_0__13169_ gnd vdd FILL
XFILL_0__9756_ gnd vdd FILL
XSFILL109560x47050 gnd vdd FILL
X_7315_ _7315_/A _7366_/B _7314_/Y gnd _7315_/Y vdd OAI21X1
XFILL_4__14639_ gnd vdd FILL
XFILL_0__6968_ gnd vdd FILL
XFILL_3__16068_ gnd vdd FILL
XFILL_2__15818_ gnd vdd FILL
XFILL_3__9465_ gnd vdd FILL
X_8295_ _8233_/A _8551_/CLK _9064_/R vdd _8295_/D gnd vdd DFFSR
XFILL_1__14459_ gnd vdd FILL
XSFILL38840x79050 gnd vdd FILL
XFILL_1__7500_ gnd vdd FILL
XFILL_0__8707_ gnd vdd FILL
XFILL_5__15929_ gnd vdd FILL
XFILL_3__15019_ gnd vdd FILL
X_7246_ _7168_/A _8654_/B gnd _7247_/C vdd NAND2X1
XFILL_1__8480_ gnd vdd FILL
XSFILL54120x27050 gnd vdd FILL
XFILL_0__6899_ gnd vdd FILL
XFILL_3__9396_ gnd vdd FILL
XFILL_2__15749_ gnd vdd FILL
XFILL_0__8638_ gnd vdd FILL
XFILL_4__16309_ gnd vdd FILL
XFILL_1__7431_ gnd vdd FILL
X_7177_ _7184_/B _7177_/B gnd _7177_/Y vdd NAND2X1
XFILL_3__8347_ gnd vdd FILL
XFILL_1__16129_ gnd vdd FILL
XSFILL64440x5050 gnd vdd FILL
XFILL_6__8056_ gnd vdd FILL
XSFILL13720x1050 gnd vdd FILL
XFILL_1__7362_ gnd vdd FILL
XFILL_0__8569_ gnd vdd FILL
XFILL_4__7071_ gnd vdd FILL
XFILL_1__9101_ gnd vdd FILL
XFILL_2_BUFX2_insert229 gnd vdd FILL
XSFILL18760x46050 gnd vdd FILL
XFILL_3__7229_ gnd vdd FILL
XSFILL8600x56050 gnd vdd FILL
XFILL_1__7293_ gnd vdd FILL
XSFILL44040x79050 gnd vdd FILL
XFILL_1__9032_ gnd vdd FILL
XFILL_1_BUFX2_insert907 gnd vdd FILL
XFILL_1_BUFX2_insert918 gnd vdd FILL
X_9818_ _9818_/Q _9818_/CLK _9441_/R vdd _9818_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert929 gnd vdd FILL
XSFILL23880x37050 gnd vdd FILL
X_10700_ _10700_/A _10700_/B _10699_/Y gnd _10700_/Y vdd OAI21X1
XFILL_4__7973_ gnd vdd FILL
X_11680_ _11062_/Y _11748_/A _11366_/B _11280_/Y gnd _11680_/Y vdd OAI22X1
XSFILL108600x63050 gnd vdd FILL
X_9749_ _9813_/B _7317_/B gnd _9750_/C vdd NAND2X1
XSFILL38920x59050 gnd vdd FILL
XFILL_4__6924_ gnd vdd FILL
XFILL112440x66050 gnd vdd FILL
X_10631_ _10629_/Y _10619_/B _10631_/C gnd _10715_/D vdd OAI21X1
XBUFX2_insert228 _12432_/Y gnd _8526_/B vdd BUFX2
XFILL_1__9934_ gnd vdd FILL
XBUFX2_insert239 _15065_/Y gnd _16151_/B vdd BUFX2
XFILL_4__6855_ gnd vdd FILL
XFILL_4__9643_ gnd vdd FILL
X_13350_ _13209_/Y _13359_/A _13350_/C gnd _13351_/A vdd OAI21X1
XSFILL79160x11050 gnd vdd FILL
XSFILL39000x68050 gnd vdd FILL
X_10562_ _10548_/B _9794_/B gnd _10562_/Y vdd NAND2X1
XFILL_1__9865_ gnd vdd FILL
XFILL_5_CLKBUF1_insert118 gnd vdd FILL
XFILL_5_BUFX2_insert840 gnd vdd FILL
XFILL_5_BUFX2_insert851 gnd vdd FILL
X_12301_ _6891_/A _12301_/B _12301_/C _11885_/B gnd _12302_/C vdd AOI22X1
XFILL_5_CLKBUF1_insert129 gnd vdd FILL
XFILL_5_BUFX2_insert862 gnd vdd FILL
X_13281_ _13230_/Y _13281_/B _13294_/A gnd _13282_/B vdd OAI21X1
XFILL_5_BUFX2_insert873 gnd vdd FILL
X_10493_ _10539_/B _9597_/B gnd _10494_/C vdd NAND2X1
XFILL_5_BUFX2_insert884 gnd vdd FILL
XFILL_1__9796_ gnd vdd FILL
XFILL_4__8525_ gnd vdd FILL
XFILL_5_BUFX2_insert895 gnd vdd FILL
X_15020_ _12770_/A _12813_/Q _12812_/Q gnd _15020_/Y vdd NOR3X1
X_12232_ _12272_/A _12707_/A _12272_/C gnd _12234_/B vdd NAND3X1
XBUFX2_insert1070 _13327_/Y gnd _8916_/A vdd BUFX2
XSFILL18840x26050 gnd vdd FILL
XSFILL114600x82050 gnd vdd FILL
XBUFX2_insert1092 rst gnd BUFX2_insert600/A vdd BUFX2
XFILL_1__8747_ gnd vdd FILL
XFILL_4__8456_ gnd vdd FILL
XSFILL59720x38050 gnd vdd FILL
X_12163_ _11935_/A gnd _12165_/A vdd INVX1
XSFILL99320x24050 gnd vdd FILL
XSFILL69080x63050 gnd vdd FILL
XFILL_2__7471_ gnd vdd FILL
XFILL_5__7180_ gnd vdd FILL
XFILL_4__8387_ gnd vdd FILL
X_11114_ _12298_/Y gnd _11115_/B vdd INVX1
XFILL_2__9210_ gnd vdd FILL
XFILL_1__7629_ gnd vdd FILL
X_12094_ _12094_/A _12094_/B _12093_/Y gnd _13158_/B vdd NAND3X1
XSFILL99480x3050 gnd vdd FILL
XSFILL104280x72050 gnd vdd FILL
XFILL_4__7338_ gnd vdd FILL
X_15922_ _14478_/Y _15981_/B _15922_/C _15922_/D gnd _15923_/A vdd OAI22X1
XFILL_4__10320_ gnd vdd FILL
X_11045_ _12270_/Y _12156_/Y gnd _11045_/Y vdd XOR2X1
XFILL_2__9141_ gnd vdd FILL
XSFILL88920x4050 gnd vdd FILL
XFILL_1__10140_ gnd vdd FILL
XFILL_0__10870_ gnd vdd FILL
XFILL_5__11610_ gnd vdd FILL
XSFILL23800x81050 gnd vdd FILL
XFILL_4__10251_ gnd vdd FILL
X_15853_ _15652_/A _9578_/Q _9650_/A _15652_/D gnd _15856_/B vdd AOI22X1
XFILL_5__12590_ gnd vdd FILL
XFILL_4__9008_ gnd vdd FILL
XFILL_2__11430_ gnd vdd FILL
XSFILL89240x76050 gnd vdd FILL
XFILL_3__10981_ gnd vdd FILL
XFILL_2_BUFX2_insert730 gnd vdd FILL
XFILL_2_BUFX2_insert741 gnd vdd FILL
X_14804_ _9034_/A gnd _14804_/Y vdd INVX1
XFILL_2_BUFX2_insert752 gnd vdd FILL
XFILL_3__12720_ gnd vdd FILL
XFILL_2_BUFX2_insert763 gnd vdd FILL
XFILL_5__11541_ gnd vdd FILL
X_12996_ _6885_/A gnd _12996_/Y vdd INVX1
XFILL_4__10182_ gnd vdd FILL
X_15784_ _15784_/A _15784_/B gnd _15785_/C vdd NOR2X1
XSFILL13880x7050 gnd vdd FILL
XFILL_2_BUFX2_insert774 gnd vdd FILL
XSFILL3720x79050 gnd vdd FILL
XFILL_2__11361_ gnd vdd FILL
XFILL_2_BUFX2_insert785 gnd vdd FILL
XFILL_6__12831_ gnd vdd FILL
XFILL_2_BUFX2_insert796 gnd vdd FILL
XFILL_5__14260_ gnd vdd FILL
XFILL_2__13100_ gnd vdd FILL
X_14735_ _7236_/A gnd _14735_/Y vdd INVX1
X_11947_ _11947_/A gnd _11949_/A vdd INVX1
XFILL_3__12651_ gnd vdd FILL
XFILL_2__10312_ gnd vdd FILL
XFILL_5__11472_ gnd vdd FILL
XFILL_1__13830_ gnd vdd FILL
XFILL_4__14990_ gnd vdd FILL
XFILL_2__14080_ gnd vdd FILL
XSFILL94360x67050 gnd vdd FILL
XFILL_0__12471_ gnd vdd FILL
XFILL_2__11292_ gnd vdd FILL
XFILL_5__13211_ gnd vdd FILL
XFILL_5__9752_ gnd vdd FILL
XFILL_5__10423_ gnd vdd FILL
XFILL_3__11602_ gnd vdd FILL
XFILL_5__6964_ gnd vdd FILL
X_14666_ _14665_/Y _14666_/B gnd _14666_/Y vdd NOR2X1
X_11878_ _12809_/Q gnd _11880_/A vdd INVX1
XFILL_3__15370_ gnd vdd FILL
XFILL_5__14191_ gnd vdd FILL
XFILL_2__13031_ gnd vdd FILL
XFILL_4__13941_ gnd vdd FILL
XFILL_0__14210_ gnd vdd FILL
XFILL_3__12582_ gnd vdd FILL
XFILL_2__10243_ gnd vdd FILL
XFILL_0__11422_ gnd vdd FILL
XFILL_5__8703_ gnd vdd FILL
XFILL_2__9974_ gnd vdd FILL
XFILL_1__13761_ gnd vdd FILL
XFILL_1__10973_ gnd vdd FILL
X_13617_ _13843_/C _13616_/Y _13615_/Y _13617_/D gnd _13618_/A vdd OAI22X1
XFILL_0__15190_ gnd vdd FILL
X_16405_ _14816_/A gnd _16407_/A vdd INVX1
XSFILL69160x43050 gnd vdd FILL
X_10829_ _10867_/Q gnd _10831_/A vdd INVX1
XFILL_5__13142_ gnd vdd FILL
XFILL_5__9683_ gnd vdd FILL
XFILL_3__14321_ gnd vdd FILL
XFILL_5__6895_ gnd vdd FILL
X_14597_ _14597_/A _14570_/Y _14597_/C gnd _13021_/B vdd AOI21X1
XFILL_1__15500_ gnd vdd FILL
XFILL_3__11533_ gnd vdd FILL
XFILL_4__13872_ gnd vdd FILL
XFILL_1__12712_ gnd vdd FILL
XFILL_2__10174_ gnd vdd FILL
XFILL_0__14141_ gnd vdd FILL
XBUFX2_insert740 _12402_/Y gnd _9008_/B vdd BUFX2
XFILL_0__11353_ gnd vdd FILL
XBUFX2_insert751 _13344_/Y gnd _9789_/B vdd BUFX2
XFILL_5__8634_ gnd vdd FILL
XFILL_1__13692_ gnd vdd FILL
XFILL_0__7940_ gnd vdd FILL
XFILL_4__15611_ gnd vdd FILL
X_13548_ _16419_/Q gnd _15145_/B vdd INVX1
X_16336_ _15275_/A gnd _16336_/Y vdd INVX1
XFILL_3__14252_ gnd vdd FILL
XSFILL104360x52050 gnd vdd FILL
XFILL_4__12823_ gnd vdd FILL
XBUFX2_insert762 _13412_/Y gnd _14051_/C vdd BUFX2
XFILL_5__10285_ gnd vdd FILL
XBUFX2_insert773 _13301_/Y gnd _7872_/B vdd BUFX2
XFILL_0__10304_ gnd vdd FILL
XFILL_1__15431_ gnd vdd FILL
XFILL_3__11464_ gnd vdd FILL
XFILL_1__12643_ gnd vdd FILL
XFILL_2__8856_ gnd vdd FILL
XFILL_2__14982_ gnd vdd FILL
XFILL_0__14072_ gnd vdd FILL
XSFILL88440x28050 gnd vdd FILL
XBUFX2_insert784 _10911_/Y gnd _12122_/A vdd BUFX2
XBUFX2_insert795 _13334_/Y gnd _9356_/A vdd BUFX2
XFILL_0__11284_ gnd vdd FILL
XFILL_5__12024_ gnd vdd FILL
XSFILL74280x34050 gnd vdd FILL
X_16267_ _16260_/Y _16267_/B _16267_/C gnd _16282_/A vdd NAND3X1
XFILL_0__7871_ gnd vdd FILL
XFILL_4__15542_ gnd vdd FILL
XFILL_3__10415_ gnd vdd FILL
X_13479_ _13479_/A _13868_/B _13479_/C _13479_/D gnd _13483_/B vdd OAI22X1
XFILL_2__7807_ gnd vdd FILL
XFILL_4__12754_ gnd vdd FILL
XFILL_3__14183_ gnd vdd FILL
XFILL_0__13023_ gnd vdd FILL
XFILL_2__13933_ gnd vdd FILL
XFILL_1__15362_ gnd vdd FILL
XFILL_3__7580_ gnd vdd FILL
XFILL_3__11395_ gnd vdd FILL
XFILL_0__10235_ gnd vdd FILL
XFILL_2__8787_ gnd vdd FILL
XFILL_0__9610_ gnd vdd FILL
XFILL_1__12574_ gnd vdd FILL
X_15218_ _9306_/Q _15892_/B _15380_/C _9946_/Q gnd _15218_/Y vdd AOI22X1
XFILL_5__8496_ gnd vdd FILL
X_16198_ _9162_/A gnd _16198_/Y vdd INVX1
XSFILL89320x56050 gnd vdd FILL
XFILL_3__13134_ gnd vdd FILL
XFILL_4__11705_ gnd vdd FILL
XSFILL49080x10050 gnd vdd FILL
XFILL_2__7738_ gnd vdd FILL
XFILL_1__14313_ gnd vdd FILL
XFILL_4__15473_ gnd vdd FILL
XFILL_2__13864_ gnd vdd FILL
XFILL_1__11525_ gnd vdd FILL
XFILL_0__10166_ gnd vdd FILL
XFILL_5__7447_ gnd vdd FILL
XFILL_1__15293_ gnd vdd FILL
X_7100_ _7100_/A _7868_/B gnd _7101_/C vdd NAND2X1
XFILL_0__9541_ gnd vdd FILL
X_15149_ _15149_/A _15792_/B _15761_/D _15149_/D gnd _15149_/Y vdd OAI22X1
X_8080_ _8078_/Y _8079_/A _8080_/C gnd _8158_/D vdd OAI21X1
XFILL_4__14424_ gnd vdd FILL
XFILL_3__9250_ gnd vdd FILL
XFILL_4__11636_ gnd vdd FILL
XFILL_2__15603_ gnd vdd FILL
XFILL_5__13975_ gnd vdd FILL
XFILL_3__10277_ gnd vdd FILL
XFILL_1__14244_ gnd vdd FILL
XFILL_2__13795_ gnd vdd FILL
XFILL_1__11456_ gnd vdd FILL
XFILL_5__15714_ gnd vdd FILL
X_7031_ _8823_/A _7068_/B gnd _7032_/C vdd NAND2X1
XFILL_0__14974_ gnd vdd FILL
XFILL_5__7378_ gnd vdd FILL
XFILL_0__9472_ gnd vdd FILL
XFILL_3__12016_ gnd vdd FILL
XFILL_3__8201_ gnd vdd FILL
XFILL_2__9408_ gnd vdd FILL
XSFILL94440x47050 gnd vdd FILL
XFILL_2__15534_ gnd vdd FILL
XFILL_4__14355_ gnd vdd FILL
XFILL_6__10388_ gnd vdd FILL
XFILL_4__11567_ gnd vdd FILL
XFILL_1__10407_ gnd vdd FILL
XFILL_2__12746_ gnd vdd FILL
XFILL_1__14175_ gnd vdd FILL
XFILL_5__9117_ gnd vdd FILL
XFILL_0__13925_ gnd vdd FILL
XFILL_1__11387_ gnd vdd FILL
XFILL_4__13306_ gnd vdd FILL
XFILL_5__15645_ gnd vdd FILL
XFILL_4__10518_ gnd vdd FILL
XFILL_5__12857_ gnd vdd FILL
XFILL_3__8132_ gnd vdd FILL
XFILL_2__9339_ gnd vdd FILL
XFILL_1__13126_ gnd vdd FILL
XFILL_4__11498_ gnd vdd FILL
XFILL_2__15465_ gnd vdd FILL
XFILL_4__14286_ gnd vdd FILL
XFILL_0__13856_ gnd vdd FILL
XFILL_4__16025_ gnd vdd FILL
XFILL_0__8354_ gnd vdd FILL
XFILL_5__11808_ gnd vdd FILL
XFILL_4__13237_ gnd vdd FILL
XFILL_4__10449_ gnd vdd FILL
XFILL_5__15576_ gnd vdd FILL
XFILL_2__14416_ gnd vdd FILL
XFILL_5__12788_ gnd vdd FILL
XFILL_3__8063_ gnd vdd FILL
X_8982_ _8982_/A _9011_/A _8981_/Y gnd _8982_/Y vdd OAI21X1
XFILL_2__11628_ gnd vdd FILL
XFILL_2__15396_ gnd vdd FILL
XFILL_1__10269_ gnd vdd FILL
XFILL_3__13967_ gnd vdd FILL
XFILL_0__7305_ gnd vdd FILL
XSFILL104440x32050 gnd vdd FILL
XFILL_0__13787_ gnd vdd FILL
XFILL_5__14527_ gnd vdd FILL
XFILL_4__13168_ gnd vdd FILL
XFILL_3__15706_ gnd vdd FILL
X_7933_ _7931_/B _9597_/B gnd _7933_/Y vdd NAND2X1
XFILL_5__11739_ gnd vdd FILL
XFILL_0__10999_ gnd vdd FILL
XFILL_1__12008_ gnd vdd FILL
XFILL_2__14347_ gnd vdd FILL
XFILL_3__12918_ gnd vdd FILL
XSFILL8680x30050 gnd vdd FILL
XFILL_0__15526_ gnd vdd FILL
XFILL_2__11559_ gnd vdd FILL
XFILL_0__12738_ gnd vdd FILL
XSFILL98680x52050 gnd vdd FILL
XFILL_3__13898_ gnd vdd FILL
XFILL_0__7236_ gnd vdd FILL
XFILL_6__9792_ gnd vdd FILL
XFILL_5__14458_ gnd vdd FILL
XFILL_4__12119_ gnd vdd FILL
XFILL_3__15637_ gnd vdd FILL
XFILL_4__13099_ gnd vdd FILL
X_7864_ _7916_/Q gnd _7866_/A vdd INVX1
XFILL_3__12849_ gnd vdd FILL
XFILL_2__14278_ gnd vdd FILL
XSFILL59160x75050 gnd vdd FILL
XFILL_0__15457_ gnd vdd FILL
X_9603_ _9613_/B _9475_/B gnd _9603_/Y vdd NAND2X1
XFILL_6__8743_ gnd vdd FILL
XFILL_5__13409_ gnd vdd FILL
XFILL_0__7167_ gnd vdd FILL
XFILL_2__16017_ gnd vdd FILL
XSFILL99560x80050 gnd vdd FILL
XFILL_2__13229_ gnd vdd FILL
XFILL_5__14389_ gnd vdd FILL
X_7795_ _7757_/A _8051_/CLK _8038_/R vdd _7759_/Y gnd vdd DFFSR
XFILL_3__15568_ gnd vdd FILL
XFILL_0__14408_ gnd vdd FILL
XFILL_3__8965_ gnd vdd FILL
XFILL_1__13959_ gnd vdd FILL
XFILL_0__15388_ gnd vdd FILL
XFILL_5__16128_ gnd vdd FILL
XFILL_6__15679_ gnd vdd FILL
X_9534_ _9534_/A gnd _9534_/Y vdd INVX1
XFILL_3__14519_ gnd vdd FILL
XFILL_0__7098_ gnd vdd FILL
XFILL_1__7980_ gnd vdd FILL
XFILL_5_BUFX2_insert103 gnd vdd FILL
XFILL_3__15499_ gnd vdd FILL
XFILL_0__14339_ gnd vdd FILL
XFILL_3__8896_ gnd vdd FILL
XSFILL13640x31050 gnd vdd FILL
XFILL_4__15809_ gnd vdd FILL
XFILL_1__6931_ gnd vdd FILL
XFILL_5__16059_ gnd vdd FILL
X_9465_ _9465_/A gnd _9467_/A vdd INVX1
XFILL_1__15629_ gnd vdd FILL
XFILL_3__7847_ gnd vdd FILL
XSFILL78840x81050 gnd vdd FILL
X_8416_ _8340_/A _9568_/CLK _7648_/R vdd _8342_/Y gnd vdd DFFSR
XFILL_1__9650_ gnd vdd FILL
XFILL_1__6862_ gnd vdd FILL
XFILL_0__16009_ gnd vdd FILL
X_9396_ _9394_/Y _9401_/A _9395_/Y gnd _9450_/D vdd OAI21X1
XFILL_4_BUFX2_insert803 gnd vdd FILL
XFILL_4_BUFX2_insert814 gnd vdd FILL
XFILL_1__8601_ gnd vdd FILL
XFILL_4_BUFX2_insert825 gnd vdd FILL
XFILL_6__7487_ gnd vdd FILL
XFILL_0__9808_ gnd vdd FILL
XFILL_4__8310_ gnd vdd FILL
X_8347_ _8356_/A _7451_/B gnd _8348_/C vdd NAND2X1
XFILL_4_BUFX2_insert836 gnd vdd FILL
XFILL_3__9517_ gnd vdd FILL
XSFILL104520x12050 gnd vdd FILL
XFILL_4__9290_ gnd vdd FILL
XFILL_4_BUFX2_insert847 gnd vdd FILL
XFILL_4_BUFX2_insert858 gnd vdd FILL
XSFILL83960x72050 gnd vdd FILL
XFILL_1__8532_ gnd vdd FILL
XFILL_4_BUFX2_insert869 gnd vdd FILL
XSFILL8760x10050 gnd vdd FILL
XFILL_0__9739_ gnd vdd FILL
X_8278_ _8278_/Q _8818_/CLK _8278_/R vdd _8278_/D gnd vdd DFFSR
XFILL_4__8241_ gnd vdd FILL
XSFILL99240x39050 gnd vdd FILL
XFILL_1__8463_ gnd vdd FILL
X_7229_ _7227_/Y _7168_/A _7229_/C gnd _7229_/Y vdd OAI21X1
XFILL_3__9379_ gnd vdd FILL
XFILL_6__8108_ gnd vdd FILL
XFILL_1__7414_ gnd vdd FILL
XFILL_1__8394_ gnd vdd FILL
XFILL_4__7123_ gnd vdd FILL
XFILL_1__7345_ gnd vdd FILL
XSFILL13720x11050 gnd vdd FILL
XFILL_4__7054_ gnd vdd FILL
XFILL112360x6050 gnd vdd FILL
X_12850_ _12928_/Q gnd _12850_/Y vdd INVX1
XFILL112040x63050 gnd vdd FILL
XFILL_5_BUFX2_insert3 gnd vdd FILL
XSFILL79400x68050 gnd vdd FILL
X_11801_ _11249_/Y _11801_/B gnd _11802_/C vdd NAND2X1
XFILL_1__9015_ gnd vdd FILL
XFILL_1_BUFX2_insert704 gnd vdd FILL
X_12781_ _12779_/Y _12777_/A _12781_/C gnd _12819_/D vdd OAI21X1
XFILL_1_BUFX2_insert715 gnd vdd FILL
XFILL_1_BUFX2_insert726 gnd vdd FILL
XSFILL69240x1050 gnd vdd FILL
X_14520_ _8120_/A gnd _14520_/Y vdd INVX1
XFILL_1_BUFX2_insert737 gnd vdd FILL
XSFILL79000x70050 gnd vdd FILL
XFILL_1_BUFX2_insert748 gnd vdd FILL
XSFILL113640x8050 gnd vdd FILL
X_11732_ _11732_/A _11732_/B gnd _11733_/C vdd NAND2X1
XFILL_1_BUFX2_insert759 gnd vdd FILL
X_14451_ _8683_/Q gnd _14451_/Y vdd INVX1
XFILL_4__7956_ gnd vdd FILL
X_11663_ _11684_/B _11067_/Y _11663_/C gnd _11664_/B vdd OAI21X1
XFILL_2__6971_ gnd vdd FILL
X_13402_ _9942_/Q gnd _13402_/Y vdd INVX1
XFILL_4__6907_ gnd vdd FILL
X_10614_ _15002_/C gnd _10616_/A vdd INVX1
XFILL_4_BUFX2_insert19 gnd vdd FILL
XFILL_4__7887_ gnd vdd FILL
X_14382_ _8041_/Q gnd _15841_/D vdd INVX1
XFILL_1__9917_ gnd vdd FILL
XFILL_2__8710_ gnd vdd FILL
X_11594_ _11593_/Y _11304_/Y _11582_/C gnd _11595_/C vdd OAI21X1
X_16121_ _16121_/A _16121_/B gnd _16122_/B vdd NOR2X1
XFILL_4__9626_ gnd vdd FILL
X_13333_ _13259_/C _13332_/Y gnd _13333_/Y vdd NOR2X1
XFILL_4__6838_ gnd vdd FILL
X_10545_ _10545_/A _10500_/B _10544_/Y gnd _10545_/Y vdd OAI21X1
XFILL_2__8641_ gnd vdd FILL
XFILL_5_BUFX2_insert670 gnd vdd FILL
XFILL_1__9848_ gnd vdd FILL
XSFILL23560x14050 gnd vdd FILL
XFILL_5_BUFX2_insert681 gnd vdd FILL
XFILL_5__8350_ gnd vdd FILL
XFILL_4__9557_ gnd vdd FILL
X_16052_ _16051_/Y _15848_/A gnd _16052_/Y vdd NOR2X1
XFILL_5_BUFX2_insert692 gnd vdd FILL
X_13264_ _13297_/A _13263_/Y gnd _13265_/B vdd OR2X2
XSFILL23800x76050 gnd vdd FILL
X_10476_ _15931_/A _7916_/CLK _9580_/R vdd _10476_/D gnd vdd DFFSR
XFILL_2__10930_ gnd vdd FILL
XFILL_0__10020_ gnd vdd FILL
XFILL_2__8572_ gnd vdd FILL
XFILL_3__11180_ gnd vdd FILL
XFILL_5__7301_ gnd vdd FILL
XFILL_4__8508_ gnd vdd FILL
X_15003_ _14986_/A _16035_/B _15024_/C gnd _15003_/Y vdd NAND3X1
XFILL_1__9779_ gnd vdd FILL
X_12215_ _12239_/A _12248_/A gnd _12215_/Y vdd NOR2X1
XFILL_4__9488_ gnd vdd FILL
X_13195_ _11947_/A _13201_/CLK _13201_/R vdd _13195_/D gnd vdd DFFSR
XFILL_4__12470_ gnd vdd FILL
XFILL_3__10131_ gnd vdd FILL
XFILL_1__11310_ gnd vdd FILL
XFILL_5__7232_ gnd vdd FILL
XFILL_4__8439_ gnd vdd FILL
XFILL_1__12290_ gnd vdd FILL
XSFILL29000x4050 gnd vdd FILL
X_12146_ _12122_/A _12929_/Q gnd _12146_/Y vdd NAND2X1
XFILL_4__11421_ gnd vdd FILL
XFILL_2__12600_ gnd vdd FILL
XFILL_5__13760_ gnd vdd FILL
XFILL_3__10062_ gnd vdd FILL
XFILL_5__10972_ gnd vdd FILL
XFILL_2__7454_ gnd vdd FILL
XFILL_2__13580_ gnd vdd FILL
XFILL_1__11241_ gnd vdd FILL
XFILL_2__10792_ gnd vdd FILL
XSFILL43720x27050 gnd vdd FILL
XFILL_5__7163_ gnd vdd FILL
XFILL_5__12711_ gnd vdd FILL
XFILL_0__11971_ gnd vdd FILL
X_12077_ _12077_/A _12073_/B _12073_/C gnd gnd _12077_/Y vdd AOI22X1
XFILL_4__14140_ gnd vdd FILL
XFILL_4__11352_ gnd vdd FILL
XSFILL53880x71050 gnd vdd FILL
XFILL_2__12531_ gnd vdd FILL
XFILL_5__13691_ gnd vdd FILL
XFILL_3__14870_ gnd vdd FILL
XFILL_0__13710_ gnd vdd FILL
XFILL_1__11172_ gnd vdd FILL
XFILL_0__10922_ gnd vdd FILL
XFILL_4__10303_ gnd vdd FILL
XFILL_5__7094_ gnd vdd FILL
X_15905_ _15351_/A _14485_/Y _14488_/Y _15351_/D gnd _15905_/Y vdd OAI22X1
XSFILL69160x38050 gnd vdd FILL
XFILL_5__15430_ gnd vdd FILL
XFILL_0__14690_ gnd vdd FILL
X_11028_ _11006_/Y _11016_/Y _11028_/C gnd _11028_/Y vdd AOI21X1
XFILL_2__9124_ gnd vdd FILL
XFILL_5__12642_ gnd vdd FILL
XFILL_4__14071_ gnd vdd FILL
XFILL_3__13821_ gnd vdd FILL
XFILL_1__10123_ gnd vdd FILL
XFILL_2__15250_ gnd vdd FILL
XSFILL3640x3050 gnd vdd FILL
XFILL_4__11283_ gnd vdd FILL
XFILL_2__12462_ gnd vdd FILL
XFILL_1__15980_ gnd vdd FILL
XFILL_0__13641_ gnd vdd FILL
XFILL_4__13022_ gnd vdd FILL
XSFILL84200x41050 gnd vdd FILL
XFILL_2__14201_ gnd vdd FILL
XFILL_5__15361_ gnd vdd FILL
X_15836_ _15836_/A _15595_/B _15836_/C gnd _15839_/A vdd OAI21X1
XFILL_0_BUFX2_insert1006 gnd vdd FILL
XFILL_4__10234_ gnd vdd FILL
XFILL_5__12573_ gnd vdd FILL
XSFILL104360x47050 gnd vdd FILL
XFILL_0_BUFX2_insert1017 gnd vdd FILL
XFILL_2__11413_ gnd vdd FILL
XFILL_3__10964_ gnd vdd FILL
XFILL_2__15181_ gnd vdd FILL
XFILL_3__13752_ gnd vdd FILL
XFILL_0_BUFX2_insert1028 gnd vdd FILL
XFILL_1__10054_ gnd vdd FILL
XFILL_1__14931_ gnd vdd FILL
XFILL_2_BUFX2_insert560 gnd vdd FILL
XFILL_0_BUFX2_insert1039 gnd vdd FILL
XFILL_2__12393_ gnd vdd FILL
XFILL_2_BUFX2_insert571 gnd vdd FILL
XFILL_0__16360_ gnd vdd FILL
XFILL_2_BUFX2_insert582 gnd vdd FILL
XFILL_0__10784_ gnd vdd FILL
XFILL_0__13572_ gnd vdd FILL
XFILL_5__14312_ gnd vdd FILL
XFILL_6__13863_ gnd vdd FILL
XFILL_2_BUFX2_insert593 gnd vdd FILL
XFILL_2__8006_ gnd vdd FILL
XSFILL74280x29050 gnd vdd FILL
XFILL_5__11524_ gnd vdd FILL
XFILL_0__8070_ gnd vdd FILL
XFILL_4__10165_ gnd vdd FILL
XFILL_3__12703_ gnd vdd FILL
XFILL_2__14132_ gnd vdd FILL
X_15767_ _15765_/Y _15767_/B gnd _15767_/Y vdd NOR2X1
XFILL_5__15292_ gnd vdd FILL
X_12979_ vdd _12979_/B gnd _12980_/C vdd NAND2X1
XFILL_0__15311_ gnd vdd FILL
XFILL_3__13683_ gnd vdd FILL
XFILL_2__11344_ gnd vdd FILL
XFILL_6_BUFX2_insert909 gnd vdd FILL
XFILL_1__14862_ gnd vdd FILL
XFILL_0__12523_ gnd vdd FILL
XFILL_5__9804_ gnd vdd FILL
XFILL_3__10895_ gnd vdd FILL
XFILL_0__16291_ gnd vdd FILL
XFILL_5__14243_ gnd vdd FILL
X_14718_ _14718_/A _14718_/B _14718_/C _14718_/D gnd _14722_/B vdd OAI22X1
XFILL_3__12634_ gnd vdd FILL
XFILL_5__7996_ gnd vdd FILL
XFILL_5__11455_ gnd vdd FILL
XFILL_3__15422_ gnd vdd FILL
XFILL_1__13813_ gnd vdd FILL
X_15698_ _10406_/A gnd _15698_/Y vdd INVX1
XFILL_2__14063_ gnd vdd FILL
XFILL_4__14973_ gnd vdd FILL
XFILL_0__15242_ gnd vdd FILL
XFILL_2__11275_ gnd vdd FILL
XFILL_1__14793_ gnd vdd FILL
XFILL_0__12454_ gnd vdd FILL
XFILL_5__9735_ gnd vdd FILL
XFILL_5__10406_ gnd vdd FILL
XFILL_5__6947_ gnd vdd FILL
XFILL_2__13014_ gnd vdd FILL
XFILL_5__14174_ gnd vdd FILL
X_14649_ _7105_/A gnd _14650_/D vdd INVX1
XFILL_4__13924_ gnd vdd FILL
XFILL_3__15353_ gnd vdd FILL
X_7580_ _7578_/Y _7562_/B _7579_/Y gnd _7650_/D vdd OAI21X1
XFILL_5__11386_ gnd vdd FILL
XFILL_1__13744_ gnd vdd FILL
XFILL_3__8750_ gnd vdd FILL
XFILL_0__11405_ gnd vdd FILL
XFILL_1__10956_ gnd vdd FILL
XFILL_0__12385_ gnd vdd FILL
XFILL_0__15173_ gnd vdd FILL
XFILL_5__13125_ gnd vdd FILL
XFILL_5__9666_ gnd vdd FILL
XFILL_0__8972_ gnd vdd FILL
XFILL_3__11516_ gnd vdd FILL
XFILL_3__14304_ gnd vdd FILL
XFILL_5__6878_ gnd vdd FILL
XFILL_4__13855_ gnd vdd FILL
XFILL_2__8908_ gnd vdd FILL
XFILL_3__7701_ gnd vdd FILL
XSFILL18680x3050 gnd vdd FILL
XFILL_3__15284_ gnd vdd FILL
XBUFX2_insert570 BUFX2_insert570/A gnd _12809_/R vdd BUFX2
XFILL_0__14124_ gnd vdd FILL
XFILL_3__12496_ gnd vdd FILL
XFILL_2__10157_ gnd vdd FILL
XFILL_0__11336_ gnd vdd FILL
XFILL_5__8617_ gnd vdd FILL
XFILL_1__13675_ gnd vdd FILL
XFILL_2__9888_ gnd vdd FILL
XBUFX2_insert581 BUFX2_insert559/A gnd _9561_/R vdd BUFX2
XSFILL93400x78050 gnd vdd FILL
XSFILL53960x51050 gnd vdd FILL
XFILL_1__10887_ gnd vdd FILL
X_16319_ _16308_/Y _16297_/Y _16318_/Y gnd _16319_/Y vdd NOR3X1
XBUFX2_insert592 BUFX2_insert559/A gnd _8542_/R vdd BUFX2
X_9250_ _9250_/A _9228_/A _9249_/Y gnd _9316_/D vdd OAI21X1
XFILL_3__14235_ gnd vdd FILL
XFILL_5__9597_ gnd vdd FILL
XSFILL109480x80050 gnd vdd FILL
XFILL_1__15414_ gnd vdd FILL
XFILL_5__10268_ gnd vdd FILL
XFILL_3__11447_ gnd vdd FILL
XFILL_3__7632_ gnd vdd FILL
XFILL_1__12626_ gnd vdd FILL
XFILL_4__13786_ gnd vdd FILL
XFILL_2__8839_ gnd vdd FILL
XSFILL69240x18050 gnd vdd FILL
XFILL_0__14055_ gnd vdd FILL
XFILL_2__14965_ gnd vdd FILL
XFILL_0__11267_ gnd vdd FILL
XFILL_1__16394_ gnd vdd FILL
XFILL_4__10998_ gnd vdd FILL
X_8201_ _8232_/B _9353_/B gnd _8202_/C vdd NAND2X1
XFILL_5__12007_ gnd vdd FILL
XFILL_4__15525_ gnd vdd FILL
XFILL_0__7854_ gnd vdd FILL
XFILL_6__11558_ gnd vdd FILL
X_9181_ _9099_/A _8051_/CLK _8051_/R vdd _9101_/Y gnd vdd DFFSR
XFILL_4__12737_ gnd vdd FILL
XFILL_3__14166_ gnd vdd FILL
XFILL_3__7563_ gnd vdd FILL
XFILL_1__15345_ gnd vdd FILL
XFILL_0__13006_ gnd vdd FILL
XFILL_2__13916_ gnd vdd FILL
XFILL_3__11378_ gnd vdd FILL
XFILL_2__14896_ gnd vdd FILL
XFILL_0__11198_ gnd vdd FILL
XFILL_3__13117_ gnd vdd FILL
X_8132_ _8132_/A gnd _8134_/A vdd INVX1
XFILL_5__8479_ gnd vdd FILL
XFILL_4__15456_ gnd vdd FILL
XFILL_2__13847_ gnd vdd FILL
XFILL_1__11508_ gnd vdd FILL
XFILL_3__14097_ gnd vdd FILL
XSFILL8680x25050 gnd vdd FILL
XFILL_0__10149_ gnd vdd FILL
XFILL_3__7494_ gnd vdd FILL
XFILL_1__15276_ gnd vdd FILL
XFILL_1__12488_ gnd vdd FILL
XFILL_0__9524_ gnd vdd FILL
XFILL_4__14407_ gnd vdd FILL
X_8063_ _8153_/Q gnd _8065_/A vdd INVX1
XFILL_5__13958_ gnd vdd FILL
XFILL_3__9233_ gnd vdd FILL
XFILL_4__11619_ gnd vdd FILL
XFILL_4__15387_ gnd vdd FILL
XFILL_1__14227_ gnd vdd FILL
XFILL_2__13778_ gnd vdd FILL
XFILL_4__12599_ gnd vdd FILL
XFILL_1__11439_ gnd vdd FILL
XFILL_0__14957_ gnd vdd FILL
X_7014_ _7014_/Q _8947_/CLK _9069_/R vdd _7014_/D gnd vdd DFFSR
XFILL_5__12909_ gnd vdd FILL
XFILL_4__14338_ gnd vdd FILL
XFILL_2__12729_ gnd vdd FILL
XFILL_3__9164_ gnd vdd FILL
XFILL_2__15517_ gnd vdd FILL
XFILL_5__13889_ gnd vdd FILL
XFILL_1__14158_ gnd vdd FILL
XFILL_0__13908_ gnd vdd FILL
XSFILL74200x73050 gnd vdd FILL
XFILL111880x69050 gnd vdd FILL
XFILL_5__15628_ gnd vdd FILL
XFILL_0__14888_ gnd vdd FILL
XSFILL89800x52050 gnd vdd FILL
XFILL_0__9386_ gnd vdd FILL
XFILL_3__8115_ gnd vdd FILL
XFILL_1__13109_ gnd vdd FILL
XFILL_4__14269_ gnd vdd FILL
XFILL_3__9095_ gnd vdd FILL
XFILL_2__15448_ gnd vdd FILL
XFILL_0__13839_ gnd vdd FILL
XSFILL109960x58050 gnd vdd FILL
XFILL_3__14999_ gnd vdd FILL
XFILL_1__14089_ gnd vdd FILL
XFILL_4__16008_ gnd vdd FILL
XFILL_0__8337_ gnd vdd FILL
XSFILL13640x26050 gnd vdd FILL
XFILL_5__15559_ gnd vdd FILL
X_8965_ _9051_/Q gnd _8965_/Y vdd INVX1
XFILL_2__15379_ gnd vdd FILL
XSFILL109560x60050 gnd vdd FILL
XFILL_0__8268_ gnd vdd FILL
X_7916_ _7916_/Q _7916_/CLK _7276_/R vdd _7866_/Y gnd vdd DFFSR
XFILL_1__7061_ gnd vdd FILL
X_8896_ _8894_/Y _8896_/B _8895_/Y gnd _8942_/D vdd OAI21X1
XFILL_0__15509_ gnd vdd FILL
XFILL_0__7219_ gnd vdd FILL
XSFILL54120x40050 gnd vdd FILL
X_7847_ _7872_/B _7847_/B gnd _7847_/Y vdd NAND2X1
XFILL_0__8199_ gnd vdd FILL
XFILL_4__7810_ gnd vdd FILL
XSFILL33800x5050 gnd vdd FILL
XFILL_0_CLKBUF1_insert115 gnd vdd FILL
XFILL_3__9997_ gnd vdd FILL
XFILL_0_CLKBUF1_insert126 gnd vdd FILL
XFILL_0_CLKBUF1_insert137 gnd vdd FILL
X_7778_ _7706_/A _7778_/CLK _8418_/R vdd _7778_/D gnd vdd DFFSR
XFILL_0_CLKBUF1_insert148 gnd vdd FILL
XFILL_4__7741_ gnd vdd FILL
XFILL_0_CLKBUF1_insert159 gnd vdd FILL
XSFILL43960x83050 gnd vdd FILL
X_9517_ _9535_/A _9517_/B gnd _9518_/C vdd NAND2X1
XSFILL58760x43050 gnd vdd FILL
XFILL_1__7963_ gnd vdd FILL
XFILL_4__7672_ gnd vdd FILL
XFILL_3__8879_ gnd vdd FILL
XFILL_1__6914_ gnd vdd FILL
XSFILL19240x66050 gnd vdd FILL
X_9448_ _9448_/Q _7010_/CLK _7413_/R vdd _9390_/Y gnd vdd DFFSR
XFILL_4__9411_ gnd vdd FILL
XFILL111960x49050 gnd vdd FILL
X_10330_ _13679_/A _9188_/CLK _9306_/R vdd _10244_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert600 gnd vdd FILL
XSFILL23480x29050 gnd vdd FILL
XFILL_1__6845_ gnd vdd FILL
XFILL_1__9633_ gnd vdd FILL
XFILL_4_BUFX2_insert611 gnd vdd FILL
X_9379_ _9379_/A gnd _9381_/A vdd INVX1
XFILL_4_BUFX2_insert622 gnd vdd FILL
XFILL_4_BUFX2_insert633 gnd vdd FILL
XFILL_4__9342_ gnd vdd FILL
XFILL_4_BUFX2_insert644 gnd vdd FILL
X_10261_ _10271_/B _6933_/B gnd _10261_/Y vdd NAND2X1
XFILL112040x58050 gnd vdd FILL
XFILL_4_BUFX2_insert655 gnd vdd FILL
XFILL_4_BUFX2_insert666 gnd vdd FILL
X_12000_ _12084_/A _12792_/Q _12084_/C gnd _12000_/Y vdd NAND3X1
XFILL_4__9273_ gnd vdd FILL
XFILL_4_BUFX2_insert677 gnd vdd FILL
XFILL_4_BUFX2_insert688 gnd vdd FILL
XFILL_6__9209_ gnd vdd FILL
XSFILL64760x62050 gnd vdd FILL
XFILL_1__8515_ gnd vdd FILL
XFILL_4_BUFX2_insert699 gnd vdd FILL
X_10192_ _10192_/A gnd _10194_/A vdd INVX1
XSFILL38920x72050 gnd vdd FILL
XFILL_1__9495_ gnd vdd FILL
XFILL_4__8224_ gnd vdd FILL
XSFILL54200x20050 gnd vdd FILL
XFILL_1__8446_ gnd vdd FILL
X_13951_ _9440_/Q _13883_/B _14214_/C _15475_/A gnd _13952_/B vdd AOI22X1
XFILL_1__8377_ gnd vdd FILL
XFILL_2__7170_ gnd vdd FILL
XFILL_4__7106_ gnd vdd FILL
XFILL_4__8086_ gnd vdd FILL
X_12902_ vdd _12902_/B gnd _12903_/C vdd NAND2X1
X_13882_ _13881_/Y _13882_/B gnd _13883_/C vdd NOR2X1
XFILL_1__7328_ gnd vdd FILL
XFILL_4__7037_ gnd vdd FILL
X_12833_ vdd _12833_/B gnd _12834_/C vdd NAND2X1
X_15621_ _14146_/B gnd _15621_/Y vdd INVX1
XFILL_1_BUFX2_insert501 gnd vdd FILL
XFILL_1_BUFX2_insert512 gnd vdd FILL
XFILL_1_BUFX2_insert523 gnd vdd FILL
XFILL_1_BUFX2_insert534 gnd vdd FILL
XFILL_5__7850_ gnd vdd FILL
X_12764_ _12764_/A gnd _12764_/Y vdd INVX1
X_15552_ _9954_/Q gnd _15554_/D vdd INVX1
XSFILL104680x83050 gnd vdd FILL
XFILL_1_BUFX2_insert545 gnd vdd FILL
XFILL_1_BUFX2_insert556 gnd vdd FILL
XFILL_3__10680_ gnd vdd FILL
XFILL_1_BUFX2_insert567 gnd vdd FILL
XFILL_1_BUFX2_insert578 gnd vdd FILL
X_14503_ _13587_/A _14502_/Y _13587_/C _14501_/Y gnd _14507_/A vdd OAI22X1
XFILL112120x38050 gnd vdd FILL
X_11715_ _11713_/Y _11074_/C _11751_/C gnd _11716_/B vdd OAI21X1
XFILL_4__8988_ gnd vdd FILL
XFILL_1_BUFX2_insert589 gnd vdd FILL
X_15483_ _7060_/A gnd _15485_/D vdd INVX1
XFILL_5__11240_ gnd vdd FILL
X_12695_ _12695_/A gnd _12695_/Y vdd INVX1
XFILL_6__10791_ gnd vdd FILL
XFILL_2__9811_ gnd vdd FILL
XFILL_4__11970_ gnd vdd FILL
XFILL_1__10810_ gnd vdd FILL
XFILL_2__11060_ gnd vdd FILL
XFILL_5__9520_ gnd vdd FILL
XSFILL64040x23050 gnd vdd FILL
XFILL_4__7939_ gnd vdd FILL
XFILL_6__12530_ gnd vdd FILL
XFILL_1__11790_ gnd vdd FILL
X_11646_ _11646_/A _11366_/B _11646_/C gnd _11648_/C vdd OAI21X1
XFILL_5__11171_ gnd vdd FILL
X_14434_ _10162_/A gnd _14436_/D vdd INVX1
XFILL_4__10921_ gnd vdd FILL
XFILL_3__12350_ gnd vdd FILL
XFILL_2__10011_ gnd vdd FILL
XFILL_2__9742_ gnd vdd FILL
XFILL_2__6954_ gnd vdd FILL
XFILL_0__12170_ gnd vdd FILL
XFILL_5__10122_ gnd vdd FILL
X_14365_ _14365_/A _14479_/B _14200_/C _14365_/D gnd _14366_/A vdd OAI22X1
XFILL_3__11301_ gnd vdd FILL
XFILL_4__13640_ gnd vdd FILL
X_11577_ _11551_/A _11577_/B _11553_/C gnd _11578_/B vdd OAI21X1
XSFILL53880x66050 gnd vdd FILL
XFILL_3__12281_ gnd vdd FILL
XFILL_0__11121_ gnd vdd FILL
XFILL_4__9609_ gnd vdd FILL
XFILL_2__6885_ gnd vdd FILL
XFILL_1__13460_ gnd vdd FILL
XFILL_2__9673_ gnd vdd FILL
XFILL_5__8402_ gnd vdd FILL
X_13316_ _13248_/A _13316_/B gnd _13316_/Y vdd NOR2X1
X_16104_ _15524_/A _16104_/B _14733_/D _15521_/C gnd _16104_/Y vdd OAI22X1
XFILL_1__10672_ gnd vdd FILL
XFILL_5__9382_ gnd vdd FILL
X_10528_ _10596_/Q gnd _10528_/Y vdd INVX1
XFILL_3__14020_ gnd vdd FILL
XFILL_5__14930_ gnd vdd FILL
XFILL_5__10053_ gnd vdd FILL
XFILL_6__12392_ gnd vdd FILL
XFILL_3__11232_ gnd vdd FILL
X_14296_ _14294_/Y _14946_/A _14456_/C _15766_/B gnd _14296_/Y vdd OAI22X1
XFILL_1__12411_ gnd vdd FILL
XFILL_2__14750_ gnd vdd FILL
XFILL_2__8624_ gnd vdd FILL
XFILL_4__10783_ gnd vdd FILL
XFILL_4__13571_ gnd vdd FILL
XFILL_2__11962_ gnd vdd FILL
XFILL_0__11052_ gnd vdd FILL
XFILL_5__8333_ gnd vdd FILL
XFILL_1__13391_ gnd vdd FILL
X_13247_ _13289_/B _13310_/A gnd _13248_/A vdd NOR2X1
X_16035_ _9918_/A _16035_/B _16037_/C gnd _16036_/C vdd NAND3X1
XFILL_4__15310_ gnd vdd FILL
XFILL_5__14861_ gnd vdd FILL
XFILL_4__12522_ gnd vdd FILL
X_10459_ _15261_/A _8151_/CLK _9048_/R vdd _10375_/Y gnd vdd DFFSR
XFILL_2__13701_ gnd vdd FILL
XFILL_2__10913_ gnd vdd FILL
XFILL_4__16290_ gnd vdd FILL
XFILL_3__11163_ gnd vdd FILL
XFILL_0__10003_ gnd vdd FILL
XFILL_1__15130_ gnd vdd FILL
XSFILL94360x80050 gnd vdd FILL
XFILL_1__12342_ gnd vdd FILL
XFILL_2__14681_ gnd vdd FILL
XFILL_2__11893_ gnd vdd FILL
XFILL_5__8264_ gnd vdd FILL
XFILL_0__15860_ gnd vdd FILL
XFILL_5__13812_ gnd vdd FILL
X_13178_ _11896_/A _12669_/CLK _9050_/R vdd _13090_/Y gnd vdd DFFSR
XFILL_3__10114_ gnd vdd FILL
XFILL_4__15241_ gnd vdd FILL
XFILL_0__7570_ gnd vdd FILL
XFILL_2__7506_ gnd vdd FILL
XFILL_2__13632_ gnd vdd FILL
XFILL_5__14792_ gnd vdd FILL
XFILL_4__12453_ gnd vdd FILL
XFILL_3__15971_ gnd vdd FILL
XFILL_2__8486_ gnd vdd FILL
XFILL_0__14811_ gnd vdd FILL
XFILL_1__15061_ gnd vdd FILL
XFILL_3__11094_ gnd vdd FILL
XFILL_5__7215_ gnd vdd FILL
XFILL_1__12273_ gnd vdd FILL
XFILL_5__8195_ gnd vdd FILL
X_12129_ _12127_/Y _12134_/A _12129_/C gnd _12129_/Y vdd OAI21X1
XFILL_0__15791_ gnd vdd FILL
XFILL_5__13743_ gnd vdd FILL
XFILL_4__11404_ gnd vdd FILL
XFILL_2__7437_ gnd vdd FILL
XFILL_5__10955_ gnd vdd FILL
XFILL_3__10045_ gnd vdd FILL
XFILL_1__14012_ gnd vdd FILL
XFILL_4__12384_ gnd vdd FILL
XFILL_2__16351_ gnd vdd FILL
XFILL_4__15172_ gnd vdd FILL
XFILL_3__14922_ gnd vdd FILL
XFILL_2__13563_ gnd vdd FILL
XFILL112200x18050 gnd vdd FILL
XFILL_1__11224_ gnd vdd FILL
XFILL_2__10775_ gnd vdd FILL
XFILL_0__14742_ gnd vdd FILL
XFILL_0__11954_ gnd vdd FILL
XFILL_0__9240_ gnd vdd FILL
XFILL_4__14123_ gnd vdd FILL
XFILL_2__15302_ gnd vdd FILL
XFILL_5__13674_ gnd vdd FILL
XFILL_2__12514_ gnd vdd FILL
XFILL_4__11335_ gnd vdd FILL
XFILL_3__14853_ gnd vdd FILL
XSFILL88440x41050 gnd vdd FILL
XFILL_2__7368_ gnd vdd FILL
XFILL_5__10886_ gnd vdd FILL
XFILL_0_BUFX2_insert17 gnd vdd FILL
XFILL_2__16282_ gnd vdd FILL
XFILL_0__10905_ gnd vdd FILL
XFILL_0_BUFX2_insert28 gnd vdd FILL
XFILL_2__13494_ gnd vdd FILL
XFILL_1__11155_ gnd vdd FILL
XFILL_5__7077_ gnd vdd FILL
XFILL_5__15413_ gnd vdd FILL
XFILL_0__14673_ gnd vdd FILL
XFILL_0_BUFX2_insert39 gnd vdd FILL
XFILL_0__11885_ gnd vdd FILL
XFILL_5__12625_ gnd vdd FILL
XFILL_0__9171_ gnd vdd FILL
XFILL_3__13804_ gnd vdd FILL
XFILL_5__16393_ gnd vdd FILL
XFILL_2__15233_ gnd vdd FILL
XFILL_4__14054_ gnd vdd FILL
XFILL_2__9107_ gnd vdd FILL
XFILL_4__11266_ gnd vdd FILL
XFILL_2__12445_ gnd vdd FILL
XFILL_1__10106_ gnd vdd FILL
XFILL_0__16412_ gnd vdd FILL
XFILL_0__13624_ gnd vdd FILL
XFILL_2__7299_ gnd vdd FILL
XFILL_3__11996_ gnd vdd FILL
XFILL_1__15963_ gnd vdd FILL
XFILL_3__14784_ gnd vdd FILL
XFILL_0__8122_ gnd vdd FILL
XFILL_1__11086_ gnd vdd FILL
XFILL_0__10836_ gnd vdd FILL
XFILL_5__15344_ gnd vdd FILL
XSFILL53960x46050 gnd vdd FILL
X_15819_ _15819_/A _15818_/Y _15816_/Y gnd _15819_/Y vdd NAND3X1
XFILL_4__13005_ gnd vdd FILL
XFILL_2__9038_ gnd vdd FILL
X_8750_ _8748_/Y _8695_/B _8750_/C gnd _8808_/D vdd OAI21X1
XSFILL3560x10050 gnd vdd FILL
XFILL_6__7890_ gnd vdd FILL
XFILL_3__9920_ gnd vdd FILL
XFILL_2_BUFX2_insert390 gnd vdd FILL
XFILL_2__15164_ gnd vdd FILL
XFILL_3__13735_ gnd vdd FILL
XFILL_4__11197_ gnd vdd FILL
XFILL_3__10947_ gnd vdd FILL
XSFILL109480x75050 gnd vdd FILL
XFILL_1__10037_ gnd vdd FILL
XFILL_0__16343_ gnd vdd FILL
XFILL_2__12376_ gnd vdd FILL
XFILL_1__14914_ gnd vdd FILL
XFILL_1__15894_ gnd vdd FILL
XFILL_0__13555_ gnd vdd FILL
XFILL_0__10767_ gnd vdd FILL
X_7701_ _7753_/B _6933_/B gnd _7702_/C vdd NAND2X1
XFILL_5__11507_ gnd vdd FILL
XFILL_4__10148_ gnd vdd FILL
XFILL_2__14115_ gnd vdd FILL
XFILL_5__15275_ gnd vdd FILL
XSFILL28760x22050 gnd vdd FILL
XFILL_5__12487_ gnd vdd FILL
X_8681_ _8681_/Q _7664_/CLK _7920_/R vdd _8681_/D gnd vdd DFFSR
XFILL_2__11327_ gnd vdd FILL
XFILL_1__14845_ gnd vdd FILL
XSFILL54040x55050 gnd vdd FILL
XFILL_0__12506_ gnd vdd FILL
XFILL_3__13666_ gnd vdd FILL
XFILL_3__10878_ gnd vdd FILL
XFILL_3__9851_ gnd vdd FILL
XFILL_2__15095_ gnd vdd FILL
XFILL_0__16274_ gnd vdd FILL
XFILL_5__14226_ gnd vdd FILL
XFILL_0__13486_ gnd vdd FILL
XFILL_3__15405_ gnd vdd FILL
XFILL_0__10698_ gnd vdd FILL
XSFILL94440x60050 gnd vdd FILL
XFILL_5__11438_ gnd vdd FILL
XFILL_5__7979_ gnd vdd FILL
X_7632_ _7632_/A gnd _7632_/Y vdd INVX1
XFILL_3__12617_ gnd vdd FILL
XFILL_2__14046_ gnd vdd FILL
XFILL_4__14956_ gnd vdd FILL
XFILL_3__16385_ gnd vdd FILL
XFILL_0__15225_ gnd vdd FILL
XFILL_2__11258_ gnd vdd FILL
XFILL_3__13597_ gnd vdd FILL
XFILL_3__9782_ gnd vdd FILL
XFILL_0__12437_ gnd vdd FILL
XFILL_5__9718_ gnd vdd FILL
XFILL_1__14776_ gnd vdd FILL
XFILL_3__6994_ gnd vdd FILL
XFILL_6__15516_ gnd vdd FILL
XFILL_1__11988_ gnd vdd FILL
XFILL_5__14157_ gnd vdd FILL
XFILL_4__13907_ gnd vdd FILL
X_7563_ _7645_/Q gnd _7563_/Y vdd INVX1
XFILL_3__15336_ gnd vdd FILL
XFILL_5__11369_ gnd vdd FILL
XFILL_3__8733_ gnd vdd FILL
XFILL_1__13727_ gnd vdd FILL
XFILL_4__14887_ gnd vdd FILL
XFILL_1__10939_ gnd vdd FILL
XFILL_0__15156_ gnd vdd FILL
XFILL_2__11189_ gnd vdd FILL
XFILL_0__12368_ gnd vdd FILL
X_9302_ _9302_/Q _6998_/CLK _9430_/R vdd _9302_/D gnd vdd DFFSR
XFILL_5__13108_ gnd vdd FILL
XFILL_5__9649_ gnd vdd FILL
XFILL_4__13838_ gnd vdd FILL
XFILL_0__8955_ gnd vdd FILL
XFILL_5__14088_ gnd vdd FILL
XSFILL18680x74050 gnd vdd FILL
X_7494_ _7492_/Y _7457_/A _7493_/Y gnd _7494_/Y vdd OAI21X1
XFILL_3__12479_ gnd vdd FILL
XFILL_0__14107_ gnd vdd FILL
XFILL_3__15267_ gnd vdd FILL
XFILL_1__13658_ gnd vdd FILL
XFILL_0__11319_ gnd vdd FILL
XSFILL74200x68050 gnd vdd FILL
XFILL_2__15997_ gnd vdd FILL
XFILL_0__15087_ gnd vdd FILL
XFILL_6__15378_ gnd vdd FILL
XFILL_5__13039_ gnd vdd FILL
XFILL_0__12299_ gnd vdd FILL
X_9233_ _9311_/Q gnd _9233_/Y vdd INVX1
XFILL_3__14218_ gnd vdd FILL
XFILL_0__8886_ gnd vdd FILL
XFILL_1__12609_ gnd vdd FILL
XFILL_3__7615_ gnd vdd FILL
XFILL_4__13769_ gnd vdd FILL
XSFILL9160x50050 gnd vdd FILL
XFILL_3__15198_ gnd vdd FILL
XFILL_0__14038_ gnd vdd FILL
XFILL_2__14948_ gnd vdd FILL
XFILL_1__16377_ gnd vdd FILL
XFILL_3__8595_ gnd vdd FILL
XFILL_1__13589_ gnd vdd FILL
XFILL_6__14329_ gnd vdd FILL
XFILL_4__15508_ gnd vdd FILL
XSFILL49000x44050 gnd vdd FILL
XFILL_0__7837_ gnd vdd FILL
X_9164_ _9164_/A _9164_/B _9164_/C gnd _9202_/D vdd OAI21X1
XFILL_3__14149_ gnd vdd FILL
XFILL_1__15328_ gnd vdd FILL
XFILL_3__7546_ gnd vdd FILL
XFILL_2__14879_ gnd vdd FILL
XSFILL109560x55050 gnd vdd FILL
X_8115_ _8133_/A _9267_/B gnd _8116_/C vdd NAND2X1
XFILL_3_BUFX2_insert607 gnd vdd FILL
XFILL_4__15439_ gnd vdd FILL
X_9095_ _9093_/Y _9086_/B _9095_/C gnd _9095_/Y vdd OAI21X1
XFILL_3_BUFX2_insert618 gnd vdd FILL
XFILL_3__7477_ gnd vdd FILL
XFILL_1__15259_ gnd vdd FILL
XFILL_3_BUFX2_insert629 gnd vdd FILL
XFILL_0__9507_ gnd vdd FILL
XFILL_0__15989_ gnd vdd FILL
XFILL_1__9280_ gnd vdd FILL
X_8046_ _8046_/Q _8046_/CLK _8670_/R vdd _8046_/D gnd vdd DFFSR
XSFILL54120x35050 gnd vdd FILL
XFILL_3__9216_ gnd vdd FILL
XFILL_0__7699_ gnd vdd FILL
XSFILL39480x53050 gnd vdd FILL
XFILL_1__8231_ gnd vdd FILL
XFILL_3__9147_ gnd vdd FILL
XSFILL43960x78050 gnd vdd FILL
XFILL_0__9369_ gnd vdd FILL
X_9997_ _9995_/Y _9996_/A _9997_/C gnd _9997_/Y vdd OAI21X1
XFILL_3__9078_ gnd vdd FILL
XFILL_1__7113_ gnd vdd FILL
XSFILL18760x54050 gnd vdd FILL
XSFILL8600x64050 gnd vdd FILL
XFILL_1__8093_ gnd vdd FILL
X_8948_ _8912_/A _8180_/CLK _8937_/R vdd _8948_/D gnd vdd DFFSR
XFILL_4__8911_ gnd vdd FILL
XFILL_4__9891_ gnd vdd FILL
XFILL_1__7044_ gnd vdd FILL
X_8879_ _8879_/A gnd _8881_/A vdd INVX1
XFILL_4__8842_ gnd vdd FILL
XSFILL43960x6050 gnd vdd FILL
XSFILL23880x45050 gnd vdd FILL
XFILL_0_BUFX2_insert508 gnd vdd FILL
XFILL_0_BUFX2_insert519 gnd vdd FILL
X_11500_ _11494_/A _11186_/Y _11500_/C gnd _11500_/Y vdd NAND3X1
XFILL_4__8773_ gnd vdd FILL
X_12480_ _12480_/A vdd _12479_/Y gnd _12548_/D vdd OAI21X1
XFILL112440x74050 gnd vdd FILL
XFILL_1__8995_ gnd vdd FILL
XFILL_4__7724_ gnd vdd FILL
X_11431_ _11431_/A _11431_/B _11431_/C gnd _11431_/Y vdd AOI21X1
XFILL_1__7946_ gnd vdd FILL
X_14150_ _7328_/A gnd _14152_/A vdd INVX1
XSFILL39000x76050 gnd vdd FILL
X_11362_ _11201_/Y gnd _11362_/Y vdd INVX1
XFILL_1__7877_ gnd vdd FILL
X_13101_ _13153_/B _13101_/B gnd _13101_/Y vdd NAND2X1
XFILL_4__7586_ gnd vdd FILL
X_10313_ _10313_/A _10280_/B _10312_/Y gnd _10353_/D vdd OAI21X1
X_14081_ _14081_/A gnd _14083_/D vdd INVX1
XFILL_4_BUFX2_insert430 gnd vdd FILL
XFILL_1__9616_ gnd vdd FILL
X_11293_ _11521_/C _11527_/C gnd _11313_/B vdd NOR2X1
XFILL_4_BUFX2_insert441 gnd vdd FILL
XFILL_4_BUFX2_insert452 gnd vdd FILL
XFILL_4_BUFX2_insert463 gnd vdd FILL
XSFILL18840x34050 gnd vdd FILL
X_13032_ _6897_/A gnd _13032_/Y vdd INVX1
XCLKBUF1_insert209 CLKBUF1_insert220/A gnd _9205_/CLK vdd CLKBUF1
X_10244_ _10244_/A _10294_/A _10243_/Y gnd _10244_/Y vdd OAI21X1
XFILL_4_BUFX2_insert474 gnd vdd FILL
XSFILL44120x67050 gnd vdd FILL
XFILL_2__8340_ gnd vdd FILL
XFILL_4_BUFX2_insert485 gnd vdd FILL
XFILL_4_BUFX2_insert496 gnd vdd FILL
XFILL_1__9547_ gnd vdd FILL
XSFILL59720x46050 gnd vdd FILL
XFILL_4__9256_ gnd vdd FILL
XSFILL69080x71050 gnd vdd FILL
X_10175_ _10127_/A _8511_/B gnd _10176_/C vdd NAND2X1
XSFILL99320x32050 gnd vdd FILL
XFILL_2__8271_ gnd vdd FILL
XFILL_1__9478_ gnd vdd FILL
XFILL_4__8207_ gnd vdd FILL
XFILL_2__7222_ gnd vdd FILL
X_14983_ _14983_/A _14982_/Y _14981_/Y gnd _14983_/Y vdd NAND3X1
XFILL_2__10560_ gnd vdd FILL
XFILL_4__8138_ gnd vdd FILL
XSFILL64040x18050 gnd vdd FILL
XFILL_4__11120_ gnd vdd FILL
XFILL_3_CLKBUF1_insert121 gnd vdd FILL
X_13934_ _15482_/A _14344_/B _13933_/Y gnd _13934_/Y vdd AOI21X1
XFILL_5__10671_ gnd vdd FILL
XFILL_3__11850_ gnd vdd FILL
XFILL_5_CLKBUF1_insert1081 gnd vdd FILL
XFILL_3_CLKBUF1_insert132 gnd vdd FILL
XFILL_3_CLKBUF1_insert143 gnd vdd FILL
XFILL_2__10491_ gnd vdd FILL
XFILL_4__8069_ gnd vdd FILL
XFILL_5__12410_ gnd vdd FILL
XFILL_5__8951_ gnd vdd FILL
XFILL_0__11670_ gnd vdd FILL
XFILL_3_CLKBUF1_insert154 gnd vdd FILL
XFILL_3_CLKBUF1_insert165 gnd vdd FILL
XFILL_4__11051_ gnd vdd FILL
X_13865_ _7902_/Q _13865_/B _13865_/C _7694_/A gnd _13873_/B vdd AOI22X1
XFILL_5__13390_ gnd vdd FILL
XFILL_3_CLKBUF1_insert176 gnd vdd FILL
XFILL_2__12230_ gnd vdd FILL
XFILL_3__10801_ gnd vdd FILL
XFILL_2__7084_ gnd vdd FILL
XFILL_3__11781_ gnd vdd FILL
XFILL_3_CLKBUF1_insert187 gnd vdd FILL
XFILL_1__12960_ gnd vdd FILL
XFILL_0__10621_ gnd vdd FILL
XFILL_3_CLKBUF1_insert198 gnd vdd FILL
XFILL_4__10002_ gnd vdd FILL
XFILL_6__13700_ gnd vdd FILL
X_15604_ _14098_/C gnd _15604_/Y vdd INVX1
XFILL_1_BUFX2_insert320 gnd vdd FILL
X_12816_ _12816_/Q _9050_/CLK _9050_/R vdd _12816_/D gnd vdd DFFSR
XFILL_5__12341_ gnd vdd FILL
XFILL_5__8882_ gnd vdd FILL
XFILL_3__13520_ gnd vdd FILL
XFILL_1_BUFX2_insert331 gnd vdd FILL
X_13796_ _13796_/A _13792_/Y gnd _13805_/B vdd NOR2X1
XFILL_1__11911_ gnd vdd FILL
XFILL_2__12161_ gnd vdd FILL
XFILL_1_BUFX2_insert342 gnd vdd FILL
XFILL_1_BUFX2_insert353 gnd vdd FILL
XFILL_0__13340_ gnd vdd FILL
XFILL_5__7833_ gnd vdd FILL
XFILL_0__10552_ gnd vdd FILL
XFILL_1__12891_ gnd vdd FILL
XFILL_1_BUFX2_insert364 gnd vdd FILL
XFILL_4__14810_ gnd vdd FILL
XFILL_5__15060_ gnd vdd FILL
X_15535_ _15535_/A _15535_/B _15534_/Y gnd _15535_/Y vdd NOR3X1
X_12747_ _12762_/A memoryOutData[17] gnd _12748_/C vdd NAND2X1
XFILL_1_BUFX2_insert375 gnd vdd FILL
XFILL_5__12272_ gnd vdd FILL
XFILL_2__11112_ gnd vdd FILL
XFILL_1__14630_ gnd vdd FILL
XFILL_3__10663_ gnd vdd FILL
XFILL_1_BUFX2_insert386 gnd vdd FILL
XFILL_3__13451_ gnd vdd FILL
XFILL_4__15790_ gnd vdd FILL
XSFILL114440x1050 gnd vdd FILL
XFILL_1_BUFX2_insert397 gnd vdd FILL
XSFILL94360x75050 gnd vdd FILL
XFILL_2__12092_ gnd vdd FILL
XFILL_1__11842_ gnd vdd FILL
XFILL_0__13271_ gnd vdd FILL
XFILL_5__14011_ gnd vdd FILL
XFILL_5__7764_ gnd vdd FILL
XFILL_6__16350_ gnd vdd FILL
XFILL_5__11223_ gnd vdd FILL
XSFILL29560x65050 gnd vdd FILL
X_12678_ _12612_/A _12538_/CLK _12689_/R vdd _12678_/D gnd vdd DFFSR
XFILL_3__12402_ gnd vdd FILL
XFILL_4__14741_ gnd vdd FILL
X_15466_ _15466_/A _15466_/B _15466_/C gnd _15473_/B vdd NAND3X1
XFILL_2__15920_ gnd vdd FILL
XFILL_3__16170_ gnd vdd FILL
XFILL_4__11953_ gnd vdd FILL
XFILL_3__13382_ gnd vdd FILL
XFILL_0__15010_ gnd vdd FILL
XFILL_2__11043_ gnd vdd FILL
XFILL_1__14561_ gnd vdd FILL
XFILL_5__9503_ gnd vdd FILL
XFILL_0__12222_ gnd vdd FILL
XSFILL69960x70050 gnd vdd FILL
XFILL_6__15301_ gnd vdd FILL
XSFILL69160x51050 gnd vdd FILL
XFILL_1__11773_ gnd vdd FILL
XSFILL99400x12050 gnd vdd FILL
XFILL_2__7986_ gnd vdd FILL
X_11629_ _11629_/A gnd _12057_/A vdd INVX1
X_14417_ _13879_/B _14415_/Y _14744_/B _15869_/B gnd _14417_/Y vdd OAI22X1
XFILL_5__7695_ gnd vdd FILL
XFILL_4__10904_ gnd vdd FILL
XFILL_1__16300_ gnd vdd FILL
XFILL_3__12333_ gnd vdd FILL
XFILL_5__11154_ gnd vdd FILL
XFILL_3__15121_ gnd vdd FILL
X_15397_ _10334_/Q _15178_/C _15397_/C gnd _15398_/C vdd AOI21X1
XFILL_2__9725_ gnd vdd FILL
XFILL_4__14672_ gnd vdd FILL
XFILL_1__13512_ gnd vdd FILL
XFILL_4__11884_ gnd vdd FILL
XFILL_2__6937_ gnd vdd FILL
XFILL_2__15851_ gnd vdd FILL
XFILL_1__14492_ gnd vdd FILL
XFILL_0__12153_ gnd vdd FILL
XFILL_0__8740_ gnd vdd FILL
XFILL_4__16411_ gnd vdd FILL
XFILL_5__10105_ gnd vdd FILL
XFILL_4__13623_ gnd vdd FILL
X_14348_ _14346_/Y _14636_/C _14555_/C _14348_/D gnd _14352_/B vdd OAI22X1
XFILL_1__16231_ gnd vdd FILL
XFILL_2__14802_ gnd vdd FILL
XFILL_5__15962_ gnd vdd FILL
XFILL_3__15052_ gnd vdd FILL
XFILL_3__12264_ gnd vdd FILL
XFILL_5__11085_ gnd vdd FILL
XFILL_4__10835_ gnd vdd FILL
XFILL_1__13443_ gnd vdd FILL
XFILL_2__9656_ gnd vdd FILL
XFILL_0__11104_ gnd vdd FILL
XFILL_0__12084_ gnd vdd FILL
XFILL_2__12994_ gnd vdd FILL
XFILL_2__6868_ gnd vdd FILL
XFILL_2__15782_ gnd vdd FILL
XFILL_1__10655_ gnd vdd FILL
XSFILL78440x6050 gnd vdd FILL
XFILL_5__9365_ gnd vdd FILL
XFILL_6__15163_ gnd vdd FILL
XFILL_4__16342_ gnd vdd FILL
XFILL_3__14003_ gnd vdd FILL
XFILL_5__10036_ gnd vdd FILL
XFILL_5__14913_ gnd vdd FILL
X_14279_ _9575_/Q gnd _14279_/Y vdd INVX1
XFILL_3__11215_ gnd vdd FILL
XFILL_5__15893_ gnd vdd FILL
XFILL_2__8607_ gnd vdd FILL
XFILL_4__13554_ gnd vdd FILL
XFILL_4__10766_ gnd vdd FILL
XFILL_3__8380_ gnd vdd FILL
XFILL_0__15912_ gnd vdd FILL
XFILL_2__11945_ gnd vdd FILL
XFILL_2__14733_ gnd vdd FILL
XFILL_3__12195_ gnd vdd FILL
XFILL_1__16162_ gnd vdd FILL
XFILL_0__11035_ gnd vdd FILL
XFILL_1__13374_ gnd vdd FILL
XFILL_5__8316_ gnd vdd FILL
XFILL_6__14114_ gnd vdd FILL
X_16018_ _16018_/A _15407_/B _16018_/C _14642_/Y gnd _16018_/Y vdd OAI22X1
XFILL_0__7622_ gnd vdd FILL
XFILL_5__14844_ gnd vdd FILL
XSFILL89320x64050 gnd vdd FILL
XFILL_4__12505_ gnd vdd FILL
XFILL_5__9296_ gnd vdd FILL
XFILL_3__7331_ gnd vdd FILL
XFILL_3__11146_ gnd vdd FILL
XFILL_1__15113_ gnd vdd FILL
XFILL_4__16273_ gnd vdd FILL
XFILL_4__13485_ gnd vdd FILL
XFILL_1__12325_ gnd vdd FILL
XFILL_2__11876_ gnd vdd FILL
XFILL_1__16093_ gnd vdd FILL
XFILL_0__15843_ gnd vdd FILL
XFILL_2__14664_ gnd vdd FILL
XFILL_4__10697_ gnd vdd FILL
XFILL_5__8247_ gnd vdd FILL
XFILL_0__7553_ gnd vdd FILL
XFILL_4__15224_ gnd vdd FILL
XFILL_6__11257_ gnd vdd FILL
XFILL_4__12436_ gnd vdd FILL
XFILL_2__16403_ gnd vdd FILL
XFILL_5__14775_ gnd vdd FILL
XFILL_2__13615_ gnd vdd FILL
XFILL_2__10827_ gnd vdd FILL
XFILL_5__11987_ gnd vdd FILL
XFILL_1__15044_ gnd vdd FILL
XFILL_3__15954_ gnd vdd FILL
XFILL_3__11077_ gnd vdd FILL
XFILL_2__14595_ gnd vdd FILL
XFILL_1__12256_ gnd vdd FILL
XFILL_2__8469_ gnd vdd FILL
XFILL_0__15774_ gnd vdd FILL
X_9920_ _9918_/Y _9920_/B _9920_/C gnd _9966_/D vdd OAI21X1
XFILL_0__12986_ gnd vdd FILL
XFILL_5__13726_ gnd vdd FILL
XFILL_5__10938_ gnd vdd FILL
XFILL_0__7484_ gnd vdd FILL
XSFILL94440x55050 gnd vdd FILL
XFILL_3__10028_ gnd vdd FILL
XFILL_4__15155_ gnd vdd FILL
XFILL_3__14905_ gnd vdd FILL
XFILL_3__9001_ gnd vdd FILL
XFILL_4__12367_ gnd vdd FILL
XFILL_2__16334_ gnd vdd FILL
XFILL_2__13546_ gnd vdd FILL
XFILL_1__11207_ gnd vdd FILL
XFILL_3__7193_ gnd vdd FILL
XFILL_0__14725_ gnd vdd FILL
XFILL_2__10758_ gnd vdd FILL
XFILL_3__15885_ gnd vdd FILL
XFILL_1__12187_ gnd vdd FILL
XFILL_0__11937_ gnd vdd FILL
XFILL_0__9223_ gnd vdd FILL
XFILL_4__14106_ gnd vdd FILL
XSFILL95080x21050 gnd vdd FILL
XFILL_5__13657_ gnd vdd FILL
XFILL_4__11318_ gnd vdd FILL
X_9851_ _9851_/A _9941_/B _9851_/C gnd _9851_/Y vdd OAI21X1
XFILL_6__8991_ gnd vdd FILL
XFILL_3__14836_ gnd vdd FILL
XFILL_4__15086_ gnd vdd FILL
XSFILL69240x31050 gnd vdd FILL
XSFILL53960x1050 gnd vdd FILL
XFILL_1__11138_ gnd vdd FILL
XFILL_2__13477_ gnd vdd FILL
XFILL_2__16265_ gnd vdd FILL
XFILL_4__12298_ gnd vdd FILL
XFILL_0__14656_ gnd vdd FILL
XFILL_2__10689_ gnd vdd FILL
XFILL_5__12608_ gnd vdd FILL
X_8802_ _8802_/Q _7778_/CLK _8418_/R vdd _8732_/Y gnd vdd DFFSR
XFILL_0__11868_ gnd vdd FILL
XFILL_6__7942_ gnd vdd FILL
XFILL_0__9154_ gnd vdd FILL
XFILL_4__14037_ gnd vdd FILL
XFILL_5__16376_ gnd vdd FILL
X_9782_ _9789_/B _9782_/B gnd _9783_/C vdd NAND2X1
XFILL_5__13588_ gnd vdd FILL
XFILL_2__12428_ gnd vdd FILL
XFILL_2__15216_ gnd vdd FILL
XFILL_4__11249_ gnd vdd FILL
XFILL_0__13607_ gnd vdd FILL
XFILL_2__16196_ gnd vdd FILL
XFILL_3__14767_ gnd vdd FILL
X_6994_ _6994_/A _6982_/B _6994_/C gnd _7028_/D vdd OAI21X1
XSFILL104440x40050 gnd vdd FILL
XFILL_1__15946_ gnd vdd FILL
XFILL_3__11979_ gnd vdd FILL
XFILL_0__10819_ gnd vdd FILL
XFILL_1__11069_ gnd vdd FILL
XFILL_0__8105_ gnd vdd FILL
XFILL_0__14587_ gnd vdd FILL
XFILL_5__15327_ gnd vdd FILL
X_8733_ _8733_/A gnd _8735_/A vdd INVX1
XFILL_0__11799_ gnd vdd FILL
XFILL_0__9085_ gnd vdd FILL
XFILL_3__13718_ gnd vdd FILL
XFILL_3__9903_ gnd vdd FILL
XFILL_2__15147_ gnd vdd FILL
XFILL_2__12359_ gnd vdd FILL
XFILL_0__16326_ gnd vdd FILL
XFILL_6__9612_ gnd vdd FILL
XFILL_3__14698_ gnd vdd FILL
XFILL_0__13538_ gnd vdd FILL
XFILL_6_BUFX2_insert536 gnd vdd FILL
XFILL_1__15877_ gnd vdd FILL
XFILL_5__15258_ gnd vdd FILL
XSFILL49000x39050 gnd vdd FILL
X_8664_ _8572_/A _8663_/CLK _8664_/R vdd _8664_/D gnd vdd DFFSR
XFILL_4__15988_ gnd vdd FILL
XFILL_3__13649_ gnd vdd FILL
XFILL_2__15078_ gnd vdd FILL
XSFILL59160x83050 gnd vdd FILL
XFILL_1__14828_ gnd vdd FILL
XSFILL89400x44050 gnd vdd FILL
XFILL_0__16257_ gnd vdd FILL
XFILL_5__14209_ gnd vdd FILL
XFILL_0__13469_ gnd vdd FILL
X_7615_ _7568_/B _7359_/B gnd _7615_/Y vdd NAND2X1
XFILL_5__15189_ gnd vdd FILL
XFILL_2__14029_ gnd vdd FILL
XFILL_4__14939_ gnd vdd FILL
XFILL_0__15208_ gnd vdd FILL
X_8595_ _8593_/Y _8657_/A _8595_/C gnd _8595_/Y vdd OAI21X1
XFILL_3__16368_ gnd vdd FILL
XFILL_3__9765_ gnd vdd FILL
XFILL_1__14759_ gnd vdd FILL
XFILL_0__16188_ gnd vdd FILL
XFILL_3__6977_ gnd vdd FILL
XFILL_1__7800_ gnd vdd FILL
XFILL_3__15319_ gnd vdd FILL
XFILL_1__8780_ gnd vdd FILL
X_7546_ _7624_/A _8314_/B gnd _7547_/C vdd NAND2X1
XFILL_3__8716_ gnd vdd FILL
XFILL_0__9987_ gnd vdd FILL
XFILL_3__16299_ gnd vdd FILL
XFILL_0__15139_ gnd vdd FILL
XFILL_1__7731_ gnd vdd FILL
XFILL_4__7440_ gnd vdd FILL
X_7477_ _7531_/Q gnd _7479_/A vdd INVX1
XSFILL64440x8050 gnd vdd FILL
XFILL_3__8647_ gnd vdd FILL
XSFILL113640x77050 gnd vdd FILL
XSFILL13720x4050 gnd vdd FILL
X_9216_ _9232_/B _7424_/B gnd _9217_/C vdd NAND2X1
XFILL_6__8356_ gnd vdd FILL
XFILL_0__8869_ gnd vdd FILL
XFILL_4__7371_ gnd vdd FILL
XFILL_6__7307_ gnd vdd FILL
XFILL_3__8578_ gnd vdd FILL
XFILL_1__9401_ gnd vdd FILL
X_9147_ _9197_/Q gnd _9147_/Y vdd INVX1
XSFILL18760x49050 gnd vdd FILL
XFILL_3_BUFX2_insert404 gnd vdd FILL
XSFILL8600x59050 gnd vdd FILL
XFILL_1__7593_ gnd vdd FILL
XFILL_4__9110_ gnd vdd FILL
XSFILL104520x20050 gnd vdd FILL
XFILL_3_BUFX2_insert415 gnd vdd FILL
XFILL_3_BUFX2_insert426 gnd vdd FILL
XFILL_3_BUFX2_insert437 gnd vdd FILL
X_9078_ _9078_/A gnd _9078_/Y vdd INVX1
XFILL_3_BUFX2_insert448 gnd vdd FILL
XSFILL99240x47050 gnd vdd FILL
XFILL_4__9041_ gnd vdd FILL
XFILL_3_BUFX2_insert459 gnd vdd FILL
X_8029_ _7947_/A _7915_/CLK _7915_/R vdd _8029_/D gnd vdd DFFSR
XFILL_1__9263_ gnd vdd FILL
XFILL_1__8214_ gnd vdd FILL
X_11980_ _13172_/A gnd _11980_/Y vdd INVX1
XSFILL108600x66050 gnd vdd FILL
XFILL111960x62050 gnd vdd FILL
XFILL112440x69050 gnd vdd FILL
X_10931_ _10930_/Y gnd _10935_/A vdd INVX1
XFILL_1__8145_ gnd vdd FILL
XFILL_0_BUFX2_insert9 gnd vdd FILL
XSFILL79160x14050 gnd vdd FILL
X_10862_ _10862_/Q _7790_/CLK _9566_/R vdd _10862_/D gnd vdd DFFSR
XFILL112040x71050 gnd vdd FILL
X_13650_ _7938_/A gnd _15226_/B vdd INVX1
XFILL_1__8076_ gnd vdd FILL
XFILL_4_CLKBUF1_insert205 gnd vdd FILL
XFILL_4_CLKBUF1_insert216 gnd vdd FILL
X_12601_ vdd memoryOutData[11] gnd _12602_/C vdd NAND2X1
XFILL_4__9874_ gnd vdd FILL
X_13581_ _7804_/A _13865_/B _14037_/C _6908_/A gnd _13582_/B vdd AOI22X1
X_10793_ _14289_/D gnd _10795_/A vdd INVX1
XFILL_0_BUFX2_insert305 gnd vdd FILL
XFILL_4__8825_ gnd vdd FILL
X_15320_ _9820_/Q gnd _15321_/B vdd INVX1
XFILL_0_BUFX2_insert316 gnd vdd FILL
X_12532_ _12436_/A gnd _12534_/A vdd INVX1
XSFILL18840x29050 gnd vdd FILL
XFILL_0_BUFX2_insert327 gnd vdd FILL
XFILL_0_BUFX2_insert338 gnd vdd FILL
XFILL_2__7840_ gnd vdd FILL
XFILL_0_BUFX2_insert349 gnd vdd FILL
XFILL_4__8756_ gnd vdd FILL
X_15251_ _8410_/Q gnd _15251_/Y vdd INVX1
X_12463_ _11912_/B gnd _12465_/A vdd INVX1
XSFILL69080x66050 gnd vdd FILL
XSFILL99320x27050 gnd vdd FILL
XFILL_4__7707_ gnd vdd FILL
XFILL_1__8978_ gnd vdd FILL
X_14202_ _9507_/A gnd _14203_/D vdd INVX1
XFILL_5__7480_ gnd vdd FILL
X_11414_ _11414_/A _11369_/Y _11414_/C gnd _11414_/Y vdd NAND3X1
X_15182_ _13615_/Y _15683_/B _15407_/C _15182_/D gnd _15183_/A vdd OAI22X1
XFILL_2__9510_ gnd vdd FILL
X_12394_ _12055_/B gnd _12394_/Y vdd INVX1
XSFILL99480x6050 gnd vdd FILL
XFILL_1__7929_ gnd vdd FILL
X_14133_ _14133_/A _14132_/Y _14133_/C gnd _14144_/B vdd NAND3X1
X_11345_ _11343_/Y _10997_/Y _11415_/C gnd _11346_/C vdd OAI21X1
XFILL_4__10620_ gnd vdd FILL
XFILL_1__10440_ gnd vdd FILL
XFILL_5__9150_ gnd vdd FILL
XFILL_5__11910_ gnd vdd FILL
X_14064_ _13621_/B _15537_/B _7578_/A _14185_/B gnd _14073_/A vdd AOI22X1
XFILL_4__7569_ gnd vdd FILL
XFILL_4_BUFX2_insert260 gnd vdd FILL
XFILL_3__11000_ gnd vdd FILL
XSFILL23000x65050 gnd vdd FILL
XFILL_4_BUFX2_insert271 gnd vdd FILL
X_11276_ _11263_/B _11271_/Y _11275_/Y gnd _11653_/A vdd OAI21X1
XFILL_4__10551_ gnd vdd FILL
XFILL_4_BUFX2_insert282 gnd vdd FILL
XFILL_5__12890_ gnd vdd FILL
XFILL_2__9372_ gnd vdd FILL
XFILL_2__11730_ gnd vdd FILL
XFILL_5__8101_ gnd vdd FILL
XFILL_4_BUFX2_insert293 gnd vdd FILL
X_13015_ vdd _13015_/B gnd _13016_/C vdd NAND2X1
XFILL112120x51050 gnd vdd FILL
XFILL_1__10371_ gnd vdd FILL
XFILL_5_BUFX2_insert1006 gnd vdd FILL
X_10227_ _10189_/A _8038_/CLK _8038_/R vdd _10227_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert1017 gnd vdd FILL
XFILL_5__9081_ gnd vdd FILL
XFILL_5_BUFX2_insert1028 gnd vdd FILL
XFILL_5__11841_ gnd vdd FILL
XFILL_4__13270_ gnd vdd FILL
XFILL_5_BUFX2_insert1039 gnd vdd FILL
XFILL_2__8323_ gnd vdd FILL
XFILL_1__12110_ gnd vdd FILL
XFILL_2__11661_ gnd vdd FILL
XFILL_1__13090_ gnd vdd FILL
XFILL_4__9239_ gnd vdd FILL
XFILL_0__12840_ gnd vdd FILL
XFILL_3_BUFX2_insert960 gnd vdd FILL
XFILL_6__11042_ gnd vdd FILL
XFILL_5__14560_ gnd vdd FILL
XFILL_2__13400_ gnd vdd FILL
X_10158_ _10158_/A _10140_/B _10158_/C gnd _10158_/Y vdd OAI21X1
XFILL_4__12221_ gnd vdd FILL
XFILL_2__8254_ gnd vdd FILL
XFILL_3_BUFX2_insert971 gnd vdd FILL
XFILL_5__11772_ gnd vdd FILL
XSFILL4360x48050 gnd vdd FILL
XFILL_3_BUFX2_insert982 gnd vdd FILL
XFILL_1__12041_ gnd vdd FILL
XFILL_3__12951_ gnd vdd FILL
XFILL_2__14380_ gnd vdd FILL
XFILL_3_BUFX2_insert993 gnd vdd FILL
XFILL_2__11592_ gnd vdd FILL
XFILL_0__12771_ gnd vdd FILL
XFILL_5__13511_ gnd vdd FILL
XFILL_2__7205_ gnd vdd FILL
XFILL_2__13331_ gnd vdd FILL
XFILL_5__14491_ gnd vdd FILL
XFILL_3__11902_ gnd vdd FILL
XFILL_4__12152_ gnd vdd FILL
X_14966_ _8147_/A gnd _14967_/A vdd INVX1
X_10089_ _15846_/A _9705_/CLK _9964_/R vdd _10089_/D gnd vdd DFFSR
XFILL_3__15670_ gnd vdd FILL
XFILL_0__14510_ gnd vdd FILL
XFILL_2__10543_ gnd vdd FILL
XFILL_2__8185_ gnd vdd FILL
XFILL_3__12882_ gnd vdd FILL
XFILL_0__11722_ gnd vdd FILL
XFILL_5__16230_ gnd vdd FILL
XSFILL69160x46050 gnd vdd FILL
XFILL_0__15490_ gnd vdd FILL
XFILL_5__9983_ gnd vdd FILL
XFILL_5__13442_ gnd vdd FILL
XFILL_4__11103_ gnd vdd FILL
X_13917_ _13917_/A _13917_/B gnd _13918_/C vdd NOR2X1
XFILL_3__14621_ gnd vdd FILL
XFILL_4__12083_ gnd vdd FILL
XFILL_5__10654_ gnd vdd FILL
XFILL_2__16050_ gnd vdd FILL
XFILL_2__13262_ gnd vdd FILL
XFILL_3_BUFX2_insert1010 gnd vdd FILL
XFILL_1__15800_ gnd vdd FILL
XFILL_3__11833_ gnd vdd FILL
X_14897_ _13879_/B _14895_/Y _16264_/A _14897_/D gnd _14897_/Y vdd OAI22X1
XFILL_3_BUFX2_insert1021 gnd vdd FILL
XFILL_0__14441_ gnd vdd FILL
XFILL_3_BUFX2_insert1032 gnd vdd FILL
XFILL_1__13992_ gnd vdd FILL
XFILL_0__11653_ gnd vdd FILL
XFILL_3_BUFX2_insert1043 gnd vdd FILL
XFILL_4__15911_ gnd vdd FILL
XFILL_2__15001_ gnd vdd FILL
XFILL_5__16161_ gnd vdd FILL
XFILL_4__11034_ gnd vdd FILL
X_13848_ _8414_/Q _13848_/B _13848_/C _7646_/Q gnd _13852_/A vdd AOI22X1
XFILL_2__12213_ gnd vdd FILL
XFILL_5__13373_ gnd vdd FILL
XFILL_3__14552_ gnd vdd FILL
XFILL_3_BUFX2_insert1054 gnd vdd FILL
XSFILL104360x55050 gnd vdd FILL
XFILL_2__7067_ gnd vdd FILL
XFILL_1__15731_ gnd vdd FILL
XFILL_3_BUFX2_insert1065 gnd vdd FILL
XFILL_3__11764_ gnd vdd FILL
XFILL_0__14372_ gnd vdd FILL
XFILL_5__15112_ gnd vdd FILL
XFILL_3_BUFX2_insert1087 gnd vdd FILL
XFILL_5__8865_ gnd vdd FILL
XSFILL74280x37050 gnd vdd FILL
XFILL_5__12324_ gnd vdd FILL
XFILL_0__11584_ gnd vdd FILL
XFILL_5__16092_ gnd vdd FILL
XFILL_4__15842_ gnd vdd FILL
XFILL_3__13503_ gnd vdd FILL
X_13779_ _13779_/A _13778_/Y gnd _13787_/B vdd NOR2X1
XFILL_0__16111_ gnd vdd FILL
XFILL_2__12144_ gnd vdd FILL
XFILL_3__6900_ gnd vdd FILL
XFILL_0__13323_ gnd vdd FILL
XFILL_3__14483_ gnd vdd FILL
XFILL_1__15662_ gnd vdd FILL
XFILL_3__11695_ gnd vdd FILL
XFILL_0__10535_ gnd vdd FILL
XFILL_5__7816_ gnd vdd FILL
XFILL_1__12874_ gnd vdd FILL
XFILL_3__7880_ gnd vdd FILL
XFILL_0__9910_ gnd vdd FILL
XFILL_5__15043_ gnd vdd FILL
X_15518_ _15518_/A _15518_/B gnd _15523_/A vdd NOR2X1
XFILL_3__16222_ gnd vdd FILL
XSFILL89320x59050 gnd vdd FILL
XFILL_5__12255_ gnd vdd FILL
XSFILL49080x13050 gnd vdd FILL
XFILL_1__14613_ gnd vdd FILL
XFILL_3__13434_ gnd vdd FILL
XFILL112200x31050 gnd vdd FILL
XFILL_4__15773_ gnd vdd FILL
XFILL_3__10646_ gnd vdd FILL
XFILL_0__16042_ gnd vdd FILL
XFILL_2__12075_ gnd vdd FILL
XFILL_4__12985_ gnd vdd FILL
XFILL_1__11825_ gnd vdd FILL
XFILL_0__13254_ gnd vdd FILL
XFILL_1__15593_ gnd vdd FILL
X_7400_ _7400_/Q _7400_/CLK _9704_/R vdd _7400_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert850 gnd vdd FILL
XFILL_5__7747_ gnd vdd FILL
XFILL_5__11206_ gnd vdd FILL
XFILL_4__14724_ gnd vdd FILL
X_15449_ _15449_/A _15527_/C _15449_/C _15448_/Y gnd _15449_/Y vdd OAI22X1
XFILL_0_BUFX2_insert861 gnd vdd FILL
X_8380_ _8360_/B _9532_/B gnd _8380_/Y vdd NAND2X1
XFILL_2__15903_ gnd vdd FILL
XFILL_5__12186_ gnd vdd FILL
XFILL_4__11936_ gnd vdd FILL
XFILL_2__11026_ gnd vdd FILL
XFILL_3__16153_ gnd vdd FILL
XFILL_3__9550_ gnd vdd FILL
XFILL_3__13365_ gnd vdd FILL
XFILL_1__14544_ gnd vdd FILL
XFILL_0_BUFX2_insert872 gnd vdd FILL
XFILL_0__12205_ gnd vdd FILL
XFILL_3__10577_ gnd vdd FILL
XFILL_2__7969_ gnd vdd FILL
XFILL_0_BUFX2_insert883 gnd vdd FILL
XFILL_1__11756_ gnd vdd FILL
XFILL_0_BUFX2_insert894 gnd vdd FILL
XFILL_0__10397_ gnd vdd FILL
XFILL_3_BUFX2_insert10 gnd vdd FILL
X_7331_ _7397_/Q gnd _7331_/Y vdd INVX1
XFILL_5__7678_ gnd vdd FILL
XFILL_5__11137_ gnd vdd FILL
XFILL_3__15104_ gnd vdd FILL
XFILL_0__9772_ gnd vdd FILL
XFILL_3__8501_ gnd vdd FILL
XFILL_3__12316_ gnd vdd FILL
XFILL112200x3050 gnd vdd FILL
XFILL_4__14655_ gnd vdd FILL
XFILL_0__6984_ gnd vdd FILL
XFILL_3__13296_ gnd vdd FILL
XFILL_3_BUFX2_insert21 gnd vdd FILL
XFILL_2__15834_ gnd vdd FILL
XFILL_4__11867_ gnd vdd FILL
XFILL_1__10707_ gnd vdd FILL
XFILL_3__16084_ gnd vdd FILL
XFILL_1__14475_ gnd vdd FILL
XFILL_0__12136_ gnd vdd FILL
XFILL_3__9481_ gnd vdd FILL
XFILL_5__9417_ gnd vdd FILL
XFILL_1_BUFX2_insert1091 gnd vdd FILL
XFILL_3_BUFX2_insert32 gnd vdd FILL
XFILL_3_BUFX2_insert43 gnd vdd FILL
XFILL_1__11687_ gnd vdd FILL
XFILL_4__13606_ gnd vdd FILL
XFILL_0__8723_ gnd vdd FILL
XFILL_3_BUFX2_insert54 gnd vdd FILL
X_7262_ _7262_/Q _8025_/CLK _7262_/R vdd _7184_/Y gnd vdd DFFSR
XFILL_1__16214_ gnd vdd FILL
XFILL_3__15035_ gnd vdd FILL
XFILL_5__15945_ gnd vdd FILL
XFILL_3_BUFX2_insert65 gnd vdd FILL
XFILL_3__12247_ gnd vdd FILL
XFILL_4__10818_ gnd vdd FILL
XFILL_5__11068_ gnd vdd FILL
XFILL_2__9639_ gnd vdd FILL
XFILL_4__14586_ gnd vdd FILL
XFILL_1__13426_ gnd vdd FILL
XSFILL69240x26050 gnd vdd FILL
XFILL_1__10638_ gnd vdd FILL
XFILL_3_BUFX2_insert76 gnd vdd FILL
XFILL_2__15765_ gnd vdd FILL
XFILL_4__11798_ gnd vdd FILL
XFILL_2__12977_ gnd vdd FILL
XFILL_5__9348_ gnd vdd FILL
XFILL_3_BUFX2_insert87 gnd vdd FILL
XFILL_0__12067_ gnd vdd FILL
X_9001_ _9063_/Q gnd _9001_/Y vdd INVX1
XFILL_5__10019_ gnd vdd FILL
XFILL_3_BUFX2_insert98 gnd vdd FILL
XFILL_4__16325_ gnd vdd FILL
XFILL_0__8654_ gnd vdd FILL
XSFILL29240x42050 gnd vdd FILL
XFILL_4__13537_ gnd vdd FILL
XFILL_3__12178_ gnd vdd FILL
X_7193_ _7191_/Y _7202_/B _7193_/C gnd _7265_/D vdd OAI21X1
XFILL_2__14716_ gnd vdd FILL
XFILL_4__10749_ gnd vdd FILL
XFILL_1__16145_ gnd vdd FILL
XFILL_5__15876_ gnd vdd FILL
XFILL_1__13357_ gnd vdd FILL
XFILL_2__11928_ gnd vdd FILL
XFILL_3__8363_ gnd vdd FILL
XFILL_0__11018_ gnd vdd FILL
XFILL_2__15696_ gnd vdd FILL
XSFILL104440x35050 gnd vdd FILL
XFILL_1__10569_ gnd vdd FILL
XFILL_5__9279_ gnd vdd FILL
XFILL_0__7605_ gnd vdd FILL
XFILL_6__8072_ gnd vdd FILL
XFILL_0__8585_ gnd vdd FILL
XFILL_5__14827_ gnd vdd FILL
XFILL_3__11129_ gnd vdd FILL
XFILL_4__16256_ gnd vdd FILL
XFILL_4__13468_ gnd vdd FILL
XSFILL8680x33050 gnd vdd FILL
XFILL_1__12308_ gnd vdd FILL
XFILL_3__7314_ gnd vdd FILL
XSFILL33720x67050 gnd vdd FILL
XFILL_2__14647_ gnd vdd FILL
XFILL_0__15826_ gnd vdd FILL
XFILL_2__11859_ gnd vdd FILL
XFILL_1__16076_ gnd vdd FILL
XFILL_1__13288_ gnd vdd FILL
XFILL_6_CLKBUF1_insert193 gnd vdd FILL
XFILL_4__15207_ gnd vdd FILL
XFILL_4__12419_ gnd vdd FILL
XFILL_5__14758_ gnd vdd FILL
XFILL_3__7245_ gnd vdd FILL
XFILL_4__16187_ gnd vdd FILL
XFILL_1__15027_ gnd vdd FILL
XFILL_3__15937_ gnd vdd FILL
XFILL_4__13399_ gnd vdd FILL
XFILL_1__12239_ gnd vdd FILL
XSFILL59160x78050 gnd vdd FILL
XFILL_2__14578_ gnd vdd FILL
XFILL_0__15757_ gnd vdd FILL
XFILL_0__12969_ gnd vdd FILL
X_9903_ _9961_/Q gnd _9903_/Y vdd INVX1
XFILL_0__7467_ gnd vdd FILL
XFILL_5__13709_ gnd vdd FILL
XFILL_4__15138_ gnd vdd FILL
XFILL_2__16317_ gnd vdd FILL
XFILL_5__14689_ gnd vdd FILL
XFILL_3__7176_ gnd vdd FILL
XFILL_0__14708_ gnd vdd FILL
XFILL_3__15868_ gnd vdd FILL
XFILL_2__13529_ gnd vdd FILL
XSFILL74200x81050 gnd vdd FILL
XFILL_0__15688_ gnd vdd FILL
XFILL_0__9206_ gnd vdd FILL
X_9834_ _9778_/A _9834_/CLK _7153_/R vdd _9834_/D gnd vdd DFFSR
XFILL_3__14819_ gnd vdd FILL
XFILL_4__15069_ gnd vdd FILL
XFILL_2__16248_ gnd vdd FILL
XFILL_0__14639_ gnd vdd FILL
XFILL_3__15799_ gnd vdd FILL
XSFILL13640x34050 gnd vdd FILL
XFILL_0__9137_ gnd vdd FILL
XFILL_5__16359_ gnd vdd FILL
X_9765_ _9763_/Y _9764_/A _9765_/C gnd _9765_/Y vdd OAI21X1
X_6977_ _7023_/Q gnd _6979_/A vdd INVX1
XFILL_1__15929_ gnd vdd FILL
XFILL_2__16179_ gnd vdd FILL
XFILL_4__6940_ gnd vdd FILL
XFILL_6_BUFX2_insert311 gnd vdd FILL
X_8716_ _8759_/B _6924_/B gnd _8716_/Y vdd NAND2X1
XFILL_0__16309_ gnd vdd FILL
X_9696_ _9696_/Q _9578_/CLK _7793_/R vdd _9622_/Y gnd vdd DFFSR
XFILL_0__8019_ gnd vdd FILL
XFILL_4__6871_ gnd vdd FILL
XFILL_6_BUFX2_insert377 gnd vdd FILL
XFILL_1__8901_ gnd vdd FILL
XFILL_6_BUFX2_insert388 gnd vdd FILL
X_8647_ _8647_/A gnd _8647_/Y vdd INVX1
XFILL_4__8610_ gnd vdd FILL
XFILL_1__9881_ gnd vdd FILL
XSFILL104520x15050 gnd vdd FILL
XFILL_4__9590_ gnd vdd FILL
XSFILL8760x13050 gnd vdd FILL
XFILL_1__8832_ gnd vdd FILL
XSFILL33800x47050 gnd vdd FILL
X_8578_ _8666_/Q gnd _8580_/A vdd INVX1
XFILL_3__9748_ gnd vdd FILL
X_7529_ _7471_/A _9705_/CLK _7914_/R vdd _7473_/Y gnd vdd DFFSR
XFILL_1__8763_ gnd vdd FILL
XSFILL59240x58050 gnd vdd FILL
XFILL_3__9679_ gnd vdd FILL
XFILL_4__8472_ gnd vdd FILL
XFILL_1__7714_ gnd vdd FILL
XFILL_4__7423_ gnd vdd FILL
XFILL111960x57050 gnd vdd FILL
XFILL_1__8694_ gnd vdd FILL
X_11130_ _11120_/Y _11130_/B _11129_/Y gnd _11140_/B vdd OAI21X1
XSFILL13720x14050 gnd vdd FILL
XFILL_4__7354_ gnd vdd FILL
X_11061_ _11059_/Y _11060_/Y _11061_/C gnd _11096_/B vdd OAI21X1
XFILL112040x66050 gnd vdd FILL
XFILL_1__7576_ gnd vdd FILL
XFILL_3_BUFX2_insert234 gnd vdd FILL
XFILL_3_BUFX2_insert245 gnd vdd FILL
X_10012_ _10010_/Y _9993_/A _10012_/C gnd _10082_/D vdd OAI21X1
XFILL_3_BUFX2_insert256 gnd vdd FILL
XFILL_3_BUFX2_insert267 gnd vdd FILL
XSFILL38920x80050 gnd vdd FILL
XFILL_3_BUFX2_insert278 gnd vdd FILL
XFILL_3_BUFX2_insert289 gnd vdd FILL
XFILL_4__9024_ gnd vdd FILL
XFILL_2_BUFX2_insert901 gnd vdd FILL
X_14820_ _13865_/C _7794_/Q _7626_/A _14185_/B gnd _14820_/Y vdd AOI22X1
XFILL_2_BUFX2_insert912 gnd vdd FILL
XFILL_2_BUFX2_insert923 gnd vdd FILL
XFILL_1__9246_ gnd vdd FILL
XFILL_2_BUFX2_insert934 gnd vdd FILL
XFILL_2_BUFX2_insert945 gnd vdd FILL
XFILL_2_BUFX2_insert956 gnd vdd FILL
XFILL_2_BUFX2_insert967 gnd vdd FILL
X_14751_ _8177_/Q gnd _14751_/Y vdd INVX1
X_11963_ _11895_/B _12418_/A gnd _11964_/C vdd NAND2X1
XFILL_2_BUFX2_insert978 gnd vdd FILL
XFILL_2_BUFX2_insert989 gnd vdd FILL
X_13702_ _13702_/A gnd _13704_/B vdd INVX1
XFILL_1__8128_ gnd vdd FILL
X_10914_ _10906_/A _10987_/Q gnd _10915_/A vdd NAND2X1
XFILL_5__6980_ gnd vdd FILL
X_11894_ _11955_/B _12349_/A gnd _11895_/C vdd NAND2X1
X_14682_ _8303_/Q gnd _14683_/A vdd INVX1
XFILL_4__9926_ gnd vdd FILL
XFILL_2__9990_ gnd vdd FILL
X_16421_ _15246_/A _7642_/CLK _7258_/R vdd _16421_/D gnd vdd DFFSR
X_10845_ _10763_/A _9963_/CLK _9963_/R vdd _10845_/D gnd vdd DFFSR
X_13633_ _13632_/Y _13882_/B _13633_/C _13631_/Y gnd _13633_/Y vdd OAI22X1
XFILL_5__10370_ gnd vdd FILL
XFILL_1__8059_ gnd vdd FILL
XFILL_2__10190_ gnd vdd FILL
XBUFX2_insert900 _15072_/Y gnd _15322_/D vdd BUFX2
XFILL_4__9857_ gnd vdd FILL
XFILL_5__8650_ gnd vdd FILL
XFILL_3__10500_ gnd vdd FILL
XFILL_0_BUFX2_insert102 gnd vdd FILL
X_16352_ gnd gnd gnd _16352_/Y vdd NAND2X1
XBUFX2_insert911 _12360_/Y gnd _7558_/B vdd BUFX2
XSFILL23800x79050 gnd vdd FILL
XBUFX2_insert922 _13370_/Y gnd _14878_/C vdd BUFX2
X_10776_ _10792_/B _6936_/B gnd _10777_/C vdd NAND2X1
X_13564_ _9304_/Q gnd _13564_/Y vdd INVX1
XFILL_3__11480_ gnd vdd FILL
XBUFX2_insert933 _12435_/Y gnd _9041_/B vdd BUFX2
XFILL_2__8872_ gnd vdd FILL
XFILL_0__10320_ gnd vdd FILL
XBUFX2_insert944 _12426_/Y gnd _8008_/B vdd BUFX2
XFILL_5__7601_ gnd vdd FILL
XBUFX2_insert955 _13365_/Y gnd _10831_/B vdd BUFX2
X_15303_ _15297_/Y _15298_/Y _15303_/C gnd _15303_/Y vdd NAND3X1
XFILL112120x46050 gnd vdd FILL
XFILL_4__9788_ gnd vdd FILL
X_12515_ vdd _12089_/A gnd _12515_/Y vdd NAND2X1
XFILL_5__12040_ gnd vdd FILL
XFILL_5__8581_ gnd vdd FILL
XBUFX2_insert966 _12417_/Y gnd _8255_/B vdd BUFX2
XFILL_3__10431_ gnd vdd FILL
X_13495_ _14762_/B _7161_/A _8407_/Q _14037_/B gnd _13503_/B vdd AOI22X1
X_16283_ _16283_/A _16283_/B _14402_/C gnd _16283_/Y vdd AOI21X1
XFILL_2__7823_ gnd vdd FILL
XFILL_4__12770_ gnd vdd FILL
XBUFX2_insert977 _16451_/Y gnd _13099_/B vdd BUFX2
XFILL_1__11610_ gnd vdd FILL
XBUFX2_insert988 _13351_/Y gnd _9985_/B vdd BUFX2
XFILL_0__10251_ gnd vdd FILL
XSFILL64040x31050 gnd vdd FILL
XFILL_1__12590_ gnd vdd FILL
XFILL_4__8739_ gnd vdd FILL
XBUFX2_insert999 _14998_/Y gnd _15681_/C vdd BUFX2
X_15234_ _15234_/A _15175_/B _15234_/C gnd _15234_/Y vdd AOI21X1
X_12446_ vdd _11997_/A gnd _12446_/Y vdd NAND2X1
XFILL_3__13150_ gnd vdd FILL
XFILL_4__11721_ gnd vdd FILL
XFILL_3__10362_ gnd vdd FILL
XFILL_2__12900_ gnd vdd FILL
XFILL_2__7754_ gnd vdd FILL
XFILL_1__11541_ gnd vdd FILL
XFILL_2__13880_ gnd vdd FILL
XFILL_0__10182_ gnd vdd FILL
XFILL_5__7463_ gnd vdd FILL
XFILL_3__12101_ gnd vdd FILL
X_12377_ _12371_/A _12600_/A gnd _12378_/C vdd NAND2X1
X_15165_ _15164_/Y _15165_/B gnd _15165_/Y vdd NAND2X1
XFILL_4__14440_ gnd vdd FILL
XFILL_3__13081_ gnd vdd FILL
XFILL_5__13991_ gnd vdd FILL
XFILL_4__11652_ gnd vdd FILL
XFILL_3__10293_ gnd vdd FILL
XFILL_1__14260_ gnd vdd FILL
XFILL_2__12831_ gnd vdd FILL
XFILL_1__11472_ gnd vdd FILL
XFILL_2__7685_ gnd vdd FILL
XFILL_0__14990_ gnd vdd FILL
X_11328_ _11327_/Y gnd _11472_/B vdd INVX1
X_14116_ _15583_/A gnd _14118_/A vdd INVX1
XFILL_5__15730_ gnd vdd FILL
XFILL_3__12032_ gnd vdd FILL
X_15096_ _7161_/A _15177_/B _15095_/Y gnd _15102_/A vdd AOI21X1
XFILL_1__13211_ gnd vdd FILL
XFILL_4__14371_ gnd vdd FILL
XSFILL3640x6050 gnd vdd FILL
XFILL_2__9424_ gnd vdd FILL
XFILL_1__10423_ gnd vdd FILL
XFILL_2__12762_ gnd vdd FILL
XFILL_2__15550_ gnd vdd FILL
XFILL_4__11583_ gnd vdd FILL
XFILL_1__14191_ gnd vdd FILL
XFILL_5__9133_ gnd vdd FILL
XFILL_0__13941_ gnd vdd FILL
XSFILL84200x44050 gnd vdd FILL
XFILL_4__16110_ gnd vdd FILL
XFILL_4__13322_ gnd vdd FILL
XFILL_5__15661_ gnd vdd FILL
X_14047_ _14037_/Y _14047_/B _14046_/Y gnd _14047_/Y vdd NAND3X1
X_11259_ _11045_/Y _11046_/Y gnd _11259_/Y vdd NAND2X1
XFILL_4__10534_ gnd vdd FILL
XFILL_2__14501_ gnd vdd FILL
XFILL_5__12873_ gnd vdd FILL
XFILL_2__11713_ gnd vdd FILL
XFILL_2__9355_ gnd vdd FILL
XFILL_1__13142_ gnd vdd FILL
XFILL_2__15481_ gnd vdd FILL
XFILL_0__13872_ gnd vdd FILL
XFILL_5__14612_ gnd vdd FILL
XFILL_4__16041_ gnd vdd FILL
XFILL_5__11824_ gnd vdd FILL
XFILL_0__8370_ gnd vdd FILL
XSFILL59000x20050 gnd vdd FILL
XFILL_4__13253_ gnd vdd FILL
XFILL_5__15592_ gnd vdd FILL
XFILL_0__15611_ gnd vdd FILL
XFILL_2__11644_ gnd vdd FILL
XFILL_2__14432_ gnd vdd FILL
XFILL_5__8015_ gnd vdd FILL
XFILL_3__13983_ gnd vdd FILL
XFILL_0__12823_ gnd vdd FILL
XFILL_2__9286_ gnd vdd FILL
XFILL_0__7321_ gnd vdd FILL
XFILL_1__10285_ gnd vdd FILL
XFILL_3_BUFX2_insert790 gnd vdd FILL
XFILL_4__12204_ gnd vdd FILL
XFILL_5__14543_ gnd vdd FILL
XFILL_3__15722_ gnd vdd FILL
XFILL_3__7030_ gnd vdd FILL
XSFILL23960x50 gnd vdd FILL
XFILL_5__11755_ gnd vdd FILL
X_15998_ _15998_/A _15997_/Y gnd _15998_/Y vdd NOR2X1
XFILL_1__12024_ gnd vdd FILL
XFILL_4__10396_ gnd vdd FILL
XFILL_2__8237_ gnd vdd FILL
XFILL_2__14363_ gnd vdd FILL
XFILL112200x26050 gnd vdd FILL
XFILL_0__15542_ gnd vdd FILL
XFILL_2__11575_ gnd vdd FILL
XFILL_0__12754_ gnd vdd FILL
XFILL_6__15833_ gnd vdd FILL
XFILL_5__10706_ gnd vdd FILL
X_6900_ _6900_/A gnd memoryWriteData[30] vdd BUFX2
XFILL_0__7252_ gnd vdd FILL
XFILL_5__14474_ gnd vdd FILL
XFILL_4__12135_ gnd vdd FILL
XFILL_2__16102_ gnd vdd FILL
X_14949_ _14947_/Y _13420_/B _14949_/C _14949_/D gnd _14950_/B vdd OAI22X1
XSFILL64120x11050 gnd vdd FILL
XFILL_2__13314_ gnd vdd FILL
XFILL_3__15653_ gnd vdd FILL
XFILL_5__11686_ gnd vdd FILL
XFILL_2__10526_ gnd vdd FILL
X_7880_ _7892_/A _7752_/B gnd _7880_/Y vdd NAND2X1
XFILL_3__12865_ gnd vdd FILL
XFILL_2__14294_ gnd vdd FILL
XFILL_0__11705_ gnd vdd FILL
XFILL_0__15473_ gnd vdd FILL
XFILL_5__16213_ gnd vdd FILL
XFILL_5__13425_ gnd vdd FILL
XFILL_0__7183_ gnd vdd FILL
XFILL_5__10637_ gnd vdd FILL
XFILL_3__14604_ gnd vdd FILL
XFILL_2__13245_ gnd vdd FILL
XFILL_2__7119_ gnd vdd FILL
XFILL_6__12976_ gnd vdd FILL
XFILL_2__16033_ gnd vdd FILL
XFILL_4__12066_ gnd vdd FILL
XSFILL18680x6050 gnd vdd FILL
XFILL_3__11816_ gnd vdd FILL
XFILL_2__8099_ gnd vdd FILL
XFILL_3__15584_ gnd vdd FILL
XFILL_0__14424_ gnd vdd FILL
XFILL_0__11636_ gnd vdd FILL
XFILL_3__8981_ gnd vdd FILL
XFILL_6__7710_ gnd vdd FILL
XFILL_1__13975_ gnd vdd FILL
XFILL_5__8917_ gnd vdd FILL
XSFILL53960x54050 gnd vdd FILL
XFILL_5__16144_ gnd vdd FILL
X_9550_ _9551_/B _8014_/B gnd _9550_/Y vdd NAND2X1
XFILL_5__13356_ gnd vdd FILL
XFILL_6__11927_ gnd vdd FILL
XFILL_4__11017_ gnd vdd FILL
XFILL_5__9897_ gnd vdd FILL
XFILL_6__15695_ gnd vdd FILL
XFILL_3__14535_ gnd vdd FILL
XFILL_5__10568_ gnd vdd FILL
XSFILL109480x83050 gnd vdd FILL
XFILL_1__15714_ gnd vdd FILL
XFILL_3__7932_ gnd vdd FILL
XFILL_3__11747_ gnd vdd FILL
XFILL_0__14355_ gnd vdd FILL
XFILL_2__10388_ gnd vdd FILL
XFILL_5__8848_ gnd vdd FILL
X_8501_ _8555_/Q gnd _8503_/A vdd INVX1
XFILL_5__12307_ gnd vdd FILL
XFILL_0__11567_ gnd vdd FILL
XFILL_6__14646_ gnd vdd FILL
XSFILL28760x30050 gnd vdd FILL
XFILL_5__16075_ gnd vdd FILL
XFILL_5__13287_ gnd vdd FILL
X_9481_ _9535_/A _9993_/B gnd _9482_/C vdd NAND2X1
XFILL_2__12127_ gnd vdd FILL
XFILL_4__15825_ gnd vdd FILL
XFILL_0__13306_ gnd vdd FILL
XFILL_3__14466_ gnd vdd FILL
XSFILL54040x63050 gnd vdd FILL
XFILL_5__10499_ gnd vdd FILL
XFILL_3__7863_ gnd vdd FILL
XFILL_1__15645_ gnd vdd FILL
XFILL_1__12857_ gnd vdd FILL
XFILL_5_BUFX2_insert307 gnd vdd FILL
XFILL_3__11678_ gnd vdd FILL
XFILL_0__10518_ gnd vdd FILL
XFILL_5__15026_ gnd vdd FILL
XFILL_5_BUFX2_insert318 gnd vdd FILL
XFILL_0__14286_ gnd vdd FILL
XFILL_3__16205_ gnd vdd FILL
XFILL_5__8779_ gnd vdd FILL
X_8432_ _8432_/Q _8289_/CLK _7649_/R vdd _8432_/D gnd vdd DFFSR
XFILL_5__12238_ gnd vdd FILL
XFILL_0__11498_ gnd vdd FILL
XFILL_5_BUFX2_insert329 gnd vdd FILL
XFILL_3__9602_ gnd vdd FILL
XFILL_3__13417_ gnd vdd FILL
XBUFX2_insert19 _13443_/Y gnd _14768_/D vdd BUFX2
XFILL_6__11789_ gnd vdd FILL
XFILL_4__15756_ gnd vdd FILL
XFILL_0__16025_ gnd vdd FILL
XFILL_2__12058_ gnd vdd FILL
XFILL_3__10629_ gnd vdd FILL
XFILL_1__11808_ gnd vdd FILL
XFILL_4__12968_ gnd vdd FILL
XFILL_0__13237_ gnd vdd FILL
XFILL_3__14397_ gnd vdd FILL
XFILL_1__15576_ gnd vdd FILL
XFILL_1__12788_ gnd vdd FILL
XFILL_0_BUFX2_insert680 gnd vdd FILL
XFILL_0__10449_ gnd vdd FILL
XFILL_4__14707_ gnd vdd FILL
XFILL_4__11919_ gnd vdd FILL
XFILL_5__12169_ gnd vdd FILL
X_8363_ _8361_/Y _8365_/A _8362_/Y gnd _8423_/D vdd OAI21X1
XSFILL33880x21050 gnd vdd FILL
XFILL_3__16136_ gnd vdd FILL
XFILL_0_BUFX2_insert691 gnd vdd FILL
XFILL_2__11009_ gnd vdd FILL
XFILL_3__9533_ gnd vdd FILL
XFILL_3__13348_ gnd vdd FILL
XFILL_4__15687_ gnd vdd FILL
XFILL_1__14527_ gnd vdd FILL
XFILL_1__11739_ gnd vdd FILL
XFILL_4__12899_ gnd vdd FILL
XFILL_0__13168_ gnd vdd FILL
X_7314_ _7366_/B _7314_/B gnd _7314_/Y vdd NAND2X1
XFILL_6__16247_ gnd vdd FILL
XFILL_4__14638_ gnd vdd FILL
XFILL_6__13459_ gnd vdd FILL
XFILL_0__9755_ gnd vdd FILL
XFILL_0__6967_ gnd vdd FILL
X_8294_ _8230_/A _7282_/CLK _8166_/R vdd _8232_/Y gnd vdd DFFSR
XSFILL48920x43050 gnd vdd FILL
XFILL_2__15817_ gnd vdd FILL
XFILL_3__16067_ gnd vdd FILL
XFILL_3__13279_ gnd vdd FILL
XFILL_1__14458_ gnd vdd FILL
XFILL_3__9464_ gnd vdd FILL
XFILL_0__12119_ gnd vdd FILL
XFILL_0__8706_ gnd vdd FILL
XFILL_0__13099_ gnd vdd FILL
X_7245_ _7245_/A gnd _7245_/Y vdd INVX1
XFILL_5__15928_ gnd vdd FILL
XFILL_3__15018_ gnd vdd FILL
XFILL_4__14569_ gnd vdd FILL
XFILL_1__13409_ gnd vdd FILL
XFILL_0__6898_ gnd vdd FILL
XFILL_2__15748_ gnd vdd FILL
XFILL_3__9395_ gnd vdd FILL
XFILL_1__14389_ gnd vdd FILL
XSFILL49000x52050 gnd vdd FILL
XFILL_4__16308_ gnd vdd FILL
XSFILL13640x29050 gnd vdd FILL
XFILL_1__7430_ gnd vdd FILL
XFILL_0__8637_ gnd vdd FILL
X_7176_ _7260_/Q gnd _7178_/A vdd INVX1
XFILL_5__15859_ gnd vdd FILL
XFILL_3__8346_ gnd vdd FILL
XFILL_1__16128_ gnd vdd FILL
XFILL_2__15679_ gnd vdd FILL
XFILL_4__16239_ gnd vdd FILL
XFILL_1__7361_ gnd vdd FILL
XFILL_0__8568_ gnd vdd FILL
XFILL_4__7070_ gnd vdd FILL
XFILL_1__16059_ gnd vdd FILL
XFILL_0__15809_ gnd vdd FILL
XFILL_3__8277_ gnd vdd FILL
XSFILL28840x10050 gnd vdd FILL
XFILL_1__9100_ gnd vdd FILL
XSFILL29320x17050 gnd vdd FILL
XSFILL54120x43050 gnd vdd FILL
XFILL_1__7292_ gnd vdd FILL
XFILL_0__8499_ gnd vdd FILL
XFILL_3__7228_ gnd vdd FILL
XSFILL33800x8050 gnd vdd FILL
XFILL_1__9031_ gnd vdd FILL
XFILL_3__7159_ gnd vdd FILL
XFILL_1_BUFX2_insert908 gnd vdd FILL
XFILL_1_BUFX2_insert919 gnd vdd FILL
X_9817_ _9817_/Q _9817_/CLK _8942_/R vdd _9817_/D gnd vdd DFFSR
XSFILL33400x44050 gnd vdd FILL
XFILL_4__7972_ gnd vdd FILL
XFILL_6__8888_ gnd vdd FILL
X_9748_ _9748_/A gnd _9750_/A vdd INVX1
XFILL_4__6923_ gnd vdd FILL
XSFILL39000x2050 gnd vdd FILL
X_10630_ _10619_/B _6918_/B gnd _10631_/C vdd NAND2X1
XFILL_6__7839_ gnd vdd FILL
XBUFX2_insert229 _12432_/Y gnd _8014_/B vdd BUFX2
XFILL_1__9933_ gnd vdd FILL
X_9679_ _9677_/Y _9639_/A _9678_/Y gnd _9715_/D vdd OAI21X1
XFILL_4__9642_ gnd vdd FILL
XFILL_4__6854_ gnd vdd FILL
X_10561_ _16072_/A gnd _10563_/A vdd INVX1
XSFILL23880x53050 gnd vdd FILL
XFILL_1__9864_ gnd vdd FILL
XFILL_5_BUFX2_insert830 gnd vdd FILL
X_12300_ _12216_/B _12340_/B _12300_/C gnd _12300_/Y vdd NAND3X1
XFILL_5_BUFX2_insert841 gnd vdd FILL
XFILL_5_CLKBUF1_insert119 gnd vdd FILL
X_13280_ _13297_/C _13280_/B gnd _13280_/Y vdd NOR2X1
XFILL_5_BUFX2_insert852 gnd vdd FILL
XFILL_5_BUFX2_insert863 gnd vdd FILL
X_10492_ _13552_/A gnd _10494_/A vdd INVX1
XSFILL38920x75050 gnd vdd FILL
XFILL_5_BUFX2_insert874 gnd vdd FILL
XFILL112440x82050 gnd vdd FILL
XFILL_4__8524_ gnd vdd FILL
XFILL_5_BUFX2_insert885 gnd vdd FILL
XFILL_1__9795_ gnd vdd FILL
XFILL_5_BUFX2_insert896 gnd vdd FILL
XBUFX2_insert1060 _15051_/Y gnd _16148_/C vdd BUFX2
X_12231_ _12239_/A gnd _12239_/C gnd _12231_/Y vdd NAND3X1
XSFILL54200x23050 gnd vdd FILL
XBUFX2_insert1071 _13327_/Y gnd _8845_/B vdd BUFX2
XFILL_1__8746_ gnd vdd FILL
XBUFX2_insert1093 rst gnd BUFX2_insert520/A vdd BUFX2
XFILL_4__8455_ gnd vdd FILL
X_12162_ _12162_/A _12137_/A _12162_/C gnd _12162_/Y vdd OAI21X1
XFILL_2__7470_ gnd vdd FILL
X_11113_ _12177_/Y gnd _11113_/Y vdd INVX1
XFILL_4__8386_ gnd vdd FILL
X_12093_ _12093_/A _12093_/B _12073_/C gnd gnd _12093_/Y vdd AOI22X1
XFILL_1__7628_ gnd vdd FILL
XSFILL18840x42050 gnd vdd FILL
XFILL_4__7337_ gnd vdd FILL
X_15921_ _7787_/Q gnd _15922_/D vdd INVX1
X_11044_ _11044_/A _11641_/C gnd _11048_/A vdd NOR2X1
XFILL_2__9140_ gnd vdd FILL
XSFILL59720x54050 gnd vdd FILL
XFILL_1__7559_ gnd vdd FILL
XFILL_4__10250_ gnd vdd FILL
XSFILL99320x40050 gnd vdd FILL
X_15852_ _15825_/Y _15852_/B _15651_/C gnd _12881_/B vdd AOI21X1
XSFILL28680x1050 gnd vdd FILL
XFILL_4__9007_ gnd vdd FILL
XFILL_2_BUFX2_insert720 gnd vdd FILL
XFILL_3__10980_ gnd vdd FILL
XFILL_2_BUFX2_insert731 gnd vdd FILL
XSFILL68840x6050 gnd vdd FILL
X_14803_ _13621_/B _10354_/Q _9162_/A _14868_/D gnd _14803_/Y vdd AOI22X1
XFILL_2_BUFX2_insert742 gnd vdd FILL
XFILL_5__11540_ gnd vdd FILL
XFILL_4__7199_ gnd vdd FILL
XFILL_1__9229_ gnd vdd FILL
XFILL_4__10181_ gnd vdd FILL
X_15783_ _15782_/Y _15025_/B _16018_/C _15781_/Y gnd _15784_/A vdd OAI22X1
XFILL_2_BUFX2_insert753 gnd vdd FILL
XFILL_2_BUFX2_insert764 gnd vdd FILL
X_12995_ _12993_/Y vdd _12995_/C gnd _13061_/D vdd OAI21X1
XFILL_2__11360_ gnd vdd FILL
XFILL_2_BUFX2_insert775 gnd vdd FILL
XSFILL64040x26050 gnd vdd FILL
XFILL_2_BUFX2_insert786 gnd vdd FILL
X_14734_ _14734_/A gnd _16104_/B vdd INVX1
X_11946_ _11946_/A _11895_/B _11946_/C gnd _6857_/A vdd OAI21X1
XFILL_2__10311_ gnd vdd FILL
XFILL_5__11471_ gnd vdd FILL
XFILL_2_BUFX2_insert797 gnd vdd FILL
XFILL_3__12650_ gnd vdd FILL
XFILL_2__11291_ gnd vdd FILL
XFILL_5__13210_ gnd vdd FILL
XFILL_5__9751_ gnd vdd FILL
XFILL_0__12470_ gnd vdd FILL
XFILL_5__10422_ gnd vdd FILL
XFILL_5__6963_ gnd vdd FILL
XFILL_5__14190_ gnd vdd FILL
XFILL_2__13030_ gnd vdd FILL
XFILL_3__11601_ gnd vdd FILL
X_14665_ _14725_/A _14665_/B _16062_/C _14752_/C gnd _14665_/Y vdd OAI22X1
XFILL_4__13940_ gnd vdd FILL
X_11877_ _11877_/A _11874_/B _11876_/Y gnd _13220_/A vdd OAI21X1
XFILL_2__10242_ gnd vdd FILL
XFILL_4__9909_ gnd vdd FILL
XFILL_3__12581_ gnd vdd FILL
XFILL_1__13760_ gnd vdd FILL
XFILL_5__8702_ gnd vdd FILL
XSFILL114840x14050 gnd vdd FILL
XFILL_0__11421_ gnd vdd FILL
XFILL_1__10972_ gnd vdd FILL
X_16404_ _16402_/Y gnd _16404_/C gnd _16404_/Y vdd OAI21X1
X_13616_ _7295_/A gnd _13616_/Y vdd INVX1
XFILL_5__13141_ gnd vdd FILL
XFILL_6__11712_ gnd vdd FILL
XFILL_5__9682_ gnd vdd FILL
X_10828_ _10826_/Y _10762_/B _10828_/C gnd _10828_/Y vdd OAI21X1
XFILL_5__6894_ gnd vdd FILL
XFILL_3__14320_ gnd vdd FILL
XFILL_6__15480_ gnd vdd FILL
X_14596_ _14596_/A _14596_/B gnd _14597_/A vdd NOR2X1
XFILL_4__13871_ gnd vdd FILL
XFILL_1__12711_ gnd vdd FILL
XFILL_3__11532_ gnd vdd FILL
XFILL_2__10173_ gnd vdd FILL
XFILL_0__14140_ gnd vdd FILL
XFILL_5__8633_ gnd vdd FILL
XBUFX2_insert730 _12411_/Y gnd _9017_/B vdd BUFX2
XFILL_0__11352_ gnd vdd FILL
XFILL_1__13691_ gnd vdd FILL
X_16335_ _16335_/A gnd _16335_/C gnd _16421_/D vdd OAI21X1
XSFILL84200x39050 gnd vdd FILL
XBUFX2_insert741 _12402_/Y gnd _6960_/B vdd BUFX2
XFILL_4__15610_ gnd vdd FILL
XFILL_6__14431_ gnd vdd FILL
XBUFX2_insert752 _13344_/Y gnd _9741_/B vdd BUFX2
X_13547_ _14030_/A _15141_/D _13461_/C _15157_/C gnd _13547_/Y vdd OAI22X1
XFILL_3__14251_ gnd vdd FILL
XBUFX2_insert763 _13412_/Y gnd _14489_/C vdd BUFX2
XFILL_5__10284_ gnd vdd FILL
X_10759_ _10759_/A _10809_/A _10759_/C gnd _10759_/Y vdd OAI21X1
XFILL_1__15430_ gnd vdd FILL
XSFILL94360x83050 gnd vdd FILL
XBUFX2_insert774 _13301_/Y gnd _7887_/B vdd BUFX2
XFILL_0__10303_ gnd vdd FILL
XFILL_1__12642_ gnd vdd FILL
XFILL_2__8855_ gnd vdd FILL
XFILL_3__11463_ gnd vdd FILL
XFILL_2__14981_ gnd vdd FILL
XFILL_0__14071_ gnd vdd FILL
XFILL_5__12023_ gnd vdd FILL
XBUFX2_insert785 _13486_/Y gnd _14481_/C vdd BUFX2
XFILL_0__11283_ gnd vdd FILL
XFILL_4__15541_ gnd vdd FILL
XFILL_6__11574_ gnd vdd FILL
XBUFX2_insert796 _13334_/Y gnd _9339_/B vdd BUFX2
X_16266_ _16266_/A _16265_/Y _16264_/Y gnd _16267_/B vdd NOR3X1
XFILL_0__7870_ gnd vdd FILL
XFILL_4__12753_ gnd vdd FILL
XFILL_3__10414_ gnd vdd FILL
XFILL_2__7806_ gnd vdd FILL
X_13478_ _8185_/A gnd _13479_/A vdd INVX1
XFILL_0__13022_ gnd vdd FILL
XFILL_3__14182_ gnd vdd FILL
XFILL_1__15361_ gnd vdd FILL
XFILL_3__11394_ gnd vdd FILL
XFILL_2__13932_ gnd vdd FILL
XFILL_1__12573_ gnd vdd FILL
XFILL_0__10234_ gnd vdd FILL
XFILL_2__8786_ gnd vdd FILL
XSFILL99400x20050 gnd vdd FILL
X_15217_ _15203_/B gnd _15892_/B vdd INVX4
X_12429_ _12427_/Y _12422_/A _12429_/C gnd _12429_/Y vdd OAI21X1
XFILL_5__8495_ gnd vdd FILL
XFILL_4__11704_ gnd vdd FILL
XFILL_6__14293_ gnd vdd FILL
X_16197_ _10098_/Q gnd _16199_/D vdd INVX1
XFILL_3__13133_ gnd vdd FILL
XFILL_4__15472_ gnd vdd FILL
XFILL111720x14050 gnd vdd FILL
XFILL_1__14312_ gnd vdd FILL
XFILL_2__7737_ gnd vdd FILL
XFILL_1__11524_ gnd vdd FILL
XFILL_2__13863_ gnd vdd FILL
XFILL_1__15292_ gnd vdd FILL
XFILL_6__13244_ gnd vdd FILL
XFILL_0__10165_ gnd vdd FILL
XFILL_6__16032_ gnd vdd FILL
XFILL_5__7446_ gnd vdd FILL
XFILL_0__9540_ gnd vdd FILL
X_15148_ _6908_/A gnd _15149_/D vdd INVX1
XFILL_4__14423_ gnd vdd FILL
XFILL_1_CLKBUF1_insert190 gnd vdd FILL
XFILL_4__11635_ gnd vdd FILL
XFILL_2__15602_ gnd vdd FILL
XFILL_3__10276_ gnd vdd FILL
XFILL_1__14243_ gnd vdd FILL
XFILL_5__13974_ gnd vdd FILL
XFILL_2_BUFX2_insert0 gnd vdd FILL
XFILL_1__11455_ gnd vdd FILL
XFILL_2__13794_ gnd vdd FILL
XSFILL74280x50050 gnd vdd FILL
XFILL_0__14973_ gnd vdd FILL
XFILL_5__15713_ gnd vdd FILL
X_7030_ _7030_/A gnd _7030_/Y vdd INVX1
XFILL_5__7377_ gnd vdd FILL
XFILL_0__9471_ gnd vdd FILL
XFILL_2__9407_ gnd vdd FILL
XFILL_3__12015_ gnd vdd FILL
XFILL_3__8200_ gnd vdd FILL
XFILL_4__14354_ gnd vdd FILL
X_15079_ _16314_/D gnd _15079_/Y vdd INVX1
XFILL_1__10406_ gnd vdd FILL
XFILL_2__15533_ gnd vdd FILL
XFILL_4__11566_ gnd vdd FILL
XFILL_2__12745_ gnd vdd FILL
XFILL_1__14174_ gnd vdd FILL
XFILL_5__9116_ gnd vdd FILL
XFILL_0__13924_ gnd vdd FILL
XFILL_6__12126_ gnd vdd FILL
XFILL_1__11386_ gnd vdd FILL
XFILL_2__7599_ gnd vdd FILL
XFILL_4__13305_ gnd vdd FILL
XSFILL89320x72050 gnd vdd FILL
XSFILL53960x49050 gnd vdd FILL
XFILL_5__15644_ gnd vdd FILL
XFILL_5__12856_ gnd vdd FILL
XFILL_4__10517_ gnd vdd FILL
XFILL_1__13125_ gnd vdd FILL
XFILL_3__8131_ gnd vdd FILL
XSFILL3560x13050 gnd vdd FILL
XFILL_2__9338_ gnd vdd FILL
XFILL_4__14285_ gnd vdd FILL
XSFILL109480x78050 gnd vdd FILL
XFILL_2__15464_ gnd vdd FILL
XFILL_4__11497_ gnd vdd FILL
XFILL_0__13855_ gnd vdd FILL
XFILL_4__16024_ gnd vdd FILL
XFILL_0__8353_ gnd vdd FILL
XFILL_5__11807_ gnd vdd FILL
XFILL_4__13236_ gnd vdd FILL
XFILL_5__12787_ gnd vdd FILL
XFILL_3__8062_ gnd vdd FILL
XFILL_4__10448_ gnd vdd FILL
X_8981_ _9011_/A _7445_/B gnd _8981_/Y vdd NAND2X1
XFILL_5__15575_ gnd vdd FILL
XFILL_2__14415_ gnd vdd FILL
XFILL_2__9269_ gnd vdd FILL
XSFILL54040x58050 gnd vdd FILL
XFILL_2__11627_ gnd vdd FILL
XFILL_3__13966_ gnd vdd FILL
XFILL_2__15395_ gnd vdd FILL
XFILL_0__7304_ gnd vdd FILL
XFILL_1__10268_ gnd vdd FILL
XFILL_6__9860_ gnd vdd FILL
XFILL_0__13786_ gnd vdd FILL
XSFILL94440x63050 gnd vdd FILL
XFILL_3__15705_ gnd vdd FILL
XFILL_5__14526_ gnd vdd FILL
X_7932_ _8024_/Q gnd _7934_/A vdd INVX1
XFILL_5__11738_ gnd vdd FILL
XFILL_0__10998_ gnd vdd FILL
XFILL_4__13167_ gnd vdd FILL
XFILL_1__12007_ gnd vdd FILL
XFILL_3__12917_ gnd vdd FILL
XFILL_4__10379_ gnd vdd FILL
XFILL_0__15525_ gnd vdd FILL
XFILL_2__14346_ gnd vdd FILL
XFILL_2__11558_ gnd vdd FILL
XFILL_0__12737_ gnd vdd FILL
XFILL_3__13897_ gnd vdd FILL
XFILL_0__7235_ gnd vdd FILL
XFILL_5__14457_ gnd vdd FILL
XFILL_4__12118_ gnd vdd FILL
X_7863_ _7861_/Y _7887_/B _7863_/C gnd _7915_/D vdd OAI21X1
XFILL_2__10509_ gnd vdd FILL
XFILL_3__15636_ gnd vdd FILL
XFILL_5__11669_ gnd vdd FILL
XSFILL33880x16050 gnd vdd FILL
XFILL_3__12848_ gnd vdd FILL
XFILL_4__13098_ gnd vdd FILL
XFILL_2__11489_ gnd vdd FILL
XFILL_0__15456_ gnd vdd FILL
XFILL_2__14277_ gnd vdd FILL
XFILL_5__13408_ gnd vdd FILL
X_9602_ _9602_/A gnd _9602_/Y vdd INVX1
XFILL_0__7166_ gnd vdd FILL
XFILL_2__16016_ gnd vdd FILL
XFILL_4__12049_ gnd vdd FILL
XFILL_5__14388_ gnd vdd FILL
XFILL_2__13228_ gnd vdd FILL
X_7794_ _7794_/Q _7662_/CLK _8166_/R vdd _7756_/Y gnd vdd DFFSR
XFILL_3__15567_ gnd vdd FILL
XSFILL48920x38050 gnd vdd FILL
XFILL_0__14407_ gnd vdd FILL
XFILL_3__12779_ gnd vdd FILL
XSFILL18680x77050 gnd vdd FILL
XFILL_3__8964_ gnd vdd FILL
XSFILL104440x9050 gnd vdd FILL
XFILL_0__11619_ gnd vdd FILL
XFILL_0__15387_ gnd vdd FILL
XFILL_6_BUFX2_insert91 gnd vdd FILL
XFILL_1__13958_ gnd vdd FILL
XFILL_5__13339_ gnd vdd FILL
X_9533_ _9533_/A _9533_/B _9532_/Y gnd _9533_/Y vdd OAI21X1
XFILL_0__12599_ gnd vdd FILL
XFILL_5__16127_ gnd vdd FILL
XFILL_3__14518_ gnd vdd FILL
XFILL_0__7097_ gnd vdd FILL
XFILL_2__13159_ gnd vdd FILL
XFILL_3__15498_ gnd vdd FILL
XFILL_1__12909_ gnd vdd FILL
XFILL_0__14338_ gnd vdd FILL
XFILL_3__8895_ gnd vdd FILL
XFILL_5_BUFX2_insert104 gnd vdd FILL
XSFILL48520x40050 gnd vdd FILL
XSFILL49000x47050 gnd vdd FILL
XFILL_5__16058_ gnd vdd FILL
XFILL_1__13889_ gnd vdd FILL
X_9464_ _9464_/A _9535_/A _9463_/Y gnd _9558_/D vdd OAI21X1
XFILL_4__15808_ gnd vdd FILL
XFILL_1__6930_ gnd vdd FILL
XFILL_3__14449_ gnd vdd FILL
XFILL_3__7846_ gnd vdd FILL
XFILL_1__15628_ gnd vdd FILL
XFILL_5__15009_ gnd vdd FILL
XFILL_0__14269_ gnd vdd FILL
XFILL_6__7555_ gnd vdd FILL
XSFILL80040x3050 gnd vdd FILL
X_8415_ _8415_/Q _9568_/CLK _8431_/R vdd _8415_/D gnd vdd DFFSR
XFILL_0__16008_ gnd vdd FILL
XFILL_1__6861_ gnd vdd FILL
X_9395_ _9401_/A _9907_/B gnd _9395_/Y vdd NAND2X1
XFILL_4__15739_ gnd vdd FILL
XFILL_1__15559_ gnd vdd FILL
XFILL_0__9807_ gnd vdd FILL
XFILL_1__8600_ gnd vdd FILL
XSFILL53640x31050 gnd vdd FILL
XFILL_4_BUFX2_insert804 gnd vdd FILL
XFILL_3__16119_ gnd vdd FILL
X_8346_ _8418_/Q gnd _8346_/Y vdd INVX1
XFILL_4_BUFX2_insert815 gnd vdd FILL
XFILL_3__9516_ gnd vdd FILL
XFILL_4_BUFX2_insert826 gnd vdd FILL
XFILL_0__7999_ gnd vdd FILL
XFILL_4_BUFX2_insert837 gnd vdd FILL
XFILL_4_BUFX2_insert848 gnd vdd FILL
XSFILL64280x82050 gnd vdd FILL
XFILL_0__9738_ gnd vdd FILL
XFILL_1__8531_ gnd vdd FILL
XFILL_4_BUFX2_insert859 gnd vdd FILL
XSFILL89800x50 gnd vdd FILL
X_8277_ _8275_/Y _8237_/A _8277_/C gnd _8309_/D vdd OAI21X1
XFILL_4__8240_ gnd vdd FILL
XFILL_6__9156_ gnd vdd FILL
X_7228_ _7168_/A _8636_/B gnd _7229_/C vdd NAND2X1
XFILL_1__8462_ gnd vdd FILL
XFILL_0__9669_ gnd vdd FILL
XSFILL83640x8050 gnd vdd FILL
XFILL_3__9378_ gnd vdd FILL
XSFILL18760x57050 gnd vdd FILL
X_7159_ _6903_/A _7207_/A gnd _7160_/C vdd NAND2X1
XFILL_1__8393_ gnd vdd FILL
XSFILL8600x67050 gnd vdd FILL
XFILL_3__8329_ gnd vdd FILL
XFILL_4__7122_ gnd vdd FILL
XFILL_1__7344_ gnd vdd FILL
XFILL_4__7053_ gnd vdd FILL
XSFILL43960x9050 gnd vdd FILL
XSFILL23880x48050 gnd vdd FILL
XFILL_5_BUFX2_insert4 gnd vdd FILL
X_11800_ _11800_/A gnd _12009_/A vdd INVX1
XFILL_1__9014_ gnd vdd FILL
X_12780_ _12777_/A memoryOutData[28] gnd _12781_/C vdd NAND2X1
XFILL_1_BUFX2_insert705 gnd vdd FILL
XFILL_6__9989_ gnd vdd FILL
XFILL_1_BUFX2_insert716 gnd vdd FILL
XFILL_1_BUFX2_insert727 gnd vdd FILL
XFILL112440x77050 gnd vdd FILL
XFILL_1_BUFX2_insert738 gnd vdd FILL
XSFILL54200x18050 gnd vdd FILL
X_11731_ _11729_/Y _11731_/B _11751_/C gnd _11741_/B vdd OAI21X1
XFILL_1_BUFX2_insert749 gnd vdd FILL
XFILL_4__7955_ gnd vdd FILL
XSFILL79160x22050 gnd vdd FILL
X_14450_ _14450_/A _14450_/B _14402_/C gnd _13012_/B vdd AOI21X1
X_11662_ _11086_/Y _11639_/Y gnd _11684_/B vdd NOR2X1
XFILL_2__6970_ gnd vdd FILL
XFILL_4__6906_ gnd vdd FILL
X_13401_ _13374_/Y _13401_/B _13401_/C gnd _13401_/Y vdd NAND3X1
XFILL_4__7886_ gnd vdd FILL
X_10613_ _16305_/A _9205_/CLK _7285_/R vdd _10581_/Y gnd vdd DFFSR
XFILL_1__9916_ gnd vdd FILL
X_14381_ _8169_/Q gnd _14383_/A vdd INVX1
X_11593_ _11289_/C _11449_/Y _11451_/B gnd _11593_/Y vdd AOI21X1
XFILL_4__9625_ gnd vdd FILL
XFILL_4__6837_ gnd vdd FILL
X_16120_ _15369_/A _16119_/Y _16118_/Y _15369_/D gnd _16121_/B vdd OAI22X1
XSFILL18840x37050 gnd vdd FILL
X_13332_ _13235_/C _13218_/A gnd _13332_/Y vdd NAND2X1
X_10544_ _10500_/B _7856_/B gnd _10544_/Y vdd NAND2X1
XSFILL84280x13050 gnd vdd FILL
XFILL_2__8640_ gnd vdd FILL
XFILL_5_BUFX2_insert660 gnd vdd FILL
XFILL_1__9847_ gnd vdd FILL
XFILL_5_BUFX2_insert671 gnd vdd FILL
XSFILL49640x9050 gnd vdd FILL
XFILL_4__9556_ gnd vdd FILL
XFILL_5_BUFX2_insert682 gnd vdd FILL
X_16051_ _9199_/Q gnd _16051_/Y vdd INVX1
X_10475_ _10475_/Q _9195_/CLK _7915_/R vdd _10475_/D gnd vdd DFFSR
X_13263_ _13278_/B _13263_/B _13263_/C gnd _13263_/Y vdd NAND3X1
XFILL_5_BUFX2_insert693 gnd vdd FILL
XSFILL99320x35050 gnd vdd FILL
XSFILL69080x74050 gnd vdd FILL
XFILL_4__8507_ gnd vdd FILL
XFILL_5__7300_ gnd vdd FILL
XFILL_2__8571_ gnd vdd FILL
XFILL_1__9778_ gnd vdd FILL
X_15002_ _16293_/A _7030_/A _15002_/C _15916_/B gnd _15008_/A vdd AOI22X1
XFILL_6__10310_ gnd vdd FILL
XFILL_4__9487_ gnd vdd FILL
X_12214_ _12216_/B _12695_/A _12300_/C gnd _12214_/Y vdd NAND3X1
X_13194_ _13194_/Q _13201_/CLK _13201_/R vdd _13194_/D gnd vdd DFFSR
XFILL_3__10130_ gnd vdd FILL
XFILL_1__8729_ gnd vdd FILL
XFILL_5__7231_ gnd vdd FILL
XFILL_4__8438_ gnd vdd FILL
X_12145_ _13185_/Q gnd _12147_/A vdd INVX1
XFILL_4__11420_ gnd vdd FILL
XFILL_5__10971_ gnd vdd FILL
XFILL_3__10061_ gnd vdd FILL
XFILL_2__7453_ gnd vdd FILL
XFILL_1__11240_ gnd vdd FILL
XFILL_2__10791_ gnd vdd FILL
XSFILL109320x20050 gnd vdd FILL
XFILL_5__12710_ gnd vdd FILL
XFILL_0__11970_ gnd vdd FILL
XFILL_4__8369_ gnd vdd FILL
XFILL_5__7162_ gnd vdd FILL
X_12076_ _12072_/A _11884_/A _12072_/C gnd _12078_/B vdd NAND3X1
XFILL_5__13690_ gnd vdd FILL
XFILL_4__11351_ gnd vdd FILL
XFILL_2__12530_ gnd vdd FILL
XFILL_0__10921_ gnd vdd FILL
XFILL_1__11171_ gnd vdd FILL
X_15904_ _15383_/A _7605_/A _7531_/Q _15383_/D gnd _15909_/B vdd AOI22X1
XSFILL3480x28050 gnd vdd FILL
X_11027_ _11021_/Y _11027_/B gnd _11028_/C vdd OR2X2
XFILL_4__10302_ gnd vdd FILL
XFILL_5__7093_ gnd vdd FILL
XFILL_5__12641_ gnd vdd FILL
XFILL_3__13820_ gnd vdd FILL
XFILL_2__9123_ gnd vdd FILL
XFILL_4__14070_ gnd vdd FILL
XFILL_1__10122_ gnd vdd FILL
XFILL_2__12461_ gnd vdd FILL
XFILL_4__11282_ gnd vdd FILL
XFILL_0__13640_ gnd vdd FILL
XSFILL114440x11050 gnd vdd FILL
XFILL_4__13021_ gnd vdd FILL
XFILL_5__15360_ gnd vdd FILL
X_15835_ _9449_/Q _15945_/C _16148_/C gnd _15836_/C vdd NAND3X1
XFILL_2__14200_ gnd vdd FILL
XFILL_5__12572_ gnd vdd FILL
XFILL_0_BUFX2_insert1007 gnd vdd FILL
XFILL_4__10233_ gnd vdd FILL
XFILL_2__11412_ gnd vdd FILL
XFILL_3__13751_ gnd vdd FILL
XFILL_2_BUFX2_insert550 gnd vdd FILL
XFILL_2__15180_ gnd vdd FILL
XFILL_2__12392_ gnd vdd FILL
XFILL_3__10963_ gnd vdd FILL
XFILL_0_BUFX2_insert1018 gnd vdd FILL
XFILL_1__14930_ gnd vdd FILL
XFILL_1__10053_ gnd vdd FILL
XFILL_2_BUFX2_insert561 gnd vdd FILL
XFILL_0_BUFX2_insert1029 gnd vdd FILL
XFILL_5__14311_ gnd vdd FILL
XFILL_0__13571_ gnd vdd FILL
XFILL_2_BUFX2_insert572 gnd vdd FILL
XFILL_5__11523_ gnd vdd FILL
XFILL_0__10783_ gnd vdd FILL
XFILL_2_BUFX2_insert583 gnd vdd FILL
XFILL_3__12702_ gnd vdd FILL
XFILL_2__8005_ gnd vdd FILL
X_15766_ _16306_/A _15766_/B _15558_/D _14307_/Y gnd _15767_/B vdd OAI22X1
XFILL_5__15291_ gnd vdd FILL
XFILL_2_BUFX2_insert594 gnd vdd FILL
XFILL_2__14131_ gnd vdd FILL
XFILL_0__15310_ gnd vdd FILL
XFILL_4__10164_ gnd vdd FILL
X_12978_ _6879_/A gnd _12978_/Y vdd INVX1
XFILL_2__11343_ gnd vdd FILL
XFILL_3__13682_ gnd vdd FILL
XFILL_5__9803_ gnd vdd FILL
XFILL_0__12522_ gnd vdd FILL
XFILL_1__14861_ gnd vdd FILL
XSFILL69160x54050 gnd vdd FILL
XFILL_0__16290_ gnd vdd FILL
XFILL_3__10894_ gnd vdd FILL
XSFILL99400x15050 gnd vdd FILL
XFILL_5__14242_ gnd vdd FILL
X_14717_ _9584_/Q gnd _14718_/A vdd INVX1
XFILL_5__7995_ gnd vdd FILL
X_11929_ _11929_/A gnd _11931_/A vdd INVX1
XFILL_5__11454_ gnd vdd FILL
XFILL_3__15421_ gnd vdd FILL
XFILL_3__12633_ gnd vdd FILL
X_15697_ _15697_/A _15696_/Y _15694_/Y gnd _15697_/Y vdd NAND3X1
XFILL_2__14062_ gnd vdd FILL
XFILL_4__14972_ gnd vdd FILL
XFILL_1__13812_ gnd vdd FILL
XFILL_0__15241_ gnd vdd FILL
XFILL_2__11274_ gnd vdd FILL
XFILL_0__12453_ gnd vdd FILL
XFILL_5__9734_ gnd vdd FILL
XFILL_5__10405_ gnd vdd FILL
XFILL_1__14792_ gnd vdd FILL
XFILL_5__6946_ gnd vdd FILL
XFILL_5__14173_ gnd vdd FILL
XFILL_4__13923_ gnd vdd FILL
X_14648_ _7361_/A gnd _14650_/A vdd INVX1
XFILL_2__13013_ gnd vdd FILL
XFILL_3__15352_ gnd vdd FILL
XFILL_5__11385_ gnd vdd FILL
XFILL_0__11404_ gnd vdd FILL
XFILL_1__10955_ gnd vdd FILL
XFILL_1__13743_ gnd vdd FILL
XFILL_0__15172_ gnd vdd FILL
XFILL_5__13124_ gnd vdd FILL
XFILL_0__12384_ gnd vdd FILL
XFILL_5__9665_ gnd vdd FILL
XFILL_5__6877_ gnd vdd FILL
XSFILL74280x45050 gnd vdd FILL
XFILL_3__14303_ gnd vdd FILL
XFILL_4__13854_ gnd vdd FILL
X_14579_ _14579_/A _14575_/Y gnd _14579_/Y vdd NOR2X1
XFILL_0__8971_ gnd vdd FILL
XFILL_2__8907_ gnd vdd FILL
XFILL_3__7700_ gnd vdd FILL
XFILL_3__11515_ gnd vdd FILL
XSFILL89880x24050 gnd vdd FILL
XFILL_0__14123_ gnd vdd FILL
XFILL_2__10156_ gnd vdd FILL
XFILL_3__15283_ gnd vdd FILL
XFILL_5__8616_ gnd vdd FILL
XFILL_1__13674_ gnd vdd FILL
XFILL_3__12495_ gnd vdd FILL
XFILL_2__9887_ gnd vdd FILL
XBUFX2_insert560 BUFX2_insert520/A gnd _7391_/R vdd BUFX2
XFILL_0__11335_ gnd vdd FILL
XFILL_1__10886_ gnd vdd FILL
X_16318_ _16317_/Y _16312_/Y gnd _16318_/Y vdd NAND2X1
XBUFX2_insert571 BUFX2_insert494/A gnd _7153_/R vdd BUFX2
XBUFX2_insert582 BUFX2_insert496/A gnd _9959_/R vdd BUFX2
XSFILL89320x67050 gnd vdd FILL
XFILL_5__9596_ gnd vdd FILL
XSFILL49080x21050 gnd vdd FILL
XFILL_3__14234_ gnd vdd FILL
XBUFX2_insert593 BUFX2_insert600/A gnd _9313_/R vdd BUFX2
XFILL_5__10267_ gnd vdd FILL
XFILL_3__7631_ gnd vdd FILL
XFILL_1__15413_ gnd vdd FILL
XFILL_1__12625_ gnd vdd FILL
XFILL_4__13785_ gnd vdd FILL
XFILL_2__8838_ gnd vdd FILL
XFILL_3__11446_ gnd vdd FILL
XFILL_0__14054_ gnd vdd FILL
XFILL_2__14964_ gnd vdd FILL
XFILL_4__10997_ gnd vdd FILL
XFILL_1__16393_ gnd vdd FILL
X_8200_ _8200_/A gnd _8202_/A vdd INVX1
XFILL_5__12006_ gnd vdd FILL
XFILL_0__11266_ gnd vdd FILL
XFILL_4__15524_ gnd vdd FILL
X_16249_ _16249_/A _16247_/Y gnd _16251_/C vdd NOR2X1
XFILL_4__12736_ gnd vdd FILL
X_9180_ _9180_/Q _7534_/CLK _8156_/R vdd _9098_/Y gnd vdd DFFSR
XFILL_0__7853_ gnd vdd FILL
XFILL_3__14165_ gnd vdd FILL
XFILL_0__13005_ gnd vdd FILL
XFILL_2__13915_ gnd vdd FILL
XFILL_1__15344_ gnd vdd FILL
XFILL_3__7562_ gnd vdd FILL
XFILL_2__8769_ gnd vdd FILL
XFILL_3__11377_ gnd vdd FILL
XFILL_2__14895_ gnd vdd FILL
XFILL_5__8478_ gnd vdd FILL
X_8131_ _8131_/A _8082_/A _8131_/C gnd _8175_/D vdd OAI21X1
XFILL_0__11197_ gnd vdd FILL
XFILL_3__13116_ gnd vdd FILL
XFILL_3__9301_ gnd vdd FILL
XFILL_4__15455_ gnd vdd FILL
XSFILL94440x58050 gnd vdd FILL
XFILL_1__11507_ gnd vdd FILL
XSFILL3400x72050 gnd vdd FILL
XFILL_2__13846_ gnd vdd FILL
XFILL_3__14096_ gnd vdd FILL
XFILL_1__15275_ gnd vdd FILL
XFILL_0__10148_ gnd vdd FILL
XFILL_1__12487_ gnd vdd FILL
XFILL_3__7493_ gnd vdd FILL
XFILL_5__7429_ gnd vdd FILL
XFILL_0__9523_ gnd vdd FILL
XFILL_6__10439_ gnd vdd FILL
XFILL_4__14406_ gnd vdd FILL
X_8062_ _8062_/A _8107_/B _8062_/C gnd _8152_/D vdd OAI21X1
XFILL_4__11618_ gnd vdd FILL
XFILL_3__9232_ gnd vdd FILL
XFILL_4__15386_ gnd vdd FILL
XFILL_1__14226_ gnd vdd FILL
XSFILL69240x34050 gnd vdd FILL
XFILL_3__10259_ gnd vdd FILL
XFILL_5__13957_ gnd vdd FILL
XFILL_4__12598_ gnd vdd FILL
XSFILL53960x4050 gnd vdd FILL
XFILL_1__11438_ gnd vdd FILL
XFILL_2__13777_ gnd vdd FILL
X_7013_ _6947_/A _7534_/CLK _8156_/R vdd _7013_/D gnd vdd DFFSR
XFILL_2__10989_ gnd vdd FILL
XFILL_0__14956_ gnd vdd FILL
XFILL_5__12908_ gnd vdd FILL
XFILL_4__14337_ gnd vdd FILL
XFILL_2__15516_ gnd vdd FILL
XFILL_4__11549_ gnd vdd FILL
XFILL_2__12728_ gnd vdd FILL
XFILL_3__9163_ gnd vdd FILL
XFILL_1__14157_ gnd vdd FILL
XFILL_5__13888_ gnd vdd FILL
XFILL_0__13907_ gnd vdd FILL
XFILL_1__11369_ gnd vdd FILL
XSFILL104440x43050 gnd vdd FILL
XFILL_0__8405_ gnd vdd FILL
XFILL_0__14887_ gnd vdd FILL
XFILL_5__15627_ gnd vdd FILL
XFILL_1__13108_ gnd vdd FILL
XFILL_3__8114_ gnd vdd FILL
XFILL_0__9385_ gnd vdd FILL
XFILL_5__12839_ gnd vdd FILL
XFILL_4__14268_ gnd vdd FILL
XSFILL33720x75050 gnd vdd FILL
XSFILL8680x41050 gnd vdd FILL
XFILL_2__15447_ gnd vdd FILL
XFILL_2__12659_ gnd vdd FILL
XFILL_0__13838_ gnd vdd FILL
XFILL_3__14998_ gnd vdd FILL
XFILL_3__9094_ gnd vdd FILL
XFILL_1__14088_ gnd vdd FILL
XFILL_4__16007_ gnd vdd FILL
XSFILL48520x35050 gnd vdd FILL
XFILL_4__13219_ gnd vdd FILL
XFILL_0__8336_ gnd vdd FILL
XFILL_5__15558_ gnd vdd FILL
XFILL_4__14199_ gnd vdd FILL
X_8964_ _8964_/A _9014_/A _8964_/C gnd _8964_/Y vdd OAI21X1
XFILL_1__13039_ gnd vdd FILL
XFILL_3__13949_ gnd vdd FILL
XFILL_2__15378_ gnd vdd FILL
XFILL_0__13769_ gnd vdd FILL
XFILL_5__14509_ gnd vdd FILL
XFILL_1__7060_ gnd vdd FILL
X_7915_ _7915_/Q _7915_/CLK _7915_/R vdd _7915_/D gnd vdd DFFSR
XFILL_0__8267_ gnd vdd FILL
X_8895_ _8896_/B _7743_/B gnd _8895_/Y vdd NAND2X1
XFILL_5__15489_ gnd vdd FILL
XFILL_2__14329_ gnd vdd FILL
XFILL_0__15508_ gnd vdd FILL
XFILL_0__7218_ gnd vdd FILL
X_7846_ _7910_/Q gnd _7848_/A vdd INVX1
XFILL_6__6986_ gnd vdd FILL
XFILL_3__15619_ gnd vdd FILL
XFILL_0__8198_ gnd vdd FILL
XFILL_0__15439_ gnd vdd FILL
XFILL_3__9996_ gnd vdd FILL
XSFILL13640x42050 gnd vdd FILL
XFILL_0_CLKBUF1_insert116 gnd vdd FILL
XFILL_0_CLKBUF1_insert127 gnd vdd FILL
X_7777_ _7703_/A _9188_/CLK _8929_/R vdd _7777_/D gnd vdd DFFSR
XFILL_0_CLKBUF1_insert138 gnd vdd FILL
XFILL_4__7740_ gnd vdd FILL
XFILL_0_CLKBUF1_insert149 gnd vdd FILL
XSFILL13720x7050 gnd vdd FILL
XSFILL94120x40050 gnd vdd FILL
X_9516_ _9516_/A gnd _9516_/Y vdd INVX1
XFILL_1__7962_ gnd vdd FILL
XFILL_4__7671_ gnd vdd FILL
XFILL_3__8878_ gnd vdd FILL
XFILL_1__6913_ gnd vdd FILL
X_9447_ _9385_/A _9447_/CLK _9447_/R vdd _9447_/D gnd vdd DFFSR
XFILL_4__9410_ gnd vdd FILL
XFILL_1__7893_ gnd vdd FILL
XFILL_3__7829_ gnd vdd FILL
XFILL_1__9632_ gnd vdd FILL
XFILL_4_BUFX2_insert601 gnd vdd FILL
XSFILL8760x21050 gnd vdd FILL
X_9378_ _9378_/A _9398_/A _9377_/Y gnd _9444_/D vdd OAI21X1
XFILL_1__6844_ gnd vdd FILL
XFILL_4_BUFX2_insert612 gnd vdd FILL
XFILL_4__9341_ gnd vdd FILL
XSFILL43160x80050 gnd vdd FILL
XFILL_4_BUFX2_insert623 gnd vdd FILL
XFILL_4_BUFX2_insert634 gnd vdd FILL
X_10260_ _15474_/A gnd _10262_/A vdd INVX1
X_8329_ _8356_/A _6921_/B gnd _8329_/Y vdd NAND2X1
XFILL_4_BUFX2_insert645 gnd vdd FILL
XFILL_4_BUFX2_insert656 gnd vdd FILL
XFILL_4_BUFX2_insert667 gnd vdd FILL
XFILL_4__9272_ gnd vdd FILL
XFILL_4_BUFX2_insert678 gnd vdd FILL
X_10191_ _10189_/Y _10191_/B _10191_/C gnd _10227_/D vdd OAI21X1
XFILL_4_BUFX2_insert689 gnd vdd FILL
XFILL_1__8514_ gnd vdd FILL
XFILL_1__9494_ gnd vdd FILL
XFILL_4__8223_ gnd vdd FILL
XFILL111960x65050 gnd vdd FILL
XFILL_1__8445_ gnd vdd FILL
XSFILL13720x22050 gnd vdd FILL
X_13950_ _9312_/Q _13854_/B _13621_/B _15474_/A gnd _13952_/A vdd AOI22X1
XFILL_1__8376_ gnd vdd FILL
XFILL_4__7105_ gnd vdd FILL
X_12901_ _12901_/A gnd _12901_/Y vdd INVX1
XFILL_4__8085_ gnd vdd FILL
X_13881_ _8030_/Q gnd _13881_/Y vdd INVX1
XFILL_1__7327_ gnd vdd FILL
XFILL_4__7036_ gnd vdd FILL
X_15620_ _15652_/A _9572_/Q _9700_/Q _15652_/D gnd _15628_/B vdd AOI22X1
X_12832_ _12125_/B gnd _12832_/Y vdd INVX1
XFILL_1_BUFX2_insert502 gnd vdd FILL
XFILL_1_BUFX2_insert513 gnd vdd FILL
X_15551_ _14041_/Y _15197_/B _15045_/D _14026_/Y gnd _15555_/A vdd OAI22X1
XFILL_1_BUFX2_insert524 gnd vdd FILL
XFILL_1_BUFX2_insert535 gnd vdd FILL
X_12763_ _12761_/Y _12762_/A _12763_/C gnd _12813_/D vdd OAI21X1
XFILL_1_BUFX2_insert546 gnd vdd FILL
XFILL_1__7189_ gnd vdd FILL
XFILL_1_BUFX2_insert557 gnd vdd FILL
X_14502_ _7736_/A gnd _14502_/Y vdd INVX1
XFILL_1_BUFX2_insert568 gnd vdd FILL
XFILL_4__8987_ gnd vdd FILL
X_11714_ _11713_/Y _11074_/C gnd _11716_/A vdd AND2X2
XSFILL84120x72050 gnd vdd FILL
XFILL_1_BUFX2_insert579 gnd vdd FILL
X_15482_ _15482_/A _15680_/B _15680_/C gnd _15482_/Y vdd NAND3X1
XFILL_2__9810_ gnd vdd FILL
X_12694_ _12694_/Q _12692_/CLK _12692_/R vdd _12694_/D gnd vdd DFFSR
XSFILL99480x9050 gnd vdd FILL
XFILL_4__7938_ gnd vdd FILL
X_14433_ _14433_/A _14725_/A _14815_/C _14431_/Y gnd _14437_/B vdd OAI22X1
XFILL_4__10920_ gnd vdd FILL
XFILL_2__10010_ gnd vdd FILL
X_11645_ _11658_/A _11681_/B gnd _11646_/C vdd NAND2X1
XFILL_5__11170_ gnd vdd FILL
XFILL_2__9741_ gnd vdd FILL
XFILL_2__6953_ gnd vdd FILL
XFILL_4__7869_ gnd vdd FILL
XFILL_5__10121_ gnd vdd FILL
X_14364_ _7145_/Q gnd _14365_/D vdd INVX1
XFILL_3__11300_ gnd vdd FILL
X_11576_ _11551_/A _11577_/B gnd _11576_/Y vdd AND2X2
XFILL_4__9608_ gnd vdd FILL
XFILL_2__9672_ gnd vdd FILL
XFILL_3__12280_ gnd vdd FILL
XFILL_0__11120_ gnd vdd FILL
XFILL_5__8401_ gnd vdd FILL
XFILL112120x54050 gnd vdd FILL
XFILL_2__6884_ gnd vdd FILL
X_16103_ _9796_/A _15390_/B gnd _16111_/A vdd NAND2X1
XFILL_1__10671_ gnd vdd FILL
X_13315_ _13299_/A _13245_/B gnd _13316_/B vdd NAND2X1
XFILL_5__9381_ gnd vdd FILL
XFILL_5__10052_ gnd vdd FILL
X_10527_ _10525_/Y _10581_/B _10526_/Y gnd _10527_/Y vdd OAI21X1
XFILL_1__12410_ gnd vdd FILL
XFILL_5_BUFX2_insert490 gnd vdd FILL
XFILL_2__8623_ gnd vdd FILL
XFILL_4__13570_ gnd vdd FILL
XSFILL39240x13050 gnd vdd FILL
X_14295_ _14295_/A gnd _15766_/B vdd INVX1
XFILL_3__11231_ gnd vdd FILL
XFILL_4__10782_ gnd vdd FILL
XFILL_5__8332_ gnd vdd FILL
XFILL_2__11961_ gnd vdd FILL
XFILL_1__13390_ gnd vdd FILL
XFILL_4__9539_ gnd vdd FILL
XFILL_0__11051_ gnd vdd FILL
X_16034_ _9838_/Q gnd _16036_/B vdd INVX1
X_13246_ _13246_/A _13246_/B gnd _13310_/A vdd NAND2X1
X_10458_ _15234_/A _9818_/CLK _8676_/R vdd _10372_/Y gnd vdd DFFSR
XFILL_4__12521_ gnd vdd FILL
XFILL_5__14860_ gnd vdd FILL
XFILL_3__11162_ gnd vdd FILL
XFILL_2__13700_ gnd vdd FILL
XFILL_2__10912_ gnd vdd FILL
XFILL_1__12341_ gnd vdd FILL
XFILL_0__10002_ gnd vdd FILL
XFILL_2__14680_ gnd vdd FILL
XFILL_2__11892_ gnd vdd FILL
XFILL_5__8263_ gnd vdd FILL
XFILL_3__10113_ gnd vdd FILL
XFILL_5__13811_ gnd vdd FILL
XFILL_4__15240_ gnd vdd FILL
XFILL_4__12452_ gnd vdd FILL
X_13177_ _13085_/A _13201_/CLK _13201_/R vdd _13087_/Y gnd vdd DFFSR
X_10389_ _10450_/B _7445_/B gnd _10389_/Y vdd NAND2X1
XFILL_2__7505_ gnd vdd FILL
XFILL_3__15970_ gnd vdd FILL
XFILL_2__13631_ gnd vdd FILL
XFILL_1__15060_ gnd vdd FILL
XFILL_3__11093_ gnd vdd FILL
XFILL_5__14791_ gnd vdd FILL
XFILL_2__8485_ gnd vdd FILL
XFILL_0__14810_ gnd vdd FILL
XFILL_5__7214_ gnd vdd FILL
XFILL_1__12272_ gnd vdd FILL
XFILL_0__15790_ gnd vdd FILL
XFILL_5__8194_ gnd vdd FILL
XSFILL69160x49050 gnd vdd FILL
X_12128_ _12134_/A _12923_/Q gnd _12129_/C vdd NAND2X1
XFILL_4__11403_ gnd vdd FILL
XFILL_5__10954_ gnd vdd FILL
XFILL_3__10044_ gnd vdd FILL
XFILL_4__15171_ gnd vdd FILL
XFILL_5__13742_ gnd vdd FILL
XFILL_1__14011_ gnd vdd FILL
XFILL_3__14921_ gnd vdd FILL
XFILL_2__7436_ gnd vdd FILL
XFILL_4__12383_ gnd vdd FILL
XFILL_2__16350_ gnd vdd FILL
XFILL_1__11223_ gnd vdd FILL
XFILL_0__14741_ gnd vdd FILL
XFILL_2__13562_ gnd vdd FILL
XFILL_2__10774_ gnd vdd FILL
XFILL_0__11953_ gnd vdd FILL
X_12059_ _11987_/A _12553_/Q _12059_/C gnd _12062_/A vdd NAND3X1
XFILL_6__10155_ gnd vdd FILL
XFILL_4__14122_ gnd vdd FILL
XFILL_2__15301_ gnd vdd FILL
XFILL_5__13673_ gnd vdd FILL
XFILL_4__11334_ gnd vdd FILL
XFILL_3__14852_ gnd vdd FILL
XFILL_2__12513_ gnd vdd FILL
XSFILL104360x58050 gnd vdd FILL
XFILL_5__10885_ gnd vdd FILL
XFILL_0__10904_ gnd vdd FILL
XFILL_0_BUFX2_insert18 gnd vdd FILL
XFILL_2__7367_ gnd vdd FILL
XFILL_1__11154_ gnd vdd FILL
XFILL_2__16281_ gnd vdd FILL
XFILL_0__14672_ gnd vdd FILL
XFILL_2__13493_ gnd vdd FILL
XFILL_5__7076_ gnd vdd FILL
XFILL_5__15412_ gnd vdd FILL
XFILL_0_BUFX2_insert29 gnd vdd FILL
XFILL_0__11884_ gnd vdd FILL
XFILL_5__12624_ gnd vdd FILL
XFILL_0__9170_ gnd vdd FILL
XFILL_3__13803_ gnd vdd FILL
XFILL_4__14053_ gnd vdd FILL
XFILL_6__14963_ gnd vdd FILL
XFILL_2__9106_ gnd vdd FILL
XFILL_2__15232_ gnd vdd FILL
XFILL_1__10105_ gnd vdd FILL
XFILL_5__16392_ gnd vdd FILL
XFILL_4__11265_ gnd vdd FILL
XFILL_0__13623_ gnd vdd FILL
XFILL_2__12444_ gnd vdd FILL
XFILL_0__16411_ gnd vdd FILL
XFILL_3__14783_ gnd vdd FILL
XFILL_2__7298_ gnd vdd FILL
XFILL_3__11995_ gnd vdd FILL
XFILL_1__15962_ gnd vdd FILL
XFILL_1__11085_ gnd vdd FILL
XFILL_0__10835_ gnd vdd FILL
XFILL_0__8121_ gnd vdd FILL
X_15818_ _8367_/A _15978_/B _16212_/A _8681_/Q gnd _15818_/Y vdd AOI22X1
XFILL_6__13914_ gnd vdd FILL
XFILL_4__13004_ gnd vdd FILL
XFILL_5__15343_ gnd vdd FILL
XFILL_2__9037_ gnd vdd FILL
XFILL112200x34050 gnd vdd FILL
XFILL_2_BUFX2_insert380 gnd vdd FILL
XSFILL49080x16050 gnd vdd FILL
XFILL_3__13734_ gnd vdd FILL
XFILL_3__10946_ gnd vdd FILL
XFILL_0__16342_ gnd vdd FILL
XFILL_2__12375_ gnd vdd FILL
XFILL_1__10036_ gnd vdd FILL
XFILL_2__15163_ gnd vdd FILL
XFILL_4__11196_ gnd vdd FILL
XFILL_1__14913_ gnd vdd FILL
XFILL_2_BUFX2_insert391 gnd vdd FILL
XSFILL23720x2050 gnd vdd FILL
XFILL_0__13554_ gnd vdd FILL
XFILL_0__10766_ gnd vdd FILL
XFILL_1__15893_ gnd vdd FILL
X_7700_ _7700_/A gnd _7700_/Y vdd INVX1
XFILL_5__11506_ gnd vdd FILL
XFILL_5__15274_ gnd vdd FILL
X_15749_ _9897_/A gnd _15749_/Y vdd INVX1
XFILL_5__12486_ gnd vdd FILL
XFILL_4__10147_ gnd vdd FILL
X_8680_ _8620_/A _8680_/CLK _8034_/R vdd _8680_/D gnd vdd DFFSR
XFILL_2__14114_ gnd vdd FILL
XFILL_2__11326_ gnd vdd FILL
XFILL_3__13665_ gnd vdd FILL
XFILL_0__12505_ gnd vdd FILL
XFILL_3__9850_ gnd vdd FILL
XFILL_1__14844_ gnd vdd FILL
XFILL_3__10877_ gnd vdd FILL
XFILL_2__15094_ gnd vdd FILL
XFILL_0__16273_ gnd vdd FILL
XFILL_0__13485_ gnd vdd FILL
X_7631_ _7631_/A _7592_/B _7631_/C gnd _7667_/D vdd OAI21X1
XFILL_3__15404_ gnd vdd FILL
XFILL_5__14225_ gnd vdd FILL
XFILL_5__11437_ gnd vdd FILL
XFILL_5__7978_ gnd vdd FILL
XFILL_0__10697_ gnd vdd FILL
XFILL_3__12616_ gnd vdd FILL
XFILL_6__13776_ gnd vdd FILL
XFILL112200x6050 gnd vdd FILL
XFILL_3__16384_ gnd vdd FILL
XFILL_2__14045_ gnd vdd FILL
XFILL_0__15224_ gnd vdd FILL
XFILL_4__14955_ gnd vdd FILL
XFILL_2__11257_ gnd vdd FILL
XFILL_3__9781_ gnd vdd FILL
XFILL_3__13596_ gnd vdd FILL
XSFILL3400x67050 gnd vdd FILL
XFILL_6__8510_ gnd vdd FILL
XFILL_0__12436_ gnd vdd FILL
XSFILL53960x62050 gnd vdd FILL
XFILL_1__11987_ gnd vdd FILL
XFILL_5__6929_ gnd vdd FILL
XFILL_3__6993_ gnd vdd FILL
XFILL_1__14775_ gnd vdd FILL
XFILL_6__12727_ gnd vdd FILL
XFILL_5__14156_ gnd vdd FILL
XFILL_3__15335_ gnd vdd FILL
X_7562_ _7560_/Y _7562_/B _7561_/Y gnd _7562_/Y vdd OAI21X1
XFILL_4__13906_ gnd vdd FILL
XFILL_5__11368_ gnd vdd FILL
XFILL_3__8732_ gnd vdd FILL
XFILL_2__9939_ gnd vdd FILL
XFILL_4__14886_ gnd vdd FILL
XFILL_1__10938_ gnd vdd FILL
XFILL_0__15155_ gnd vdd FILL
XFILL_2__11188_ gnd vdd FILL
XFILL_1__13726_ gnd vdd FILL
XFILL_0__12367_ gnd vdd FILL
XFILL_5__13107_ gnd vdd FILL
X_9301_ _9299_/Y _9301_/B _9301_/C gnd _9333_/D vdd OAI21X1
XFILL_5__9648_ gnd vdd FILL
XFILL_5__10319_ gnd vdd FILL
XFILL_0__8954_ gnd vdd FILL
XFILL_5__14087_ gnd vdd FILL
XSFILL54040x71050 gnd vdd FILL
XFILL_4__13837_ gnd vdd FILL
X_7493_ _7457_/A _8005_/B gnd _7493_/Y vdd NAND2X1
XFILL_2__10139_ gnd vdd FILL
XFILL_0__14106_ gnd vdd FILL
XFILL_5__11299_ gnd vdd FILL
XFILL_3__15266_ gnd vdd FILL
XBUFX2_insert390 _12387_/Y gnd _8225_/B vdd BUFX2
XFILL_3__12478_ gnd vdd FILL
XFILL_0__11318_ gnd vdd FILL
XFILL_2__15996_ gnd vdd FILL
XFILL_1__13657_ gnd vdd FILL
XFILL_0__15086_ gnd vdd FILL
X_9232_ _9232_/A _9232_/B _9231_/Y gnd _9310_/D vdd OAI21X1
XFILL_5__13038_ gnd vdd FILL
XSFILL104440x38050 gnd vdd FILL
XFILL_0__12298_ gnd vdd FILL
XFILL_3__14217_ gnd vdd FILL
XFILL_0__8885_ gnd vdd FILL
XFILL_3__7614_ gnd vdd FILL
XFILL_4__13768_ gnd vdd FILL
XFILL_3__11429_ gnd vdd FILL
XFILL_3__15197_ gnd vdd FILL
XFILL_1__12608_ gnd vdd FILL
XFILL_0__14037_ gnd vdd FILL
XSFILL8680x36050 gnd vdd FILL
XFILL_2__14947_ gnd vdd FILL
XFILL_1__13588_ gnd vdd FILL
XFILL_1__16376_ gnd vdd FILL
XFILL_3__8594_ gnd vdd FILL
XFILL_0__11249_ gnd vdd FILL
XFILL_4__12719_ gnd vdd FILL
X_9163_ _9163_/A _7243_/B gnd _9164_/C vdd NAND2X1
XFILL_4__15507_ gnd vdd FILL
XFILL_0__7836_ gnd vdd FILL
XFILL_3__14148_ gnd vdd FILL
XFILL_1__15327_ gnd vdd FILL
XFILL_4__13699_ gnd vdd FILL
XFILL_3__7545_ gnd vdd FILL
XFILL_2__14878_ gnd vdd FILL
X_8114_ _8170_/Q gnd _8116_/A vdd INVX1
XFILL_3_BUFX2_insert608 gnd vdd FILL
X_9094_ _9086_/B _9094_/B gnd _9095_/C vdd NAND2X1
XFILL_4__15438_ gnd vdd FILL
XFILL_2__13829_ gnd vdd FILL
XFILL_5__14989_ gnd vdd FILL
XFILL_3_BUFX2_insert619 gnd vdd FILL
XFILL_3__14079_ gnd vdd FILL
XFILL_1__15258_ gnd vdd FILL
XFILL_3__7476_ gnd vdd FILL
XFILL_0__9506_ gnd vdd FILL
XFILL_0__15988_ gnd vdd FILL
X_8045_ _8045_/Q _7411_/CLK _7411_/R vdd _8045_/D gnd vdd DFFSR
XFILL_3__9215_ gnd vdd FILL
XFILL_4__15369_ gnd vdd FILL
XFILL_1__14209_ gnd vdd FILL
XFILL_0__7698_ gnd vdd FILL
XFILL_1__15189_ gnd vdd FILL
XSFILL49000x60050 gnd vdd FILL
XSFILL13640x37050 gnd vdd FILL
XFILL_0__14939_ gnd vdd FILL
XFILL_1__8230_ gnd vdd FILL
XFILL_3__9146_ gnd vdd FILL
XSFILL109560x71050 gnd vdd FILL
XFILL_0__9368_ gnd vdd FILL
X_9996_ _9996_/A _7948_/B gnd _9997_/C vdd NAND2X1
XFILL_0__8319_ gnd vdd FILL
XSFILL54120x51050 gnd vdd FILL
XFILL_1__7112_ gnd vdd FILL
XFILL_1__8092_ gnd vdd FILL
X_8947_ _8909_/A _8947_/CLK _9069_/R vdd _8947_/D gnd vdd DFFSR
XFILL_4__8910_ gnd vdd FILL
XFILL_0__9299_ gnd vdd FILL
XSFILL104520x18050 gnd vdd FILL
XFILL_4__9890_ gnd vdd FILL
XFILL_1__7043_ gnd vdd FILL
XSFILL8760x16050 gnd vdd FILL
XFILL_4__8841_ gnd vdd FILL
X_8878_ _8878_/A _8859_/A _8877_/Y gnd _8936_/D vdd OAI21X1
X_7829_ _7892_/A _8853_/B gnd _7830_/C vdd NAND2X1
XFILL_0_BUFX2_insert509 gnd vdd FILL
XFILL_4__8772_ gnd vdd FILL
XFILL_3__9979_ gnd vdd FILL
XSFILL23880x8050 gnd vdd FILL
XFILL_1__8994_ gnd vdd FILL
XFILL_4__7723_ gnd vdd FILL
X_11430_ _11256_/Y gnd _11431_/A vdd INVX1
XFILL_1__7945_ gnd vdd FILL
XSFILL13720x17050 gnd vdd FILL
X_11361_ _11778_/B gnd _11764_/A vdd INVX4
XFILL112040x69050 gnd vdd FILL
XSFILL23880x61050 gnd vdd FILL
XFILL_1__7876_ gnd vdd FILL
X_13100_ _13182_/Q gnd _13100_/Y vdd INVX1
X_10312_ _10280_/B _8136_/B gnd _10312_/Y vdd NAND2X1
XFILL_4__7585_ gnd vdd FILL
XFILL_4_BUFX2_insert420 gnd vdd FILL
XFILL_1__9615_ gnd vdd FILL
XFILL_4_BUFX2_insert431 gnd vdd FILL
X_11292_ _11529_/A _11105_/Y gnd _11527_/C vdd OR2X2
X_14080_ _14078_/Y _14441_/B _14744_/B _15589_/B gnd _14084_/B vdd OAI22X1
XSFILL38920x83050 gnd vdd FILL
XFILL_4_BUFX2_insert442 gnd vdd FILL
XFILL_4_BUFX2_insert453 gnd vdd FILL
XSFILL69240x7050 gnd vdd FILL
X_10243_ _10294_/A _7555_/B gnd _10243_/Y vdd NAND2X1
X_13031_ _13029_/Y vdd _13031_/C gnd _13073_/D vdd OAI21X1
XFILL_4_BUFX2_insert464 gnd vdd FILL
XFILL_4_BUFX2_insert475 gnd vdd FILL
XFILL_1__9546_ gnd vdd FILL
XFILL_4_BUFX2_insert486 gnd vdd FILL
XFILL_4__9255_ gnd vdd FILL
XFILL_4_BUFX2_insert497 gnd vdd FILL
X_10174_ _10222_/Q gnd _10174_/Y vdd INVX1
XFILL_4__8206_ gnd vdd FILL
XFILL_2__8270_ gnd vdd FILL
XFILL_1__9477_ gnd vdd FILL
XFILL_2__7221_ gnd vdd FILL
X_14982_ _12767_/A _12764_/A gnd _14982_/Y vdd AND2X2
XSFILL18840x50050 gnd vdd FILL
XFILL_4__8137_ gnd vdd FILL
X_13933_ _15476_/C _14377_/B gnd _13933_/Y vdd NOR2X1
XFILL_5__10670_ gnd vdd FILL
XFILL_3_CLKBUF1_insert111 gnd vdd FILL
XFILL_1__8359_ gnd vdd FILL
XFILL_3_CLKBUF1_insert122 gnd vdd FILL
XFILL_3_CLKBUF1_insert133 gnd vdd FILL
XFILL_2__10490_ gnd vdd FILL
XFILL_5__8950_ gnd vdd FILL
XFILL_3_CLKBUF1_insert144 gnd vdd FILL
XFILL_4__8068_ gnd vdd FILL
XFILL_5_CLKBUF1_insert1082 gnd vdd FILL
X_13864_ _8670_/Q _13864_/B _13864_/C _8542_/Q gnd _13864_/Y vdd AOI22X1
XFILL_3__10800_ gnd vdd FILL
XFILL_3_CLKBUF1_insert155 gnd vdd FILL
XFILL_4__11050_ gnd vdd FILL
XFILL_3_CLKBUF1_insert166 gnd vdd FILL
XFILL_2__7083_ gnd vdd FILL
XFILL_3_CLKBUF1_insert177 gnd vdd FILL
XFILL_0__10620_ gnd vdd FILL
XFILL_3__11780_ gnd vdd FILL
XFILL_3_CLKBUF1_insert188 gnd vdd FILL
XSFILL84920x7050 gnd vdd FILL
X_15603_ _15449_/C _14091_/A _14118_/D _16314_/A gnd _15603_/Y vdd OAI22X1
X_12815_ _12767_/A _8171_/CLK _12795_/R vdd _12815_/D gnd vdd DFFSR
XFILL112120x49050 gnd vdd FILL
XFILL_5__12340_ gnd vdd FILL
XFILL_4__10001_ gnd vdd FILL
XFILL_1_BUFX2_insert310 gnd vdd FILL
XFILL_5__8881_ gnd vdd FILL
XFILL_3_CLKBUF1_insert199 gnd vdd FILL
XFILL_1_BUFX2_insert321 gnd vdd FILL
X_13795_ _13794_/Y _13795_/B _13876_/C _13793_/Y gnd _13796_/A vdd OAI22X1
XFILL_2__12160_ gnd vdd FILL
XFILL_6__11891_ gnd vdd FILL
XFILL_1_BUFX2_insert332 gnd vdd FILL
XFILL_1__11910_ gnd vdd FILL
XFILL_0__10551_ gnd vdd FILL
XFILL_5__7832_ gnd vdd FILL
XFILL_1__12890_ gnd vdd FILL
XFILL_1_BUFX2_insert343 gnd vdd FILL
XFILL_1_BUFX2_insert354 gnd vdd FILL
X_15534_ _15533_/Y _15528_/Y gnd _15534_/Y vdd NAND2X1
X_12746_ _12808_/Q gnd _12748_/A vdd INVX1
XFILL_1_BUFX2_insert365 gnd vdd FILL
XFILL_5__12271_ gnd vdd FILL
XFILL_2__11111_ gnd vdd FILL
XFILL_3__13450_ gnd vdd FILL
XFILL_1_BUFX2_insert376 gnd vdd FILL
XFILL_3__10662_ gnd vdd FILL
XFILL_2__12091_ gnd vdd FILL
XFILL_1__11841_ gnd vdd FILL
XFILL_0__13270_ gnd vdd FILL
XFILL_5__14010_ gnd vdd FILL
XFILL_1_BUFX2_insert387 gnd vdd FILL
XFILL_1_BUFX2_insert398 gnd vdd FILL
XFILL_5__7763_ gnd vdd FILL
XFILL_5__11222_ gnd vdd FILL
XFILL_3__12401_ gnd vdd FILL
XFILL_4__14740_ gnd vdd FILL
XFILL_6__13561_ gnd vdd FILL
X_15465_ _15463_/Y _15464_/Y gnd _15466_/B vdd NOR2X1
X_12677_ _12609_/A _8171_/CLK _12795_/R vdd _12677_/D gnd vdd DFFSR
XFILL_4__11952_ gnd vdd FILL
XFILL_2__11042_ gnd vdd FILL
XFILL_3__13381_ gnd vdd FILL
XFILL_5__9502_ gnd vdd FILL
XFILL_0__12221_ gnd vdd FILL
XFILL_1__14560_ gnd vdd FILL
XFILL_2__7985_ gnd vdd FILL
XFILL_1__11772_ gnd vdd FILL
X_14416_ _7530_/Q gnd _15869_/B vdd INVX1
XFILL_5__7694_ gnd vdd FILL
XFILL_4__10903_ gnd vdd FILL
XFILL_5__11153_ gnd vdd FILL
X_11628_ _11628_/A _11619_/Y _11627_/Y gnd _11629_/A vdd AOI21X1
XFILL_3__15120_ gnd vdd FILL
X_15396_ _15677_/A _13855_/Y _13844_/Y _15677_/D gnd _15397_/C vdd OAI22X1
XFILL_3__12332_ gnd vdd FILL
XFILL_2__9724_ gnd vdd FILL
XSFILL3640x9050 gnd vdd FILL
XFILL_4__14671_ gnd vdd FILL
XFILL_4__11883_ gnd vdd FILL
XFILL_2__6936_ gnd vdd FILL
XFILL_2__15850_ gnd vdd FILL
XFILL_1__13511_ gnd vdd FILL
XFILL_1__14491_ gnd vdd FILL
XFILL_0__12152_ gnd vdd FILL
XSFILL84200x47050 gnd vdd FILL
XFILL_5__10104_ gnd vdd FILL
XFILL_4__13622_ gnd vdd FILL
XFILL_4__16410_ gnd vdd FILL
X_14347_ _6956_/A gnd _14348_/D vdd INVX1
XFILL_6__12443_ gnd vdd FILL
XFILL_2__14801_ gnd vdd FILL
XFILL_3__15051_ gnd vdd FILL
XFILL_5__15961_ gnd vdd FILL
XFILL_5__11084_ gnd vdd FILL
X_11559_ _11157_/Y gnd _11559_/Y vdd INVX1
XFILL_4__10834_ gnd vdd FILL
XFILL_2__9655_ gnd vdd FILL
XFILL_1__16230_ gnd vdd FILL
XFILL_1__13442_ gnd vdd FILL
XFILL_3__12263_ gnd vdd FILL
XFILL_0__11103_ gnd vdd FILL
XFILL_2__6867_ gnd vdd FILL
XFILL_2__15781_ gnd vdd FILL
XFILL_1__10654_ gnd vdd FILL
XFILL_0__12083_ gnd vdd FILL
XFILL_2__12993_ gnd vdd FILL
XFILL_5__9364_ gnd vdd FILL
XFILL_4__16341_ gnd vdd FILL
XFILL_3__14002_ gnd vdd FILL
XFILL_5__10035_ gnd vdd FILL
XFILL_5__14912_ gnd vdd FILL
XSFILL59000x23050 gnd vdd FILL
XFILL_2__8606_ gnd vdd FILL
XFILL_4__13553_ gnd vdd FILL
X_14278_ _14030_/A _14278_/B _13461_/C _14278_/D gnd _14278_/Y vdd OAI22X1
XFILL_3__11214_ gnd vdd FILL
XFILL_4__10765_ gnd vdd FILL
XFILL_5__15892_ gnd vdd FILL
XFILL_2__14732_ gnd vdd FILL
XFILL_0__15911_ gnd vdd FILL
XFILL_2__11944_ gnd vdd FILL
XFILL_3__12194_ gnd vdd FILL
XFILL_1__13373_ gnd vdd FILL
XFILL_5__8315_ gnd vdd FILL
XFILL_1__16161_ gnd vdd FILL
XFILL_0__11034_ gnd vdd FILL
X_16017_ _8430_/Q gnd _16018_/A vdd INVX1
X_13229_ _13246_/A _13246_/B gnd _13288_/B vdd NOR2X1
XFILL_5__9295_ gnd vdd FILL
XFILL_4__12504_ gnd vdd FILL
XFILL_0__7621_ gnd vdd FILL
XFILL_5__14843_ gnd vdd FILL
XFILL_4__16272_ gnd vdd FILL
XFILL_3__7330_ gnd vdd FILL
XFILL_4__13484_ gnd vdd FILL
XFILL_1__12324_ gnd vdd FILL
XFILL_3__11145_ gnd vdd FILL
XFILL_1__15112_ gnd vdd FILL
XSFILL74680x56050 gnd vdd FILL
XFILL_1__16092_ gnd vdd FILL
XFILL112200x29050 gnd vdd FILL
XFILL_2__14663_ gnd vdd FILL
XFILL_4__10696_ gnd vdd FILL
XFILL_2__11875_ gnd vdd FILL
XFILL_5__8246_ gnd vdd FILL
XFILL_0__15842_ gnd vdd FILL
XFILL_4__15223_ gnd vdd FILL
XSFILL89480x16050 gnd vdd FILL
XFILL_0__7552_ gnd vdd FILL
XFILL_4__12435_ gnd vdd FILL
XFILL_2__16402_ gnd vdd FILL
XSFILL64120x14050 gnd vdd FILL
XFILL_2__13614_ gnd vdd FILL
XFILL_3__15953_ gnd vdd FILL
XFILL_5__14774_ gnd vdd FILL
XFILL_2__10826_ gnd vdd FILL
XFILL_5__11986_ gnd vdd FILL
XFILL_1__15043_ gnd vdd FILL
XFILL_1__12255_ gnd vdd FILL
XFILL_3__11076_ gnd vdd FILL
XFILL_2__8468_ gnd vdd FILL
XFILL_2__14594_ gnd vdd FILL
XFILL_0__12985_ gnd vdd FILL
XFILL_0__15773_ gnd vdd FILL
XFILL_3__9000_ gnd vdd FILL
XFILL_4__15154_ gnd vdd FILL
XFILL_5__13725_ gnd vdd FILL
XFILL_5__10937_ gnd vdd FILL
XFILL_4__12366_ gnd vdd FILL
XFILL_0__7483_ gnd vdd FILL
XFILL_2__16333_ gnd vdd FILL
XFILL_2__7419_ gnd vdd FILL
XFILL_1__11206_ gnd vdd FILL
XFILL_3__14904_ gnd vdd FILL
XFILL_3__10027_ gnd vdd FILL
XFILL_2__13545_ gnd vdd FILL
XFILL_3__15884_ gnd vdd FILL
XFILL_2__8399_ gnd vdd FILL
XFILL_1__12186_ gnd vdd FILL
XFILL_0__11936_ gnd vdd FILL
XFILL_3__7192_ gnd vdd FILL
XFILL_0__14724_ gnd vdd FILL
XFILL_2__10757_ gnd vdd FILL
XSFILL89320x80050 gnd vdd FILL
XFILL_4__14105_ gnd vdd FILL
XFILL_0__9222_ gnd vdd FILL
XFILL_4__11317_ gnd vdd FILL
XFILL_3__14835_ gnd vdd FILL
XFILL_5__13656_ gnd vdd FILL
X_9850_ _9941_/B _8314_/B gnd _9851_/C vdd NAND2X1
XFILL_4__15085_ gnd vdd FILL
XSFILL3560x21050 gnd vdd FILL
XFILL_1__11137_ gnd vdd FILL
XFILL_2__16264_ gnd vdd FILL
XFILL_4__12297_ gnd vdd FILL
XFILL_2__13476_ gnd vdd FILL
XFILL_0__14655_ gnd vdd FILL
XFILL_2__10688_ gnd vdd FILL
XFILL_0__11867_ gnd vdd FILL
XFILL_5__7059_ gnd vdd FILL
XFILL_5__12607_ gnd vdd FILL
X_8801_ _8801_/Q _7411_/CLK _8801_/R vdd _8801_/D gnd vdd DFFSR
XFILL_4__14036_ gnd vdd FILL
XSFILL28760x33050 gnd vdd FILL
XFILL_0__9153_ gnd vdd FILL
XFILL_2__15215_ gnd vdd FILL
XFILL_5__16375_ gnd vdd FILL
XFILL_4__11248_ gnd vdd FILL
X_9781_ _9835_/Q gnd _9781_/Y vdd INVX1
XFILL_5__13587_ gnd vdd FILL
XFILL_2__12427_ gnd vdd FILL
XFILL_5__10799_ gnd vdd FILL
XFILL_3__14766_ gnd vdd FILL
X_6993_ _6982_/B _8401_/B gnd _6994_/C vdd NAND2X1
XSFILL54040x66050 gnd vdd FILL
XFILL_0__13606_ gnd vdd FILL
XFILL_2__16195_ gnd vdd FILL
XFILL_1__15945_ gnd vdd FILL
XFILL_3__11978_ gnd vdd FILL
XFILL_0__10818_ gnd vdd FILL
XFILL_1__11068_ gnd vdd FILL
XFILL_0__8104_ gnd vdd FILL
XFILL_0__14586_ gnd vdd FILL
XSFILL94440x71050 gnd vdd FILL
XFILL_5__15326_ gnd vdd FILL
XFILL_0__11798_ gnd vdd FILL
X_8732_ _8730_/Y _8695_/B _8731_/Y gnd _8732_/Y vdd OAI21X1
XFILL_3__13717_ gnd vdd FILL
XFILL_0__9084_ gnd vdd FILL
XFILL_3__9902_ gnd vdd FILL
XFILL_1__10019_ gnd vdd FILL
XFILL_3__10929_ gnd vdd FILL
XFILL_4__11179_ gnd vdd FILL
XFILL_2__15146_ gnd vdd FILL
XFILL_6_BUFX2_insert515 gnd vdd FILL
XFILL_2__12358_ gnd vdd FILL
XFILL_3__14697_ gnd vdd FILL
XFILL_0__16325_ gnd vdd FILL
XFILL_0__13537_ gnd vdd FILL
XFILL_0__10749_ gnd vdd FILL
XFILL_6_BUFX2_insert526 gnd vdd FILL
XFILL_1__15876_ gnd vdd FILL
XFILL_5__15257_ gnd vdd FILL
XFILL_5__12469_ gnd vdd FILL
X_8663_ _8663_/Q _8663_/CLK _7131_/R vdd _8663_/D gnd vdd DFFSR
XFILL_3__13648_ gnd vdd FILL
XFILL_2__11309_ gnd vdd FILL
XSFILL33880x24050 gnd vdd FILL
XFILL_4__15987_ gnd vdd FILL
XFILL_1__14827_ gnd vdd FILL
XFILL_2__15077_ gnd vdd FILL
XFILL_0__13468_ gnd vdd FILL
XFILL_2__12289_ gnd vdd FILL
XFILL_0__16256_ gnd vdd FILL
XFILL_5__14208_ gnd vdd FILL
X_7614_ _7662_/Q gnd _7614_/Y vdd INVX1
XSFILL74760x36050 gnd vdd FILL
XFILL_3__16367_ gnd vdd FILL
XFILL_5__15188_ gnd vdd FILL
XSFILL48920x46050 gnd vdd FILL
XFILL_2__14028_ gnd vdd FILL
XFILL_4__14938_ gnd vdd FILL
X_8594_ _8657_/A _8466_/B gnd _8595_/C vdd NAND2X1
XFILL_3__9764_ gnd vdd FILL
XFILL_0__15207_ gnd vdd FILL
XFILL_0__12419_ gnd vdd FILL
XFILL_3__13579_ gnd vdd FILL
XFILL_3__6976_ gnd vdd FILL
XFILL_0__16187_ gnd vdd FILL
XFILL_1__14758_ gnd vdd FILL
XSFILL74200x79050 gnd vdd FILL
XFILL_0__13399_ gnd vdd FILL
XFILL_3__15318_ gnd vdd FILL
XFILL_5__14139_ gnd vdd FILL
X_7545_ _7639_/Q gnd _7547_/A vdd INVX1
XFILL_3__8715_ gnd vdd FILL
XFILL_0__9986_ gnd vdd FILL
XSFILL79240x2050 gnd vdd FILL
XFILL_4__14869_ gnd vdd FILL
XFILL_3__16298_ gnd vdd FILL
XFILL_1__13709_ gnd vdd FILL
XFILL_0__15138_ gnd vdd FILL
XSFILL49000x55050 gnd vdd FILL
XFILL_6__15429_ gnd vdd FILL
XFILL_1__14689_ gnd vdd FILL
XFILL_1__7730_ gnd vdd FILL
XFILL_3__15249_ gnd vdd FILL
X_7476_ _7476_/A _7430_/A _7476_/C gnd _7530_/D vdd OAI21X1
XSFILL89400x60050 gnd vdd FILL
XFILL_3__8646_ gnd vdd FILL
XFILL_2__15979_ gnd vdd FILL
XFILL_0__15069_ gnd vdd FILL
X_9215_ _9215_/A gnd _9217_/A vdd INVX1
XFILL_0__8868_ gnd vdd FILL
XFILL_1__16359_ gnd vdd FILL
XFILL_3__8577_ gnd vdd FILL
XFILL_4__7370_ gnd vdd FILL
XSFILL28840x13050 gnd vdd FILL
XFILL_1__9400_ gnd vdd FILL
XFILL_0__7819_ gnd vdd FILL
X_9146_ _9144_/Y _9164_/B _9146_/C gnd _9196_/D vdd OAI21X1
XSFILL79720x8050 gnd vdd FILL
XSFILL54120x46050 gnd vdd FILL
XFILL_1__7592_ gnd vdd FILL
XFILL_3_BUFX2_insert405 gnd vdd FILL
XFILL_3_BUFX2_insert416 gnd vdd FILL
XFILL_3_BUFX2_insert427 gnd vdd FILL
XFILL_3_BUFX2_insert438 gnd vdd FILL
X_9077_ _9043_/A _9077_/CLK _8433_/R vdd _9077_/D gnd vdd DFFSR
XFILL_4__9040_ gnd vdd FILL
XFILL_3__7459_ gnd vdd FILL
XFILL_3_BUFX2_insert449 gnd vdd FILL
X_8028_ _7944_/A _8926_/CLK _7262_/R vdd _8028_/D gnd vdd DFFSR
XFILL_1__9262_ gnd vdd FILL
XFILL_1__8213_ gnd vdd FILL
XFILL_6__7099_ gnd vdd FILL
XSFILL18760x65050 gnd vdd FILL
XSFILL34040x13050 gnd vdd FILL
XFILL_3__9129_ gnd vdd FILL
XSFILL39000x5050 gnd vdd FILL
X_10930_ _12785_/A _12788_/A gnd _10930_/Y vdd NOR2X1
XFILL_1__8144_ gnd vdd FILL
X_9979_ _9979_/A _9979_/B _9978_/Y gnd _9979_/Y vdd OAI21X1
X_10861_ _10861_/Q _8429_/CLK _9203_/R vdd _10813_/Y gnd vdd DFFSR
XFILL_1__8075_ gnd vdd FILL
XFILL_4_CLKBUF1_insert206 gnd vdd FILL
X_12600_ _12600_/A gnd _12602_/A vdd INVX1
XFILL_4__9873_ gnd vdd FILL
XFILL_4_CLKBUF1_insert217 gnd vdd FILL
X_13580_ _13420_/C gnd _13865_/B vdd INVX8
X_10792_ _10792_/A _10792_/B _10791_/Y gnd _10854_/D vdd OAI21X1
XFILL_4__8824_ gnd vdd FILL
XSFILL54200x26050 gnd vdd FILL
XFILL_0_BUFX2_insert306 gnd vdd FILL
X_12531_ _12529_/Y vdd _12531_/C gnd _12565_/D vdd OAI21X1
XFILL_0_BUFX2_insert317 gnd vdd FILL
XFILL_0_BUFX2_insert328 gnd vdd FILL
XFILL_0_BUFX2_insert339 gnd vdd FILL
XSFILL79160x30050 gnd vdd FILL
XFILL_4__8755_ gnd vdd FILL
X_15250_ _15249_/Y _15247_/Y gnd _15250_/Y vdd NOR2X1
X_12462_ _12462_/A vdd _12461_/Y gnd _12542_/D vdd OAI21X1
XFILL_4__7706_ gnd vdd FILL
XFILL_1__8977_ gnd vdd FILL
X_14201_ _9701_/Q gnd _14203_/A vdd INVX1
X_11413_ _11411_/Y _11412_/Y _11334_/A gnd _11414_/C vdd OAI21X1
X_15181_ _8191_/A gnd _15182_/D vdd INVX1
X_12393_ _12391_/Y _12422_/A _12393_/C gnd _12393_/Y vdd OAI21X1
XFILL_1__7928_ gnd vdd FILL
XFILL_4__7637_ gnd vdd FILL
X_14132_ _8864_/A _14482_/B _13854_/B _9248_/A gnd _14132_/Y vdd AOI22X1
XSFILL18840x45050 gnd vdd FILL
X_11344_ _11762_/B gnd _11344_/Y vdd INVX8
XFILL_1__7859_ gnd vdd FILL
XFILL_4__7568_ gnd vdd FILL
XFILL_4_BUFX2_insert250 gnd vdd FILL
XSFILL99320x43050 gnd vdd FILL
X_14063_ _14063_/A _14055_/Y gnd _14074_/A vdd NAND2X1
XFILL_4_BUFX2_insert261 gnd vdd FILL
XSFILL69080x82050 gnd vdd FILL
XFILL_4__10550_ gnd vdd FILL
X_11275_ _11275_/A _11713_/C _11709_/A gnd _11275_/Y vdd AOI21X1
XFILL_5__8100_ gnd vdd FILL
XFILL_2__9371_ gnd vdd FILL
XFILL_4_BUFX2_insert272 gnd vdd FILL
XFILL_1__10370_ gnd vdd FILL
XFILL_4_BUFX2_insert283 gnd vdd FILL
X_13014_ _6891_/A gnd _13014_/Y vdd INVX1
XFILL_5__9080_ gnd vdd FILL
XFILL_4_BUFX2_insert294 gnd vdd FILL
XFILL_5_BUFX2_insert1007 gnd vdd FILL
XFILL_4__7499_ gnd vdd FILL
X_10226_ _10186_/A _7282_/CLK _7411_/R vdd _10226_/D gnd vdd DFFSR
XFILL_6__12090_ gnd vdd FILL
XFILL_2__8322_ gnd vdd FILL
XFILL_5_BUFX2_insert1018 gnd vdd FILL
XFILL_1__9529_ gnd vdd FILL
XFILL_5__11840_ gnd vdd FILL
XFILL_5_BUFX2_insert1029 gnd vdd FILL
XSFILL63560x22050 gnd vdd FILL
XFILL_2__11660_ gnd vdd FILL
XFILL_4__9238_ gnd vdd FILL
XSFILL64040x29050 gnd vdd FILL
XFILL_4__12220_ gnd vdd FILL
XFILL_3_BUFX2_insert950 gnd vdd FILL
X_10157_ _10140_/B _9517_/B gnd _10158_/C vdd NAND2X1
XFILL_3_BUFX2_insert961 gnd vdd FILL
XFILL_5__11771_ gnd vdd FILL
XFILL_2__8253_ gnd vdd FILL
XFILL_3_BUFX2_insert972 gnd vdd FILL
XFILL_1__12040_ gnd vdd FILL
XFILL_3_BUFX2_insert983 gnd vdd FILL
XFILL_2__11591_ gnd vdd FILL
XFILL_0__12770_ gnd vdd FILL
XFILL_4__9169_ gnd vdd FILL
XFILL_3_BUFX2_insert994 gnd vdd FILL
XFILL_5__13510_ gnd vdd FILL
XFILL_2__7204_ gnd vdd FILL
XFILL_5__14490_ gnd vdd FILL
XFILL_3__11901_ gnd vdd FILL
XFILL_4__12151_ gnd vdd FILL
X_10088_ _15797_/A _7400_/CLK _9704_/R vdd _10088_/D gnd vdd DFFSR
X_14965_ _8275_/A _14323_/B _14065_/C _16305_/A gnd _14976_/A vdd AOI22X1
XFILL_2__13330_ gnd vdd FILL
XFILL_2__8184_ gnd vdd FILL
XFILL_2__10542_ gnd vdd FILL
XFILL_3__12881_ gnd vdd FILL
XFILL_0__11721_ gnd vdd FILL
XFILL_6__14800_ gnd vdd FILL
XFILL_4__11102_ gnd vdd FILL
XFILL_5__9982_ gnd vdd FILL
X_13916_ _14700_/A _15445_/D _14711_/B _13915_/Y gnd _13917_/A vdd OAI22X1
XFILL_3__14620_ gnd vdd FILL
XFILL_5__13441_ gnd vdd FILL
XFILL_5__10653_ gnd vdd FILL
XFILL_4__12082_ gnd vdd FILL
XFILL_3_BUFX2_insert1000 gnd vdd FILL
X_14896_ _9204_/Q gnd _16264_/A vdd INVX1
XFILL_3__11832_ gnd vdd FILL
XFILL_2__13261_ gnd vdd FILL
XFILL_3_BUFX2_insert1011 gnd vdd FILL
XFILL_0__14440_ gnd vdd FILL
XFILL_0__11652_ gnd vdd FILL
XSFILL53480x74050 gnd vdd FILL
XFILL_3_BUFX2_insert1022 gnd vdd FILL
XFILL_1__13991_ gnd vdd FILL
XFILL_3_BUFX2_insert1033 gnd vdd FILL
X_13847_ _13847_/A _13846_/Y gnd _13852_/C vdd NOR2X1
XFILL_4__15910_ gnd vdd FILL
XFILL_5__13372_ gnd vdd FILL
XFILL_2__15000_ gnd vdd FILL
XFILL_5__16160_ gnd vdd FILL
XFILL_4__11033_ gnd vdd FILL
XFILL_3_BUFX2_insert1044 gnd vdd FILL
XFILL_3__14551_ gnd vdd FILL
XFILL_2__12212_ gnd vdd FILL
XFILL_1__15730_ gnd vdd FILL
XFILL_3_BUFX2_insert1055 gnd vdd FILL
XFILL_2__7066_ gnd vdd FILL
XFILL_3__11763_ gnd vdd FILL
XFILL_3_BUFX2_insert1066 gnd vdd FILL
XFILL_0__14371_ gnd vdd FILL
XFILL_5__8864_ gnd vdd FILL
XFILL_5__12323_ gnd vdd FILL
XFILL_0__11583_ gnd vdd FILL
XFILL_5__15111_ gnd vdd FILL
XFILL_3__13502_ gnd vdd FILL
XSFILL59000x18050 gnd vdd FILL
X_13778_ _13777_/Y _13857_/B _13633_/C _13776_/Y gnd _13778_/Y vdd OAI22X1
XFILL_3_BUFX2_insert1088 gnd vdd FILL
XFILL_5__16091_ gnd vdd FILL
XFILL_4__15841_ gnd vdd FILL
XFILL_0__13322_ gnd vdd FILL
XFILL_3__14482_ gnd vdd FILL
XFILL_0__16110_ gnd vdd FILL
XFILL_2__12143_ gnd vdd FILL
XFILL_0__10534_ gnd vdd FILL
XFILL_1__15661_ gnd vdd FILL
XFILL_6__16401_ gnd vdd FILL
XFILL_3__11694_ gnd vdd FILL
XFILL_5__7815_ gnd vdd FILL
XSFILL99400x23050 gnd vdd FILL
XFILL_6__13613_ gnd vdd FILL
XSFILL69160x62050 gnd vdd FILL
X_15517_ _16235_/A _15517_/B _15516_/Y _15633_/D gnd _15518_/B vdd OAI22X1
XFILL_1__12873_ gnd vdd FILL
X_12729_ _12762_/A memoryOutData[11] gnd _12730_/C vdd NAND2X1
XFILL_3__16221_ gnd vdd FILL
XFILL_5__15042_ gnd vdd FILL
XFILL_5__12254_ gnd vdd FILL
XFILL_3__13433_ gnd vdd FILL
XFILL_1__14612_ gnd vdd FILL
XFILL_0__16041_ gnd vdd FILL
XFILL_2__12074_ gnd vdd FILL
XFILL_4__12984_ gnd vdd FILL
XFILL_4__15772_ gnd vdd FILL
XFILL_3__10645_ gnd vdd FILL
XFILL_0__13253_ gnd vdd FILL
XFILL_1__11824_ gnd vdd FILL
XFILL_5__7746_ gnd vdd FILL
XFILL_5__11205_ gnd vdd FILL
XFILL_1__15592_ gnd vdd FILL
X_15448_ _8209_/A gnd _15448_/Y vdd INVX1
XFILL_0_BUFX2_insert840 gnd vdd FILL
XSFILL104360x71050 gnd vdd FILL
XFILL_2__15902_ gnd vdd FILL
XFILL_5__12185_ gnd vdd FILL
XFILL_4__11935_ gnd vdd FILL
XFILL_0_BUFX2_insert851 gnd vdd FILL
XFILL_4__14723_ gnd vdd FILL
XFILL_2__11025_ gnd vdd FILL
XFILL_3__16152_ gnd vdd FILL
XFILL_3__13364_ gnd vdd FILL
XFILL_0_BUFX2_insert862 gnd vdd FILL
XFILL_0__12204_ gnd vdd FILL
XFILL_2__7968_ gnd vdd FILL
XFILL_1__14543_ gnd vdd FILL
XFILL_0_BUFX2_insert873 gnd vdd FILL
XFILL_3__10576_ gnd vdd FILL
XFILL_1__11755_ gnd vdd FILL
XSFILL74280x53050 gnd vdd FILL
X_7330_ _7330_/A _7308_/A _7329_/Y gnd _7396_/D vdd OAI21X1
XFILL_6__16263_ gnd vdd FILL
XFILL_0__10396_ gnd vdd FILL
XFILL_0_BUFX2_insert884 gnd vdd FILL
XFILL_5__7677_ gnd vdd FILL
XFILL_5__11136_ gnd vdd FILL
XFILL_3__15103_ gnd vdd FILL
X_15379_ _15379_/A _15378_/Y _15379_/C gnd _15381_/C vdd NOR3X1
XFILL_0_BUFX2_insert895 gnd vdd FILL
XFILL_3__12315_ gnd vdd FILL
XFILL_0__9771_ gnd vdd FILL
XFILL_3__8500_ gnd vdd FILL
XFILL_6__10687_ gnd vdd FILL
XFILL_3_BUFX2_insert11 gnd vdd FILL
XFILL_2__15833_ gnd vdd FILL
XFILL_4__11866_ gnd vdd FILL
XFILL_2__6919_ gnd vdd FILL
XFILL_1_BUFX2_insert1070 gnd vdd FILL
XFILL_4__14654_ gnd vdd FILL
XFILL_3__16083_ gnd vdd FILL
XFILL_0__6983_ gnd vdd FILL
XFILL_3__13295_ gnd vdd FILL
XFILL_3__9480_ gnd vdd FILL
XFILL_0__12135_ gnd vdd FILL
XFILL_5__9416_ gnd vdd FILL
XFILL_3_BUFX2_insert22 gnd vdd FILL
XFILL_1__10706_ gnd vdd FILL
XFILL_1__14474_ gnd vdd FILL
XFILL_6__15214_ gnd vdd FILL
XFILL_1__11686_ gnd vdd FILL
XFILL_3_BUFX2_insert33 gnd vdd FILL
XFILL_1_BUFX2_insert1092 gnd vdd FILL
XFILL_0__8722_ gnd vdd FILL
X_7261_ _7261_/Q _7261_/CLK _8669_/R vdd _7261_/D gnd vdd DFFSR
XFILL_4__13605_ gnd vdd FILL
XFILL_5__15944_ gnd vdd FILL
XFILL_3__15034_ gnd vdd FILL
XFILL_3_BUFX2_insert44 gnd vdd FILL
XFILL_4__10817_ gnd vdd FILL
XFILL_5__11067_ gnd vdd FILL
XFILL_2__9638_ gnd vdd FILL
XFILL_1__16213_ gnd vdd FILL
XFILL_3_BUFX2_insert55 gnd vdd FILL
XFILL_4__14585_ gnd vdd FILL
XFILL_3__12246_ gnd vdd FILL
XSFILL3560x16050 gnd vdd FILL
XFILL_1__10637_ gnd vdd FILL
XFILL_1__13425_ gnd vdd FILL
XFILL_3_BUFX2_insert66 gnd vdd FILL
XFILL_2__15764_ gnd vdd FILL
XFILL_4__11797_ gnd vdd FILL
X_9000_ _8998_/Y _8961_/B _9000_/C gnd _9062_/D vdd OAI21X1
XFILL_2__12976_ gnd vdd FILL
XFILL_5__9347_ gnd vdd FILL
XFILL_3_BUFX2_insert77 gnd vdd FILL
XFILL_0__12066_ gnd vdd FILL
XFILL_5__10018_ gnd vdd FILL
XFILL_3_BUFX2_insert88 gnd vdd FILL
XSFILL3800x78050 gnd vdd FILL
XFILL_0__8653_ gnd vdd FILL
XFILL_6__12357_ gnd vdd FILL
XFILL_4__16324_ gnd vdd FILL
XFILL_4__13536_ gnd vdd FILL
X_7192_ _7202_/B _6936_/B gnd _7193_/C vdd NAND2X1
XFILL_3_BUFX2_insert99 gnd vdd FILL
XFILL_2__14715_ gnd vdd FILL
XSFILL28760x28050 gnd vdd FILL
XFILL_4__10748_ gnd vdd FILL
XFILL_5__15875_ gnd vdd FILL
XFILL_2__11927_ gnd vdd FILL
XFILL_3__8362_ gnd vdd FILL
XFILL_3__12177_ gnd vdd FILL
XFILL_0__11017_ gnd vdd FILL
XFILL_1__16144_ gnd vdd FILL
XFILL_1__13356_ gnd vdd FILL
XFILL_2__15695_ gnd vdd FILL
XFILL_1__10568_ gnd vdd FILL
XFILL_5__9278_ gnd vdd FILL
XFILL_6__11308_ gnd vdd FILL
XFILL_0__7604_ gnd vdd FILL
XFILL_5__14826_ gnd vdd FILL
XFILL_6__15076_ gnd vdd FILL
XSFILL43800x31050 gnd vdd FILL
XFILL_0__8584_ gnd vdd FILL
XSFILL94440x66050 gnd vdd FILL
XFILL_4__13467_ gnd vdd FILL
XFILL_3__11128_ gnd vdd FILL
XFILL_3__7313_ gnd vdd FILL
XFILL_4__16255_ gnd vdd FILL
XFILL_4__10679_ gnd vdd FILL
XSFILL68600x76050 gnd vdd FILL
XFILL_2__14646_ gnd vdd FILL
XFILL_1__12307_ gnd vdd FILL
XFILL_5__8229_ gnd vdd FILL
XFILL_1__13287_ gnd vdd FILL
XFILL_0__15825_ gnd vdd FILL
XFILL_1__16075_ gnd vdd FILL
XFILL_2__11858_ gnd vdd FILL
XFILL_1__10499_ gnd vdd FILL
XFILL_6__14027_ gnd vdd FILL
XFILL_6_CLKBUF1_insert183 gnd vdd FILL
XFILL_4__15206_ gnd vdd FILL
XFILL_4__12418_ gnd vdd FILL
XFILL_4__16186_ gnd vdd FILL
XSFILL69240x42050 gnd vdd FILL
XFILL_5__14757_ gnd vdd FILL
XFILL_3__7244_ gnd vdd FILL
XFILL_4__13398_ gnd vdd FILL
XFILL_1__15026_ gnd vdd FILL
XFILL_3__15936_ gnd vdd FILL
XFILL_5__11969_ gnd vdd FILL
XFILL_2__10809_ gnd vdd FILL
XFILL_1__12238_ gnd vdd FILL
XFILL_3__11059_ gnd vdd FILL
XSFILL33880x19050 gnd vdd FILL
XFILL_2__14577_ gnd vdd FILL
XFILL_2__11789_ gnd vdd FILL
XFILL_0__15756_ gnd vdd FILL
XFILL_5__13708_ gnd vdd FILL
XFILL_4__15137_ gnd vdd FILL
XFILL_0__12968_ gnd vdd FILL
X_9902_ _9900_/Y _9902_/B _9901_/Y gnd _9902_/Y vdd OAI21X1
XFILL_4__12349_ gnd vdd FILL
XFILL_2__16316_ gnd vdd FILL
XFILL_0__7466_ gnd vdd FILL
XFILL_5__14688_ gnd vdd FILL
XFILL_2__13528_ gnd vdd FILL
XFILL_0__14707_ gnd vdd FILL
XFILL_1__12169_ gnd vdd FILL
XFILL_3__15867_ gnd vdd FILL
XFILL_3__7175_ gnd vdd FILL
XSFILL104440x51050 gnd vdd FILL
XFILL_0__11919_ gnd vdd FILL
XFILL_0__15687_ gnd vdd FILL
XFILL_0__12899_ gnd vdd FILL
XFILL_5__13639_ gnd vdd FILL
XFILL_4__15068_ gnd vdd FILL
X_9833_ _9833_/Q _7664_/CLK _7920_/R vdd _9777_/Y gnd vdd DFFSR
XFILL_3__14818_ gnd vdd FILL
XFILL_2__16247_ gnd vdd FILL
XFILL_2__13459_ gnd vdd FILL
XFILL_3__15798_ gnd vdd FILL
XFILL_0__14638_ gnd vdd FILL
XFILL_4__14019_ gnd vdd FILL
XFILL_0__9136_ gnd vdd FILL
XFILL_5__16358_ gnd vdd FILL
X_9764_ _9764_/A _8228_/B gnd _9765_/C vdd NAND2X1
XFILL_3__14749_ gnd vdd FILL
X_6976_ _6974_/Y _6988_/B _6976_/C gnd _7022_/D vdd OAI21X1
XFILL_6_BUFX2_insert301 gnd vdd FILL
XFILL_1__15928_ gnd vdd FILL
XFILL_2__16178_ gnd vdd FILL
XFILL_0__14569_ gnd vdd FILL
XFILL_5__15309_ gnd vdd FILL
X_8715_ _8715_/A gnd _8717_/A vdd INVX1
XFILL_5__16289_ gnd vdd FILL
XFILL_2__15129_ gnd vdd FILL
XFILL_0__16308_ gnd vdd FILL
X_9695_ _9695_/Q _9716_/CLK _8682_/R vdd _9695_/D gnd vdd DFFSR
XFILL_4__6870_ gnd vdd FILL
XFILL_1__15859_ gnd vdd FILL
XFILL_6_BUFX2_insert367 gnd vdd FILL
XFILL_1__8900_ gnd vdd FILL
XFILL_0__8018_ gnd vdd FILL
XFILL_1__9880_ gnd vdd FILL
X_8646_ _8646_/A _8609_/A _8646_/C gnd _8646_/Y vdd OAI21X1
XFILL_0__16239_ gnd vdd FILL
XSFILL13640x50050 gnd vdd FILL
XFILL_1__8831_ gnd vdd FILL
XSFILL79880x64050 gnd vdd FILL
X_8577_ _8575_/Y _8577_/B _8576_/Y gnd _8577_/Y vdd OAI21X1
XFILL_3__9747_ gnd vdd FILL
XFILL_3__6959_ gnd vdd FILL
XFILL_1__8762_ gnd vdd FILL
X_7528_ _7468_/A _7527_/CLK _8935_/R vdd _7528_/D gnd vdd DFFSR
XFILL_3__9678_ gnd vdd FILL
XFILL_4__8471_ gnd vdd FILL
XFILL_1__7713_ gnd vdd FILL
X_7459_ _7459_/A gnd _7461_/A vdd INVX1
XFILL_3__8629_ gnd vdd FILL
XSFILL104520x31050 gnd vdd FILL
XFILL_4__7422_ gnd vdd FILL
XSFILL89880x9050 gnd vdd FILL
XFILL_4__7353_ gnd vdd FILL
X_11060_ _12274_/Y _12159_/Y gnd _11060_/Y vdd NOR2X1
X_9129_ _9191_/Q gnd _9129_/Y vdd INVX1
XFILL_1__7575_ gnd vdd FILL
X_10011_ _9993_/A _8987_/B gnd _10012_/C vdd NAND2X1
XFILL_3_BUFX2_insert235 gnd vdd FILL
XFILL_3_BUFX2_insert246 gnd vdd FILL
XFILL_3_BUFX2_insert257 gnd vdd FILL
XFILL_4__9023_ gnd vdd FILL
XFILL_3_BUFX2_insert268 gnd vdd FILL
XFILL111960x73050 gnd vdd FILL
XFILL_3_BUFX2_insert279 gnd vdd FILL
XFILL_2_BUFX2_insert902 gnd vdd FILL
XFILL_1__9245_ gnd vdd FILL
XFILL_2_BUFX2_insert913 gnd vdd FILL
XFILL_2_BUFX2_insert924 gnd vdd FILL
XSFILL13720x30050 gnd vdd FILL
XFILL_2_BUFX2_insert935 gnd vdd FILL
XFILL_2_BUFX2_insert946 gnd vdd FILL
X_14750_ _10311_/A gnd _14750_/Y vdd INVX1
XSFILL79160x25050 gnd vdd FILL
X_11962_ _13200_/Q gnd _11962_/Y vdd INVX1
XFILL_2_BUFX2_insert957 gnd vdd FILL
XFILL_2_BUFX2_insert968 gnd vdd FILL
XFILL_2_BUFX2_insert979 gnd vdd FILL
X_13701_ _14887_/B _13701_/B _13574_/C _15283_/D gnd _13705_/A vdd OAI22X1
X_10913_ _10920_/B _10938_/B gnd _10913_/Y vdd NOR2X1
XFILL_1__8127_ gnd vdd FILL
X_14681_ _8559_/Q gnd _16083_/B vdd INVX1
X_11893_ _13085_/A gnd _11895_/A vdd INVX1
X_16420_ _13594_/A _8537_/CLK _9054_/R vdd _16332_/Y gnd vdd DFFSR
XFILL_4__9925_ gnd vdd FILL
X_13632_ _8025_/Q gnd _13632_/Y vdd INVX1
X_10844_ _10844_/Q _9436_/CLK _8156_/R vdd _10844_/D gnd vdd DFFSR
XSFILL84280x16050 gnd vdd FILL
XFILL_1__8058_ gnd vdd FILL
XFILL_4__9856_ gnd vdd FILL
X_16351_ _15482_/A gnd _16353_/A vdd INVX1
XBUFX2_insert901 _15072_/Y gnd _16261_/D vdd BUFX2
XFILL_0_BUFX2_insert103 gnd vdd FILL
XBUFX2_insert912 _12360_/Y gnd _9478_/B vdd BUFX2
XSFILL53800x1050 gnd vdd FILL
X_13563_ _15149_/A _14071_/B _14897_/D _13562_/Y gnd _13567_/A vdd OAI22X1
X_10775_ _15509_/A gnd _10777_/A vdd INVX1
XSFILL99320x38050 gnd vdd FILL
XBUFX2_insert923 _13370_/Y gnd _14065_/C vdd BUFX2
XFILL_2__8871_ gnd vdd FILL
XFILL_5__7600_ gnd vdd FILL
X_15302_ _15302_/A _15302_/B gnd _15303_/C vdd NOR2X1
XBUFX2_insert934 _12435_/Y gnd _7889_/B vdd BUFX2
XFILL_4__9787_ gnd vdd FILL
XFILL_5__8580_ gnd vdd FILL
X_12514_ _12418_/A gnd _12516_/A vdd INVX1
XBUFX2_insert945 _11987_/Y gnd _12025_/B vdd BUFX2
XBUFX2_insert956 _13365_/Y gnd _10792_/B vdd BUFX2
X_16282_ _16282_/A _16281_/Y gnd _16283_/B vdd NOR2X1
XFILL_2__7822_ gnd vdd FILL
XBUFX2_insert967 _12417_/Y gnd _7359_/B vdd BUFX2
XFILL_3__10430_ gnd vdd FILL
X_13494_ _14865_/B gnd _13494_/Y vdd INVX8
XBUFX2_insert978 _16451_/Y gnd _13173_/A vdd BUFX2
XFILL_0__10250_ gnd vdd FILL
XFILL_4__8738_ gnd vdd FILL
X_15233_ _16002_/C _15232_/Y _15233_/C _15912_/D gnd _15234_/C vdd OAI22X1
XBUFX2_insert989 _13351_/Y gnd _10024_/B vdd BUFX2
X_12445_ _12349_/A gnd _12447_/A vdd INVX1
XFILL_4__11720_ gnd vdd FILL
XFILL_3__10361_ gnd vdd FILL
XFILL_1__11540_ gnd vdd FILL
XFILL_2__7753_ gnd vdd FILL
XFILL_5__7462_ gnd vdd FILL
XFILL_0__10181_ gnd vdd FILL
XFILL_6__13260_ gnd vdd FILL
XFILL_3__12100_ gnd vdd FILL
XSFILL13800x10050 gnd vdd FILL
X_15164_ _15162_/Y _15164_/B gnd _15164_/Y vdd NOR2X1
X_12376_ _12031_/B gnd _12376_/Y vdd INVX1
XFILL_4__11651_ gnd vdd FILL
XFILL_3__13080_ gnd vdd FILL
XFILL_5__13990_ gnd vdd FILL
XFILL_2__12830_ gnd vdd FILL
XFILL_2__7684_ gnd vdd FILL
XFILL_1__11471_ gnd vdd FILL
XFILL_3__10292_ gnd vdd FILL
XFILL112120x62050 gnd vdd FILL
X_14115_ _14115_/A _14768_/D _14342_/B _14115_/D gnd _14115_/Y vdd OAI22X1
X_11327_ _11181_/Y _11494_/A _11175_/Y gnd _11327_/Y vdd AOI21X1
XFILL_2__9423_ gnd vdd FILL
XFILL_3__12031_ gnd vdd FILL
XFILL_4__14370_ gnd vdd FILL
X_15095_ _15095_/A _15565_/B _15569_/C _15095_/D gnd _15095_/Y vdd OAI22X1
XFILL_1__10422_ gnd vdd FILL
XFILL_1__13210_ gnd vdd FILL
XFILL_4__11582_ gnd vdd FILL
XFILL_2__12761_ gnd vdd FILL
XFILL_1__14190_ gnd vdd FILL
XFILL_5__9132_ gnd vdd FILL
XFILL_0__13940_ gnd vdd FILL
XFILL_4__13321_ gnd vdd FILL
X_14046_ _14046_/A _14046_/B _14040_/Y gnd _14046_/Y vdd NOR3X1
XFILL_6__12142_ gnd vdd FILL
XFILL_4__10533_ gnd vdd FILL
XFILL_2__14500_ gnd vdd FILL
XFILL_5__15660_ gnd vdd FILL
X_11258_ _11044_/A _11641_/C gnd _11258_/Y vdd NAND2X1
XSFILL4360x59050 gnd vdd FILL
XFILL_2__9354_ gnd vdd FILL
XFILL_5__12872_ gnd vdd FILL
XFILL_1__13141_ gnd vdd FILL
XFILL_2__11712_ gnd vdd FILL
XFILL_2__15480_ gnd vdd FILL
XSFILL43720x46050 gnd vdd FILL
XFILL_0__13871_ gnd vdd FILL
XFILL_4__16040_ gnd vdd FILL
XFILL_5__14611_ gnd vdd FILL
X_10209_ _13994_/A _8560_/CLK _9313_/R vdd _10209_/D gnd vdd DFFSR
XFILL_4__13252_ gnd vdd FILL
XFILL_5__11823_ gnd vdd FILL
XFILL_5__15591_ gnd vdd FILL
X_11189_ _11494_/A _11186_/Y _11189_/C gnd _11189_/Y vdd OAI21X1
XFILL_2__14431_ gnd vdd FILL
XFILL_5__8014_ gnd vdd FILL
XFILL_3__13982_ gnd vdd FILL
XFILL_2__9285_ gnd vdd FILL
XFILL_2__11643_ gnd vdd FILL
XFILL_0__15610_ gnd vdd FILL
XFILL_1__10284_ gnd vdd FILL
XSFILL99400x18050 gnd vdd FILL
XSFILL69160x57050 gnd vdd FILL
XFILL_4__12203_ gnd vdd FILL
XFILL_0__7320_ gnd vdd FILL
XFILL_3_BUFX2_insert780 gnd vdd FILL
XFILL_5__14542_ gnd vdd FILL
XFILL_3_BUFX2_insert791 gnd vdd FILL
X_15997_ _15920_/C _14577_/Y _15997_/C _15915_/C gnd _15997_/Y vdd OAI22X1
XFILL_3__15721_ gnd vdd FILL
XFILL_5__11754_ gnd vdd FILL
XFILL_1__12023_ gnd vdd FILL
XFILL_2__8236_ gnd vdd FILL
XFILL_4__10395_ gnd vdd FILL
XFILL_2__14362_ gnd vdd FILL
XFILL_0__12753_ gnd vdd FILL
XSFILL84200x60050 gnd vdd FILL
XFILL_0__15541_ gnd vdd FILL
XFILL_2__11574_ gnd vdd FILL
XFILL_4__12134_ gnd vdd FILL
XFILL_2__16101_ gnd vdd FILL
X_14948_ _8019_/A gnd _14949_/D vdd INVX1
XFILL_5__10705_ gnd vdd FILL
XFILL_0__7251_ gnd vdd FILL
XFILL_2__13313_ gnd vdd FILL
XFILL_3__15652_ gnd vdd FILL
XFILL_5__14473_ gnd vdd FILL
XSFILL104360x66050 gnd vdd FILL
XFILL_5__11685_ gnd vdd FILL
XFILL_0__11704_ gnd vdd FILL
XFILL_2__10525_ gnd vdd FILL
XFILL_3__12864_ gnd vdd FILL
XFILL_2__14293_ gnd vdd FILL
XFILL_5__16212_ gnd vdd FILL
XFILL_0__15472_ gnd vdd FILL
XFILL_0__7182_ gnd vdd FILL
XFILL_5__10636_ gnd vdd FILL
XFILL_3__14603_ gnd vdd FILL
XFILL_5__13424_ gnd vdd FILL
XFILL_2__7118_ gnd vdd FILL
X_14879_ _14877_/Y _14879_/B _14879_/C gnd _14879_/Y vdd NAND3X1
XFILL_2__16032_ gnd vdd FILL
XFILL_4__12065_ gnd vdd FILL
XFILL_3__11815_ gnd vdd FILL
XFILL_2__13244_ gnd vdd FILL
XFILL_3__15583_ gnd vdd FILL
XFILL_2__8098_ gnd vdd FILL
XFILL_3__8980_ gnd vdd FILL
XFILL_0__11635_ gnd vdd FILL
XFILL_0__14423_ gnd vdd FILL
XFILL_1__13974_ gnd vdd FILL
XFILL_5__8916_ gnd vdd FILL
XFILL_5__16143_ gnd vdd FILL
XFILL_4__11016_ gnd vdd FILL
XFILL_5__13355_ gnd vdd FILL
XFILL_5__9896_ gnd vdd FILL
XFILL_3__14534_ gnd vdd FILL
XFILL_5__10567_ gnd vdd FILL
XFILL_1__15713_ gnd vdd FILL
XFILL_2__7049_ gnd vdd FILL
XFILL112200x42050 gnd vdd FILL
XFILL_3__11746_ gnd vdd FILL
XFILL_3__7931_ gnd vdd FILL
XFILL_0__14354_ gnd vdd FILL
XFILL_2__10387_ gnd vdd FILL
XFILL_0__11566_ gnd vdd FILL
XFILL_5__8847_ gnd vdd FILL
XFILL_5__12306_ gnd vdd FILL
X_8500_ _8500_/A _8496_/A _8500_/C gnd _8554_/D vdd OAI21X1
XFILL_5__13286_ gnd vdd FILL
XFILL_4__15824_ gnd vdd FILL
XFILL_5__16074_ gnd vdd FILL
XFILL_0__13305_ gnd vdd FILL
XFILL_3__14465_ gnd vdd FILL
XFILL_2__12126_ gnd vdd FILL
X_9480_ _9564_/Q gnd _9482_/A vdd INVX1
XFILL_5__10498_ gnd vdd FILL
XFILL_3__7862_ gnd vdd FILL
XFILL_1__15644_ gnd vdd FILL
XFILL_3__11677_ gnd vdd FILL
XFILL_0__10517_ gnd vdd FILL
XFILL_5_BUFX2_insert308 gnd vdd FILL
XFILL_1__12856_ gnd vdd FILL
XFILL_0__14285_ gnd vdd FILL
XFILL_3__16204_ gnd vdd FILL
XFILL_5__8778_ gnd vdd FILL
XFILL_5__15025_ gnd vdd FILL
XFILL_5_BUFX2_insert319 gnd vdd FILL
XFILL_5__12237_ gnd vdd FILL
XFILL_0__11497_ gnd vdd FILL
XFILL_3__9601_ gnd vdd FILL
XFILL_3__13416_ gnd vdd FILL
X_8431_ _8385_/A _9716_/CLK _8431_/R vdd _8387_/Y gnd vdd DFFSR
XSFILL43800x26050 gnd vdd FILL
XFILL_3__10628_ gnd vdd FILL
XFILL_4__15755_ gnd vdd FILL
XFILL_0__13236_ gnd vdd FILL
XFILL_0__16024_ gnd vdd FILL
XFILL_2__12057_ gnd vdd FILL
XFILL_3__14396_ gnd vdd FILL
XFILL_1__11807_ gnd vdd FILL
XFILL_4__12967_ gnd vdd FILL
XFILL_5__7729_ gnd vdd FILL
XFILL_0__10448_ gnd vdd FILL
XFILL_1__15575_ gnd vdd FILL
XFILL_1__12787_ gnd vdd FILL
XSFILL53960x70050 gnd vdd FILL
XFILL_0_BUFX2_insert670 gnd vdd FILL
XFILL_4__14706_ gnd vdd FILL
XFILL_5__12168_ gnd vdd FILL
XFILL_0_BUFX2_insert681 gnd vdd FILL
X_8362_ _8365_/A _7594_/B gnd _8362_/Y vdd NAND2X1
XFILL_3__16135_ gnd vdd FILL
XFILL_3__9532_ gnd vdd FILL
XFILL_3__13347_ gnd vdd FILL
XFILL_4__11918_ gnd vdd FILL
XFILL_0_BUFX2_insert692 gnd vdd FILL
XFILL_2__11008_ gnd vdd FILL
XFILL_3__10559_ gnd vdd FILL
XFILL_4__15686_ gnd vdd FILL
XFILL_1__14526_ gnd vdd FILL
XSFILL69240x37050 gnd vdd FILL
XFILL_4__12898_ gnd vdd FILL
XFILL_0__13167_ gnd vdd FILL
XFILL_1__11738_ gnd vdd FILL
XFILL_0__10379_ gnd vdd FILL
XFILL_5__11119_ gnd vdd FILL
X_7313_ _7391_/Q gnd _7315_/A vdd INVX1
XFILL_0__9754_ gnd vdd FILL
X_8293_ _8293_/Q _8025_/CLK _8025_/R vdd _8229_/Y gnd vdd DFFSR
XFILL_0__6966_ gnd vdd FILL
XFILL_4__14637_ gnd vdd FILL
XFILL_5__12099_ gnd vdd FILL
XFILL_2__15816_ gnd vdd FILL
XFILL_3__16066_ gnd vdd FILL
XFILL_4__11849_ gnd vdd FILL
XFILL_3__13278_ gnd vdd FILL
XFILL_3__9463_ gnd vdd FILL
XFILL_0__12118_ gnd vdd FILL
XFILL_1__14457_ gnd vdd FILL
XFILL_0__8705_ gnd vdd FILL
XFILL_0__13098_ gnd vdd FILL
XFILL_1__11669_ gnd vdd FILL
XFILL_6__9172_ gnd vdd FILL
X_7244_ _7242_/Y _7168_/A _7244_/C gnd _7244_/Y vdd OAI21X1
XFILL_5__15927_ gnd vdd FILL
XFILL_3__15017_ gnd vdd FILL
XFILL_0__9685_ gnd vdd FILL
XFILL_3__12229_ gnd vdd FILL
XFILL_4__14568_ gnd vdd FILL
XFILL_1__13408_ gnd vdd FILL
XSFILL8680x44050 gnd vdd FILL
XFILL_2__15747_ gnd vdd FILL
XFILL_0__6897_ gnd vdd FILL
XFILL_6__8123_ gnd vdd FILL
XFILL_0__12049_ gnd vdd FILL
XFILL_3__9394_ gnd vdd FILL
XFILL_2__12959_ gnd vdd FILL
XFILL_1__14388_ gnd vdd FILL
XFILL_0__8636_ gnd vdd FILL
XFILL_4__16307_ gnd vdd FILL
X_7175_ _7173_/Y _7166_/B _7175_/C gnd _7259_/D vdd OAI21X1
XFILL_4__13519_ gnd vdd FILL
XFILL_5__15858_ gnd vdd FILL
XFILL_4__14499_ gnd vdd FILL
XFILL_3__8345_ gnd vdd FILL
XFILL_1__16127_ gnd vdd FILL
XFILL_1__13339_ gnd vdd FILL
XFILL_2__15678_ gnd vdd FILL
XFILL_5__14809_ gnd vdd FILL
XFILL_0__8567_ gnd vdd FILL
XFILL_1__7360_ gnd vdd FILL
XFILL_4__16238_ gnd vdd FILL
XFILL_2__14629_ gnd vdd FILL
XFILL_5__15789_ gnd vdd FILL
XFILL_0__15808_ gnd vdd FILL
XFILL_3__8276_ gnd vdd FILL
XFILL_1__16058_ gnd vdd FILL
XFILL_3__7227_ gnd vdd FILL
XFILL_3__15919_ gnd vdd FILL
XFILL_4__16169_ gnd vdd FILL
XFILL_1__15009_ gnd vdd FILL
XFILL_0__8498_ gnd vdd FILL
XFILL_1__7291_ gnd vdd FILL
XFILL_0__15739_ gnd vdd FILL
XSFILL13640x45050 gnd vdd FILL
XFILL_1__9030_ gnd vdd FILL
XFILL_0__7449_ gnd vdd FILL
XFILL_3__7158_ gnd vdd FILL
XSFILL54520x57050 gnd vdd FILL
XFILL_1_BUFX2_insert909 gnd vdd FILL
X_9816_ _9816_/Q _7515_/CLK _7515_/R vdd _9816_/D gnd vdd DFFSR
XFILL_6__8956_ gnd vdd FILL
XFILL_4__7971_ gnd vdd FILL
XFILL_3__7089_ gnd vdd FILL
XFILL_0__9119_ gnd vdd FILL
X_9747_ _9745_/Y _9798_/B _9747_/C gnd _9823_/D vdd OAI21X1
XFILL_4__6922_ gnd vdd FILL
X_6959_ _6959_/A gnd _6959_/Y vdd INVX1
XSFILL104520x26050 gnd vdd FILL
XSFILL114680x70050 gnd vdd FILL
XFILL_1__9932_ gnd vdd FILL
XSFILL33800x58050 gnd vdd FILL
X_9678_ _9639_/A _8654_/B gnd _9678_/Y vdd NAND2X1
XFILL_4__9641_ gnd vdd FILL
XFILL_4__6853_ gnd vdd FILL
X_10560_ _10560_/A _10511_/A _10560_/C gnd _10606_/D vdd OAI21X1
X_8629_ _8683_/Q gnd _8631_/A vdd INVX1
XFILL_1__9863_ gnd vdd FILL
XSFILL33400x60050 gnd vdd FILL
XFILL_5_BUFX2_insert820 gnd vdd FILL
XFILL_5_BUFX2_insert831 gnd vdd FILL
XFILL_6__9508_ gnd vdd FILL
XFILL_5_BUFX2_insert842 gnd vdd FILL
XFILL_5_BUFX2_insert853 gnd vdd FILL
XFILL_5_BUFX2_insert864 gnd vdd FILL
X_10491_ _10489_/Y _10539_/B _10491_/C gnd _10583_/D vdd OAI21X1
XFILL_4__8523_ gnd vdd FILL
XFILL_1__9794_ gnd vdd FILL
XFILL111960x68050 gnd vdd FILL
XFILL_5_BUFX2_insert875 gnd vdd FILL
XFILL_5_BUFX2_insert886 gnd vdd FILL
X_12230_ _12227_/Y _12228_/Y _12230_/C gnd _12230_/Y vdd NAND3X1
XBUFX2_insert1050 _12806_/Q gnd _12340_/B vdd BUFX2
XFILL_5_BUFX2_insert897 gnd vdd FILL
XBUFX2_insert1061 _15051_/Y gnd _15071_/C vdd BUFX2
XBUFX2_insert1072 _13327_/Y gnd _8896_/B vdd BUFX2
XSFILL109240x38050 gnd vdd FILL
XFILL_1__8745_ gnd vdd FILL
XFILL_4__8454_ gnd vdd FILL
XSFILL13720x25050 gnd vdd FILL
X_12161_ _12137_/A _12934_/Q gnd _12162_/C vdd NAND2X1
XFILL_4__8385_ gnd vdd FILL
X_11112_ _11111_/Y _11110_/Y gnd _11553_/B vdd NOR2X1
XSFILL94200x23050 gnd vdd FILL
X_12092_ _12072_/A _12767_/A _12072_/C gnd _12094_/B vdd NAND3X1
XFILL_1__7627_ gnd vdd FILL
XSFILL114360x29050 gnd vdd FILL
XFILL_4__7336_ gnd vdd FILL
X_15920_ _15920_/A _15920_/B _15920_/C _14475_/Y gnd _15923_/B vdd OAI22X1
X_11043_ _12274_/Y _12159_/Y gnd _11641_/C vdd XOR2X1
XSFILL34600x4050 gnd vdd FILL
XFILL_1__7558_ gnd vdd FILL
X_15851_ _15851_/A _15851_/B _15850_/Y gnd _15852_/B vdd NOR3X1
XFILL_2_BUFX2_insert710 gnd vdd FILL
XFILL_4__9006_ gnd vdd FILL
XFILL_1__7489_ gnd vdd FILL
X_14802_ _9802_/A _13751_/B _13751_/C _9970_/Q gnd _14802_/Y vdd AOI22X1
XFILL_2_BUFX2_insert721 gnd vdd FILL
XFILL_2_BUFX2_insert732 gnd vdd FILL
XFILL_4__7198_ gnd vdd FILL
XFILL_1__9228_ gnd vdd FILL
X_15782_ _8424_/Q gnd _15782_/Y vdd INVX1
XFILL_2__8021_ gnd vdd FILL
XFILL_2_BUFX2_insert743 gnd vdd FILL
X_12994_ vdd _12994_/B gnd _12995_/C vdd NAND2X1
XFILL_4__10180_ gnd vdd FILL
XFILL_2_BUFX2_insert754 gnd vdd FILL
XFILL_2_BUFX2_insert765 gnd vdd FILL
XFILL_2_BUFX2_insert776 gnd vdd FILL
X_14733_ _14731_/Y _13680_/B _14466_/C _14733_/D gnd _14737_/A vdd OAI22X1
X_11945_ _11895_/B _12496_/A gnd _11946_/C vdd NAND2X1
XFILL_2_BUFX2_insert787 gnd vdd FILL
XFILL_5__11470_ gnd vdd FILL
XFILL_2_BUFX2_insert798 gnd vdd FILL
XFILL_2__10310_ gnd vdd FILL
XFILL_1__9159_ gnd vdd FILL
XFILL_2__11290_ gnd vdd FILL
XFILL_5__10421_ gnd vdd FILL
XFILL_5__9750_ gnd vdd FILL
XFILL_5__6962_ gnd vdd FILL
XFILL_3__11600_ gnd vdd FILL
X_14664_ _8129_/A gnd _16062_/C vdd INVX1
XFILL_2__10241_ gnd vdd FILL
X_11876_ _11874_/B _11876_/B gnd _11876_/Y vdd NAND2X1
XFILL_3__12580_ gnd vdd FILL
XFILL_0__11420_ gnd vdd FILL
XFILL_4__9908_ gnd vdd FILL
XFILL_5__8701_ gnd vdd FILL
X_16403_ gnd gnd gnd _16404_/C vdd NAND2X1
X_13615_ _7807_/A gnd _13615_/Y vdd INVX1
XFILL_1__10971_ gnd vdd FILL
XFILL112120x57050 gnd vdd FILL
XFILL_5__13140_ gnd vdd FILL
XFILL_5__9681_ gnd vdd FILL
XFILL_5__6893_ gnd vdd FILL
X_10827_ _10762_/B _7883_/B gnd _10828_/C vdd NAND2X1
X_14595_ _14595_/A _14587_/Y gnd _14596_/A vdd NAND2X1
XFILL_3__11531_ gnd vdd FILL
XFILL_2__10172_ gnd vdd FILL
XFILL_4__13870_ gnd vdd FILL
XFILL_1__12710_ gnd vdd FILL
XFILL_5__8632_ gnd vdd FILL
XSFILL64040x42050 gnd vdd FILL
XBUFX2_insert720 _13352_/Y gnd _10193_/A vdd BUFX2
XFILL_0__11351_ gnd vdd FILL
XBUFX2_insert731 _12411_/Y gnd _8377_/B vdd BUFX2
X_16334_ gnd gnd gnd _16335_/C vdd NAND2X1
XFILL_1__13690_ gnd vdd FILL
XBUFX2_insert742 _15055_/Y gnd _15342_/B vdd BUFX2
X_13546_ _8024_/Q gnd _15157_/C vdd INVX1
XFILL_3__14250_ gnd vdd FILL
XFILL_5__10283_ gnd vdd FILL
X_10758_ _10809_/A _6918_/B gnd _10759_/C vdd NAND2X1
XFILL_0__10302_ gnd vdd FILL
XBUFX2_insert753 _13344_/Y gnd _9785_/A vdd BUFX2
XFILL_2__8854_ gnd vdd FILL
XFILL112280x1050 gnd vdd FILL
XFILL_3__11462_ gnd vdd FILL
XBUFX2_insert764 _12393_/Y gnd _7847_/B vdd BUFX2
XFILL_1__12641_ gnd vdd FILL
XFILL_2__14980_ gnd vdd FILL
XFILL_0__14070_ gnd vdd FILL
XFILL_5__12022_ gnd vdd FILL
XFILL_0__11282_ gnd vdd FILL
XBUFX2_insert775 _13301_/Y gnd _7892_/A vdd BUFX2
XBUFX2_insert786 _13486_/Y gnd _14926_/C vdd BUFX2
X_16265_ _14894_/D _15656_/B _15656_/C gnd _16265_/Y vdd NOR3X1
XFILL_4__12752_ gnd vdd FILL
XFILL_4__15540_ gnd vdd FILL
XFILL_3__10413_ gnd vdd FILL
XFILL_2__7805_ gnd vdd FILL
X_13477_ _9047_/Q gnd _13479_/D vdd INVX1
XBUFX2_insert797 _13334_/Y gnd _9425_/A vdd BUFX2
XFILL_0__13021_ gnd vdd FILL
XFILL_3__14181_ gnd vdd FILL
XFILL_2__13931_ gnd vdd FILL
X_10689_ _14689_/B gnd _10691_/A vdd INVX1
XFILL_1__15360_ gnd vdd FILL
XFILL_3__11393_ gnd vdd FILL
XFILL_0__10233_ gnd vdd FILL
XFILL_2__8785_ gnd vdd FILL
XFILL_1__12572_ gnd vdd FILL
X_15216_ _15321_/C gnd _15380_/C vdd INVX4
X_12428_ _12368_/A _12428_/B gnd _12429_/C vdd NAND2X1
XFILL_5__8494_ gnd vdd FILL
XFILL_4__11703_ gnd vdd FILL
X_16196_ _15407_/C _14805_/Y _14804_/Y _15169_/A gnd _16200_/A vdd OAI22X1
XFILL_3__13132_ gnd vdd FILL
XFILL_2__7736_ gnd vdd FILL
XFILL_1__14311_ gnd vdd FILL
XFILL_4__15471_ gnd vdd FILL
XFILL_2__13862_ gnd vdd FILL
XFILL_1__11523_ gnd vdd FILL
XFILL_0__10164_ gnd vdd FILL
XFILL_5__7445_ gnd vdd FILL
XFILL_1__15291_ gnd vdd FILL
XSFILL84200x55050 gnd vdd FILL
X_15147_ _15760_/A _13576_/Y _15147_/C gnd _15150_/A vdd OAI21X1
X_12359_ _12359_/A _12668_/Q gnd _12360_/C vdd NAND2X1
XFILL_4__11634_ gnd vdd FILL
XFILL_2__15601_ gnd vdd FILL
XFILL_4__14422_ gnd vdd FILL
XFILL_1_CLKBUF1_insert180 gnd vdd FILL
XFILL_5__13973_ gnd vdd FILL
XFILL_1_CLKBUF1_insert191 gnd vdd FILL
XFILL_3__10275_ gnd vdd FILL
XFILL_1__14242_ gnd vdd FILL
XFILL_1__11454_ gnd vdd FILL
XFILL_2__13793_ gnd vdd FILL
XFILL_5__15712_ gnd vdd FILL
XFILL_2_BUFX2_insert1 gnd vdd FILL
XFILL_5__7376_ gnd vdd FILL
XFILL_0__14972_ gnd vdd FILL
XFILL_2__9406_ gnd vdd FILL
XFILL_3__12014_ gnd vdd FILL
XFILL_4__14353_ gnd vdd FILL
XFILL_0__9470_ gnd vdd FILL
X_15078_ _16314_/A gnd _15078_/Y vdd INVX1
XFILL_2__15532_ gnd vdd FILL
XFILL_4__11565_ gnd vdd FILL
XFILL_2__12744_ gnd vdd FILL
XFILL_1__10405_ gnd vdd FILL
XFILL_5__9115_ gnd vdd FILL
XFILL_1__14173_ gnd vdd FILL
XFILL_2__7598_ gnd vdd FILL
XFILL_0__13923_ gnd vdd FILL
XFILL_1__11385_ gnd vdd FILL
X_14029_ _8602_/A gnd _14029_/Y vdd INVX1
XFILL_4__13304_ gnd vdd FILL
XFILL_5__15643_ gnd vdd FILL
XFILL_4__10516_ gnd vdd FILL
XFILL_3__8130_ gnd vdd FILL
XFILL_5__12855_ gnd vdd FILL
XFILL_2__9337_ gnd vdd FILL
XFILL_4__14284_ gnd vdd FILL
XFILL_1__13124_ gnd vdd FILL
XFILL112200x37050 gnd vdd FILL
XFILL_2__15463_ gnd vdd FILL
XFILL_4__11496_ gnd vdd FILL
XSFILL23720x5050 gnd vdd FILL
XFILL_0__13854_ gnd vdd FILL
XFILL_4__13235_ gnd vdd FILL
XFILL_4__16023_ gnd vdd FILL
XFILL_0__8352_ gnd vdd FILL
XFILL_5__11806_ gnd vdd FILL
XFILL_4__10447_ gnd vdd FILL
XFILL_5__15574_ gnd vdd FILL
XFILL_2__14414_ gnd vdd FILL
XFILL_5__12786_ gnd vdd FILL
XFILL_2__9268_ gnd vdd FILL
XFILL_3__8061_ gnd vdd FILL
X_8980_ _8980_/A gnd _8982_/A vdd INVX1
XFILL_2__11626_ gnd vdd FILL
XFILL_3__13965_ gnd vdd FILL
XFILL_2__15394_ gnd vdd FILL
XFILL_1__10267_ gnd vdd FILL
XFILL_0__7303_ gnd vdd FILL
XFILL_0__13785_ gnd vdd FILL
XFILL_5__14525_ gnd vdd FILL
XFILL_0__10997_ gnd vdd FILL
XFILL_4__13166_ gnd vdd FILL
XFILL_3__15704_ gnd vdd FILL
XFILL_2__8219_ gnd vdd FILL
XFILL_5__11737_ gnd vdd FILL
X_7931_ _7929_/Y _7931_/B _7930_/Y gnd _8023_/D vdd OAI21X1
XFILL_4__10378_ gnd vdd FILL
XFILL_1__12006_ gnd vdd FILL
XFILL_2__14345_ gnd vdd FILL
XFILL_3__12916_ gnd vdd FILL
XFILL_0__15524_ gnd vdd FILL
XFILL_3__13896_ gnd vdd FILL
XFILL_2__11557_ gnd vdd FILL
XFILL_0__12736_ gnd vdd FILL
XSFILL53960x65050 gnd vdd FILL
XFILL_4__12117_ gnd vdd FILL
XFILL_0__7234_ gnd vdd FILL
XFILL_5__14456_ gnd vdd FILL
X_7862_ _7887_/B _7990_/B gnd _7863_/C vdd NAND2X1
XFILL_2__10508_ gnd vdd FILL
XFILL_3__15635_ gnd vdd FILL
XFILL_3__12847_ gnd vdd FILL
XFILL_4__13097_ gnd vdd FILL
XFILL_5__11668_ gnd vdd FILL
XFILL_2__14276_ gnd vdd FILL
XFILL_0__15455_ gnd vdd FILL
XFILL_2__11488_ gnd vdd FILL
X_9601_ _9599_/Y _9639_/A _9600_/Y gnd _9601_/Y vdd OAI21X1
XFILL_5__13407_ gnd vdd FILL
XFILL_6__15746_ gnd vdd FILL
XFILL_2__16015_ gnd vdd FILL
XFILL_4__12048_ gnd vdd FILL
XSFILL28760x41050 gnd vdd FILL
XFILL_5__10619_ gnd vdd FILL
XFILL_0__7165_ gnd vdd FILL
XFILL_2__13227_ gnd vdd FILL
XFILL_3__15566_ gnd vdd FILL
XFILL_5__14387_ gnd vdd FILL
XFILL_3__12778_ gnd vdd FILL
XFILL_3__8963_ gnd vdd FILL
XFILL_6_BUFX2_insert70 gnd vdd FILL
XFILL_2__10439_ gnd vdd FILL
XFILL_5__11599_ gnd vdd FILL
XFILL_0__14406_ gnd vdd FILL
X_7793_ _7751_/A _9834_/CLK _7793_/R vdd _7753_/Y gnd vdd DFFSR
XFILL_6_BUFX2_insert81 gnd vdd FILL
XFILL_1__13957_ gnd vdd FILL
XFILL_0__11618_ gnd vdd FILL
XFILL_0__15386_ gnd vdd FILL
XFILL_0__12598_ gnd vdd FILL
XFILL_5__16126_ gnd vdd FILL
XFILL_5__13338_ gnd vdd FILL
X_9532_ _9533_/B _9532_/B gnd _9532_/Y vdd NAND2X1
XFILL_5__9879_ gnd vdd FILL
XFILL_0__7096_ gnd vdd FILL
XFILL_3__14517_ gnd vdd FILL
XFILL_3__11729_ gnd vdd FILL
XFILL_1__12908_ gnd vdd FILL
XFILL_2__13158_ gnd vdd FILL
XFILL_3__15497_ gnd vdd FILL
XFILL_3__8894_ gnd vdd FILL
XFILL_0__14337_ gnd vdd FILL
XFILL_0__11549_ gnd vdd FILL
XFILL_1__13888_ gnd vdd FILL
XFILL_5_BUFX2_insert105 gnd vdd FILL
XFILL_4__15807_ gnd vdd FILL
XFILL_5__16057_ gnd vdd FILL
XFILL_5__13269_ gnd vdd FILL
X_9463_ _8951_/A _9535_/A gnd _9463_/Y vdd NAND2X1
XFILL_2__12109_ gnd vdd FILL
XSFILL33880x32050 gnd vdd FILL
XFILL_3__14448_ gnd vdd FILL
XFILL_3__7845_ gnd vdd FILL
XFILL_1__15627_ gnd vdd FILL
XFILL_2__13089_ gnd vdd FILL
XFILL_4__13999_ gnd vdd FILL
XFILL_1__12839_ gnd vdd FILL
XFILL_5__15008_ gnd vdd FILL
XFILL_0__14268_ gnd vdd FILL
X_8414_ _8414_/Q _7902_/CLK _7150_/R vdd _8414_/D gnd vdd DFFSR
XFILL_6__14559_ gnd vdd FILL
XFILL_1__6860_ gnd vdd FILL
XFILL_4__15738_ gnd vdd FILL
XFILL_0__16007_ gnd vdd FILL
XSFILL48920x54050 gnd vdd FILL
XFILL_3__14379_ gnd vdd FILL
X_9394_ _9394_/A gnd _9394_/Y vdd INVX1
XSFILL73720x80050 gnd vdd FILL
XFILL_0__13219_ gnd vdd FILL
XFILL_1__15558_ gnd vdd FILL
XFILL_0__9806_ gnd vdd FILL
XFILL_0__14199_ gnd vdd FILL
XFILL_4_BUFX2_insert805 gnd vdd FILL
XFILL_4_BUFX2_insert816 gnd vdd FILL
XFILL_3__16118_ gnd vdd FILL
X_8345_ _8343_/Y _8345_/B _8344_/Y gnd _8417_/D vdd OAI21X1
XFILL_3__9515_ gnd vdd FILL
XFILL_0__7998_ gnd vdd FILL
XFILL_4__15669_ gnd vdd FILL
XFILL_1__14509_ gnd vdd FILL
XFILL_4_BUFX2_insert827 gnd vdd FILL
XFILL_6__9224_ gnd vdd FILL
XFILL_4_BUFX2_insert838 gnd vdd FILL
XFILL_1__15489_ gnd vdd FILL
XSFILL49000x63050 gnd vdd FILL
XFILL_0__9737_ gnd vdd FILL
XFILL_1__8530_ gnd vdd FILL
XFILL_4_BUFX2_insert849 gnd vdd FILL
XFILL_0__6949_ gnd vdd FILL
X_8276_ _8237_/A _7380_/B gnd _8277_/C vdd NAND2X1
XFILL_3__16049_ gnd vdd FILL
XSFILL109560x74050 gnd vdd FILL
X_7227_ _7277_/Q gnd _7227_/Y vdd INVX1
XFILL_1__8461_ gnd vdd FILL
XFILL_0__9668_ gnd vdd FILL
XFILL_3__9377_ gnd vdd FILL
XSFILL28840x21050 gnd vdd FILL
XFILL_0__8619_ gnd vdd FILL
XSFILL54120x54050 gnd vdd FILL
X_7158_ _7158_/A gnd _7160_/A vdd INVX1
XFILL_0__9599_ gnd vdd FILL
XFILL_3__8328_ gnd vdd FILL
XFILL_4__7121_ gnd vdd FILL
XFILL_1__8392_ gnd vdd FILL
XCLKBUF1_insert190 CLKBUF1_insert192/A gnd _7902_/CLK vdd CLKBUF1
XFILL_1__7343_ gnd vdd FILL
X_7089_ _7087_/Y _7124_/A _7089_/C gnd _7089_/Y vdd OAI21X1
XFILL_4__7052_ gnd vdd FILL
XFILL_3__8259_ gnd vdd FILL
XSFILL33960x12050 gnd vdd FILL
XFILL_1__9013_ gnd vdd FILL
XFILL_5_BUFX2_insert5 gnd vdd FILL
XSFILL18760x73050 gnd vdd FILL
XSFILL8600x83050 gnd vdd FILL
XFILL_1_BUFX2_insert706 gnd vdd FILL
XFILL_1_BUFX2_insert717 gnd vdd FILL
XFILL_1_BUFX2_insert728 gnd vdd FILL
X_11730_ _11729_/Y _11731_/B gnd _11741_/A vdd AND2X2
XFILL_1_BUFX2_insert739 gnd vdd FILL
XSFILL108760x26050 gnd vdd FILL
XSFILL99240x71050 gnd vdd FILL
XFILL_4__7954_ gnd vdd FILL
X_11661_ _11661_/A _11661_/B _11660_/Y gnd _12485_/B vdd NAND3X1
XSFILL23880x64050 gnd vdd FILL
XFILL_4__6905_ gnd vdd FILL
X_13400_ _13394_/Y _13399_/Y gnd _13401_/C vdd NOR2X1
XFILL_4__7885_ gnd vdd FILL
X_10612_ _16246_/A _8297_/CLK _7796_/R vdd _10578_/Y gnd vdd DFFSR
X_14380_ _14380_/A _14380_/B gnd _14402_/A vdd NOR2X1
XFILL_1__9915_ gnd vdd FILL
X_11592_ _11592_/A _11592_/B gnd _11600_/B vdd NOR2X1
XFILL_4__6836_ gnd vdd FILL
XFILL_4__9624_ gnd vdd FILL
X_13331_ _13273_/A _13337_/B gnd _13331_/Y vdd AND2X2
XSFILL54200x34050 gnd vdd FILL
X_10543_ _15837_/A gnd _10545_/A vdd INVX1
XFILL_1__9846_ gnd vdd FILL
XFILL_5_BUFX2_insert650 gnd vdd FILL
XFILL_5_BUFX2_insert661 gnd vdd FILL
XFILL_4__9555_ gnd vdd FILL
XFILL_5_BUFX2_insert672 gnd vdd FILL
X_16050_ _16049_/Y _15656_/B _15656_/C gnd _16053_/B vdd NOR3X1
X_13262_ _13209_/B _13262_/B gnd _13263_/B vdd NAND2X1
XFILL_5_BUFX2_insert683 gnd vdd FILL
X_10474_ _10418_/A _9194_/CLK _7914_/R vdd _10474_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert694 gnd vdd FILL
XFILL_1__9777_ gnd vdd FILL
XFILL_2__8570_ gnd vdd FILL
XFILL_1__6989_ gnd vdd FILL
X_15001_ _16235_/A gnd _15916_/B vdd INVX4
XFILL_4__8506_ gnd vdd FILL
XFILL_4__9486_ gnd vdd FILL
X_12213_ _12216_/A gnd _12213_/Y vdd INVX8
XFILL_1__8728_ gnd vdd FILL
X_13193_ _13133_/A _13201_/CLK _13201_/R vdd _13193_/D gnd vdd DFFSR
XFILL_5__7230_ gnd vdd FILL
XSFILL18840x53050 gnd vdd FILL
X_12144_ _12144_/A _12122_/A _12143_/Y gnd _12144_/Y vdd OAI21X1
XFILL_5__10970_ gnd vdd FILL
XFILL_3__10060_ gnd vdd FILL
XFILL_2__7452_ gnd vdd FILL
XFILL_1__8659_ gnd vdd FILL
XFILL_2_CLKBUF1_insert220 gnd vdd FILL
XFILL_2__10790_ gnd vdd FILL
XFILL_4__8368_ gnd vdd FILL
XFILL_5__7161_ gnd vdd FILL
XSFILL99320x51050 gnd vdd FILL
X_12075_ _11987_/A _12409_/A _12011_/C gnd _12078_/A vdd NAND3X1
XFILL_4__11350_ gnd vdd FILL
XFILL_0__10920_ gnd vdd FILL
XFILL_4__7319_ gnd vdd FILL
XFILL_1__11170_ gnd vdd FILL
XFILL_4__10301_ gnd vdd FILL
X_15903_ _7019_/Q _15382_/B _16096_/C _7403_/Q gnd _15903_/Y vdd AOI22X1
XFILL_5__7092_ gnd vdd FILL
X_11026_ _11026_/A _11026_/B _11026_/C _11025_/Y gnd _11027_/B vdd OAI22X1
XFILL_5__12640_ gnd vdd FILL
XFILL_2__9122_ gnd vdd FILL
XFILL_1__10121_ gnd vdd FILL
XFILL_4__11281_ gnd vdd FILL
XFILL_2__12460_ gnd vdd FILL
XFILL112280x11050 gnd vdd FILL
XSFILL64040x37050 gnd vdd FILL
XFILL_4__13020_ gnd vdd FILL
XFILL_6__13930_ gnd vdd FILL
XFILL_4__10232_ gnd vdd FILL
X_15834_ _9321_/Q gnd _15836_/A vdd INVX1
XFILL_5__12571_ gnd vdd FILL
XFILL_3__13750_ gnd vdd FILL
XFILL_2__11411_ gnd vdd FILL
XFILL_3__10962_ gnd vdd FILL
XFILL_1__10052_ gnd vdd FILL
XFILL_0_BUFX2_insert1008 gnd vdd FILL
XFILL_2_BUFX2_insert540 gnd vdd FILL
XFILL_2__12391_ gnd vdd FILL
XFILL_0_BUFX2_insert1019 gnd vdd FILL
XFILL_2_BUFX2_insert551 gnd vdd FILL
XFILL_0__13570_ gnd vdd FILL
XFILL_2_BUFX2_insert562 gnd vdd FILL
XFILL_5__14310_ gnd vdd FILL
XFILL_0__10782_ gnd vdd FILL
XFILL_3__12701_ gnd vdd FILL
XFILL_2_BUFX2_insert573 gnd vdd FILL
XFILL_2__8004_ gnd vdd FILL
XFILL_5__11522_ gnd vdd FILL
X_12977_ _12977_/A vdd _12977_/C gnd _13055_/D vdd OAI21X1
XFILL_2__14130_ gnd vdd FILL
XFILL_4__10163_ gnd vdd FILL
X_15765_ _15765_/A _15795_/B _15765_/C gnd _15765_/Y vdd OAI21X1
XFILL_5__15290_ gnd vdd FILL
XFILL_3__13681_ gnd vdd FILL
XFILL_2_BUFX2_insert584 gnd vdd FILL
XFILL_0__12521_ gnd vdd FILL
XFILL_2__11342_ gnd vdd FILL
XFILL_1__14860_ gnd vdd FILL
XFILL_2_BUFX2_insert595 gnd vdd FILL
XFILL_5__9802_ gnd vdd FILL
XFILL_3__10893_ gnd vdd FILL
XFILL_5__14241_ gnd vdd FILL
XFILL_5__7994_ gnd vdd FILL
X_14716_ _9412_/A gnd _14718_/D vdd INVX1
X_11928_ _11926_/Y _11900_/A _11928_/C gnd _6851_/A vdd OAI21X1
XFILL_3__15420_ gnd vdd FILL
XFILL_3__12632_ gnd vdd FILL
XFILL_6__13792_ gnd vdd FILL
X_15696_ _15696_/A _14245_/A _9702_/Q _15652_/D gnd _15696_/Y vdd AOI22X1
XFILL_5__11453_ gnd vdd FILL
XFILL_1__13811_ gnd vdd FILL
XFILL_2__14061_ gnd vdd FILL
XFILL_4__14971_ gnd vdd FILL
XFILL_0__15240_ gnd vdd FILL
XFILL_0__12452_ gnd vdd FILL
XFILL_2__11273_ gnd vdd FILL
XSFILL58920x17050 gnd vdd FILL
XFILL_5__6945_ gnd vdd FILL
XFILL_6__15531_ gnd vdd FILL
XFILL_5__9733_ gnd vdd FILL
XFILL_1__14791_ gnd vdd FILL
XFILL_6__12743_ gnd vdd FILL
X_14647_ _14647_/A _14647_/B _14265_/C gnd _13024_/B vdd AOI21X1
XFILL_5__10404_ gnd vdd FILL
XFILL_5__14172_ gnd vdd FILL
XFILL_3__15351_ gnd vdd FILL
X_11859_ _11774_/A _11689_/Y _11718_/A gnd _11863_/A vdd NAND3X1
XFILL_4__13922_ gnd vdd FILL
XFILL_5__11384_ gnd vdd FILL
XFILL_2__13012_ gnd vdd FILL
XSFILL69560x68050 gnd vdd FILL
XFILL_0__11403_ gnd vdd FILL
XFILL_0__15171_ gnd vdd FILL
XFILL_1__13742_ gnd vdd FILL
XFILL_1__10954_ gnd vdd FILL
XFILL_0__12383_ gnd vdd FILL
XFILL_5__9664_ gnd vdd FILL
XFILL_5__13123_ gnd vdd FILL
XFILL_5__6876_ gnd vdd FILL
XFILL_3__14302_ gnd vdd FILL
X_14578_ _15986_/A _13843_/C _14200_/C _14577_/Y gnd _14579_/A vdd OAI22X1
XFILL_0__8970_ gnd vdd FILL
XFILL_3__11514_ gnd vdd FILL
XSFILL59000x26050 gnd vdd FILL
XFILL_4__13853_ gnd vdd FILL
XFILL_2__8906_ gnd vdd FILL
XFILL_3__15282_ gnd vdd FILL
XFILL_3__12494_ gnd vdd FILL
XFILL_2__10155_ gnd vdd FILL
XSFILL99400x31050 gnd vdd FILL
XFILL_2__9886_ gnd vdd FILL
XFILL_0__14122_ gnd vdd FILL
XBUFX2_insert550 BUFX2_insert496/A gnd _7015_/R vdd BUFX2
XFILL_0__11334_ gnd vdd FILL
XFILL_5__8615_ gnd vdd FILL
XFILL_1__13673_ gnd vdd FILL
XBUFX2_insert561 BUFX2_insert524/A gnd _7000_/R vdd BUFX2
XSFILL104760x77050 gnd vdd FILL
XFILL_1__10885_ gnd vdd FILL
X_16317_ _16314_/Y _16316_/Y gnd _16317_/Y vdd NOR2X1
XFILL_6__11625_ gnd vdd FILL
X_13529_ _14894_/B gnd _14214_/C vdd INVX8
XFILL_5__9595_ gnd vdd FILL
XBUFX2_insert572 BUFX2_insert570/A gnd _12685_/R vdd BUFX2
XFILL_6__15393_ gnd vdd FILL
XFILL_3__14233_ gnd vdd FILL
XFILL_5__10266_ gnd vdd FILL
XFILL_3__7630_ gnd vdd FILL
XBUFX2_insert583 BUFX2_insert518/A gnd _7531_/R vdd BUFX2
XFILL_1__15412_ gnd vdd FILL
XFILL111880x3050 gnd vdd FILL
XFILL_2__8837_ gnd vdd FILL
XFILL_3__11445_ gnd vdd FILL
XBUFX2_insert594 BUFX2_insert518/A gnd _9203_/R vdd BUFX2
XFILL_1__12624_ gnd vdd FILL
XFILL_4__13784_ gnd vdd FILL
XFILL_0__14053_ gnd vdd FILL
XFILL_2__14963_ gnd vdd FILL
XFILL_4__10996_ gnd vdd FILL
XFILL_1__16392_ gnd vdd FILL
XFILL_0__11265_ gnd vdd FILL
XFILL_5__12005_ gnd vdd FILL
XFILL_6__14344_ gnd vdd FILL
X_16248_ _14883_/Y _15239_/B _16106_/A _14884_/B gnd _16249_/A vdd OAI22X1
XFILL_4__15523_ gnd vdd FILL
XFILL_0__7852_ gnd vdd FILL
XFILL_4__12735_ gnd vdd FILL
XFILL_3__14164_ gnd vdd FILL
XFILL_5__10197_ gnd vdd FILL
XSFILL64120x17050 gnd vdd FILL
XFILL_2__13914_ gnd vdd FILL
XFILL_0__13004_ gnd vdd FILL
XFILL_2__8768_ gnd vdd FILL
XFILL_1__15343_ gnd vdd FILL
XFILL_3__7561_ gnd vdd FILL
XFILL_3__11376_ gnd vdd FILL
XFILL_2__14894_ gnd vdd FILL
XFILL_6__10507_ gnd vdd FILL
XSFILL74280x61050 gnd vdd FILL
XFILL_5__8477_ gnd vdd FILL
X_8130_ _8082_/A _9282_/B gnd _8131_/C vdd NAND2X1
XFILL_0__11196_ gnd vdd FILL
X_16179_ _16179_/A _16179_/B gnd _16203_/A vdd NOR2X1
XFILL_3__13115_ gnd vdd FILL
XFILL_3__9300_ gnd vdd FILL
XFILL_2__7719_ gnd vdd FILL
XSFILL48440x71050 gnd vdd FILL
XFILL_6__11487_ gnd vdd FILL
XFILL_4__15454_ gnd vdd FILL
XFILL_2__13845_ gnd vdd FILL
XFILL_1__11506_ gnd vdd FILL
XFILL_3__14095_ gnd vdd FILL
XFILL_5__7428_ gnd vdd FILL
XFILL_0__10147_ gnd vdd FILL
XFILL_3__7492_ gnd vdd FILL
XFILL_2__8699_ gnd vdd FILL
XFILL_1__15274_ gnd vdd FILL
XFILL_1__12486_ gnd vdd FILL
XFILL_0__9522_ gnd vdd FILL
XSFILL89320x83050 gnd vdd FILL
XFILL_4__14405_ gnd vdd FILL
X_8061_ _8107_/B _9981_/B gnd _8062_/C vdd NAND2X1
XFILL_3__9231_ gnd vdd FILL
XFILL_3__13046_ gnd vdd FILL
XFILL_5__13956_ gnd vdd FILL
XFILL_4__11617_ gnd vdd FILL
XSFILL3560x24050 gnd vdd FILL
XFILL_4__15385_ gnd vdd FILL
XFILL_1__14225_ gnd vdd FILL
XFILL_4__12597_ gnd vdd FILL
XFILL_3__10258_ gnd vdd FILL
XFILL_2__13776_ gnd vdd FILL
XFILL_1__11437_ gnd vdd FILL
XFILL_5__7359_ gnd vdd FILL
X_7012_ _7012_/Q _8161_/CLK _7140_/R vdd _7012_/D gnd vdd DFFSR
XFILL_2__10988_ gnd vdd FILL
XFILL_0__14955_ gnd vdd FILL
XFILL_5__12907_ gnd vdd FILL
XFILL_2__15515_ gnd vdd FILL
XFILL_4__14336_ gnd vdd FILL
XFILL_4__11548_ gnd vdd FILL
XFILL_2__12727_ gnd vdd FILL
XFILL_5__13887_ gnd vdd FILL
XFILL_3__9162_ gnd vdd FILL
XFILL_3__10189_ gnd vdd FILL
XSFILL54040x69050 gnd vdd FILL
XFILL_1__14156_ gnd vdd FILL
XFILL_0__13906_ gnd vdd FILL
XSFILL115000x14050 gnd vdd FILL
XFILL_0__8404_ gnd vdd FILL
XSFILL33880x6050 gnd vdd FILL
XFILL_1__11368_ gnd vdd FILL
XSFILL68360x22050 gnd vdd FILL
XFILL_5__15626_ gnd vdd FILL
XFILL_0__14886_ gnd vdd FILL
XFILL_0__9384_ gnd vdd FILL
XFILL_3__8113_ gnd vdd FILL
XFILL_5__12838_ gnd vdd FILL
XFILL_1__13107_ gnd vdd FILL
XFILL_2__15446_ gnd vdd FILL
XFILL_4__11479_ gnd vdd FILL
XFILL_4__14267_ gnd vdd FILL
XFILL_2__12658_ gnd vdd FILL
XFILL_1__10319_ gnd vdd FILL
XFILL_5__9029_ gnd vdd FILL
XFILL_3__9093_ gnd vdd FILL
XFILL_6__9911_ gnd vdd FILL
XFILL_0__13837_ gnd vdd FILL
XFILL_3__14997_ gnd vdd FILL
XFILL_1__14087_ gnd vdd FILL
XFILL_1__11299_ gnd vdd FILL
XFILL_0__8335_ gnd vdd FILL
XFILL_4__16006_ gnd vdd FILL
XFILL_6__12039_ gnd vdd FILL
XFILL_4__13218_ gnd vdd FILL
XFILL_5__15557_ gnd vdd FILL
XFILL_4__14198_ gnd vdd FILL
XFILL_5__12769_ gnd vdd FILL
X_8963_ _9014_/A _8195_/B gnd _8964_/C vdd NAND2X1
XSFILL69240x50050 gnd vdd FILL
XSFILL33880x27050 gnd vdd FILL
XFILL_2__11609_ gnd vdd FILL
XFILL_2__15377_ gnd vdd FILL
XFILL_1__13038_ gnd vdd FILL
XFILL_3__13948_ gnd vdd FILL
XFILL_2__12589_ gnd vdd FILL
XFILL_0__13768_ gnd vdd FILL
XFILL_5__14508_ gnd vdd FILL
XFILL_0__8266_ gnd vdd FILL
XFILL_4__13149_ gnd vdd FILL
X_7914_ _7914_/Q _9194_/CLK _7914_/R vdd _7914_/D gnd vdd DFFSR
XFILL_2__14328_ gnd vdd FILL
XFILL_5__15488_ gnd vdd FILL
X_8894_ _8894_/A gnd _8894_/Y vdd INVX1
XFILL_0__15507_ gnd vdd FILL
XSFILL48920x49050 gnd vdd FILL
XFILL_0__12719_ gnd vdd FILL
XFILL_3__13879_ gnd vdd FILL
XFILL_0__7217_ gnd vdd FILL
XSFILL58280x74050 gnd vdd FILL
XFILL_0__13699_ gnd vdd FILL
XFILL_5__14439_ gnd vdd FILL
X_7845_ _7843_/Y _7824_/B _7845_/C gnd _7909_/D vdd OAI21X1
XFILL_3__15618_ gnd vdd FILL
XSFILL79240x5050 gnd vdd FILL
XFILL_0__8197_ gnd vdd FILL
XFILL_2__14259_ gnd vdd FILL
XFILL_0__15438_ gnd vdd FILL
XFILL_3__9995_ gnd vdd FILL
XFILL_1__14989_ gnd vdd FILL
XSFILL49000x58050 gnd vdd FILL
XFILL_0_CLKBUF1_insert117 gnd vdd FILL
XFILL_0_CLKBUF1_insert128 gnd vdd FILL
XFILL_3__15549_ gnd vdd FILL
X_7776_ _7700_/A _7530_/CLK _7523_/R vdd _7702_/Y gnd vdd DFFSR
XFILL_0_CLKBUF1_insert139 gnd vdd FILL
XFILL_0__15369_ gnd vdd FILL
XFILL_5__16109_ gnd vdd FILL
XFILL_6__8655_ gnd vdd FILL
X_9515_ _9515_/A _9514_/A _9515_/C gnd _9515_/Y vdd OAI21X1
XSFILL109560x69050 gnd vdd FILL
XFILL_0__7079_ gnd vdd FILL
XFILL_1__7961_ gnd vdd FILL
XFILL_4__7670_ gnd vdd FILL
XFILL_3__8877_ gnd vdd FILL
XFILL_6__7606_ gnd vdd FILL
XFILL_1__6912_ gnd vdd FILL
X_9446_ _9382_/A _8306_/CLK _9054_/R vdd _9446_/D gnd vdd DFFSR
XSFILL54120x49050 gnd vdd FILL
XFILL_1__7892_ gnd vdd FILL
XFILL_3__7828_ gnd vdd FILL
XFILL_1__9631_ gnd vdd FILL
XFILL_1__6843_ gnd vdd FILL
X_9377_ _9398_/A _9889_/B gnd _9377_/Y vdd NAND2X1
XFILL_4__9340_ gnd vdd FILL
XFILL_4_BUFX2_insert602 gnd vdd FILL
XFILL_3__7759_ gnd vdd FILL
XFILL_4_BUFX2_insert613 gnd vdd FILL
XFILL_4_BUFX2_insert624 gnd vdd FILL
XFILL_4_BUFX2_insert635 gnd vdd FILL
X_8328_ _8328_/A gnd _8328_/Y vdd INVX1
XFILL_4_BUFX2_insert646 gnd vdd FILL
XFILL_4__9271_ gnd vdd FILL
XFILL_4_BUFX2_insert657 gnd vdd FILL
XFILL_4_BUFX2_insert668 gnd vdd FILL
X_10190_ _10191_/B _8910_/B gnd _10191_/C vdd NAND2X1
XFILL_4_BUFX2_insert679 gnd vdd FILL
XFILL_1__8513_ gnd vdd FILL
XSFILL8600x78050 gnd vdd FILL
XFILL_1__9493_ gnd vdd FILL
XFILL_4__8222_ gnd vdd FILL
X_8259_ _8257_/Y _8187_/B _8259_/C gnd _8303_/D vdd OAI21X1
XFILL_3__9429_ gnd vdd FILL
XSFILL39000x8050 gnd vdd FILL
XSFILL33800x71050 gnd vdd FILL
XFILL_1__8444_ gnd vdd FILL
XFILL_2_BUFX2_insert90 gnd vdd FILL
XFILL_1__8375_ gnd vdd FILL
XFILL_4__7104_ gnd vdd FILL
XFILL_4__8084_ gnd vdd FILL
X_12900_ _12900_/A vdd _12900_/C gnd _12900_/Y vdd OAI21X1
X_13880_ _13880_/A _13876_/Y gnd _13880_/Y vdd NOR2X1
XFILL_1__7326_ gnd vdd FILL
XFILL_4__7035_ gnd vdd FILL
X_12831_ _12831_/A vdd _12830_/Y gnd _12831_/Y vdd OAI21X1
XFILL_1_BUFX2_insert503 gnd vdd FILL
X_15550_ _15550_/A _14045_/D _15550_/C gnd _15550_/Y vdd NOR3X1
XSFILL79160x33050 gnd vdd FILL
XFILL_1_BUFX2_insert514 gnd vdd FILL
X_12762_ _12762_/A memoryOutData[22] gnd _12763_/C vdd NAND2X1
XFILL_1_BUFX2_insert525 gnd vdd FILL
XFILL_1_BUFX2_insert536 gnd vdd FILL
XFILL_1__7188_ gnd vdd FILL
XFILL_1_BUFX2_insert547 gnd vdd FILL
X_14501_ _7608_/A gnd _14501_/Y vdd INVX1
XFILL_1_BUFX2_insert558 gnd vdd FILL
X_11713_ _11713_/A _11726_/B _11713_/C gnd _11713_/Y vdd AOI21X1
XFILL_1_BUFX2_insert569 gnd vdd FILL
XFILL_4__8986_ gnd vdd FILL
X_15481_ _15481_/A _15481_/B _15477_/Y gnd _15496_/A vdd NAND3X1
X_12693_ _12693_/Q _12809_/CLK _12809_/R vdd _12693_/D gnd vdd DFFSR
XFILL_4__7937_ gnd vdd FILL
X_14432_ _8810_/Q gnd _14433_/A vdd INVX1
X_11644_ _11044_/A _11642_/Y _11644_/C gnd _11661_/A vdd OAI21X1
XSFILL84280x24050 gnd vdd FILL
XFILL_2__9740_ gnd vdd FILL
XFILL_2__6952_ gnd vdd FILL
XSFILL58440x34050 gnd vdd FILL
XFILL_5__10120_ gnd vdd FILL
XFILL_4__7868_ gnd vdd FILL
X_14363_ _7913_/Q gnd _14365_/A vdd INVX1
XSFILL99320x46050 gnd vdd FILL
X_11575_ _11561_/A _11846_/C _11575_/C gnd _11575_/Y vdd AOI21X1
XFILL_2__9671_ gnd vdd FILL
X_16102_ _16101_/Y _16102_/B gnd _16102_/Y vdd NOR2X1
XFILL_1__10670_ gnd vdd FILL
XFILL_4__9607_ gnd vdd FILL
XFILL_2__6883_ gnd vdd FILL
XFILL_5__8400_ gnd vdd FILL
X_13314_ _13313_/Y _13297_/C gnd _13314_/Y vdd NOR2X1
XFILL_5__9380_ gnd vdd FILL
XFILL_6__11410_ gnd vdd FILL
XFILL_4__7799_ gnd vdd FILL
XFILL_5__10051_ gnd vdd FILL
X_10526_ _10581_/B _7326_/B gnd _10526_/Y vdd NAND2X1
XFILL_2__8622_ gnd vdd FILL
X_14294_ _10727_/Q gnd _14294_/Y vdd INVX1
XFILL_3__11230_ gnd vdd FILL
XFILL_5_BUFX2_insert480 gnd vdd FILL
XFILL_4__10781_ gnd vdd FILL
XFILL_5__8331_ gnd vdd FILL
XFILL_2__11960_ gnd vdd FILL
XFILL_0__11050_ gnd vdd FILL
XFILL_5_BUFX2_insert491 gnd vdd FILL
X_16033_ _16032_/Y _16033_/B gnd _16045_/C vdd NAND2X1
XFILL_4__9538_ gnd vdd FILL
X_13245_ _13244_/Y _13245_/B gnd _13253_/A vdd AND2X2
X_10457_ _10457_/Q _9817_/CLK _8942_/R vdd _10457_/D gnd vdd DFFSR
XFILL_4__12520_ gnd vdd FILL
XFILL_2__10911_ gnd vdd FILL
XFILL_3__11161_ gnd vdd FILL
XFILL_0__10001_ gnd vdd FILL
XSFILL24040x48050 gnd vdd FILL
XFILL_1__12340_ gnd vdd FILL
XFILL_5__8262_ gnd vdd FILL
XFILL_2__11891_ gnd vdd FILL
XSFILL109320x31050 gnd vdd FILL
XFILL_5__13810_ gnd vdd FILL
XFILL_4__9469_ gnd vdd FILL
XFILL_3__10112_ gnd vdd FILL
XFILL_4__12451_ gnd vdd FILL
X_13176_ _11890_/A _13180_/CLK _13180_/R vdd _13176_/D gnd vdd DFFSR
XFILL_6__11272_ gnd vdd FILL
XFILL_2__7504_ gnd vdd FILL
XFILL_2__13630_ gnd vdd FILL
X_10388_ _13972_/A gnd _10390_/A vdd INVX1
XFILL_5__14790_ gnd vdd FILL
XFILL_2__8484_ gnd vdd FILL
XFILL_5__7213_ gnd vdd FILL
XFILL_3__11092_ gnd vdd FILL
XFILL_1__12271_ gnd vdd FILL
XFILL_6__13011_ gnd vdd FILL
XFILL_5__8193_ gnd vdd FILL
X_12127_ _12127_/A gnd _12127_/Y vdd INVX1
XFILL_4__11402_ gnd vdd FILL
XFILL_5__13741_ gnd vdd FILL
XFILL_5__10953_ gnd vdd FILL
XFILL_2__7435_ gnd vdd FILL
XFILL_3__10043_ gnd vdd FILL
XFILL_4__15170_ gnd vdd FILL
XFILL_1__14010_ gnd vdd FILL
XFILL_4__12382_ gnd vdd FILL
XFILL_3__14920_ gnd vdd FILL
XFILL_2__13561_ gnd vdd FILL
XFILL_1__11222_ gnd vdd FILL
XFILL_0__14740_ gnd vdd FILL
XFILL_2__10773_ gnd vdd FILL
XFILL_0__11952_ gnd vdd FILL
XSFILL114440x22050 gnd vdd FILL
XFILL_2__15300_ gnd vdd FILL
X_12058_ _12055_/Y _12056_/Y _12057_/Y gnd _13131_/B vdd NAND3X1
XFILL_4__14121_ gnd vdd FILL
XFILL_4__11333_ gnd vdd FILL
XFILL_2__12512_ gnd vdd FILL
XFILL_5__13672_ gnd vdd FILL
XFILL_3__14851_ gnd vdd FILL
XFILL_5__10884_ gnd vdd FILL
XFILL_2__7366_ gnd vdd FILL
XFILL_1__11153_ gnd vdd FILL
XFILL_2__16280_ gnd vdd FILL
XFILL_0__10903_ gnd vdd FILL
XSFILL43720x54050 gnd vdd FILL
XFILL_2__13492_ gnd vdd FILL
XFILL_5__7075_ gnd vdd FILL
XFILL_5__15411_ gnd vdd FILL
XFILL_0_BUFX2_insert19 gnd vdd FILL
XFILL_0__14671_ gnd vdd FILL
X_11009_ _12117_/Y gnd _11009_/Y vdd INVX1
XFILL_5__12623_ gnd vdd FILL
XFILL_0__11883_ gnd vdd FILL
XFILL_4__14052_ gnd vdd FILL
XFILL_2__9105_ gnd vdd FILL
XFILL_3__13802_ gnd vdd FILL
XFILL_2__15231_ gnd vdd FILL
XFILL_1__10104_ gnd vdd FILL
XFILL_5__16391_ gnd vdd FILL
XFILL_4__11264_ gnd vdd FILL
XFILL_0__16410_ gnd vdd FILL
XFILL_2__12443_ gnd vdd FILL
XFILL_2__7297_ gnd vdd FILL
XFILL_0__13622_ gnd vdd FILL
XFILL_1__15961_ gnd vdd FILL
XFILL_3__11994_ gnd vdd FILL
XFILL_1__11084_ gnd vdd FILL
XFILL_3__14782_ gnd vdd FILL
XSFILL69160x65050 gnd vdd FILL
XFILL_0__8120_ gnd vdd FILL
XSFILL99400x26050 gnd vdd FILL
XFILL_4__13003_ gnd vdd FILL
XFILL_0__10834_ gnd vdd FILL
XFILL_5__15342_ gnd vdd FILL
X_15817_ _7273_/Q _15177_/B _16293_/A _7145_/Q gnd _15819_/A vdd AOI22X1
XFILL_2__9036_ gnd vdd FILL
XFILL_3__10945_ gnd vdd FILL
XFILL_2_BUFX2_insert370 gnd vdd FILL
XFILL_1__10035_ gnd vdd FILL
XFILL_2__15162_ gnd vdd FILL
XFILL_3__13733_ gnd vdd FILL
XFILL_4__11195_ gnd vdd FILL
XFILL_1__14912_ gnd vdd FILL
XFILL_2_BUFX2_insert381 gnd vdd FILL
XFILL_0__16341_ gnd vdd FILL
XFILL_2__12374_ gnd vdd FILL
XFILL_0__10765_ gnd vdd FILL
XFILL_1__15892_ gnd vdd FILL
XFILL_2_BUFX2_insert392 gnd vdd FILL
XFILL_0__13553_ gnd vdd FILL
XFILL_5__11505_ gnd vdd FILL
XFILL_4__10146_ gnd vdd FILL
X_15748_ _15550_/A _15748_/B _15550_/C gnd _15769_/B vdd NOR3X1
XFILL_2__14113_ gnd vdd FILL
XFILL_5__15273_ gnd vdd FILL
XFILL_3__13664_ gnd vdd FILL
XFILL_5__12485_ gnd vdd FILL
XFILL_2__11325_ gnd vdd FILL
XFILL_1__14843_ gnd vdd FILL
XFILL_0__12504_ gnd vdd FILL
XFILL_3__10876_ gnd vdd FILL
XFILL_2__15093_ gnd vdd FILL
XFILL_0__16272_ gnd vdd FILL
XFILL_5__14224_ gnd vdd FILL
XFILL_0__13484_ gnd vdd FILL
XFILL_0__10696_ gnd vdd FILL
XFILL_3__12615_ gnd vdd FILL
X_7630_ _7592_/B _7502_/B gnd _7631_/C vdd NAND2X1
XFILL_3__15403_ gnd vdd FILL
XFILL_5__11436_ gnd vdd FILL
XFILL_5__7977_ gnd vdd FILL
X_15679_ _15679_/A _15675_/Y _15678_/Y gnd _15690_/A vdd NAND3X1
XFILL_2__14044_ gnd vdd FILL
XFILL_4__14954_ gnd vdd FILL
XSFILL109400x11050 gnd vdd FILL
XFILL_3__16383_ gnd vdd FILL
XFILL_3__13595_ gnd vdd FILL
XFILL_0__15223_ gnd vdd FILL
XFILL_2__11256_ gnd vdd FILL
XFILL_3__9780_ gnd vdd FILL
XFILL_0__12435_ gnd vdd FILL
XFILL_3__6992_ gnd vdd FILL
XFILL_1__14774_ gnd vdd FILL
XFILL_5__6928_ gnd vdd FILL
XFILL_1__11986_ gnd vdd FILL
XSFILL89320x78050 gnd vdd FILL
XFILL_5__14155_ gnd vdd FILL
XFILL_4__13905_ gnd vdd FILL
XFILL_3__15334_ gnd vdd FILL
X_7561_ _7562_/B _9737_/B gnd _7561_/Y vdd NAND2X1
XFILL112200x50050 gnd vdd FILL
XFILL_3__8731_ gnd vdd FILL
XSFILL3560x19050 gnd vdd FILL
XFILL_5__11367_ gnd vdd FILL
XFILL_1__13725_ gnd vdd FILL
XFILL_4__14885_ gnd vdd FILL
XFILL_2__9938_ gnd vdd FILL
XFILL_1__10937_ gnd vdd FILL
XFILL_0__12366_ gnd vdd FILL
XFILL_0__15154_ gnd vdd FILL
XFILL_2__11187_ gnd vdd FILL
XFILL_5__13106_ gnd vdd FILL
X_9300_ _9301_/B _7508_/B gnd _9301_/C vdd NAND2X1
XFILL_5__9647_ gnd vdd FILL
XFILL_5__10318_ gnd vdd FILL
XFILL_5__6859_ gnd vdd FILL
XFILL_0__8953_ gnd vdd FILL
XFILL_4__13836_ gnd vdd FILL
XFILL_5__11298_ gnd vdd FILL
XFILL_5__14086_ gnd vdd FILL
XFILL_3__15265_ gnd vdd FILL
XFILL_2__10138_ gnd vdd FILL
XFILL_3__12477_ gnd vdd FILL
X_7492_ _7536_/Q gnd _7492_/Y vdd INVX1
XBUFX2_insert380 _12211_/Y gnd _12307_/C vdd BUFX2
XFILL_0__11317_ gnd vdd FILL
XFILL_0__14105_ gnd vdd FILL
XFILL_2__9869_ gnd vdd FILL
XFILL_1__13656_ gnd vdd FILL
XFILL_2__15995_ gnd vdd FILL
XBUFX2_insert391 _12387_/Y gnd _7713_/B vdd BUFX2
XFILL_6__8371_ gnd vdd FILL
XFILL_0__15085_ gnd vdd FILL
XFILL_0__12297_ gnd vdd FILL
X_9231_ _9232_/B _9487_/B gnd _9231_/Y vdd NAND2X1
XFILL_5__10249_ gnd vdd FILL
XFILL_3__14216_ gnd vdd FILL
XFILL_5__13037_ gnd vdd FILL
XFILL_6__12588_ gnd vdd FILL
XFILL_3__7613_ gnd vdd FILL
XSFILL94440x69050 gnd vdd FILL
XSFILL43800x34050 gnd vdd FILL
XFILL_0__8884_ gnd vdd FILL
XFILL_3__11428_ gnd vdd FILL
XFILL_3__15196_ gnd vdd FILL
XFILL_4__13767_ gnd vdd FILL
XFILL_1__12607_ gnd vdd FILL
XSFILL49000x3050 gnd vdd FILL
XFILL_4__10979_ gnd vdd FILL
XFILL_6__7322_ gnd vdd FILL
XFILL_0__14036_ gnd vdd FILL
XFILL_2__10069_ gnd vdd FILL
XFILL_2__14946_ gnd vdd FILL
XFILL_1__16375_ gnd vdd FILL
XFILL_0__11248_ gnd vdd FILL
XFILL_3__8593_ gnd vdd FILL
XFILL_1__13587_ gnd vdd FILL
XFILL_5__8529_ gnd vdd FILL
XFILL_4__15506_ gnd vdd FILL
XFILL_0__7835_ gnd vdd FILL
XFILL_1__10799_ gnd vdd FILL
XFILL_4__12718_ gnd vdd FILL
XFILL_3__14147_ gnd vdd FILL
X_9162_ _9162_/A gnd _9164_/A vdd INVX1
XFILL_1__15326_ gnd vdd FILL
XSFILL69240x45050 gnd vdd FILL
XFILL_3__7544_ gnd vdd FILL
XFILL_3__11359_ gnd vdd FILL
XFILL_2__14877_ gnd vdd FILL
XFILL_4__13698_ gnd vdd FILL
XFILL_0__11179_ gnd vdd FILL
X_8113_ _8111_/Y _8133_/A _8113_/C gnd _8169_/D vdd OAI21X1
XSFILL29240x61050 gnd vdd FILL
XFILL_4__15437_ gnd vdd FILL
XFILL_4__12649_ gnd vdd FILL
XFILL_2__13828_ gnd vdd FILL
XFILL_5__14988_ gnd vdd FILL
X_9093_ _9179_/Q gnd _9093_/Y vdd INVX1
XFILL_3__14078_ gnd vdd FILL
XFILL_1__15257_ gnd vdd FILL
XFILL_3__7475_ gnd vdd FILL
XFILL_3_BUFX2_insert609 gnd vdd FILL
XFILL_0__9505_ gnd vdd FILL
XFILL_1__12469_ gnd vdd FILL
XFILL_0__15987_ gnd vdd FILL
X_8044_ _7992_/A _8560_/CLK _8033_/R vdd _8044_/D gnd vdd DFFSR
XFILL_3__13029_ gnd vdd FILL
XFILL_5__13939_ gnd vdd FILL
XFILL_3__9214_ gnd vdd FILL
XFILL_4__15368_ gnd vdd FILL
XFILL_1__14208_ gnd vdd FILL
XSFILL8680x52050 gnd vdd FILL
XFILL_0__7697_ gnd vdd FILL
XFILL_2__13759_ gnd vdd FILL
XSFILL98680x74050 gnd vdd FILL
XFILL_1__15188_ gnd vdd FILL
XFILL_0__14938_ gnd vdd FILL
XFILL_4__14319_ gnd vdd FILL
XFILL_3__9145_ gnd vdd FILL
XFILL_4__15299_ gnd vdd FILL
XFILL_1__14139_ gnd vdd FILL
XSFILL89400x58050 gnd vdd FILL
XFILL_0__14869_ gnd vdd FILL
XFILL_5__15609_ gnd vdd FILL
XFILL_0__9367_ gnd vdd FILL
XFILL_2__15429_ gnd vdd FILL
X_9995_ _9995_/A gnd _9995_/Y vdd INVX1
XFILL_1__7111_ gnd vdd FILL
XFILL_0__8318_ gnd vdd FILL
X_8946_ _8946_/Q _8562_/CLK _7270_/R vdd _8946_/D gnd vdd DFFSR
XFILL_1__8091_ gnd vdd FILL
XFILL_0__9298_ gnd vdd FILL
XFILL_0__8249_ gnd vdd FILL
XFILL_1__7042_ gnd vdd FILL
X_8877_ _8859_/A _9005_/B gnd _8877_/Y vdd NAND2X1
XFILL_4__8840_ gnd vdd FILL
XFILL_6__9756_ gnd vdd FILL
X_7828_ _7828_/A gnd _7830_/A vdd INVX1
XFILL_4__8771_ gnd vdd FILL
XFILL_6__8707_ gnd vdd FILL
XFILL_3__9978_ gnd vdd FILL
X_7759_ _7759_/A _7759_/B _7758_/Y gnd _7759_/Y vdd OAI21X1
XFILL_1__8993_ gnd vdd FILL
XSFILL104520x34050 gnd vdd FILL
XFILL_6__6899_ gnd vdd FILL
XFILL_4__7722_ gnd vdd FILL
XSFILL8760x32050 gnd vdd FILL
XFILL_1__7944_ gnd vdd FILL
X_11360_ _11359_/A _11359_/B _11360_/C gnd _11360_/Y vdd OAI21X1
X_9429_ _9427_/Y _9372_/B _9428_/Y gnd _9429_/Y vdd OAI21X1
XFILL_1__7875_ gnd vdd FILL
XFILL_4__7584_ gnd vdd FILL
XFILL_4_BUFX2_insert410 gnd vdd FILL
X_10311_ _10311_/A gnd _10313_/A vdd INVX1
XFILL_1__9614_ gnd vdd FILL
XFILL_4_BUFX2_insert421 gnd vdd FILL
X_11291_ _11099_/Y _11546_/A gnd _11521_/C vdd NAND2X1
XFILL_4_BUFX2_insert432 gnd vdd FILL
XFILL111960x76050 gnd vdd FILL
XFILL_4_BUFX2_insert443 gnd vdd FILL
XFILL_4_BUFX2_insert454 gnd vdd FILL
X_13030_ vdd _13030_/B gnd _13031_/C vdd NAND2X1
X_10242_ _13679_/A gnd _10244_/A vdd INVX1
XFILL_1__9545_ gnd vdd FILL
XFILL_4_BUFX2_insert465 gnd vdd FILL
XSFILL63880x61050 gnd vdd FILL
XFILL_4_BUFX2_insert476 gnd vdd FILL
XFILL_4__9254_ gnd vdd FILL
XSFILL13720x33050 gnd vdd FILL
XFILL_4_BUFX2_insert487 gnd vdd FILL
XFILL_4_BUFX2_insert498 gnd vdd FILL
XSFILL79160x28050 gnd vdd FILL
X_10173_ _10171_/Y _10191_/B _10173_/C gnd _10221_/D vdd OAI21X1
XFILL_1__9476_ gnd vdd FILL
XFILL_4__8205_ gnd vdd FILL
XFILL_2__7220_ gnd vdd FILL
X_14981_ _12813_/Q _14980_/Y gnd _14981_/Y vdd NOR2X1
XFILL_4__8136_ gnd vdd FILL
X_13932_ _13932_/A gnd _15476_/C vdd INVX1
XSFILL84280x19050 gnd vdd FILL
XFILL_1__8358_ gnd vdd FILL
XFILL_3_CLKBUF1_insert112 gnd vdd FILL
XSFILL103960x3050 gnd vdd FILL
XFILL_4__8067_ gnd vdd FILL
XFILL_3_CLKBUF1_insert123 gnd vdd FILL
XFILL_3_CLKBUF1_insert134 gnd vdd FILL
XFILL_5_CLKBUF1_insert1083 gnd vdd FILL
X_13863_ _13863_/A _13862_/Y gnd _13863_/Y vdd NOR2X1
XFILL_1__7309_ gnd vdd FILL
XFILL_3_CLKBUF1_insert145 gnd vdd FILL
XFILL_3_CLKBUF1_insert156 gnd vdd FILL
XFILL_3_CLKBUF1_insert167 gnd vdd FILL
XFILL_2__7082_ gnd vdd FILL
X_12814_ _12764_/A _12809_/CLK _12685_/R vdd _12814_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert300 gnd vdd FILL
XFILL_6__10910_ gnd vdd FILL
XFILL_3_CLKBUF1_insert178 gnd vdd FILL
XFILL_4__10000_ gnd vdd FILL
X_15602_ _15601_/Y _15602_/B gnd _15608_/A vdd NOR2X1
XFILL_5__8880_ gnd vdd FILL
XFILL_3_CLKBUF1_insert189 gnd vdd FILL
X_13794_ _9099_/A gnd _13794_/Y vdd INVX1
XFILL_1_BUFX2_insert311 gnd vdd FILL
XFILL_1_BUFX2_insert322 gnd vdd FILL
XFILL_0__10550_ gnd vdd FILL
XFILL_1_BUFX2_insert333 gnd vdd FILL
XFILL_5__7831_ gnd vdd FILL
XFILL_1_BUFX2_insert344 gnd vdd FILL
X_12745_ _12745_/A _12721_/B _12745_/C gnd _12745_/Y vdd OAI21X1
XFILL_1_BUFX2_insert355 gnd vdd FILL
X_15533_ _15533_/A _15532_/Y gnd _15533_/Y vdd NOR2X1
XFILL_5__12270_ gnd vdd FILL
XFILL_2__11110_ gnd vdd FILL
XFILL_3__10661_ gnd vdd FILL
XFILL_1_BUFX2_insert366 gnd vdd FILL
XFILL_2__12090_ gnd vdd FILL
XFILL_1_BUFX2_insert377 gnd vdd FILL
XFILL_1__11840_ gnd vdd FILL
XFILL_1_BUFX2_insert388 gnd vdd FILL
XFILL_4__8969_ gnd vdd FILL
XFILL_3__12400_ gnd vdd FILL
XSFILL63960x41050 gnd vdd FILL
XFILL_1_BUFX2_insert399 gnd vdd FILL
X_15464_ _16261_/A _15464_/B _15464_/C _16261_/D gnd _15464_/Y vdd OAI22X1
XFILL_5__7762_ gnd vdd FILL
XFILL_5__11221_ gnd vdd FILL
X_12676_ _12676_/Q _9050_/CLK _8171_/R vdd _12608_/Y gnd vdd DFFSR
XSFILL13800x13050 gnd vdd FILL
XFILL_4__11951_ gnd vdd FILL
XFILL_3__13380_ gnd vdd FILL
XFILL_0__12220_ gnd vdd FILL
XFILL_2__11041_ gnd vdd FILL
XFILL_2__7984_ gnd vdd FILL
XFILL_5__9501_ gnd vdd FILL
XFILL112120x65050 gnd vdd FILL
XFILL_1__11771_ gnd vdd FILL
X_14415_ _9778_/A gnd _14415_/Y vdd INVX1
XFILL_5__7693_ gnd vdd FILL
XFILL_5__11152_ gnd vdd FILL
X_11627_ _11627_/A _11626_/Y _11627_/C gnd _11627_/Y vdd OAI21X1
XFILL_4__10902_ gnd vdd FILL
X_15395_ _15395_/A _15394_/Y gnd _15395_/Y vdd NOR2X1
XFILL_3__12331_ gnd vdd FILL
XFILL_2__6935_ gnd vdd FILL
XFILL_4__14670_ gnd vdd FILL
XFILL_2__9723_ gnd vdd FILL
XFILL_1__13510_ gnd vdd FILL
XFILL_4__11882_ gnd vdd FILL
XSFILL64040x50050 gnd vdd FILL
XFILL_0__12151_ gnd vdd FILL
XFILL_1__14490_ gnd vdd FILL
XFILL_5__10103_ gnd vdd FILL
X_14346_ _10216_/Q gnd _14346_/Y vdd INVX1
XSFILL114440x17050 gnd vdd FILL
XFILL_4__13621_ gnd vdd FILL
XFILL_3__15050_ gnd vdd FILL
XFILL_5__15960_ gnd vdd FILL
XFILL_5__11083_ gnd vdd FILL
X_11558_ _11558_/A gnd _11558_/Y vdd INVX1
XFILL_2__14800_ gnd vdd FILL
XFILL_3__12262_ gnd vdd FILL
XFILL_0__11102_ gnd vdd FILL
XFILL_4__10833_ gnd vdd FILL
XFILL_2__9654_ gnd vdd FILL
XFILL_2__6866_ gnd vdd FILL
XFILL_1__13441_ gnd vdd FILL
XFILL_2__15780_ gnd vdd FILL
XFILL_0__12082_ gnd vdd FILL
XFILL_1__10653_ gnd vdd FILL
XFILL_2__12992_ gnd vdd FILL
X_10509_ _10509_/A _10535_/A _10508_/Y gnd _10509_/Y vdd OAI21X1
XFILL_3__14001_ gnd vdd FILL
XFILL_5__9363_ gnd vdd FILL
XFILL_5__10034_ gnd vdd FILL
XFILL_5__14911_ gnd vdd FILL
XFILL_4__16340_ gnd vdd FILL
X_14277_ _8039_/Q gnd _14278_/D vdd INVX1
XFILL_3__11213_ gnd vdd FILL
XFILL_4__10764_ gnd vdd FILL
XFILL_2__14731_ gnd vdd FILL
XFILL_4__13552_ gnd vdd FILL
XFILL_2__8605_ gnd vdd FILL
X_11489_ _11182_/Y gnd _11511_/A vdd INVX1
XFILL_5__15891_ gnd vdd FILL
XFILL_0__15910_ gnd vdd FILL
XFILL_2__11943_ gnd vdd FILL
XFILL_3__12193_ gnd vdd FILL
XFILL_1__16160_ gnd vdd FILL
XFILL_0__11033_ gnd vdd FILL
X_16016_ _16016_/A _15392_/B _16225_/C _14631_/Y gnd _16019_/A vdd OAI22X1
XFILL_1__13372_ gnd vdd FILL
XFILL_5__8314_ gnd vdd FILL
XFILL_5__9294_ gnd vdd FILL
X_13228_ _13215_/A gnd _13246_/B vdd INVX1
XFILL_0__7620_ gnd vdd FILL
XSFILL18520x25050 gnd vdd FILL
XFILL_5__14842_ gnd vdd FILL
XFILL_4__12503_ gnd vdd FILL
XFILL_3__11144_ gnd vdd FILL
XFILL_1__15111_ gnd vdd FILL
XFILL_4__16271_ gnd vdd FILL
XFILL_1__12323_ gnd vdd FILL
XFILL_2__14662_ gnd vdd FILL
XFILL_4__13483_ gnd vdd FILL
XFILL_4__10695_ gnd vdd FILL
XFILL_2__11874_ gnd vdd FILL
XFILL_5__8245_ gnd vdd FILL
XFILL_1__16091_ gnd vdd FILL
XFILL_0__15841_ gnd vdd FILL
XFILL_0__7551_ gnd vdd FILL
X_13159_ _13157_/Y _13149_/A _13159_/C gnd _13201_/D vdd OAI21X1
XFILL_4__15222_ gnd vdd FILL
XFILL_2__13613_ gnd vdd FILL
XFILL_4__12434_ gnd vdd FILL
XFILL_2__16401_ gnd vdd FILL
XFILL_5__14773_ gnd vdd FILL
XSFILL104360x69050 gnd vdd FILL
XFILL_5__11985_ gnd vdd FILL
XFILL_1__15042_ gnd vdd FILL
XFILL_3__15952_ gnd vdd FILL
XFILL_3__11075_ gnd vdd FILL
XFILL_2__8467_ gnd vdd FILL
XFILL_2__10825_ gnd vdd FILL
XFILL_2__14593_ gnd vdd FILL
XFILL_1__12254_ gnd vdd FILL
XFILL_0__15772_ gnd vdd FILL
XFILL_0__12984_ gnd vdd FILL
XFILL_5__13724_ gnd vdd FILL
XFILL_4__12365_ gnd vdd FILL
XFILL_5__10936_ gnd vdd FILL
XFILL_2__16332_ gnd vdd FILL
XFILL_0__7482_ gnd vdd FILL
XFILL_4__15153_ gnd vdd FILL
XFILL_2__7418_ gnd vdd FILL
XFILL_3__14903_ gnd vdd FILL
XFILL_3__10026_ gnd vdd FILL
XFILL_1__11205_ gnd vdd FILL
XFILL_2__13544_ gnd vdd FILL
XFILL_2__8398_ gnd vdd FILL
XFILL_2__10756_ gnd vdd FILL
XFILL_3__7191_ gnd vdd FILL
XFILL_0__14723_ gnd vdd FILL
XFILL_3__15883_ gnd vdd FILL
XFILL_1__12185_ gnd vdd FILL
XFILL_0__11935_ gnd vdd FILL
XFILL_0__9221_ gnd vdd FILL
XFILL_4__14104_ gnd vdd FILL
XFILL_5__13655_ gnd vdd FILL
XFILL_4__11316_ gnd vdd FILL
XFILL_2__7349_ gnd vdd FILL
XFILL_3__14834_ gnd vdd FILL
XFILL_2__16263_ gnd vdd FILL
XFILL_4__12296_ gnd vdd FILL
XFILL_4__15084_ gnd vdd FILL
XFILL_2__13475_ gnd vdd FILL
XFILL_1__11136_ gnd vdd FILL
XFILL_2__10687_ gnd vdd FILL
XFILL_0__14654_ gnd vdd FILL
XFILL_5__7058_ gnd vdd FILL
XFILL_0__9152_ gnd vdd FILL
XFILL_5__12606_ gnd vdd FILL
XFILL_0__11866_ gnd vdd FILL
X_8800_ _8724_/A _7535_/CLK _7648_/R vdd _8726_/Y gnd vdd DFFSR
XFILL_2__15214_ gnd vdd FILL
XFILL_4__14035_ gnd vdd FILL
XSFILL64120x30050 gnd vdd FILL
XFILL_5__16374_ gnd vdd FILL
XFILL_4__11247_ gnd vdd FILL
XFILL_5__13586_ gnd vdd FILL
XFILL_2__12426_ gnd vdd FILL
X_9780_ _9780_/A _9785_/A _9779_/Y gnd _9834_/D vdd OAI21X1
XFILL_0__13605_ gnd vdd FILL
XFILL_2__16194_ gnd vdd FILL
XFILL_1__15944_ gnd vdd FILL
XFILL_3__11977_ gnd vdd FILL
XFILL_5__10798_ gnd vdd FILL
XFILL_1__11067_ gnd vdd FILL
X_6992_ _6992_/A gnd _6994_/A vdd INVX1
XFILL_3__14765_ gnd vdd FILL
XFILL_0__8103_ gnd vdd FILL
XFILL_0__10817_ gnd vdd FILL
XFILL_0__14585_ gnd vdd FILL
XFILL_5__15325_ gnd vdd FILL
XFILL_2__9019_ gnd vdd FILL
XFILL_6__14876_ gnd vdd FILL
X_8731_ _8695_/B _7579_/B gnd _8731_/Y vdd NAND2X1
XFILL_0__11797_ gnd vdd FILL
XFILL_0__9083_ gnd vdd FILL
XFILL_3__10928_ gnd vdd FILL
XFILL_3__13716_ gnd vdd FILL
XFILL_4__11178_ gnd vdd FILL
XFILL_2__15145_ gnd vdd FILL
XFILL_3__9901_ gnd vdd FILL
XFILL_1__10018_ gnd vdd FILL
XFILL_2__12357_ gnd vdd FILL
XFILL_6_BUFX2_insert505 gnd vdd FILL
XFILL_0__16324_ gnd vdd FILL
XFILL_3__14696_ gnd vdd FILL
XFILL_0__13536_ gnd vdd FILL
XFILL_1__15875_ gnd vdd FILL
XSFILL53960x73050 gnd vdd FILL
XFILL_0__10748_ gnd vdd FILL
XFILL_6__13827_ gnd vdd FILL
XFILL_5__15256_ gnd vdd FILL
XSFILL99880x7050 gnd vdd FILL
XFILL_4__10129_ gnd vdd FILL
X_8662_ _8662_/Q _8022_/CLK _9046_/R vdd _8662_/D gnd vdd DFFSR
XFILL_5__12468_ gnd vdd FILL
XSFILL4040x44050 gnd vdd FILL
XFILL_2__11308_ gnd vdd FILL
XFILL_1__14826_ gnd vdd FILL
XFILL_4__15986_ gnd vdd FILL
XFILL_3__13647_ gnd vdd FILL
XFILL_2__15076_ gnd vdd FILL
XFILL_2__12288_ gnd vdd FILL
XFILL_0__16255_ gnd vdd FILL
XFILL_0__10679_ gnd vdd FILL
XFILL_5__14207_ gnd vdd FILL
XFILL_0__13467_ gnd vdd FILL
X_7613_ _7613_/A _7592_/B _7613_/C gnd _7661_/D vdd OAI21X1
XFILL_5__11419_ gnd vdd FILL
XFILL_5__15187_ gnd vdd FILL
XSFILL29240x56050 gnd vdd FILL
XFILL_2__14027_ gnd vdd FILL
XFILL_4__14937_ gnd vdd FILL
XSFILL54040x82050 gnd vdd FILL
XFILL_0__15206_ gnd vdd FILL
XFILL_5__12399_ gnd vdd FILL
XFILL_3__13578_ gnd vdd FILL
X_8593_ _8671_/Q gnd _8593_/Y vdd INVX1
XFILL_2__11239_ gnd vdd FILL
XFILL_3__16366_ gnd vdd FILL
XFILL_3__9763_ gnd vdd FILL
XFILL_3__6975_ gnd vdd FILL
XFILL_0__12418_ gnd vdd FILL
XFILL_1__14757_ gnd vdd FILL
XFILL_0__16186_ gnd vdd FILL
XFILL_1__11969_ gnd vdd FILL
XFILL_6__9472_ gnd vdd FILL
XFILL_0__13398_ gnd vdd FILL
XFILL_5__14138_ gnd vdd FILL
XSFILL104440x49050 gnd vdd FILL
XFILL_3__15317_ gnd vdd FILL
X_7544_ _7542_/Y _7562_/B _7543_/Y gnd _7544_/Y vdd OAI21X1
XFILL_6__13689_ gnd vdd FILL
XFILL_0__9985_ gnd vdd FILL
XFILL_4__14868_ gnd vdd FILL
XFILL_3__8714_ gnd vdd FILL
XFILL_3__12529_ gnd vdd FILL
XFILL_1__13708_ gnd vdd FILL
XSFILL8680x47050 gnd vdd FILL
XFILL_3__16297_ gnd vdd FILL
XFILL_0__15137_ gnd vdd FILL
XFILL_0__12349_ gnd vdd FILL
XFILL_1__14688_ gnd vdd FILL
XFILL_4__13819_ gnd vdd FILL
XFILL_5__14069_ gnd vdd FILL
XFILL_3__15248_ gnd vdd FILL
X_7475_ _7430_/A _8243_/B gnd _7476_/C vdd NAND2X1
XFILL_1__13639_ gnd vdd FILL
XFILL_4__14799_ gnd vdd FILL
XFILL_3__8645_ gnd vdd FILL
XSFILL59160x4050 gnd vdd FILL
XFILL_2__15978_ gnd vdd FILL
XFILL_0__15068_ gnd vdd FILL
X_9214_ _9212_/Y _9238_/B _9214_/C gnd _9214_/Y vdd OAI21X1
XSFILL99320x9050 gnd vdd FILL
XFILL_0__8867_ gnd vdd FILL
XSFILL48920x62050 gnd vdd FILL
XFILL_3__8576_ gnd vdd FILL
XFILL_3__15179_ gnd vdd FILL
XFILL_0__14019_ gnd vdd FILL
XFILL_1__16358_ gnd vdd FILL
XFILL_2__14929_ gnd vdd FILL
XSFILL64200x10050 gnd vdd FILL
XFILL_0__7818_ gnd vdd FILL
X_9145_ _9164_/B _8889_/B gnd _9146_/C vdd NAND2X1
XFILL_1__7591_ gnd vdd FILL
XFILL_1__15309_ gnd vdd FILL
XSFILL108680x54050 gnd vdd FILL
XFILL_3_BUFX2_insert406 gnd vdd FILL
XFILL_1__16289_ gnd vdd FILL
XFILL_3_BUFX2_insert417 gnd vdd FILL
XFILL_0__7749_ gnd vdd FILL
XFILL_3_BUFX2_insert428 gnd vdd FILL
X_9076_ _9040_/A _9328_/CLK _7152_/R vdd _9076_/D gnd vdd DFFSR
XFILL_3__7458_ gnd vdd FILL
XFILL_3_BUFX2_insert439 gnd vdd FILL
XFILL_6__7167_ gnd vdd FILL
XFILL_1__9261_ gnd vdd FILL
X_8027_ _7941_/A _8152_/CLK _9944_/R vdd _7943_/Y gnd vdd DFFSR
XFILL_0__9419_ gnd vdd FILL
XFILL_1__8212_ gnd vdd FILL
XSFILL54120x62050 gnd vdd FILL
XFILL_3__9128_ gnd vdd FILL
XFILL_1__8143_ gnd vdd FILL
X_9978_ _9979_/B _9978_/B gnd _9978_/Y vdd NAND2X1
XFILL_4__9941_ gnd vdd FILL
X_10860_ _14522_/A _7020_/CLK _8053_/R vdd _10860_/D gnd vdd DFFSR
XFILL_1__8074_ gnd vdd FILL
X_8929_ _8855_/A _9453_/CLK _8929_/R vdd _8929_/D gnd vdd DFFSR
XFILL_4_CLKBUF1_insert207 gnd vdd FILL
XFILL_4__9872_ gnd vdd FILL
XFILL_6__9808_ gnd vdd FILL
XFILL_4_CLKBUF1_insert218 gnd vdd FILL
XSFILL18760x81050 gnd vdd FILL
X_10791_ _10792_/B _9895_/B gnd _10791_/Y vdd NAND2X1
XFILL_4__8823_ gnd vdd FILL
X_12530_ vdd _12109_/A gnd _12531_/C vdd NAND2X1
XFILL_0_BUFX2_insert307 gnd vdd FILL
XFILL_0_BUFX2_insert318 gnd vdd FILL
XSFILL13720x28050 gnd vdd FILL
XFILL_0_BUFX2_insert329 gnd vdd FILL
XFILL_4__8754_ gnd vdd FILL
X_12461_ vdd _12461_/B gnd _12461_/Y vdd NAND2X1
XFILL_1__8976_ gnd vdd FILL
X_14200_ _14199_/Y _14045_/A _14200_/C _14198_/Y gnd _14204_/A vdd OAI22X1
XFILL_4__7705_ gnd vdd FILL
XSFILL28920x50 gnd vdd FILL
X_11412_ _11419_/A gnd _11412_/Y vdd INVX1
X_15180_ _13613_/Y _15407_/B _15180_/C _15179_/Y gnd _15183_/B vdd OAI22X1
X_12392_ _12380_/A _12615_/A gnd _12393_/C vdd NAND2X1
XFILL_1__7927_ gnd vdd FILL
X_14131_ _13813_/B gnd _14482_/B vdd INVX2
XSFILL54200x42050 gnd vdd FILL
XFILL_4__7636_ gnd vdd FILL
X_11343_ _11211_/Y _11212_/A gnd _11343_/Y vdd NOR2X1
XFILL_1__7858_ gnd vdd FILL
XFILL_4__7567_ gnd vdd FILL
XFILL_4_BUFX2_insert240 gnd vdd FILL
X_14062_ _14062_/A _14061_/Y gnd _14063_/A vdd NOR2X1
X_11274_ _11274_/A _11083_/Y gnd _11275_/A vdd NAND2X1
XFILL_4_BUFX2_insert251 gnd vdd FILL
XFILL_2__9370_ gnd vdd FILL
XFILL_4_BUFX2_insert262 gnd vdd FILL
XFILL_4_BUFX2_insert273 gnd vdd FILL
XSFILL84680x35050 gnd vdd FILL
XFILL_4_BUFX2_insert284 gnd vdd FILL
X_13013_ _13011_/Y vdd _13013_/C gnd _13013_/Y vdd OAI21X1
XFILL_4__7498_ gnd vdd FILL
X_10225_ _10225_/Q _7786_/CLK _7153_/R vdd _10225_/D gnd vdd DFFSR
XFILL_2__8321_ gnd vdd FILL
XFILL_4_BUFX2_insert295 gnd vdd FILL
XFILL_5_BUFX2_insert1008 gnd vdd FILL
XFILL_1__9528_ gnd vdd FILL
XFILL_5_BUFX2_insert1019 gnd vdd FILL
XSFILL18840x61050 gnd vdd FILL
XFILL_4__9237_ gnd vdd FILL
XSFILL19320x68050 gnd vdd FILL
XFILL_3_BUFX2_insert940 gnd vdd FILL
XFILL_3_BUFX2_insert951 gnd vdd FILL
X_10156_ _10216_/Q gnd _10158_/A vdd INVX1
XFILL_2__8252_ gnd vdd FILL
XFILL_5__11770_ gnd vdd FILL
XFILL_3_BUFX2_insert962 gnd vdd FILL
XFILL_3_BUFX2_insert973 gnd vdd FILL
XFILL_2__11590_ gnd vdd FILL
XFILL_4__9168_ gnd vdd FILL
XFILL_3_BUFX2_insert984 gnd vdd FILL
XFILL_3_BUFX2_insert995 gnd vdd FILL
XFILL_2__7203_ gnd vdd FILL
XFILL_4__12150_ gnd vdd FILL
XFILL_3__11900_ gnd vdd FILL
X_14964_ _14964_/A _14956_/Y _14964_/C gnd _14964_/Y vdd NAND3X1
X_10087_ _10087_/Q _7527_/CLK _8935_/R vdd _10027_/Y gnd vdd DFFSR
XFILL_2__8183_ gnd vdd FILL
XFILL_2__10541_ gnd vdd FILL
XFILL_3__12880_ gnd vdd FILL
XFILL_4__8119_ gnd vdd FILL
XFILL_0__11720_ gnd vdd FILL
XFILL_4__9099_ gnd vdd FILL
XFILL_4__11101_ gnd vdd FILL
XFILL_5__13440_ gnd vdd FILL
XFILL_5__9981_ gnd vdd FILL
X_13915_ _7441_/A gnd _13915_/Y vdd INVX1
XFILL_4__12081_ gnd vdd FILL
XFILL_5__10652_ gnd vdd FILL
XFILL_6__12991_ gnd vdd FILL
XFILL_3__11831_ gnd vdd FILL
XFILL_2__13260_ gnd vdd FILL
X_14895_ _9844_/Q gnd _14895_/Y vdd INVX1
XSFILL64040x45050 gnd vdd FILL
XFILL_3_BUFX2_insert1001 gnd vdd FILL
XFILL_3_BUFX2_insert1012 gnd vdd FILL
XFILL_1__13990_ gnd vdd FILL
XFILL_0__11651_ gnd vdd FILL
XFILL_6__11942_ gnd vdd FILL
XFILL_4__11032_ gnd vdd FILL
XFILL_3_BUFX2_insert1023 gnd vdd FILL
X_13846_ _13846_/A _13844_/Y _13846_/C _14203_/B gnd _13846_/Y vdd OAI22X1
XFILL_5__13371_ gnd vdd FILL
XFILL_3_BUFX2_insert1034 gnd vdd FILL
XFILL_2__12211_ gnd vdd FILL
XFILL_3__14550_ gnd vdd FILL
XFILL_2__7065_ gnd vdd FILL
XFILL_3__11762_ gnd vdd FILL
XSFILL78600x60050 gnd vdd FILL
XFILL_3_BUFX2_insert1045 gnd vdd FILL
XFILL_3_BUFX2_insert1056 gnd vdd FILL
XFILL_0__14370_ gnd vdd FILL
XFILL_0__11582_ gnd vdd FILL
XFILL_5__15110_ gnd vdd FILL
XFILL_5__12322_ gnd vdd FILL
XFILL_6__14661_ gnd vdd FILL
XFILL_5__8863_ gnd vdd FILL
XFILL_3_BUFX2_insert1067 gnd vdd FILL
X_13777_ _8156_/Q gnd _13777_/Y vdd INVX1
XFILL_5__16090_ gnd vdd FILL
XFILL_4__15840_ gnd vdd FILL
XFILL_3__13501_ gnd vdd FILL
XFILL_3_BUFX2_insert1089 gnd vdd FILL
XFILL_3__14481_ gnd vdd FILL
XFILL_2__12142_ gnd vdd FILL
X_10989_ _12210_/Y _10988_/B gnd _10989_/Y vdd NAND2X1
XFILL_0__13321_ gnd vdd FILL
XFILL_0__10533_ gnd vdd FILL
XFILL_1__15660_ gnd vdd FILL
XFILL_3__11693_ gnd vdd FILL
XFILL_1__12872_ gnd vdd FILL
XFILL_5__7814_ gnd vdd FILL
XFILL_5__15041_ gnd vdd FILL
X_15516_ _6935_/A gnd _15516_/Y vdd INVX1
X_12728_ _12802_/Q gnd _12728_/Y vdd INVX1
XFILL_3__16220_ gnd vdd FILL
XFILL_3__13432_ gnd vdd FILL
XFILL_5__12253_ gnd vdd FILL
XFILL_1__14611_ gnd vdd FILL
XFILL_4__15771_ gnd vdd FILL
XFILL_3__10644_ gnd vdd FILL
XFILL_0__16040_ gnd vdd FILL
XFILL_2__12073_ gnd vdd FILL
XFILL_4__12983_ gnd vdd FILL
XFILL_1__11823_ gnd vdd FILL
XFILL_0__13252_ gnd vdd FILL
XFILL_1__15591_ gnd vdd FILL
XSFILL84200x58050 gnd vdd FILL
XFILL_0_BUFX2_insert830 gnd vdd FILL
XFILL_5__7745_ gnd vdd FILL
XFILL_5__11204_ gnd vdd FILL
X_12659_ _12657_/Y vdd _12659_/C gnd _12693_/D vdd OAI21X1
XFILL_6__10755_ gnd vdd FILL
XFILL_4__14722_ gnd vdd FILL
X_15447_ _8415_/Q gnd _15449_/A vdd INVX1
XFILL_0_BUFX2_insert841 gnd vdd FILL
XFILL_3__13363_ gnd vdd FILL
XFILL_0_BUFX2_insert852 gnd vdd FILL
XFILL_2__15901_ gnd vdd FILL
XFILL_4__11934_ gnd vdd FILL
XFILL_5__12184_ gnd vdd FILL
XFILL_2__11024_ gnd vdd FILL
XFILL_3__16151_ gnd vdd FILL
XFILL_3__10575_ gnd vdd FILL
XFILL_0__12203_ gnd vdd FILL
XFILL_1__14542_ gnd vdd FILL
XFILL_1__11754_ gnd vdd FILL
XFILL_0_BUFX2_insert863 gnd vdd FILL
XFILL_2__7967_ gnd vdd FILL
XFILL_0_BUFX2_insert874 gnd vdd FILL
XFILL_0__10395_ gnd vdd FILL
XFILL_0__9770_ gnd vdd FILL
XFILL_6__13474_ gnd vdd FILL
XFILL_3__12314_ gnd vdd FILL
XFILL_0_BUFX2_insert885 gnd vdd FILL
XFILL_5__7676_ gnd vdd FILL
XFILL_5__11135_ gnd vdd FILL
XFILL_3__15102_ gnd vdd FILL
X_15378_ _15378_/A _15378_/B gnd _15378_/Y vdd NOR2X1
XFILL_0_BUFX2_insert896 gnd vdd FILL
XFILL_0__6982_ gnd vdd FILL
XFILL_4__14653_ gnd vdd FILL
XFILL_3__16082_ gnd vdd FILL
XFILL_3__13294_ gnd vdd FILL
XFILL_0__12134_ gnd vdd FILL
XFILL_1_BUFX2_insert1060 gnd vdd FILL
XFILL_2__15832_ gnd vdd FILL
XFILL_4__11865_ gnd vdd FILL
XFILL_2__6918_ gnd vdd FILL
XFILL_1__10705_ gnd vdd FILL
XFILL_1__14473_ gnd vdd FILL
XFILL_1_BUFX2_insert1071 gnd vdd FILL
XFILL_3_BUFX2_insert12 gnd vdd FILL
XFILL_5__9415_ gnd vdd FILL
XFILL_0__8721_ gnd vdd FILL
XFILL_1__11685_ gnd vdd FILL
XFILL_3_BUFX2_insert23 gnd vdd FILL
XFILL_4__13604_ gnd vdd FILL
XFILL_3_BUFX2_insert34 gnd vdd FILL
XFILL_5__15943_ gnd vdd FILL
XFILL_1_BUFX2_insert1093 gnd vdd FILL
X_14329_ _9960_/Q gnd _14330_/D vdd INVX1
X_7260_ _7260_/Q _8926_/CLK _7262_/R vdd _7260_/D gnd vdd DFFSR
XFILL_4__10816_ gnd vdd FILL
XFILL_1__16212_ gnd vdd FILL
XFILL_3__15033_ gnd vdd FILL
XFILL_3__12245_ gnd vdd FILL
XFILL_3_BUFX2_insert45 gnd vdd FILL
XFILL_5__11066_ gnd vdd FILL
XFILL_2__9637_ gnd vdd FILL
XFILL_4__14584_ gnd vdd FILL
XFILL_1__13424_ gnd vdd FILL
XFILL_2__6849_ gnd vdd FILL
XFILL_3_BUFX2_insert56 gnd vdd FILL
XFILL_1__10636_ gnd vdd FILL
XFILL_2__12975_ gnd vdd FILL
XFILL_0__12065_ gnd vdd FILL
XFILL_2__15763_ gnd vdd FILL
XFILL_4__11796_ gnd vdd FILL
XFILL_5__9346_ gnd vdd FILL
XFILL_3_BUFX2_insert67 gnd vdd FILL
XSFILL89480x27050 gnd vdd FILL
XSFILL23720x8050 gnd vdd FILL
XFILL_0__8652_ gnd vdd FILL
XFILL_5__10017_ gnd vdd FILL
XFILL_3_BUFX2_insert78 gnd vdd FILL
XFILL_4__16323_ gnd vdd FILL
XFILL_3_BUFX2_insert89 gnd vdd FILL
X_7191_ _7191_/A gnd _7191_/Y vdd INVX1
XFILL_4__13535_ gnd vdd FILL
XFILL_5__15874_ gnd vdd FILL
XSFILL64120x25050 gnd vdd FILL
XFILL_2__14714_ gnd vdd FILL
XFILL_2__11926_ gnd vdd FILL
XFILL_1__16143_ gnd vdd FILL
XFILL_3__8361_ gnd vdd FILL
XFILL_4__10747_ gnd vdd FILL
XFILL_3__12176_ gnd vdd FILL
XFILL_0__11016_ gnd vdd FILL
XFILL_1__13355_ gnd vdd FILL
XFILL_2__15694_ gnd vdd FILL
XFILL_0__7603_ gnd vdd FILL
XFILL_1__10567_ gnd vdd FILL
XFILL_5__9277_ gnd vdd FILL
XFILL_5__14825_ gnd vdd FILL
XFILL_3__7312_ gnd vdd FILL
XFILL_3__11127_ gnd vdd FILL
XFILL_0__8583_ gnd vdd FILL
XFILL_4__16254_ gnd vdd FILL
XFILL_4__13466_ gnd vdd FILL
XFILL_2__8519_ gnd vdd FILL
XFILL_1__12306_ gnd vdd FILL
XSFILL43880x50 gnd vdd FILL
XFILL_4__10678_ gnd vdd FILL
XFILL_2__14645_ gnd vdd FILL
XFILL_2__9499_ gnd vdd FILL
XFILL_0__15824_ gnd vdd FILL
XFILL_1__16074_ gnd vdd FILL
XFILL_2__11857_ gnd vdd FILL
XFILL_5__8228_ gnd vdd FILL
XFILL_1__13286_ gnd vdd FILL
XFILL_6_CLKBUF1_insert162 gnd vdd FILL
XSFILL53960x68050 gnd vdd FILL
XFILL_4__15205_ gnd vdd FILL
XFILL_6_CLKBUF1_insert173 gnd vdd FILL
XFILL_1__10498_ gnd vdd FILL
XFILL_4__12417_ gnd vdd FILL
XSFILL3560x32050 gnd vdd FILL
XFILL_5__14756_ gnd vdd FILL
XFILL_3__7243_ gnd vdd FILL
XFILL_4__16185_ gnd vdd FILL
XFILL_1__15025_ gnd vdd FILL
XFILL_3__15935_ gnd vdd FILL
XFILL_5__11968_ gnd vdd FILL
XFILL_2__10808_ gnd vdd FILL
XFILL_3__11058_ gnd vdd FILL
XFILL_2__14576_ gnd vdd FILL
XFILL_4__13397_ gnd vdd FILL
XFILL_1__12237_ gnd vdd FILL
XSFILL13160x65050 gnd vdd FILL
XFILL_2__11788_ gnd vdd FILL
XFILL_0__15755_ gnd vdd FILL
XFILL_5__13707_ gnd vdd FILL
XFILL_0__12967_ gnd vdd FILL
X_9901_ _9902_/B _9901_/B gnd _9901_/Y vdd NAND2X1
XFILL_5__10919_ gnd vdd FILL
XFILL_3__10009_ gnd vdd FILL
XFILL_0__7465_ gnd vdd FILL
XFILL_4__15136_ gnd vdd FILL
XFILL_2__13527_ gnd vdd FILL
XFILL_4__12348_ gnd vdd FILL
XFILL_2__16315_ gnd vdd FILL
XFILL_5__14687_ gnd vdd FILL
XSFILL54040x77050 gnd vdd FILL
XFILL_5__11899_ gnd vdd FILL
XFILL_0__14706_ gnd vdd FILL
XFILL_3__7174_ gnd vdd FILL
XFILL_3__15866_ gnd vdd FILL
XFILL_0__11918_ gnd vdd FILL
XFILL_1__12168_ gnd vdd FILL
XFILL_0__15686_ gnd vdd FILL
XFILL_5__13638_ gnd vdd FILL
X_9832_ _9772_/A _7527_/CLK _8935_/R vdd _9832_/D gnd vdd DFFSR
XFILL_0__12898_ gnd vdd FILL
XFILL_3__14817_ gnd vdd FILL
XFILL_4__15067_ gnd vdd FILL
XFILL_2__13458_ gnd vdd FILL
XFILL_4__12279_ gnd vdd FILL
XFILL_1__11119_ gnd vdd FILL
XFILL_2__16246_ gnd vdd FILL
XFILL_0__14637_ gnd vdd FILL
XFILL_3__15797_ gnd vdd FILL
XFILL_1__12099_ gnd vdd FILL
XFILL_0__9135_ gnd vdd FILL
XFILL_0__11849_ gnd vdd FILL
XFILL_4__14018_ gnd vdd FILL
XFILL_5__16357_ gnd vdd FILL
XSFILL3560x1050 gnd vdd FILL
X_9763_ _9829_/Q gnd _9763_/Y vdd INVX1
XFILL_2__12409_ gnd vdd FILL
XFILL_5__13569_ gnd vdd FILL
XSFILL33880x35050 gnd vdd FILL
X_6975_ _6988_/B _8255_/B gnd _6976_/C vdd NAND2X1
XFILL_2__16177_ gnd vdd FILL
XFILL_3__14748_ gnd vdd FILL
XFILL_1__15927_ gnd vdd FILL
XFILL_2__13389_ gnd vdd FILL
XFILL_0__14568_ gnd vdd FILL
XFILL_5__15308_ gnd vdd FILL
XFILL111800x13050 gnd vdd FILL
X_8714_ _8714_/A _8714_/B _8713_/Y gnd _8714_/Y vdd OAI21X1
XFILL_6__7854_ gnd vdd FILL
XFILL_5__16288_ gnd vdd FILL
XFILL_2__15128_ gnd vdd FILL
X_9694_ _9694_/Q _8926_/CLK _7262_/R vdd _9616_/Y gnd vdd DFFSR
XSFILL48920x57050 gnd vdd FILL
XFILL_0__16307_ gnd vdd FILL
XFILL_3__14679_ gnd vdd FILL
XFILL_0__13519_ gnd vdd FILL
XFILL_0__8017_ gnd vdd FILL
XFILL_1__15858_ gnd vdd FILL
XFILL_0__14499_ gnd vdd FILL
XFILL_6_BUFX2_insert357 gnd vdd FILL
XFILL_5__15239_ gnd vdd FILL
X_8645_ _8609_/A _9413_/B gnd _8646_/C vdd NAND2X1
XFILL_4__15969_ gnd vdd FILL
XFILL_2__15059_ gnd vdd FILL
XFILL_0__16238_ gnd vdd FILL
XFILL_1__14809_ gnd vdd FILL
XFILL_1__15789_ gnd vdd FILL
XFILL_6__9524_ gnd vdd FILL
XSFILL49000x66050 gnd vdd FILL
XFILL_1__8830_ gnd vdd FILL
X_8576_ _8577_/B _8576_/B gnd _8576_/Y vdd NAND2X1
XFILL_3__16349_ gnd vdd FILL
XSFILL89400x71050 gnd vdd FILL
XFILL_3__9746_ gnd vdd FILL
XFILL_0__16169_ gnd vdd FILL
XFILL_3__6958_ gnd vdd FILL
XSFILL3640x12050 gnd vdd FILL
XFILL_1__8761_ gnd vdd FILL
X_7527_ _7527_/Q _7527_/CLK _8935_/R vdd _7527_/D gnd vdd DFFSR
XFILL_4__8470_ gnd vdd FILL
XFILL_3__9677_ gnd vdd FILL
XSFILL79480x59050 gnd vdd FILL
XFILL_3__6889_ gnd vdd FILL
XFILL_1__7712_ gnd vdd FILL
X_7458_ _7456_/Y _7457_/A _7458_/C gnd _7524_/D vdd OAI21X1
XFILL_4__7421_ gnd vdd FILL
XFILL_3__8628_ gnd vdd FILL
XFILL_0__9899_ gnd vdd FILL
X_7389_ _7389_/Q _7389_/CLK _7531_/R vdd _7389_/D gnd vdd DFFSR
XFILL_4__7352_ gnd vdd FILL
X_9128_ _9126_/Y _9164_/B _9128_/C gnd _9190_/D vdd OAI21X1
XFILL_1__7574_ gnd vdd FILL
XFILL_3_BUFX2_insert225 gnd vdd FILL
X_10010_ _10082_/Q gnd _10010_/Y vdd INVX1
XFILL_3_BUFX2_insert236 gnd vdd FILL
XSFILL18760x76050 gnd vdd FILL
XFILL_3_BUFX2_insert247 gnd vdd FILL
XFILL_3_BUFX2_insert258 gnd vdd FILL
X_9059_ _9059_/Q _7651_/CLK _7011_/R vdd _8991_/Y gnd vdd DFFSR
XFILL_4__9022_ gnd vdd FILL
XFILL_3_BUFX2_insert269 gnd vdd FILL
XSFILL88600x23050 gnd vdd FILL
XFILL_2_BUFX2_insert903 gnd vdd FILL
XFILL_1__9244_ gnd vdd FILL
XFILL_2_BUFX2_insert914 gnd vdd FILL
XFILL_2_BUFX2_insert925 gnd vdd FILL
XFILL_2_BUFX2_insert936 gnd vdd FILL
X_11961_ _11961_/A _11975_/A _11961_/C gnd _6862_/A vdd OAI21X1
XFILL_2_BUFX2_insert947 gnd vdd FILL
XFILL_2_BUFX2_insert958 gnd vdd FILL
XFILL_2_BUFX2_insert969 gnd vdd FILL
XSFILL38680x27050 gnd vdd FILL
X_10912_ _10897_/Y _10910_/B gnd _10938_/B vdd NAND2X1
X_13700_ _13700_/A gnd _13701_/B vdd INVX1
XFILL_1__8126_ gnd vdd FILL
X_14680_ _14680_/A _14680_/B _14680_/C gnd _14691_/B vdd NAND3X1
X_11892_ _11892_/A _11969_/A _11891_/Y gnd _6839_/A vdd OAI21X1
XFILL_4__9924_ gnd vdd FILL
X_13631_ _9343_/A gnd _13631_/Y vdd INVX1
X_10843_ _15268_/A _7640_/CLK _7896_/R vdd _10759_/Y gnd vdd DFFSR
XFILL_1__8057_ gnd vdd FILL
XFILL_4__9855_ gnd vdd FILL
XSFILL79160x41050 gnd vdd FILL
X_13562_ _9176_/Q gnd _13562_/Y vdd INVX1
X_16350_ _16350_/A gnd _16349_/Y gnd _16426_/D vdd OAI21X1
XBUFX2_insert902 _15072_/Y gnd _15980_/C vdd BUFX2
X_10774_ _10772_/Y _10773_/A _10774_/C gnd _10774_/Y vdd OAI21X1
XFILL_0_BUFX2_insert104 gnd vdd FILL
XBUFX2_insert913 _12360_/Y gnd _8582_/B vdd BUFX2
XFILL_2__8870_ gnd vdd FILL
XBUFX2_insert924 _13370_/Y gnd _14739_/C vdd BUFX2
X_12513_ _12511_/Y vdd _12513_/C gnd _12513_/Y vdd OAI21X1
X_15301_ _15301_/A _15394_/B _16225_/C _13783_/Y gnd _15302_/A vdd OAI22X1
XBUFX2_insert935 _13423_/Y gnd _14567_/D vdd BUFX2
XBUFX2_insert946 _11987_/Y gnd _12113_/B vdd BUFX2
XFILL_4__9786_ gnd vdd FILL
X_16281_ _16273_/Y _16281_/B _16268_/Y gnd _16281_/Y vdd NAND3X1
X_13493_ _7639_/Q _14290_/C _13493_/C gnd _13493_/Y vdd AOI21X1
XFILL_2__7821_ gnd vdd FILL
XBUFX2_insert957 _13365_/Y gnd _10797_/A vdd BUFX2
XBUFX2_insert968 _12417_/Y gnd _7231_/B vdd BUFX2
XBUFX2_insert979 _13455_/Y gnd _13871_/D vdd BUFX2
XSFILL18840x56050 gnd vdd FILL
XFILL_4__8737_ gnd vdd FILL
X_15232_ _9986_/A gnd _15232_/Y vdd INVX1
X_12444_ _12442_/Y vdd _12443_/Y gnd _12444_/Y vdd OAI21X1
XFILL_3__10360_ gnd vdd FILL
XFILL_2__7752_ gnd vdd FILL
XFILL_1__8959_ gnd vdd FILL
XFILL_5__7461_ gnd vdd FILL
XFILL_0__10180_ gnd vdd FILL
X_15163_ _16306_/A _15163_/B _13562_/Y _16314_/D gnd _15164_/B vdd OAI22X1
XSFILL99320x54050 gnd vdd FILL
X_12375_ _12373_/Y _12395_/A _12375_/C gnd _12375_/Y vdd OAI21X1
XFILL_4__11650_ gnd vdd FILL
XFILL_2__7683_ gnd vdd FILL
XFILL_3__10291_ gnd vdd FILL
X_14114_ _9501_/A gnd _14115_/D vdd INVX1
XFILL_4__7619_ gnd vdd FILL
XFILL_1__11470_ gnd vdd FILL
X_11326_ _11325_/Y gnd _11331_/B vdd INVX1
XFILL_4__8599_ gnd vdd FILL
XFILL_3__12030_ gnd vdd FILL
X_15094_ _15094_/A _15094_/B _15093_/Y gnd _15094_/Y vdd NAND3X1
XFILL_2__9422_ gnd vdd FILL
XFILL_4__11581_ gnd vdd FILL
XFILL_1__10421_ gnd vdd FILL
XFILL_2__12760_ gnd vdd FILL
XFILL112280x14050 gnd vdd FILL
XFILL_5__9131_ gnd vdd FILL
X_14045_ _14045_/A _14044_/Y _13420_/B _14045_/D gnd _14046_/B vdd OAI22X1
XFILL_4__13320_ gnd vdd FILL
X_11257_ _11251_/Y _11768_/B _11256_/Y gnd _11257_/Y vdd AOI21X1
XSFILL79640x19050 gnd vdd FILL
XFILL_4__10532_ gnd vdd FILL
XFILL_2__9353_ gnd vdd FILL
XFILL_5__12871_ gnd vdd FILL
XFILL_2__11711_ gnd vdd FILL
XFILL_1__13140_ gnd vdd FILL
XFILL_0__13870_ gnd vdd FILL
XFILL_5__14610_ gnd vdd FILL
X_10208_ _13932_/A _7647_/CLK _9823_/R vdd _10134_/Y gnd vdd DFFSR
XFILL_5__11822_ gnd vdd FILL
XFILL_4__13251_ gnd vdd FILL
XFILL_5__15590_ gnd vdd FILL
X_11188_ _12192_/Y _11188_/B gnd _11189_/C vdd NAND2X1
XFILL_2__14430_ gnd vdd FILL
XFILL_2__9284_ gnd vdd FILL
XFILL_2__11642_ gnd vdd FILL
XFILL_5__8013_ gnd vdd FILL
XFILL_3__13981_ gnd vdd FILL
XFILL_1__10283_ gnd vdd FILL
XFILL_3_BUFX2_insert770 gnd vdd FILL
XFILL_5__14541_ gnd vdd FILL
XFILL_4__12202_ gnd vdd FILL
X_10139_ _10140_/B _8091_/B gnd _10139_/Y vdd NAND2X1
XFILL_3_BUFX2_insert781 gnd vdd FILL
XFILL_3__15720_ gnd vdd FILL
XSFILL39400x3050 gnd vdd FILL
XFILL_5__11753_ gnd vdd FILL
XFILL_2__8235_ gnd vdd FILL
X_15996_ _15170_/D _15996_/B _15995_/Y gnd _15998_/A vdd OAI21X1
XFILL_1__12022_ gnd vdd FILL
XFILL_3_BUFX2_insert792 gnd vdd FILL
XFILL_4__10394_ gnd vdd FILL
XFILL_2__14361_ gnd vdd FILL
XFILL_0__15540_ gnd vdd FILL
XFILL_2__11573_ gnd vdd FILL
XFILL_0__12752_ gnd vdd FILL
XSFILL114440x30050 gnd vdd FILL
XFILL_5__10704_ gnd vdd FILL
XFILL_0__7250_ gnd vdd FILL
XFILL_2__13312_ gnd vdd FILL
XFILL_5__14472_ gnd vdd FILL
XFILL_4__12133_ gnd vdd FILL
XFILL_2__16100_ gnd vdd FILL
X_14947_ _16448_/Q gnd _14947_/Y vdd INVX1
XFILL_3__15651_ gnd vdd FILL
XFILL_2__10524_ gnd vdd FILL
XFILL_5__11684_ gnd vdd FILL
XFILL_0__11703_ gnd vdd FILL
XSFILL84360x12050 gnd vdd FILL
XFILL_3__12863_ gnd vdd FILL
XFILL_2__14292_ gnd vdd FILL
XFILL_5__16211_ gnd vdd FILL
XFILL_0__15471_ gnd vdd FILL
XFILL_5__13423_ gnd vdd FILL
XFILL_2__7117_ gnd vdd FILL
XFILL_5__10635_ gnd vdd FILL
XFILL_0__7181_ gnd vdd FILL
XFILL_3__14602_ gnd vdd FILL
XFILL_2__16031_ gnd vdd FILL
XFILL_4__12064_ gnd vdd FILL
XSFILL59000x29050 gnd vdd FILL
XFILL_2__13243_ gnd vdd FILL
X_14878_ _7629_/A _13848_/C _14878_/C _10573_/A gnd _14879_/B vdd AOI22X1
XFILL_3__11814_ gnd vdd FILL
XFILL_2__8097_ gnd vdd FILL
XFILL_3__15582_ gnd vdd FILL
XFILL_0__14422_ gnd vdd FILL
XSFILL69160x73050 gnd vdd FILL
XSFILL103480x54050 gnd vdd FILL
XSFILL99400x34050 gnd vdd FILL
XFILL_0__11634_ gnd vdd FILL
XFILL_1__13973_ gnd vdd FILL
XFILL_5__8915_ gnd vdd FILL
XFILL_6__14713_ gnd vdd FILL
XFILL_5__16142_ gnd vdd FILL
XFILL_4__11015_ gnd vdd FILL
XFILL_5__13354_ gnd vdd FILL
X_13829_ _13828_/Y _14849_/B gnd _13830_/C vdd NOR2X1
XFILL_5__9895_ gnd vdd FILL
XFILL_3__14533_ gnd vdd FILL
XFILL_2__7048_ gnd vdd FILL
XFILL_5__10566_ gnd vdd FILL
XFILL_1__15712_ gnd vdd FILL
XFILL_2__13174_ gnd vdd FILL
XFILL111880x6050 gnd vdd FILL
XFILL_3__11745_ gnd vdd FILL
XFILL_3__7930_ gnd vdd FILL
XFILL_0__14353_ gnd vdd FILL
XFILL_2__10386_ gnd vdd FILL
XFILL_5__8846_ gnd vdd FILL
XFILL_5__12305_ gnd vdd FILL
XFILL_0__11565_ gnd vdd FILL
XFILL_4__15823_ gnd vdd FILL
XFILL_5__16073_ gnd vdd FILL
XSFILL104360x82050 gnd vdd FILL
XFILL_5__13285_ gnd vdd FILL
XFILL_2__12125_ gnd vdd FILL
XFILL_0__13304_ gnd vdd FILL
XFILL_5__10497_ gnd vdd FILL
XFILL_3__14464_ gnd vdd FILL
XFILL_1__15643_ gnd vdd FILL
XFILL_3__11676_ gnd vdd FILL
XFILL_3__7861_ gnd vdd FILL
XFILL_1__12855_ gnd vdd FILL
XFILL_0__10516_ gnd vdd FILL
XSFILL74280x64050 gnd vdd FILL
XFILL_5__15024_ gnd vdd FILL
XFILL_0__14284_ gnd vdd FILL
X_8430_ _8430_/Q _7406_/CLK _8430_/R vdd _8384_/Y gnd vdd DFFSR
XFILL_3__16203_ gnd vdd FILL
XFILL_5__12236_ gnd vdd FILL
XFILL_6__7570_ gnd vdd FILL
XFILL_0__11496_ gnd vdd FILL
XFILL_5_BUFX2_insert309 gnd vdd FILL
XFILL_5__8777_ gnd vdd FILL
XFILL_3__9600_ gnd vdd FILL
XFILL_3__13415_ gnd vdd FILL
XFILL_3__10627_ gnd vdd FILL
XFILL_4__15754_ gnd vdd FILL
XFILL_0__16023_ gnd vdd FILL
XFILL_2__12056_ gnd vdd FILL
XFILL_1__11806_ gnd vdd FILL
XFILL_4__12966_ gnd vdd FILL
XFILL_0__13235_ gnd vdd FILL
XFILL_3__14395_ gnd vdd FILL
XFILL_1__15574_ gnd vdd FILL
XFILL_1__12786_ gnd vdd FILL
XFILL_2__8999_ gnd vdd FILL
XFILL_0__10447_ gnd vdd FILL
XFILL_0_BUFX2_insert660 gnd vdd FILL
XFILL_5__7728_ gnd vdd FILL
XFILL_6__16314_ gnd vdd FILL
XFILL_6__13526_ gnd vdd FILL
XFILL_0_BUFX2_insert671 gnd vdd FILL
XFILL_4__14705_ gnd vdd FILL
XFILL_4__11917_ gnd vdd FILL
XFILL_5__12167_ gnd vdd FILL
X_8361_ _8423_/Q gnd _8361_/Y vdd INVX1
XFILL_2__11007_ gnd vdd FILL
XFILL_3__16134_ gnd vdd FILL
XFILL_3__9531_ gnd vdd FILL
XFILL_3__13346_ gnd vdd FILL
XFILL_3__10558_ gnd vdd FILL
XFILL_4__15685_ gnd vdd FILL
XFILL_1__14525_ gnd vdd FILL
XFILL_0_BUFX2_insert682 gnd vdd FILL
XFILL_4__12897_ gnd vdd FILL
XFILL_0_BUFX2_insert693 gnd vdd FILL
XFILL_1__11737_ gnd vdd FILL
XFILL_0__13166_ gnd vdd FILL
XFILL_0__10378_ gnd vdd FILL
XFILL_6__9240_ gnd vdd FILL
X_7312_ _7312_/A _7297_/B _7311_/Y gnd _7390_/D vdd OAI21X1
XFILL_5__11118_ gnd vdd FILL
XFILL_0__6965_ gnd vdd FILL
XFILL_4__14636_ gnd vdd FILL
XFILL_0__9753_ gnd vdd FILL
XSFILL28760x39050 gnd vdd FILL
XFILL_3__13277_ gnd vdd FILL
X_8292_ _8292_/Q _9050_/CLK _7258_/R vdd _8292_/D gnd vdd DFFSR
XFILL_5__12098_ gnd vdd FILL
XFILL_2__15815_ gnd vdd FILL
XFILL_3__16065_ gnd vdd FILL
XSFILL114520x10050 gnd vdd FILL
XFILL_4__11848_ gnd vdd FILL
XFILL_1__14456_ gnd vdd FILL
XFILL_3__9462_ gnd vdd FILL
XFILL_0__12117_ gnd vdd FILL
XFILL_3__10489_ gnd vdd FILL
XFILL_6__12408_ gnd vdd FILL
XFILL_1__11668_ gnd vdd FILL
XFILL_0__8704_ gnd vdd FILL
XFILL_6__16176_ gnd vdd FILL
XFILL_0__13097_ gnd vdd FILL
XSFILL33880x9050 gnd vdd FILL
XSFILL94440x77050 gnd vdd FILL
X_7243_ _7168_/A _7243_/B gnd _7244_/C vdd NAND2X1
XFILL_5__15926_ gnd vdd FILL
XFILL_6__13388_ gnd vdd FILL
XSFILL43800x42050 gnd vdd FILL
XFILL_0__9684_ gnd vdd FILL
XFILL_3__12228_ gnd vdd FILL
XFILL_3__15016_ gnd vdd FILL
XFILL_5__11049_ gnd vdd FILL
XFILL_4__14567_ gnd vdd FILL
XFILL_1__13407_ gnd vdd FILL
XFILL_0__6896_ gnd vdd FILL
XFILL_3__9393_ gnd vdd FILL
XFILL_2__15746_ gnd vdd FILL
XFILL_1__10619_ gnd vdd FILL
XFILL_4__11779_ gnd vdd FILL
XFILL_0__12048_ gnd vdd FILL
XFILL_1__14387_ gnd vdd FILL
XFILL_6__15127_ gnd vdd FILL
XFILL_2__12958_ gnd vdd FILL
XFILL_0__8635_ gnd vdd FILL
XFILL_4__16306_ gnd vdd FILL
XFILL_1__11599_ gnd vdd FILL
XFILL_4__13518_ gnd vdd FILL
XSFILL69240x53050 gnd vdd FILL
XFILL_3__12159_ gnd vdd FILL
XFILL_1__16126_ gnd vdd FILL
X_7174_ _7166_/B _7558_/B gnd _7175_/C vdd NAND2X1
XFILL_5__15857_ gnd vdd FILL
XFILL_1__13338_ gnd vdd FILL
XFILL_4__14498_ gnd vdd FILL
XFILL_2__11909_ gnd vdd FILL
XFILL_3__8344_ gnd vdd FILL
XFILL_2__15677_ gnd vdd FILL
XFILL_2__12889_ gnd vdd FILL
XFILL_4__16237_ gnd vdd FILL
XFILL_5__14808_ gnd vdd FILL
XFILL_0__8566_ gnd vdd FILL
XFILL_4__13449_ gnd vdd FILL
XFILL_5__15788_ gnd vdd FILL
XFILL_2__14628_ gnd vdd FILL
XFILL_0__15807_ gnd vdd FILL
XFILL_3__8275_ gnd vdd FILL
XFILL_1__16057_ gnd vdd FILL
XSFILL73720x78050 gnd vdd FILL
XFILL_1__13269_ gnd vdd FILL
XFILL_0__13999_ gnd vdd FILL
XFILL_5__14739_ gnd vdd FILL
XFILL_3__15918_ gnd vdd FILL
XFILL_4__16168_ gnd vdd FILL
XFILL_1__15008_ gnd vdd FILL
XFILL_3__7226_ gnd vdd FILL
XFILL_0__8497_ gnd vdd FILL
XFILL_1__7290_ gnd vdd FILL
XSFILL8680x60050 gnd vdd FILL
XFILL_2__14559_ gnd vdd FILL
XFILL_0__15738_ gnd vdd FILL
XFILL_0__7448_ gnd vdd FILL
XFILL_4__15119_ gnd vdd FILL
XFILL_4__16099_ gnd vdd FILL
XFILL_3__15849_ gnd vdd FILL
XSFILL89400x66050 gnd vdd FILL
XFILL_0__15669_ gnd vdd FILL
XFILL_5__16409_ gnd vdd FILL
X_9815_ _9815_/Q _8679_/CLK _9959_/R vdd _9815_/D gnd vdd DFFSR
XFILL_0__7379_ gnd vdd FILL
XFILL_2__16229_ gnd vdd FILL
XFILL_3__7088_ gnd vdd FILL
XFILL_4__7970_ gnd vdd FILL
XFILL_0__9118_ gnd vdd FILL
XSFILL28840x19050 gnd vdd FILL
X_9746_ _9798_/B _7314_/B gnd _9747_/C vdd NAND2X1
X_6958_ _6956_/Y _6948_/A _6958_/C gnd _7016_/D vdd OAI21X1
XFILL_4__6921_ gnd vdd FILL
XSFILL13640x61050 gnd vdd FILL
XSFILL94520x57050 gnd vdd FILL
XFILL_1__9931_ gnd vdd FILL
X_9677_ _9677_/A gnd _9677_/Y vdd INVX1
XFILL_4__9640_ gnd vdd FILL
X_6889_ _6889_/A gnd memoryWriteData[19] vdd BUFX2
XFILL_4__6852_ gnd vdd FILL
X_8628_ _8626_/Y _8657_/A _8628_/C gnd _8682_/D vdd OAI21X1
XFILL_1__9862_ gnd vdd FILL
XFILL_5_BUFX2_insert810 gnd vdd FILL
XFILL_5_BUFX2_insert821 gnd vdd FILL
XFILL_5_BUFX2_insert832 gnd vdd FILL
XFILL_5_BUFX2_insert843 gnd vdd FILL
X_10490_ _10539_/B _9978_/B gnd _10491_/C vdd NAND2X1
XFILL_5_BUFX2_insert854 gnd vdd FILL
XSFILL73800x58050 gnd vdd FILL
X_8559_ _8559_/Q _7651_/CLK _9711_/R vdd _8559_/D gnd vdd DFFSR
XFILL_6__7699_ gnd vdd FILL
XFILL_3__9729_ gnd vdd FILL
XFILL_4__8522_ gnd vdd FILL
XFILL_1__9793_ gnd vdd FILL
XFILL_5_BUFX2_insert865 gnd vdd FILL
XFILL_5_BUFX2_insert876 gnd vdd FILL
XBUFX2_insert1040 _13297_/Y gnd _7753_/B vdd BUFX2
XFILL_5_BUFX2_insert887 gnd vdd FILL
XSFILL8760x40050 gnd vdd FILL
XBUFX2_insert1051 _12806_/Q gnd _12313_/D vdd BUFX2
XSFILL33800x74050 gnd vdd FILL
XBUFX2_insert1062 _14992_/Y gnd _15322_/A vdd BUFX2
XFILL_5_BUFX2_insert898 gnd vdd FILL
XFILL_1__8744_ gnd vdd FILL
XBUFX2_insert1073 _13327_/Y gnd _8823_/B vdd BUFX2
XBUFX2_insert1084 rst gnd BUFX2_insert570/A vdd BUFX2
XFILL_4__8453_ gnd vdd FILL
X_12160_ _13190_/Q gnd _12162_/A vdd INVX1
XFILL_6__9369_ gnd vdd FILL
X_11111_ _12180_/Y _12302_/Y gnd _11111_/Y vdd NOR2X1
XFILL_4__8384_ gnd vdd FILL
XSFILL8840x3050 gnd vdd FILL
X_12091_ _11987_/A _12091_/B _12011_/C gnd _12094_/A vdd NAND3X1
XFILL_1__7626_ gnd vdd FILL
XSFILL54200x5050 gnd vdd FILL
XFILL_4__7335_ gnd vdd FILL
X_11042_ _12278_/Y _12162_/Y gnd _11044_/A vdd XOR2X1
XFILL_1__7557_ gnd vdd FILL
X_15850_ _15843_/Y _15850_/B gnd _15850_/Y vdd NAND2X1
XFILL_1__7488_ gnd vdd FILL
XFILL_4__9005_ gnd vdd FILL
XFILL_2_BUFX2_insert700 gnd vdd FILL
XSFILL39160x52050 gnd vdd FILL
XFILL_2_BUFX2_insert711 gnd vdd FILL
X_14801_ _14801_/A _14801_/B _14800_/Y gnd _14812_/A vdd NAND3X1
XFILL_2_BUFX2_insert722 gnd vdd FILL
XFILL_4__7197_ gnd vdd FILL
XFILL_2__8020_ gnd vdd FILL
XFILL_1__9227_ gnd vdd FILL
X_15781_ _8620_/A gnd _15781_/Y vdd INVX1
XFILL_2_BUFX2_insert733 gnd vdd FILL
X_12993_ _6884_/A gnd _12993_/Y vdd INVX1
XFILL_2_BUFX2_insert744 gnd vdd FILL
XFILL_2_BUFX2_insert755 gnd vdd FILL
XFILL_2_BUFX2_insert766 gnd vdd FILL
XFILL_2_BUFX2_insert777 gnd vdd FILL
X_14732_ _14732_/A gnd _14733_/D vdd INVX1
XSFILL84280x27050 gnd vdd FILL
X_11944_ _13194_/Q gnd _11946_/A vdd INVX1
XFILL_1__9158_ gnd vdd FILL
XFILL_2_BUFX2_insert788 gnd vdd FILL
XFILL_2_BUFX2_insert799 gnd vdd FILL
XFILL_1__8109_ gnd vdd FILL
XFILL_5__6961_ gnd vdd FILL
XFILL_5__10420_ gnd vdd FILL
X_11875_ _12808_/Q gnd _11877_/A vdd INVX1
XSFILL99320x49050 gnd vdd FILL
X_14663_ _8815_/Q gnd _14665_/B vdd INVX1
XFILL_1__9089_ gnd vdd FILL
XFILL_2__10240_ gnd vdd FILL
XFILL_4__9907_ gnd vdd FILL
XFILL_5__8700_ gnd vdd FILL
XSFILL34520x20050 gnd vdd FILL
XFILL_1__10970_ gnd vdd FILL
X_16402_ _14776_/A gnd _16402_/Y vdd INVX1
X_13614_ _13613_/Y _14865_/B _13614_/C _13612_/Y gnd _13618_/B vdd OAI22X1
X_10826_ _14793_/C gnd _10826_/Y vdd INVX1
XFILL_5__9680_ gnd vdd FILL
XFILL_5__6892_ gnd vdd FILL
XFILL_3__11530_ gnd vdd FILL
X_14594_ _14594_/A _14594_/B gnd _14595_/A vdd NOR2X1
XFILL_2__10171_ gnd vdd FILL
XBUFX2_insert710 _12816_/Q gnd _15064_/A vdd BUFX2
XFILL_5__8631_ gnd vdd FILL
XFILL_0__11350_ gnd vdd FILL
X_16333_ _15246_/A gnd _16335_/A vdd INVX1
XBUFX2_insert721 _13352_/Y gnd _10140_/B vdd BUFX2
XBUFX2_insert732 _12411_/Y gnd _8889_/B vdd BUFX2
X_10757_ _15268_/A gnd _10759_/A vdd INVX1
X_13545_ _8572_/A gnd _15141_/D vdd INVX1
XBUFX2_insert743 _15055_/Y gnd _15595_/B vdd BUFX2
XFILL_5__10282_ gnd vdd FILL
XFILL_3__11461_ gnd vdd FILL
XFILL_1__12640_ gnd vdd FILL
XFILL_0__10301_ gnd vdd FILL
XFILL_2__8853_ gnd vdd FILL
XBUFX2_insert754 _13344_/Y gnd _9770_/A vdd BUFX2
XBUFX2_insert765 _12393_/Y gnd _7079_/B vdd BUFX2
XSFILL43880x4050 gnd vdd FILL
XFILL_0__11281_ gnd vdd FILL
XFILL_5__12021_ gnd vdd FILL
XFILL_6__14360_ gnd vdd FILL
XFILL_4__9769_ gnd vdd FILL
XBUFX2_insert776 _13301_/Y gnd _7824_/B vdd BUFX2
X_13476_ _13476_/A _13476_/B _15338_/C gnd _12952_/A vdd AOI21X1
XFILL_3__10412_ gnd vdd FILL
XSFILL13800x21050 gnd vdd FILL
X_16264_ _16264_/A _15848_/A gnd _16264_/Y vdd NOR2X1
XFILL_4__12751_ gnd vdd FILL
X_10688_ _10688_/A _10661_/B _10688_/C gnd _10688_/Y vdd OAI21X1
XFILL_3__14180_ gnd vdd FILL
XBUFX2_insert787 _13486_/Y gnd _14037_/C vdd BUFX2
XFILL_2__7804_ gnd vdd FILL
XFILL_0__13020_ gnd vdd FILL
XFILL_0__10232_ gnd vdd FILL
XBUFX2_insert798 _13334_/Y gnd _9372_/B vdd BUFX2
XFILL_3__11392_ gnd vdd FILL
XFILL_2__13930_ gnd vdd FILL
XFILL_6__13311_ gnd vdd FILL
XFILL112120x73050 gnd vdd FILL
XFILL_1__12571_ gnd vdd FILL
XFILL_2__8784_ gnd vdd FILL
X_15215_ _15215_/A _15215_/B _15215_/C gnd _15219_/C vdd NOR3X1
X_12427_ _12427_/A gnd _12427_/Y vdd INVX1
XFILL_3__13131_ gnd vdd FILL
XFILL_5__8493_ gnd vdd FILL
XFILL_4__11702_ gnd vdd FILL
X_16195_ _16195_/A _16194_/Y gnd _16201_/A vdd NOR2X1
XFILL_1__14310_ gnd vdd FILL
XFILL_4__15470_ gnd vdd FILL
XFILL_2__7735_ gnd vdd FILL
XFILL_1__11522_ gnd vdd FILL
XFILL_2__13861_ gnd vdd FILL
XFILL_0__10163_ gnd vdd FILL
XFILL_1__15290_ gnd vdd FILL
XFILL_5__7444_ gnd vdd FILL
X_12358_ _12454_/A gnd _12358_/Y vdd INVX1
XFILL_4__14421_ gnd vdd FILL
X_15146_ _7292_/A _15114_/B _15114_/C gnd _15147_/C vdd NAND3X1
XSFILL114440x25050 gnd vdd FILL
XFILL_1_CLKBUF1_insert170 gnd vdd FILL
XFILL_4__11633_ gnd vdd FILL
XFILL_2__15600_ gnd vdd FILL
XFILL_5__13972_ gnd vdd FILL
XFILL_1_CLKBUF1_insert181 gnd vdd FILL
XFILL_1__14241_ gnd vdd FILL
XFILL_3__10274_ gnd vdd FILL
XFILL_1_CLKBUF1_insert192 gnd vdd FILL
XFILL_2__13792_ gnd vdd FILL
XSFILL43720x57050 gnd vdd FILL
XFILL_1__11453_ gnd vdd FILL
XFILL_0__14971_ gnd vdd FILL
X_11309_ _11550_/C gnd _11533_/A vdd INVX1
XFILL_5__15711_ gnd vdd FILL
XFILL_5__7375_ gnd vdd FILL
XFILL_3__12013_ gnd vdd FILL
X_15077_ _15077_/A _15077_/B _15338_/C gnd _12824_/A vdd AOI21X1
XFILL_2__9405_ gnd vdd FILL
XFILL_2_BUFX2_insert2 gnd vdd FILL
XFILL_4__14352_ gnd vdd FILL
X_12289_ _6888_/A _12289_/B _12289_/C _12308_/B gnd _12289_/Y vdd AOI22X1
XSFILL89240x3050 gnd vdd FILL
XFILL_2__12743_ gnd vdd FILL
XFILL_1__10404_ gnd vdd FILL
XFILL_2__15531_ gnd vdd FILL
XFILL_4__11564_ gnd vdd FILL
XFILL_1__14172_ gnd vdd FILL
XFILL_5__9114_ gnd vdd FILL
XFILL_2__7597_ gnd vdd FILL
XFILL_0__13922_ gnd vdd FILL
X_14028_ _10082_/Q gnd _14030_/D vdd INVX1
XSFILL99400x29050 gnd vdd FILL
XFILL_1__11384_ gnd vdd FILL
XFILL_4__13303_ gnd vdd FILL
XFILL_5__15642_ gnd vdd FILL
XFILL_5__12854_ gnd vdd FILL
XFILL_4__10515_ gnd vdd FILL
XFILL_2__9336_ gnd vdd FILL
XFILL_1__13123_ gnd vdd FILL
XFILL_4__14283_ gnd vdd FILL
XFILL_4__11495_ gnd vdd FILL
XFILL_2__15462_ gnd vdd FILL
XFILL_0__13853_ gnd vdd FILL
XFILL_5__9045_ gnd vdd FILL
XFILL_4__16022_ gnd vdd FILL
XFILL_6__12055_ gnd vdd FILL
XFILL_0__8351_ gnd vdd FILL
XFILL_5__11805_ gnd vdd FILL
XFILL_4__13234_ gnd vdd FILL
XFILL_5__15573_ gnd vdd FILL
XFILL_5__12785_ gnd vdd FILL
XFILL_4__10446_ gnd vdd FILL
XFILL_3__8060_ gnd vdd FILL
XFILL_2__11625_ gnd vdd FILL
XFILL_2__14413_ gnd vdd FILL
XFILL_2__15393_ gnd vdd FILL
XFILL_2__9267_ gnd vdd FILL
XFILL_3__13964_ gnd vdd FILL
XFILL_1__10266_ gnd vdd FILL
XFILL_6__11006_ gnd vdd FILL
XFILL_0__7302_ gnd vdd FILL
XFILL_0__13784_ gnd vdd FILL
XFILL_5__14524_ gnd vdd FILL
XFILL_3__15703_ gnd vdd FILL
XSFILL74280x59050 gnd vdd FILL
XFILL_0__10996_ gnd vdd FILL
XFILL_5__11736_ gnd vdd FILL
X_7930_ _7931_/B _9082_/B gnd _7930_/Y vdd NAND2X1
X_15979_ _9837_/Q gnd _15979_/Y vdd INVX1
XFILL_4__10377_ gnd vdd FILL
XFILL_4__13165_ gnd vdd FILL
XFILL_1__12005_ gnd vdd FILL
XFILL_2__8218_ gnd vdd FILL
XFILL_2__14344_ gnd vdd FILL
XFILL_3__12915_ gnd vdd FILL
XSFILL109400x14050 gnd vdd FILL
XFILL_0__15523_ gnd vdd FILL
XFILL_2__11556_ gnd vdd FILL
XFILL_0__12735_ gnd vdd FILL
XFILL_3__13895_ gnd vdd FILL
XFILL_1__10197_ gnd vdd FILL
XFILL_0__7233_ gnd vdd FILL
XFILL_5__14455_ gnd vdd FILL
XFILL_4__12116_ gnd vdd FILL
X_7861_ _7915_/Q gnd _7861_/Y vdd INVX1
XFILL_2__10507_ gnd vdd FILL
XFILL112200x53050 gnd vdd FILL
XFILL_3__15634_ gnd vdd FILL
XFILL_2__8149_ gnd vdd FILL
XFILL_5__11667_ gnd vdd FILL
XFILL_3__12846_ gnd vdd FILL
XFILL_4__13096_ gnd vdd FILL
XFILL_2__14275_ gnd vdd FILL
XFILL_2__11487_ gnd vdd FILL
XFILL_0__15454_ gnd vdd FILL
X_9600_ _9639_/A _9600_/B gnd _9600_/Y vdd NAND2X1
XFILL_5__13406_ gnd vdd FILL
XFILL_5__10618_ gnd vdd FILL
XFILL_0__7164_ gnd vdd FILL
XFILL_2__13226_ gnd vdd FILL
XFILL_2__16014_ gnd vdd FILL
XFILL_4__12047_ gnd vdd FILL
XFILL_5__14386_ gnd vdd FILL
XFILL_2__10438_ gnd vdd FILL
XFILL_3__15565_ gnd vdd FILL
XFILL_6_BUFX2_insert60 gnd vdd FILL
XFILL_0__14405_ gnd vdd FILL
X_7792_ _7748_/A _7664_/CLK _7920_/R vdd _7750_/Y gnd vdd DFFSR
XFILL_5__11598_ gnd vdd FILL
XFILL_3__12777_ gnd vdd FILL
XFILL_3__8962_ gnd vdd FILL
XFILL_1__13956_ gnd vdd FILL
XFILL_0__11617_ gnd vdd FILL
XFILL_0__15385_ gnd vdd FILL
XFILL_5__16125_ gnd vdd FILL
XFILL_5__13337_ gnd vdd FILL
X_9531_ _9581_/Q gnd _9533_/A vdd INVX1
XFILL_0__12597_ gnd vdd FILL
XFILL_5__9878_ gnd vdd FILL
XFILL_5__10549_ gnd vdd FILL
XFILL_0__7095_ gnd vdd FILL
XFILL_3__14516_ gnd vdd FILL
XFILL_2__13157_ gnd vdd FILL
XFILL_1__12907_ gnd vdd FILL
XFILL_3__11728_ gnd vdd FILL
XFILL_2__10369_ gnd vdd FILL
XFILL_0__14336_ gnd vdd FILL
XSFILL49000x6050 gnd vdd FILL
XFILL_3__15496_ gnd vdd FILL
XSFILL53960x81050 gnd vdd FILL
XFILL_1__13887_ gnd vdd FILL
XFILL_3__8893_ gnd vdd FILL
XFILL_5__8829_ gnd vdd FILL
XFILL_0__11548_ gnd vdd FILL
XFILL_4__15806_ gnd vdd FILL
XFILL_5__16056_ gnd vdd FILL
XFILL_5__13268_ gnd vdd FILL
X_9462_ _9558_/Q gnd _9464_/A vdd INVX1
XFILL_5_BUFX2_insert106 gnd vdd FILL
XFILL_2__12108_ gnd vdd FILL
XSFILL69240x48050 gnd vdd FILL
XSFILL103560x29050 gnd vdd FILL
XFILL_3__14447_ gnd vdd FILL
XFILL_3__7844_ gnd vdd FILL
XFILL_2__13088_ gnd vdd FILL
XFILL_1__15626_ gnd vdd FILL
XFILL_4__13998_ gnd vdd FILL
XFILL_3__11659_ gnd vdd FILL
XFILL_1__12838_ gnd vdd FILL
XFILL_5__15007_ gnd vdd FILL
XFILL_0__14267_ gnd vdd FILL
X_8413_ _8413_/Q _7915_/CLK _7915_/R vdd _8333_/Y gnd vdd DFFSR
XFILL_0__11479_ gnd vdd FILL
XFILL_5__12219_ gnd vdd FILL
XFILL_4__15737_ gnd vdd FILL
XFILL_0__16006_ gnd vdd FILL
XFILL_2__12039_ gnd vdd FILL
X_9393_ _9393_/A _9401_/A _9393_/C gnd _9449_/D vdd OAI21X1
XFILL_0__13218_ gnd vdd FILL
XFILL_1__15557_ gnd vdd FILL
XFILL_3__14378_ gnd vdd FILL
XFILL_1__12769_ gnd vdd FILL
XFILL_0_BUFX2_insert490 gnd vdd FILL
XFILL_0__9805_ gnd vdd FILL
XFILL_0__14198_ gnd vdd FILL
XSFILL104440x57050 gnd vdd FILL
XFILL_3__16117_ gnd vdd FILL
X_8344_ _8345_/B _8600_/B gnd _8344_/Y vdd NAND2X1
XFILL_3__13329_ gnd vdd FILL
XFILL_4__15668_ gnd vdd FILL
XFILL_1__14508_ gnd vdd FILL
XFILL_4_BUFX2_insert806 gnd vdd FILL
XFILL_3__9514_ gnd vdd FILL
XFILL_0__7997_ gnd vdd FILL
XSFILL8680x55050 gnd vdd FILL
XFILL_4_BUFX2_insert817 gnd vdd FILL
XFILL_4_BUFX2_insert828 gnd vdd FILL
XFILL_0__13149_ gnd vdd FILL
XFILL_1__15488_ gnd vdd FILL
XFILL_4_BUFX2_insert839 gnd vdd FILL
XFILL_4__14619_ gnd vdd FILL
XFILL_0__9736_ gnd vdd FILL
XFILL_0__6948_ gnd vdd FILL
X_8275_ _8275_/A gnd _8275_/Y vdd INVX1
XFILL_3__16048_ gnd vdd FILL
XFILL_4__15599_ gnd vdd FILL
XFILL_1__14439_ gnd vdd FILL
XFILL_5__15909_ gnd vdd FILL
XFILL_1__8460_ gnd vdd FILL
X_7226_ _7226_/A _7202_/B _7225_/Y gnd _7226_/Y vdd OAI21X1
XFILL_0__9667_ gnd vdd FILL
XFILL_0__6879_ gnd vdd FILL
XFILL_2__15729_ gnd vdd FILL
XFILL_3__9376_ gnd vdd FILL
XFILL_6__9085_ gnd vdd FILL
XFILL_0__8618_ gnd vdd FILL
X_7157_ _7157_/Q _9958_/CLK _8053_/R vdd _7125_/Y gnd vdd DFFSR
XFILL_4__7120_ gnd vdd FILL
XFILL_1__8391_ gnd vdd FILL
XFILL_1__16109_ gnd vdd FILL
XFILL_0__9598_ gnd vdd FILL
XFILL_3__8327_ gnd vdd FILL
XSFILL13640x56050 gnd vdd FILL
XCLKBUF1_insert180 CLKBUF1_insert216/A gnd _7781_/CLK vdd CLKBUF1
XFILL_1__7342_ gnd vdd FILL
XCLKBUF1_insert191 CLKBUF1_insert218/A gnd _9195_/CLK vdd CLKBUF1
XSFILL28440x16050 gnd vdd FILL
XFILL_4__7051_ gnd vdd FILL
X_7088_ _7124_/A _8496_/B gnd _7089_/C vdd NAND2X1
XFILL_3__8258_ gnd vdd FILL
XSFILL39080x67050 gnd vdd FILL
XFILL_3__7209_ gnd vdd FILL
XFILL_3__8189_ gnd vdd FILL
XFILL_1__9012_ gnd vdd FILL
XFILL_5_BUFX2_insert6 gnd vdd FILL
XFILL_1_BUFX2_insert707 gnd vdd FILL
XFILL_1_BUFX2_insert718 gnd vdd FILL
XFILL_1_BUFX2_insert729 gnd vdd FILL
XSFILL33800x69050 gnd vdd FILL
XSFILL8760x35050 gnd vdd FILL
XFILL_4__7953_ gnd vdd FILL
X_11660_ _11660_/A _11660_/B _11658_/Y gnd _11660_/Y vdd NAND3X1
X_9729_ _9727_/Y _9764_/A _9729_/C gnd _9817_/D vdd OAI21X1
XFILL_4__6904_ gnd vdd FILL
X_10611_ _10573_/A _8051_/CLK _7789_/R vdd _10575_/Y gnd vdd DFFSR
XFILL_4__7884_ gnd vdd FILL
XFILL_1__9914_ gnd vdd FILL
X_11591_ _11591_/A _11621_/C _11591_/C _11484_/B gnd _11592_/A vdd OAI22X1
XFILL_4__9623_ gnd vdd FILL
X_13330_ _13259_/C gnd _13337_/B vdd INVX2
X_10542_ _10540_/Y _10505_/A _10542_/C gnd _10600_/D vdd OAI21X1
XFILL_5_BUFX2_insert640 gnd vdd FILL
XFILL_5_BUFX2_insert651 gnd vdd FILL
XFILL_4__9554_ gnd vdd FILL
X_13261_ _13289_/B _13337_/A gnd _13262_/B vdd NOR2X1
XFILL_5_BUFX2_insert662 gnd vdd FILL
XFILL_5_BUFX2_insert673 gnd vdd FILL
X_10473_ _15822_/B _9705_/CLK _7914_/R vdd _10473_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert684 gnd vdd FILL
XFILL_5_BUFX2_insert695 gnd vdd FILL
XFILL_4__8505_ gnd vdd FILL
XFILL_1__9776_ gnd vdd FILL
XFILL_1__6988_ gnd vdd FILL
X_15000_ _15000_/A _14982_/Y _15024_/C gnd _15000_/Y vdd NAND3X1
X_12212_ _12227_/A gnd _12307_/C gnd _12218_/A vdd NAND3X1
XFILL_4__9485_ gnd vdd FILL
X_13192_ _13192_/Q _13180_/CLK _13180_/R vdd _13132_/Y gnd vdd DFFSR
XFILL_1__8727_ gnd vdd FILL
X_12143_ _12122_/A _12928_/Q gnd _12143_/Y vdd NAND2X1
XFILL_2__7451_ gnd vdd FILL
XSFILL104600x17050 gnd vdd FILL
XFILL_1__8658_ gnd vdd FILL
XFILL_2_CLKBUF1_insert210 gnd vdd FILL
XFILL_5__7160_ gnd vdd FILL
XFILL_4__8367_ gnd vdd FILL
XFILL_2_CLKBUF1_insert221 gnd vdd FILL
XSFILL13640x2050 gnd vdd FILL
X_12074_ _12074_/A _12072_/Y _12073_/Y gnd _13143_/B vdd NAND3X1
XFILL_6__10170_ gnd vdd FILL
XFILL_1__7609_ gnd vdd FILL
XFILL_1__8589_ gnd vdd FILL
XFILL_4__7318_ gnd vdd FILL
X_15902_ _15892_/Y _15902_/B _15902_/C gnd _15910_/B vdd NAND3X1
XFILL_5__7091_ gnd vdd FILL
X_11025_ _11025_/A _12129_/Y gnd _11025_/Y vdd NOR2X1
XFILL_4__10300_ gnd vdd FILL
XFILL_2__9121_ gnd vdd FILL
XFILL_4__11280_ gnd vdd FILL
XFILL_1__10120_ gnd vdd FILL
XFILL_4__7249_ gnd vdd FILL
XFILL_4__10231_ gnd vdd FILL
X_15833_ _15829_/Y _15833_/B gnd _15833_/Y vdd NOR2X1
XFILL_5__12570_ gnd vdd FILL
XFILL_2__11410_ gnd vdd FILL
XFILL_2_BUFX2_insert530 gnd vdd FILL
XFILL_3__10961_ gnd vdd FILL
XFILL_2__12390_ gnd vdd FILL
XFILL_1__10051_ gnd vdd FILL
XFILL_2_BUFX2_insert541 gnd vdd FILL
XSFILL108840x22050 gnd vdd FILL
XFILL_0_BUFX2_insert1009 gnd vdd FILL
XFILL_2_BUFX2_insert552 gnd vdd FILL
XFILL_5__11521_ gnd vdd FILL
XFILL_2__8003_ gnd vdd FILL
XFILL_0__10781_ gnd vdd FILL
XFILL_2_BUFX2_insert563 gnd vdd FILL
XFILL_3__12700_ gnd vdd FILL
X_15764_ _9385_/A _15794_/B _15764_/C gnd _15765_/C vdd NAND3X1
XFILL_4__10162_ gnd vdd FILL
X_12976_ vdd _12976_/B gnd _12977_/C vdd NAND2X1
XSFILL59000x1050 gnd vdd FILL
XFILL_2_BUFX2_insert574 gnd vdd FILL
XFILL_2__11341_ gnd vdd FILL
XFILL_3__13680_ gnd vdd FILL
XFILL_0__12520_ gnd vdd FILL
XFILL_3__10892_ gnd vdd FILL
XFILL_2_BUFX2_insert585 gnd vdd FILL
XFILL_5__9801_ gnd vdd FILL
XFILL_2_BUFX2_insert596 gnd vdd FILL
XFILL112120x68050 gnd vdd FILL
XFILL_5__14240_ gnd vdd FILL
X_14715_ _14715_/A _14702_/Y gnd _14742_/A vdd NOR2X1
XFILL_5__7993_ gnd vdd FILL
X_11927_ _11900_/A _12382_/A gnd _11928_/C vdd NAND2X1
XFILL_5__11452_ gnd vdd FILL
XSFILL38760x20050 gnd vdd FILL
XFILL_3__12631_ gnd vdd FILL
XFILL_1__13810_ gnd vdd FILL
X_15695_ _15652_/A _9574_/Q _10214_/Q _15695_/D gnd _15697_/A vdd AOI22X1
XFILL_2__14060_ gnd vdd FILL
XFILL_4__14970_ gnd vdd FILL
XSFILL64040x53050 gnd vdd FILL
XFILL_2__11272_ gnd vdd FILL
XSFILL94360x50 gnd vdd FILL
XFILL_5__9732_ gnd vdd FILL
XFILL_0__12451_ gnd vdd FILL
XFILL_1__14790_ gnd vdd FILL
XFILL_5__10403_ gnd vdd FILL
XFILL_5__6944_ gnd vdd FILL
X_14646_ _14645_/Y _14646_/B gnd _14647_/B vdd NOR2X1
XFILL_5__14171_ gnd vdd FILL
XFILL_4__13921_ gnd vdd FILL
XFILL_2__13011_ gnd vdd FILL
XFILL_3__15350_ gnd vdd FILL
XFILL_5__11383_ gnd vdd FILL
X_11858_ _11855_/Y _12089_/A _11857_/Y gnd _11858_/Y vdd NOR3X1
XFILL_1__13741_ gnd vdd FILL
XFILL_0__11402_ gnd vdd FILL
XFILL_1__10953_ gnd vdd FILL
XFILL_0__15170_ gnd vdd FILL
XFILL_6_BUFX2_insert1093 gnd vdd FILL
XFILL_5__9663_ gnd vdd FILL
XFILL_5__13122_ gnd vdd FILL
XFILL_0__12382_ gnd vdd FILL
X_10809_ _10809_/A _9785_/B gnd _10810_/C vdd NAND2X1
XFILL_3__14301_ gnd vdd FILL
XFILL_5__6875_ gnd vdd FILL
X_14577_ _7149_/Q gnd _14577_/Y vdd INVX1
XFILL_4__13852_ gnd vdd FILL
XFILL_2__8905_ gnd vdd FILL
XFILL_3__11513_ gnd vdd FILL
XSFILL43880x11050 gnd vdd FILL
X_11789_ _11034_/B _11789_/B gnd _11790_/C vdd NOR2X1
XFILL_3__12493_ gnd vdd FILL
XFILL_2__10154_ gnd vdd FILL
XFILL_0__14121_ gnd vdd FILL
XFILL_3__15281_ gnd vdd FILL
XFILL_5__8614_ gnd vdd FILL
XFILL_1__13672_ gnd vdd FILL
XFILL_2__9885_ gnd vdd FILL
XBUFX2_insert540 BUFX2_insert494/A gnd _7793_/R vdd BUFX2
XFILL_0__11333_ gnd vdd FILL
XFILL_1__10884_ gnd vdd FILL
X_16316_ _16316_/A _15792_/B _15726_/A _14959_/D gnd _16316_/Y vdd OAI22X1
XBUFX2_insert551 BUFX2_insert524/A gnd _7896_/R vdd BUFX2
XBUFX2_insert562 BUFX2_insert607/A gnd _8156_/R vdd BUFX2
X_13528_ _13528_/A _14389_/B _13751_/B _9815_/Q gnd _13528_/Y vdd AOI22X1
XFILL_5__9594_ gnd vdd FILL
XFILL_3__14232_ gnd vdd FILL
XFILL_1__15411_ gnd vdd FILL
XBUFX2_insert573 BUFX2_insert556/A gnd _8929_/R vdd BUFX2
XFILL_5__10265_ gnd vdd FILL
XFILL_3__11444_ gnd vdd FILL
XFILL_1__12623_ gnd vdd FILL
XFILL_4__13783_ gnd vdd FILL
XFILL_2__8836_ gnd vdd FILL
XBUFX2_insert584 BUFX2_insert607/A gnd _9430_/R vdd BUFX2
XFILL_0__14052_ gnd vdd FILL
XFILL_1__16391_ gnd vdd FILL
XFILL_2__14962_ gnd vdd FILL
XFILL_4__10995_ gnd vdd FILL
XBUFX2_insert595 BUFX2_insert559/A gnd _8670_/R vdd BUFX2
XSFILL84200x66050 gnd vdd FILL
XFILL_5__12004_ gnd vdd FILL
XFILL_0__11264_ gnd vdd FILL
XFILL_4__15522_ gnd vdd FILL
X_16247_ _16247_/A _15622_/A _16247_/C _16246_/Y gnd _16247_/Y vdd OAI22X1
XFILL_4__12734_ gnd vdd FILL
X_13459_ _13423_/A _13407_/Y _13465_/C gnd _13459_/Y vdd NAND3X1
XFILL_0__7851_ gnd vdd FILL
XFILL_1__15342_ gnd vdd FILL
XFILL_3__14163_ gnd vdd FILL
XFILL_5__10196_ gnd vdd FILL
XFILL_0__13003_ gnd vdd FILL
XFILL_2__13913_ gnd vdd FILL
XFILL_3__11375_ gnd vdd FILL
XFILL_2__8767_ gnd vdd FILL
XFILL_3__7560_ gnd vdd FILL
XFILL_0__11195_ gnd vdd FILL
XFILL_2__14893_ gnd vdd FILL
XFILL_5__8476_ gnd vdd FILL
XSFILL59000x42050 gnd vdd FILL
XSFILL23640x19050 gnd vdd FILL
X_16178_ _16178_/A _16178_/B _16178_/C gnd _16179_/A vdd NAND3X1
XFILL_3__13114_ gnd vdd FILL
XFILL_4__15453_ gnd vdd FILL
XFILL_2__7718_ gnd vdd FILL
XFILL_1__11505_ gnd vdd FILL
XFILL_3__14094_ gnd vdd FILL
XFILL_2__13844_ gnd vdd FILL
XFILL_0__10146_ gnd vdd FILL
XFILL_3__7491_ gnd vdd FILL
XFILL_1__15273_ gnd vdd FILL
XFILL_5__7427_ gnd vdd FILL
XFILL_1__12485_ gnd vdd FILL
XFILL_2__8698_ gnd vdd FILL
XFILL_0__9521_ gnd vdd FILL
X_15129_ _8700_/A _15821_/B _15969_/C _7768_/Q gnd _15136_/A vdd AOI22X1
XFILL_4__14404_ gnd vdd FILL
XFILL_3__13045_ gnd vdd FILL
XFILL_4__11616_ gnd vdd FILL
X_8060_ _8152_/Q gnd _8062_/A vdd INVX1
XFILL_5__13955_ gnd vdd FILL
XFILL_3__9230_ gnd vdd FILL
XFILL_4__15384_ gnd vdd FILL
XFILL_1__14224_ gnd vdd FILL
XFILL112200x48050 gnd vdd FILL
XFILL_3__10257_ gnd vdd FILL
XFILL_4__12596_ gnd vdd FILL
XFILL_1__11436_ gnd vdd FILL
XFILL_2__13775_ gnd vdd FILL
XFILL_0__14954_ gnd vdd FILL
XFILL_5__7358_ gnd vdd FILL
XFILL_6__13156_ gnd vdd FILL
X_7011_ _7011_/Q _6999_/CLK _7011_/R vdd _7011_/D gnd vdd DFFSR
XFILL_4__14335_ gnd vdd FILL
XSFILL64120x33050 gnd vdd FILL
XFILL_5__12906_ gnd vdd FILL
XFILL_5__13886_ gnd vdd FILL
XFILL_2__15514_ gnd vdd FILL
XFILL_4__11547_ gnd vdd FILL
XFILL_2__12726_ gnd vdd FILL
XFILL_3__10188_ gnd vdd FILL
XFILL_1__14155_ gnd vdd FILL
XFILL_0__13905_ gnd vdd FILL
XFILL_3__9161_ gnd vdd FILL
XFILL_1__11367_ gnd vdd FILL
XFILL_0__8403_ gnd vdd FILL
XFILL_0__14885_ gnd vdd FILL
XFILL_0__9383_ gnd vdd FILL
XFILL_5__15625_ gnd vdd FILL
XFILL_5__12837_ gnd vdd FILL
XFILL_5__7289_ gnd vdd FILL
XFILL_1__13106_ gnd vdd FILL
XFILL_3__8112_ gnd vdd FILL
XFILL_4__14266_ gnd vdd FILL
XFILL_3__9092_ gnd vdd FILL
XFILL_2__12657_ gnd vdd FILL
XFILL_1__10318_ gnd vdd FILL
XFILL_4__11478_ gnd vdd FILL
XFILL_2__15445_ gnd vdd FILL
XFILL_0__13836_ gnd vdd FILL
XFILL_3__14996_ gnd vdd FILL
XFILL_5__9028_ gnd vdd FILL
XFILL_1__14086_ gnd vdd FILL
XFILL_0__8334_ gnd vdd FILL
XFILL_4__16005_ gnd vdd FILL
XFILL_1__11298_ gnd vdd FILL
XSFILL53960x76050 gnd vdd FILL
XFILL_4__13217_ gnd vdd FILL
XFILL_4__10429_ gnd vdd FILL
XFILL_5__12768_ gnd vdd FILL
X_8962_ _8962_/A gnd _8964_/A vdd INVX1
XFILL_5__15556_ gnd vdd FILL
XSFILL3560x40050 gnd vdd FILL
XFILL_4__14197_ gnd vdd FILL
XFILL_1__13037_ gnd vdd FILL
XFILL_2__11608_ gnd vdd FILL
XFILL_3__13947_ gnd vdd FILL
XFILL_2__12588_ gnd vdd FILL
XFILL_1__10249_ gnd vdd FILL
XFILL_2__15376_ gnd vdd FILL
XFILL_0__13767_ gnd vdd FILL
XFILL_0__10979_ gnd vdd FILL
XSFILL28760x52050 gnd vdd FILL
XFILL_5__14507_ gnd vdd FILL
X_7913_ _7913_/Q _7664_/CLK _7920_/R vdd _7913_/D gnd vdd DFFSR
XFILL_5__11719_ gnd vdd FILL
XFILL_0__8265_ gnd vdd FILL
XFILL_4__13148_ gnd vdd FILL
XFILL_5__15487_ gnd vdd FILL
XFILL_5__12699_ gnd vdd FILL
X_8893_ _8893_/A _8893_/B _8892_/Y gnd _8893_/Y vdd OAI21X1
XFILL_0__15506_ gnd vdd FILL
XFILL_2__14327_ gnd vdd FILL
XFILL_2__11539_ gnd vdd FILL
XFILL_3__13878_ gnd vdd FILL
XFILL_0__12718_ gnd vdd FILL
XFILL_0__7216_ gnd vdd FILL
XFILL_6__9772_ gnd vdd FILL
XFILL_0__13698_ gnd vdd FILL
XFILL_5__14438_ gnd vdd FILL
X_7844_ _7824_/B _8868_/B gnd _7845_/C vdd NAND2X1
XFILL_0__8196_ gnd vdd FILL
XFILL_3__15617_ gnd vdd FILL
XFILL_4__13079_ gnd vdd FILL
XFILL_3__12829_ gnd vdd FILL
XFILL_2__14258_ gnd vdd FILL
XFILL_0__15437_ gnd vdd FILL
XFILL_0__12649_ gnd vdd FILL
XFILL_3__9994_ gnd vdd FILL
XFILL_6__8723_ gnd vdd FILL
XFILL_1__14988_ gnd vdd FILL
XSFILL33880x43050 gnd vdd FILL
XFILL_5__14369_ gnd vdd FILL
XFILL_2__13209_ gnd vdd FILL
XFILL_3__15548_ gnd vdd FILL
XFILL_0_CLKBUF1_insert118 gnd vdd FILL
X_7775_ _7697_/A _7156_/CLK _7775_/R vdd _7775_/D gnd vdd DFFSR
XFILL_2__14189_ gnd vdd FILL
XFILL_0_CLKBUF1_insert129 gnd vdd FILL
XFILL_0__15368_ gnd vdd FILL
XSFILL59160x7050 gnd vdd FILL
XFILL_1__13939_ gnd vdd FILL
XFILL111800x21050 gnd vdd FILL
XFILL_5__16108_ gnd vdd FILL
X_9514_ _9514_/A _9898_/B gnd _9515_/C vdd NAND2X1
XFILL_6__15659_ gnd vdd FILL
XFILL_0__7078_ gnd vdd FILL
XSFILL48920x65050 gnd vdd FILL
XFILL_1__7960_ gnd vdd FILL
XFILL_0__14319_ gnd vdd FILL
XFILL_3__15479_ gnd vdd FILL
XFILL_3__8876_ gnd vdd FILL
XSFILL64200x13050 gnd vdd FILL
XFILL_5__16039_ gnd vdd FILL
XFILL_0__15299_ gnd vdd FILL
XFILL_1__6911_ gnd vdd FILL
X_9445_ _9379_/A _7902_/CLK _7150_/R vdd _9445_/D gnd vdd DFFSR
XFILL_1__7891_ gnd vdd FILL
XFILL_1__15609_ gnd vdd FILL
XFILL_3__7827_ gnd vdd FILL
XFILL_1__9630_ gnd vdd FILL
X_9376_ _9376_/A gnd _9378_/A vdd INVX1
XFILL_1__6842_ gnd vdd FILL
XFILL_4_BUFX2_insert603 gnd vdd FILL
XFILL_3__7758_ gnd vdd FILL
XFILL_4_BUFX2_insert614 gnd vdd FILL
XSFILL3640x20050 gnd vdd FILL
XFILL_4_BUFX2_insert625 gnd vdd FILL
XFILL_6__7467_ gnd vdd FILL
X_8327_ _8325_/Y _8315_/B _8327_/C gnd _8411_/D vdd OAI21X1
XFILL_4_BUFX2_insert636 gnd vdd FILL
XFILL_4_BUFX2_insert647 gnd vdd FILL
XFILL_4__9270_ gnd vdd FILL
XFILL_4_BUFX2_insert658 gnd vdd FILL
XSFILL28840x32050 gnd vdd FILL
XFILL_3__7689_ gnd vdd FILL
XSFILL54120x65050 gnd vdd FILL
XFILL_1__8512_ gnd vdd FILL
XFILL_0__9719_ gnd vdd FILL
XFILL_4_BUFX2_insert669 gnd vdd FILL
XFILL112120x1050 gnd vdd FILL
X_8258_ _8187_/B _8642_/B gnd _8259_/C vdd NAND2X1
XFILL_3__9428_ gnd vdd FILL
XFILL_1__9492_ gnd vdd FILL
XFILL_4__8221_ gnd vdd FILL
X_7209_ _7271_/Q gnd _7211_/A vdd INVX1
XSFILL114680x76050 gnd vdd FILL
XFILL_1__8443_ gnd vdd FILL
X_8189_ _8187_/B _8701_/B gnd _8189_/Y vdd NAND2X1
XFILL_3__9359_ gnd vdd FILL
XFILL_2_BUFX2_insert80 gnd vdd FILL
XFILL_2_BUFX2_insert91 gnd vdd FILL
XSFILL33960x23050 gnd vdd FILL
XSFILL104920x53050 gnd vdd FILL
XFILL_1__8374_ gnd vdd FILL
XFILL_4__7103_ gnd vdd FILL
XFILL_4__8083_ gnd vdd FILL
XFILL_6__8019_ gnd vdd FILL
XFILL_1__7325_ gnd vdd FILL
XFILL_4__7034_ gnd vdd FILL
X_12830_ vdd _15167_/Y gnd _12830_/Y vdd NAND2X1
XFILL_1_BUFX2_insert504 gnd vdd FILL
XFILL_1_BUFX2_insert515 gnd vdd FILL
X_12761_ _12813_/Q gnd _12761_/Y vdd INVX1
XFILL_1__7187_ gnd vdd FILL
XFILL_1_BUFX2_insert526 gnd vdd FILL
XFILL_1_BUFX2_insert537 gnd vdd FILL
X_14500_ _14500_/A _14500_/B _14597_/C gnd _13015_/B vdd AOI21X1
XFILL_1_BUFX2_insert548 gnd vdd FILL
XFILL_4__8985_ gnd vdd FILL
X_11712_ _11257_/Y _11261_/Y _11271_/Y gnd _11726_/B vdd OAI21X1
XFILL_1_BUFX2_insert559 gnd vdd FILL
X_12692_ _12654_/A _12692_/CLK _12692_/R vdd _12692_/D gnd vdd DFFSR
X_15480_ _10720_/Q _15916_/B _15480_/C gnd _15481_/B vdd AOI21X1
XFILL_4__7936_ gnd vdd FILL
X_11643_ _11044_/A _11642_/Y _11762_/B gnd _11644_/C vdd AOI21X1
X_14431_ _9578_/Q gnd _14431_/Y vdd INVX1
XFILL_2__6951_ gnd vdd FILL
XFILL_4__7867_ gnd vdd FILL
XSFILL114760x56050 gnd vdd FILL
X_14362_ _14361_/Y _13843_/C _14506_/C _14360_/Y gnd _14366_/B vdd OAI22X1
X_11574_ _11577_/B _11574_/B _11574_/C gnd _11575_/C vdd OAI21X1
XFILL_2__9670_ gnd vdd FILL
XFILL_4__9606_ gnd vdd FILL
X_16101_ _16096_/Y _16097_/Y _16100_/Y gnd _16101_/Y vdd NAND3X1
XFILL_2__6882_ gnd vdd FILL
X_13313_ _13308_/A _13312_/Y _13253_/A gnd _13313_/Y vdd NAND3X1
X_10525_ _10595_/Q gnd _10525_/Y vdd INVX1
XFILL_4__7798_ gnd vdd FILL
XFILL_5__10050_ gnd vdd FILL
X_14293_ _14293_/A _14071_/B _13879_/B _14292_/Y gnd _14293_/Y vdd OAI22X1
XFILL_2__8621_ gnd vdd FILL
XFILL_5_BUFX2_insert470 gnd vdd FILL
XFILL_4__10780_ gnd vdd FILL
XFILL_5_BUFX2_insert481 gnd vdd FILL
XSFILL18840x64050 gnd vdd FILL
XFILL_5__8330_ gnd vdd FILL
XFILL_4__9537_ gnd vdd FILL
X_13244_ _13244_/A _13244_/B gnd _13244_/Y vdd OR2X2
X_16032_ _16032_/A _16032_/B gnd _16032_/Y vdd NOR2X1
XSFILL84280x40050 gnd vdd FILL
XFILL_5_BUFX2_insert492 gnd vdd FILL
X_10456_ _10364_/A _8792_/CLK _7896_/R vdd _10366_/Y gnd vdd DFFSR
XFILL_2__10910_ gnd vdd FILL
XFILL_0__10000_ gnd vdd FILL
XFILL_3__11160_ gnd vdd FILL
XSFILL64040x50 gnd vdd FILL
XFILL_1__9759_ gnd vdd FILL
XFILL_2__11890_ gnd vdd FILL
XFILL_5__8261_ gnd vdd FILL
XFILL_4__9468_ gnd vdd FILL
XFILL_3__10111_ gnd vdd FILL
XSFILL99320x62050 gnd vdd FILL
X_13175_ _11887_/A _13175_/CLK _13199_/R vdd _13175_/D gnd vdd DFFSR
XFILL_2__7503_ gnd vdd FILL
XFILL_4__12450_ gnd vdd FILL
X_10387_ _10387_/A _10450_/B _10386_/Y gnd _10463_/D vdd OAI21X1
XFILL_3__11091_ gnd vdd FILL
XFILL_2__8483_ gnd vdd FILL
XFILL_5__7212_ gnd vdd FILL
XFILL_1__12270_ gnd vdd FILL
X_12126_ _12126_/A _12137_/A _12126_/C gnd _12126_/Y vdd OAI21X1
XFILL_5__8192_ gnd vdd FILL
XFILL_4__9399_ gnd vdd FILL
XFILL_5__13740_ gnd vdd FILL
XFILL_4__11401_ gnd vdd FILL
XFILL_5__10952_ gnd vdd FILL
XFILL_3__10042_ gnd vdd FILL
XFILL_2__7434_ gnd vdd FILL
XFILL_4__12381_ gnd vdd FILL
XFILL_2__13560_ gnd vdd FILL
XFILL_1__11221_ gnd vdd FILL
XFILL_2__10772_ gnd vdd FILL
XFILL112280x22050 gnd vdd FILL
XFILL_0__11951_ gnd vdd FILL
XSFILL64040x48050 gnd vdd FILL
X_12057_ _12057_/A _12113_/B _12113_/C gnd gnd _12057_/Y vdd AOI22X1
XFILL_4__14120_ gnd vdd FILL
XFILL_2__12511_ gnd vdd FILL
XFILL_5__13671_ gnd vdd FILL
XFILL_4__11332_ gnd vdd FILL
XFILL_3__14850_ gnd vdd FILL
XFILL_5__10883_ gnd vdd FILL
XFILL_2__7365_ gnd vdd FILL
XFILL_0__10902_ gnd vdd FILL
XFILL_1__11152_ gnd vdd FILL
XFILL112280x7050 gnd vdd FILL
XFILL_2__13491_ gnd vdd FILL
XFILL_5__7074_ gnd vdd FILL
XFILL_0__14670_ gnd vdd FILL
X_11008_ _12222_/Y _11007_/Y gnd _11008_/Y vdd NOR2X1
XFILL_5__12622_ gnd vdd FILL
XFILL_0__11882_ gnd vdd FILL
XFILL_5__15410_ gnd vdd FILL
XFILL_2__9104_ gnd vdd FILL
XFILL_5__16390_ gnd vdd FILL
XFILL_3__13801_ gnd vdd FILL
XFILL_4__14051_ gnd vdd FILL
XFILL_2__15230_ gnd vdd FILL
XFILL_2__12442_ gnd vdd FILL
XFILL_4__11263_ gnd vdd FILL
XFILL_1__10103_ gnd vdd FILL
XFILL_2__7296_ gnd vdd FILL
XFILL_0__13621_ gnd vdd FILL
XFILL_3__14781_ gnd vdd FILL
XSFILL3480x55050 gnd vdd FILL
XFILL_1__15960_ gnd vdd FILL
XFILL_3__11993_ gnd vdd FILL
XFILL_1__11083_ gnd vdd FILL
XFILL_0__10833_ gnd vdd FILL
XFILL_5__15341_ gnd vdd FILL
X_15816_ _15813_/Y _15816_/B gnd _15816_/Y vdd NOR2X1
XFILL_4__13002_ gnd vdd FILL
XFILL_2__9035_ gnd vdd FILL
XFILL_3__13732_ gnd vdd FILL
XFILL_2_BUFX2_insert360 gnd vdd FILL
XFILL_2__15161_ gnd vdd FILL
XFILL_4__11194_ gnd vdd FILL
XFILL_6__14892_ gnd vdd FILL
XFILL_0__16340_ gnd vdd FILL
XFILL_3__10944_ gnd vdd FILL
XFILL_2__12373_ gnd vdd FILL
XSFILL69160x2050 gnd vdd FILL
XFILL_1__10034_ gnd vdd FILL
XFILL_1__14911_ gnd vdd FILL
XFILL_2_BUFX2_insert371 gnd vdd FILL
XFILL_0__13552_ gnd vdd FILL
XFILL_0__10764_ gnd vdd FILL
XFILL_5__11504_ gnd vdd FILL
XFILL_2_BUFX2_insert382 gnd vdd FILL
XFILL_1__15891_ gnd vdd FILL
XFILL_6__13843_ gnd vdd FILL
XFILL_2_BUFX2_insert393 gnd vdd FILL
X_15747_ _15747_/A gnd _15748_/B vdd INVX1
XFILL_5__15272_ gnd vdd FILL
XFILL_3__16451_ gnd vdd FILL
XFILL_5__12484_ gnd vdd FILL
XFILL_4__10145_ gnd vdd FILL
XFILL_2__11324_ gnd vdd FILL
XFILL_2__14112_ gnd vdd FILL
X_12959_ _12957_/Y vdd _12958_/Y gnd _12959_/Y vdd OAI21X1
XFILL_0__12503_ gnd vdd FILL
XFILL_3__13663_ gnd vdd FILL
XFILL_2__15092_ gnd vdd FILL
XSFILL84360x20050 gnd vdd FILL
XFILL_6_CLKBUF1_insert1078 gnd vdd FILL
XFILL_1__14842_ gnd vdd FILL
XFILL_3__10875_ gnd vdd FILL
XFILL_0__16271_ gnd vdd FILL
XFILL_5__14223_ gnd vdd FILL
XFILL_0__13483_ gnd vdd FILL
XFILL_5__7976_ gnd vdd FILL
XFILL_3__15402_ gnd vdd FILL
XSFILL59000x37050 gnd vdd FILL
XFILL_5__11435_ gnd vdd FILL
XFILL_0__10695_ gnd vdd FILL
X_15678_ _10341_/Q _15178_/C _15678_/C gnd _15678_/Y vdd AOI21X1
XFILL_3__12614_ gnd vdd FILL
XFILL_2__14043_ gnd vdd FILL
XFILL_4__14953_ gnd vdd FILL
XFILL_3__16382_ gnd vdd FILL
XFILL_0__15222_ gnd vdd FILL
XFILL_2__11255_ gnd vdd FILL
XFILL_0__12434_ gnd vdd FILL
XFILL_3__13594_ gnd vdd FILL
XSFILL99400x42050 gnd vdd FILL
XFILL_1__14773_ gnd vdd FILL
XFILL_3__6991_ gnd vdd FILL
XFILL_5__6927_ gnd vdd FILL
XFILL_1__11985_ gnd vdd FILL
X_14629_ _9326_/Q _13854_/B _14629_/C gnd _14630_/B vdd AOI21X1
XFILL_5__14154_ gnd vdd FILL
XFILL_4__13904_ gnd vdd FILL
XFILL_3__15333_ gnd vdd FILL
X_7560_ _7560_/A gnd _7560_/Y vdd INVX1
XFILL_5__11366_ gnd vdd FILL
XFILL_3__8730_ gnd vdd FILL
XFILL_2__9937_ gnd vdd FILL
XFILL_4__14884_ gnd vdd FILL
XFILL_1__10936_ gnd vdd FILL
XFILL_0__15153_ gnd vdd FILL
XFILL_2__11186_ gnd vdd FILL
XFILL_1__13724_ gnd vdd FILL
XFILL_0__12365_ gnd vdd FILL
XFILL_5__13105_ gnd vdd FILL
XFILL_5__9646_ gnd vdd FILL
XFILL_5__10317_ gnd vdd FILL
XFILL_5__6858_ gnd vdd FILL
XFILL_6__15444_ gnd vdd FILL
XFILL_4__13835_ gnd vdd FILL
XSFILL64120x28050 gnd vdd FILL
XFILL_0__8952_ gnd vdd FILL
XFILL_5__14085_ gnd vdd FILL
XFILL_2__10137_ gnd vdd FILL
XFILL_5__11297_ gnd vdd FILL
X_7491_ _7489_/Y _7430_/A _7490_/Y gnd _7535_/D vdd OAI21X1
XFILL_3__15264_ gnd vdd FILL
XFILL_0__14104_ gnd vdd FILL
XFILL_2__9868_ gnd vdd FILL
XFILL_1__13655_ gnd vdd FILL
XFILL_3__12476_ gnd vdd FILL
XBUFX2_insert370 _13338_/Y gnd _9466_/A vdd BUFX2
XFILL_0__11316_ gnd vdd FILL
XFILL_3__8661_ gnd vdd FILL
XBUFX2_insert381 _13331_/Y gnd _9163_/A vdd BUFX2
XFILL_2__15994_ gnd vdd FILL
XFILL_0__15084_ gnd vdd FILL
X_9230_ _9310_/Q gnd _9232_/A vdd INVX1
XSFILL74280x72050 gnd vdd FILL
XBUFX2_insert392 _12387_/Y gnd _7329_/B vdd BUFX2
XFILL_5__13036_ gnd vdd FILL
XFILL_0__12296_ gnd vdd FILL
XFILL_5__10248_ gnd vdd FILL
XFILL_3__14215_ gnd vdd FILL
XFILL_3__7612_ gnd vdd FILL
XFILL_1__12606_ gnd vdd FILL
XFILL_4__13766_ gnd vdd FILL
XFILL_0__8883_ gnd vdd FILL
XFILL_3__11427_ gnd vdd FILL
XFILL_4__10978_ gnd vdd FILL
XFILL_3__15195_ gnd vdd FILL
XFILL_0__14035_ gnd vdd FILL
XFILL_2__10068_ gnd vdd FILL
XFILL_2__14945_ gnd vdd FILL
XFILL_1__13586_ gnd vdd FILL
XFILL_3__8592_ gnd vdd FILL
XFILL_1__16374_ gnd vdd FILL
XFILL_5__8528_ gnd vdd FILL
XFILL_2__9799_ gnd vdd FILL
XFILL_0__11247_ gnd vdd FILL
XFILL_4__15505_ gnd vdd FILL
XFILL_1__10798_ gnd vdd FILL
XFILL_6__11538_ gnd vdd FILL
XFILL_4__12717_ gnd vdd FILL
XFILL_0__7834_ gnd vdd FILL
X_9161_ _9161_/A _9086_/B _9161_/C gnd _9161_/Y vdd OAI21X1
XFILL_3__14146_ gnd vdd FILL
XFILL_5__10179_ gnd vdd FILL
XFILL_1__15325_ gnd vdd FILL
XFILL_3__7543_ gnd vdd FILL
XFILL_4__13697_ gnd vdd FILL
XFILL_3__11358_ gnd vdd FILL
XFILL_2__14876_ gnd vdd FILL
XFILL_5__8459_ gnd vdd FILL
X_8112_ _8133_/A _9008_/B gnd _8113_/C vdd NAND2X1
XFILL_0__11178_ gnd vdd FILL
XFILL_6__14257_ gnd vdd FILL
XFILL_4__15436_ gnd vdd FILL
XFILL_4__12648_ gnd vdd FILL
X_9092_ _9090_/Y _9101_/B _9092_/C gnd _9178_/D vdd OAI21X1
XSFILL28760x47050 gnd vdd FILL
XFILL_3__10309_ gnd vdd FILL
XFILL_0__7765_ gnd vdd FILL
XFILL_2__13827_ gnd vdd FILL
XFILL_1__15256_ gnd vdd FILL
XFILL_5__14987_ gnd vdd FILL
XFILL_3__11289_ gnd vdd FILL
XFILL_3__14077_ gnd vdd FILL
XFILL_1__12468_ gnd vdd FILL
XFILL_3__7474_ gnd vdd FILL
XFILL_0__10129_ gnd vdd FILL
XFILL_6__13208_ gnd vdd FILL
XFILL_0__15986_ gnd vdd FILL
XFILL_0__9504_ gnd vdd FILL
X_8043_ _7989_/A _7915_/CLK _7915_/R vdd _8043_/D gnd vdd DFFSR
XFILL_6__7183_ gnd vdd FILL
XFILL_0__7696_ gnd vdd FILL
XFILL_4__15367_ gnd vdd FILL
XFILL_1__14207_ gnd vdd FILL
XFILL_5__13938_ gnd vdd FILL
XFILL_3__13028_ gnd vdd FILL
XFILL_3__9213_ gnd vdd FILL
XFILL_4__12579_ gnd vdd FILL
XFILL_1__11419_ gnd vdd FILL
XFILL_1__15187_ gnd vdd FILL
XFILL_2__13758_ gnd vdd FILL
XFILL_1__12399_ gnd vdd FILL
XFILL_0__14937_ gnd vdd FILL
XFILL_4__14318_ gnd vdd FILL
XSFILL3560x4050 gnd vdd FILL
XSFILL69240x61050 gnd vdd FILL
XSFILL103560x42050 gnd vdd FILL
XFILL_5__13869_ gnd vdd FILL
XFILL_2__12709_ gnd vdd FILL
XFILL_4__15298_ gnd vdd FILL
XFILL_1__14138_ gnd vdd FILL
XFILL_3__9144_ gnd vdd FILL
XSFILL33880x38050 gnd vdd FILL
XFILL_0__14868_ gnd vdd FILL
XFILL_2__13689_ gnd vdd FILL
XFILL_5__15608_ gnd vdd FILL
XFILL_4__14249_ gnd vdd FILL
XFILL_0__9366_ gnd vdd FILL
X_9994_ _9994_/A _9993_/A _9994_/C gnd _9994_/Y vdd OAI21X1
XFILL_2__15428_ gnd vdd FILL
XFILL_0__13819_ gnd vdd FILL
XFILL_3__14979_ gnd vdd FILL
XFILL_1__14069_ gnd vdd FILL
XSFILL104440x70050 gnd vdd FILL
XFILL_1__7110_ gnd vdd FILL
XFILL_0__14799_ gnd vdd FILL
XFILL_0__8317_ gnd vdd FILL
XFILL_1__8090_ gnd vdd FILL
XFILL_5__15539_ gnd vdd FILL
XFILL_0__9297_ gnd vdd FILL
X_8945_ _8945_/Q _9589_/CLK _7413_/R vdd _8945_/D gnd vdd DFFSR
XFILL_2__15359_ gnd vdd FILL
XFILL_1__7041_ gnd vdd FILL
XFILL_0__8248_ gnd vdd FILL
XSFILL49000x69050 gnd vdd FILL
X_8876_ _8936_/Q gnd _8878_/A vdd INVX1
XSFILL3640x15050 gnd vdd FILL
X_7827_ _7827_/A _7878_/B _7827_/C gnd _7903_/D vdd OAI21X1
XSFILL28840x27050 gnd vdd FILL
XFILL_4__8770_ gnd vdd FILL
XFILL_3__9977_ gnd vdd FILL
X_7758_ _7759_/B _8014_/B gnd _7758_/Y vdd NAND2X1
XFILL_1__8992_ gnd vdd FILL
XFILL_4__7721_ gnd vdd FILL
XSFILL94520x65050 gnd vdd FILL
XFILL_1__7943_ gnd vdd FILL
X_7689_ _7690_/B _7177_/B gnd _7690_/C vdd NAND2X1
XFILL_3__8859_ gnd vdd FILL
XFILL_6__8568_ gnd vdd FILL
X_9428_ _9372_/B _9556_/B gnd _9428_/Y vdd NAND2X1
XSFILL33960x18050 gnd vdd FILL
XFILL_1__7874_ gnd vdd FILL
X_10310_ _10308_/Y _10264_/A _10310_/C gnd _10352_/D vdd OAI21X1
XFILL_4__7583_ gnd vdd FILL
XFILL_4_BUFX2_insert400 gnd vdd FILL
XFILL_1__9613_ gnd vdd FILL
XFILL_4_BUFX2_insert411 gnd vdd FILL
X_11290_ _11290_/A gnd _11546_/A vdd INVX1
XSFILL18760x79050 gnd vdd FILL
X_9359_ _9359_/A _8719_/B gnd _9360_/C vdd NAND2X1
XFILL_4_BUFX2_insert422 gnd vdd FILL
XFILL_4_BUFX2_insert433 gnd vdd FILL
XSFILL104520x50050 gnd vdd FILL
X_10241_ _10239_/Y _10318_/A _10241_/C gnd _10329_/D vdd OAI21X1
XFILL_4_BUFX2_insert444 gnd vdd FILL
XSFILL33800x82050 gnd vdd FILL
XFILL_4_BUFX2_insert455 gnd vdd FILL
XFILL_4_BUFX2_insert466 gnd vdd FILL
XFILL_1__9544_ gnd vdd FILL
XFILL_4_BUFX2_insert477 gnd vdd FILL
XFILL_4__9253_ gnd vdd FILL
XFILL_4_BUFX2_insert488 gnd vdd FILL
X_10172_ _10191_/B _7868_/B gnd _10173_/C vdd NAND2X1
XFILL_4_BUFX2_insert499 gnd vdd FILL
XFILL_1__9475_ gnd vdd FILL
XFILL_4__8204_ gnd vdd FILL
X_14980_ _12812_/Q gnd _14980_/Y vdd INVX2
XFILL_4__8135_ gnd vdd FILL
XSFILL38280x32050 gnd vdd FILL
X_13931_ _7188_/A _14762_/B _14413_/A _8212_/A gnd _13931_/Y vdd AOI22X1
XFILL_1__8357_ gnd vdd FILL
XFILL_3_CLKBUF1_insert113 gnd vdd FILL
XFILL_4__8066_ gnd vdd FILL
XSFILL79160x44050 gnd vdd FILL
XFILL_3_CLKBUF1_insert124 gnd vdd FILL
XFILL_3_CLKBUF1_insert135 gnd vdd FILL
X_13862_ _13853_/Y _13854_/Y _13862_/C gnd _13862_/Y vdd NAND3X1
XFILL_1__7308_ gnd vdd FILL
XFILL_3_CLKBUF1_insert146 gnd vdd FILL
XFILL_2__7081_ gnd vdd FILL
XFILL_3_CLKBUF1_insert157 gnd vdd FILL
XSFILL69400x21050 gnd vdd FILL
XFILL_3_CLKBUF1_insert168 gnd vdd FILL
X_15601_ _14999_/A _15601_/B _14088_/D _15172_/A gnd _15601_/Y vdd OAI22X1
X_12813_ _12813_/Q _12685_/CLK _12685_/R vdd _12813_/D gnd vdd DFFSR
XFILL_3_CLKBUF1_insert179 gnd vdd FILL
XFILL_1_BUFX2_insert301 gnd vdd FILL
X_13793_ _9949_/Q gnd _13793_/Y vdd INVX1
XSFILL114360x53050 gnd vdd FILL
XFILL_1_BUFX2_insert312 gnd vdd FILL
XFILL_1__7239_ gnd vdd FILL
XFILL_1_BUFX2_insert323 gnd vdd FILL
XFILL_5__7830_ gnd vdd FILL
XSFILL18840x59050 gnd vdd FILL
X_15532_ _13995_/A _15622_/A _15726_/A _15531_/Y gnd _15532_/Y vdd OAI22X1
XFILL_1_BUFX2_insert334 gnd vdd FILL
X_12744_ _12762_/A memoryOutData[16] gnd _12745_/C vdd NAND2X1
XFILL_1_BUFX2_insert345 gnd vdd FILL
XFILL_3__10660_ gnd vdd FILL
XFILL_1_BUFX2_insert356 gnd vdd FILL
XFILL_1_BUFX2_insert367 gnd vdd FILL
XFILL_4__8968_ gnd vdd FILL
XFILL_1_BUFX2_insert378 gnd vdd FILL
XFILL_5__11220_ gnd vdd FILL
XFILL_5__7761_ gnd vdd FILL
XSFILL99320x57050 gnd vdd FILL
XFILL_1_BUFX2_insert389 gnd vdd FILL
XSFILL59080x11050 gnd vdd FILL
X_15463_ _15172_/A _13966_/A _16155_/D _13948_/D gnd _15463_/Y vdd OAI22X1
X_12675_ _12675_/Q _12685_/CLK _12799_/R vdd _12675_/D gnd vdd DFFSR
XFILL_4__11950_ gnd vdd FILL
XFILL_2__11040_ gnd vdd FILL
XFILL_5__9500_ gnd vdd FILL
XFILL_2__7983_ gnd vdd FILL
XFILL_1__11770_ gnd vdd FILL
XFILL_6__12510_ gnd vdd FILL
X_14414_ _8426_/Q _14414_/B _14868_/A _14414_/D gnd _14414_/Y vdd AOI22X1
XFILL_5__7692_ gnd vdd FILL
XFILL_4__10901_ gnd vdd FILL
XFILL_6__13490_ gnd vdd FILL
XFILL_5__11151_ gnd vdd FILL
XFILL_4__8899_ gnd vdd FILL
X_11626_ _11150_/C _11802_/A _11626_/C gnd _11626_/Y vdd NAND3X1
X_15394_ _15394_/A _15394_/B _15394_/C _13869_/Y gnd _15394_/Y vdd OAI22X1
XFILL_3__12330_ gnd vdd FILL
XFILL_2__9722_ gnd vdd FILL
XFILL_4__11881_ gnd vdd FILL
XFILL_2__6934_ gnd vdd FILL
XFILL_0__12150_ gnd vdd FILL
XFILL_5__10102_ gnd vdd FILL
XFILL_4__13620_ gnd vdd FILL
X_14345_ _14345_/A _14344_/Y _14340_/Y gnd _14345_/Y vdd NAND3X1
XFILL_5__11082_ gnd vdd FILL
X_11557_ _11554_/Y _11556_/Y gnd _11558_/A vdd AND2X2
XFILL_4__10832_ gnd vdd FILL
XFILL_2__9653_ gnd vdd FILL
XFILL_1__13440_ gnd vdd FILL
XFILL_3__12261_ gnd vdd FILL
XFILL_0__11101_ gnd vdd FILL
XFILL_1__10652_ gnd vdd FILL
XFILL_2__6865_ gnd vdd FILL
XFILL_0__12081_ gnd vdd FILL
XFILL_5__9362_ gnd vdd FILL
XFILL_2__12991_ gnd vdd FILL
X_10508_ _10535_/A _9100_/B gnd _10508_/Y vdd NAND2X1
XFILL_6__12372_ gnd vdd FILL
XFILL_3__14000_ gnd vdd FILL
XFILL_5__10033_ gnd vdd FILL
XFILL_5__14910_ gnd vdd FILL
XFILL_2__8604_ gnd vdd FILL
XFILL_4__13551_ gnd vdd FILL
X_11488_ _11485_/Y _11481_/Y _11487_/Y gnd _12093_/A vdd NAND3X1
X_14276_ _8617_/A gnd _14278_/B vdd INVX1
XFILL_3__11212_ gnd vdd FILL
XFILL_4__10763_ gnd vdd FILL
XFILL_2__14730_ gnd vdd FILL
XFILL_3__12192_ gnd vdd FILL
XSFILL79240x24050 gnd vdd FILL
XFILL_5__15890_ gnd vdd FILL
XFILL_1__13371_ gnd vdd FILL
XFILL_2__11942_ gnd vdd FILL
XFILL_5__8313_ gnd vdd FILL
XFILL_0__11032_ gnd vdd FILL
XFILL112120x81050 gnd vdd FILL
X_16015_ _10862_/Q gnd _16016_/A vdd INVX1
XFILL_6__11323_ gnd vdd FILL
X_13227_ _13220_/A _13305_/A gnd _13231_/A vdd NOR2X1
XFILL_5__9293_ gnd vdd FILL
XFILL_4__12502_ gnd vdd FILL
X_10439_ _10481_/Q gnd _10441_/A vdd INVX1
XFILL_6__15091_ gnd vdd FILL
XFILL_5__14841_ gnd vdd FILL
XFILL_3__11143_ gnd vdd FILL
XFILL_1__15110_ gnd vdd FILL
XFILL_4__16270_ gnd vdd FILL
XFILL_1__12322_ gnd vdd FILL
XFILL_4__13482_ gnd vdd FILL
XFILL_4__10694_ gnd vdd FILL
XFILL_1__16090_ gnd vdd FILL
XFILL_0__15840_ gnd vdd FILL
XFILL_2__14661_ gnd vdd FILL
XFILL_2__11873_ gnd vdd FILL
XSFILL83720x49050 gnd vdd FILL
XFILL_6__14042_ gnd vdd FILL
XFILL_5__8244_ gnd vdd FILL
XFILL_4__15221_ gnd vdd FILL
XSFILL114440x33050 gnd vdd FILL
XFILL_0__7550_ gnd vdd FILL
X_13158_ _13149_/A _13158_/B gnd _13159_/C vdd NAND2X1
XFILL_2__16400_ gnd vdd FILL
XFILL_4__12433_ gnd vdd FILL
XFILL_2__13612_ gnd vdd FILL
XFILL_5__11984_ gnd vdd FILL
XFILL_1__15041_ gnd vdd FILL
XFILL_3__15951_ gnd vdd FILL
XFILL_3__11074_ gnd vdd FILL
XFILL_5__14772_ gnd vdd FILL
XFILL_1__12253_ gnd vdd FILL
XFILL_2__8466_ gnd vdd FILL
XFILL_2__10824_ gnd vdd FILL
XFILL_2__14592_ gnd vdd FILL
XFILL_0__15771_ gnd vdd FILL
XSFILL84360x15050 gnd vdd FILL
X_12109_ _12109_/A _12113_/B _12113_/C gnd gnd _12110_/C vdd AOI22X1
XFILL_0__12983_ gnd vdd FILL
XFILL_5__10935_ gnd vdd FILL
X_13089_ _13168_/B _13089_/B gnd _13089_/Y vdd NAND2X1
XFILL_0__7481_ gnd vdd FILL
XFILL_5__13723_ gnd vdd FILL
XFILL_6__11185_ gnd vdd FILL
XFILL_4__15152_ gnd vdd FILL
XFILL_3__14902_ gnd vdd FILL
XFILL_3__10025_ gnd vdd FILL
XFILL_4__12364_ gnd vdd FILL
XFILL_2__16331_ gnd vdd FILL
XFILL_2__7417_ gnd vdd FILL
XFILL_1__11204_ gnd vdd FILL
XFILL_2__10755_ gnd vdd FILL
XFILL_0__14722_ gnd vdd FILL
XFILL_3__7190_ gnd vdd FILL
XFILL_2__13543_ gnd vdd FILL
XFILL_3__15882_ gnd vdd FILL
XFILL_2__8397_ gnd vdd FILL
XFILL_0__11934_ gnd vdd FILL
XFILL_1__12184_ gnd vdd FILL
XSFILL99400x37050 gnd vdd FILL
XFILL_0__9220_ gnd vdd FILL
XFILL_4__14103_ gnd vdd FILL
XFILL_5__13654_ gnd vdd FILL
XFILL_4__11315_ gnd vdd FILL
XFILL_3__14833_ gnd vdd FILL
XFILL_4__15083_ gnd vdd FILL
XFILL_4__12295_ gnd vdd FILL
XFILL_1__11135_ gnd vdd FILL
XFILL_2__16262_ gnd vdd FILL
XFILL_2__7348_ gnd vdd FILL
XFILL_2__10686_ gnd vdd FILL
XFILL_2__13474_ gnd vdd FILL
XFILL_0__14653_ gnd vdd FILL
XFILL_5__12605_ gnd vdd FILL
XFILL_0__9151_ gnd vdd FILL
XFILL_0__11865_ gnd vdd FILL
XFILL_5__7057_ gnd vdd FILL
XFILL_4__14034_ gnd vdd FILL
XFILL_6__10067_ gnd vdd FILL
XFILL_5__13585_ gnd vdd FILL
XFILL_2__15213_ gnd vdd FILL
XFILL_4__11246_ gnd vdd FILL
XFILL_5__16373_ gnd vdd FILL
X_6991_ _6989_/Y _6951_/A _6991_/C gnd _7027_/D vdd OAI21X1
XFILL_0__13604_ gnd vdd FILL
XFILL_2__12425_ gnd vdd FILL
XFILL_5__10797_ gnd vdd FILL
XFILL_3__14764_ gnd vdd FILL
XFILL_0__10816_ gnd vdd FILL
XFILL_3__11976_ gnd vdd FILL
XFILL_0__8102_ gnd vdd FILL
XFILL_2__16193_ gnd vdd FILL
XFILL_1__15943_ gnd vdd FILL
XFILL_1__11066_ gnd vdd FILL
XFILL_0__14584_ gnd vdd FILL
XFILL_6__7870_ gnd vdd FILL
XFILL_5__15324_ gnd vdd FILL
X_8730_ _8802_/Q gnd _8730_/Y vdd INVX1
XFILL_0__11796_ gnd vdd FILL
XFILL_0__9082_ gnd vdd FILL
XFILL_2__9018_ gnd vdd FILL
XFILL_3__13715_ gnd vdd FILL
XFILL_3__9900_ gnd vdd FILL
XFILL_3__10927_ gnd vdd FILL
XFILL_2__12356_ gnd vdd FILL
XFILL_1__10017_ gnd vdd FILL
XFILL_0__16323_ gnd vdd FILL
XFILL_2__15144_ gnd vdd FILL
XFILL_4__11177_ gnd vdd FILL
XFILL_3__14695_ gnd vdd FILL
XFILL_0__13535_ gnd vdd FILL
XFILL_0__10747_ gnd vdd FILL
XFILL_1__15874_ gnd vdd FILL
XFILL_5__15255_ gnd vdd FILL
XFILL_4__10128_ gnd vdd FILL
XFILL112200x61050 gnd vdd FILL
XSFILL49080x43050 gnd vdd FILL
XFILL_5__12467_ gnd vdd FILL
XFILL_2__11307_ gnd vdd FILL
X_8661_ _8661_/A _8607_/B _8660_/Y gnd _8661_/Y vdd OAI21X1
XFILL_3__13646_ gnd vdd FILL
XFILL_4__15985_ gnd vdd FILL
XFILL_1__14825_ gnd vdd FILL
XFILL_2__15075_ gnd vdd FILL
XFILL_2__12287_ gnd vdd FILL
XFILL_0__16254_ gnd vdd FILL
XFILL_5__14206_ gnd vdd FILL
XFILL_0__13466_ gnd vdd FILL
XFILL_0__10678_ gnd vdd FILL
X_7612_ _7592_/B _9788_/B gnd _7613_/C vdd NAND2X1
XFILL_5__7959_ gnd vdd FILL
XFILL_5__11418_ gnd vdd FILL
XFILL_5__15186_ gnd vdd FILL
X_8592_ _8590_/Y _8577_/B _8592_/C gnd _8670_/D vdd OAI21X1
XFILL_1_BUFX2_insert890 gnd vdd FILL
XFILL_5__12398_ gnd vdd FILL
XFILL_0__15205_ gnd vdd FILL
XFILL_4__10059_ gnd vdd FILL
XFILL_3__16365_ gnd vdd FILL
XFILL_2__14026_ gnd vdd FILL
XFILL_4__14936_ gnd vdd FILL
XFILL_2__11238_ gnd vdd FILL
XFILL_0__12417_ gnd vdd FILL
XFILL_3__9762_ gnd vdd FILL
XSFILL114520x13050 gnd vdd FILL
XFILL_3__13577_ gnd vdd FILL
XFILL_3__10789_ gnd vdd FILL
XFILL_3__6974_ gnd vdd FILL
XFILL_0__16185_ gnd vdd FILL
XFILL_1__11968_ gnd vdd FILL
XFILL_1__14756_ gnd vdd FILL
XFILL_0__13397_ gnd vdd FILL
XFILL_5__14137_ gnd vdd FILL
XFILL_3__15316_ gnd vdd FILL
X_7543_ _8183_/A _7562_/B gnd _7543_/Y vdd NAND2X1
XFILL_5__11349_ gnd vdd FILL
XFILL_0__9984_ gnd vdd FILL
XFILL_4__14867_ gnd vdd FILL
XFILL_3__8713_ gnd vdd FILL
XFILL_3__12528_ gnd vdd FILL
XFILL_1__10919_ gnd vdd FILL
XSFILL28360x44050 gnd vdd FILL
XFILL_3__16296_ gnd vdd FILL
XFILL_0__15136_ gnd vdd FILL
XFILL_1__13707_ gnd vdd FILL
XFILL_2__11169_ gnd vdd FILL
XFILL_0__12348_ gnd vdd FILL
XFILL_5__9629_ gnd vdd FILL
XFILL_1__11899_ gnd vdd FILL
XFILL_1__14687_ gnd vdd FILL
XFILL_6__12639_ gnd vdd FILL
XFILL_4__13818_ gnd vdd FILL
XFILL_5__14068_ gnd vdd FILL
XFILL_3__15247_ gnd vdd FILL
X_7474_ _7530_/Q gnd _7476_/A vdd INVX1
XSFILL69240x56050 gnd vdd FILL
XFILL_3__12459_ gnd vdd FILL
XFILL_4__14798_ gnd vdd FILL
XFILL_3__8644_ gnd vdd FILL
XFILL_2__15977_ gnd vdd FILL
XFILL_1__13638_ gnd vdd FILL
XFILL_0__15067_ gnd vdd FILL
XFILL_5__13019_ gnd vdd FILL
XFILL_0__12279_ gnd vdd FILL
X_9213_ _9238_/B _7293_/B gnd _9214_/C vdd NAND2X1
XFILL_4__13749_ gnd vdd FILL
XFILL_0__8866_ gnd vdd FILL
XFILL_3__15178_ gnd vdd FILL
XFILL_0__14018_ gnd vdd FILL
XFILL_2__14928_ gnd vdd FILL
XFILL_3__8575_ gnd vdd FILL
XFILL_1__13569_ gnd vdd FILL
XFILL_1__16357_ gnd vdd FILL
XSFILL104440x65050 gnd vdd FILL
XFILL_0__7817_ gnd vdd FILL
X_9144_ _9144_/A gnd _9144_/Y vdd INVX1
XFILL_1__7590_ gnd vdd FILL
XFILL_3__14129_ gnd vdd FILL
XSFILL8680x63050 gnd vdd FILL
XFILL_1__15308_ gnd vdd FILL
XSFILL23720x12050 gnd vdd FILL
XFILL_2__14859_ gnd vdd FILL
XFILL_1__16288_ gnd vdd FILL
XFILL_3_BUFX2_insert407 gnd vdd FILL
XFILL_4__15419_ gnd vdd FILL
X_9075_ _9075_/Q _8947_/CLK _9069_/R vdd _9075_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert418 gnd vdd FILL
XFILL_0__7748_ gnd vdd FILL
XFILL_3_BUFX2_insert429 gnd vdd FILL
XFILL_4__16399_ gnd vdd FILL
XFILL_3__7457_ gnd vdd FILL
XFILL_1__15239_ gnd vdd FILL
XSFILL89400x69050 gnd vdd FILL
XFILL_0__15969_ gnd vdd FILL
X_8026_ _7938_/A _9050_/CLK _7258_/R vdd _8026_/D gnd vdd DFFSR
XFILL_1__9260_ gnd vdd FILL
XFILL_0__7679_ gnd vdd FILL
XFILL_0__9418_ gnd vdd FILL
XFILL_1__8211_ gnd vdd FILL
XFILL_3__9127_ gnd vdd FILL
XSFILL109160x77050 gnd vdd FILL
XFILL_1__8142_ gnd vdd FILL
XFILL_0__9349_ gnd vdd FILL
X_9977_ _9977_/A gnd _9979_/A vdd INVX1
XFILL_4__9940_ gnd vdd FILL
XSFILL39080x75050 gnd vdd FILL
XFILL_1__8073_ gnd vdd FILL
X_8928_ _8928_/Q _7535_/CLK _8431_/R vdd _8854_/Y gnd vdd DFFSR
XFILL_3__8009_ gnd vdd FILL
XFILL_4__9871_ gnd vdd FILL
XFILL_4_CLKBUF1_insert208 gnd vdd FILL
X_10790_ _14252_/D gnd _10792_/A vdd INVX1
XFILL_6__7999_ gnd vdd FILL
XFILL_4_CLKBUF1_insert219 gnd vdd FILL
XFILL_4__8822_ gnd vdd FILL
X_8859_ _8859_/A _8091_/B gnd _8860_/C vdd NAND2X1
XSFILL8760x43050 gnd vdd FILL
XSFILL33800x77050 gnd vdd FILL
XFILL_0_BUFX2_insert308 gnd vdd FILL
XFILL_0_BUFX2_insert319 gnd vdd FILL
XFILL_4__8753_ gnd vdd FILL
X_12460_ _12364_/A gnd _12462_/A vdd INVX1
XFILL_1__8975_ gnd vdd FILL
XFILL_4__7704_ gnd vdd FILL
XSFILL104360x7050 gnd vdd FILL
X_11411_ _11411_/A _11411_/B _11411_/C gnd _11411_/Y vdd AOI21X1
X_12391_ _11936_/B gnd _12391_/Y vdd INVX1
XFILL_1__7926_ gnd vdd FILL
XFILL_4__7635_ gnd vdd FILL
X_14130_ _8420_/Q _13647_/B _14557_/C _8292_/Q gnd _14133_/A vdd AOI22X1
X_11342_ _11230_/Y _11341_/Y _11342_/C gnd _12113_/A vdd NAND3X1
XSFILL13720x44050 gnd vdd FILL
XFILL_1__7857_ gnd vdd FILL
XFILL_4__7566_ gnd vdd FILL
XSFILL8680x50 gnd vdd FILL
XFILL_4_BUFX2_insert230 gnd vdd FILL
X_14061_ _14061_/A _14830_/B _14643_/C _14060_/Y gnd _14061_/Y vdd OAI22X1
XFILL_4_BUFX2_insert241 gnd vdd FILL
X_11273_ _11274_/A _11083_/Y gnd _11709_/A vdd NOR2X1
XFILL_4_BUFX2_insert252 gnd vdd FILL
XFILL_4_BUFX2_insert263 gnd vdd FILL
XFILL_4_BUFX2_insert274 gnd vdd FILL
X_10224_ _14732_/A _7268_/CLK _9313_/R vdd _10182_/Y gnd vdd DFFSR
X_13012_ vdd _13012_/B gnd _13013_/C vdd NAND2X1
XFILL_4_BUFX2_insert285 gnd vdd FILL
XFILL_4__7497_ gnd vdd FILL
XFILL_1__9527_ gnd vdd FILL
XFILL_2__8320_ gnd vdd FILL
XFILL_4_BUFX2_insert296 gnd vdd FILL
XFILL_5_BUFX2_insert1009 gnd vdd FILL
XFILL_4__9236_ gnd vdd FILL
X_10155_ _10153_/Y _10140_/B _10155_/C gnd _10215_/D vdd OAI21X1
XFILL_3_BUFX2_insert930 gnd vdd FILL
XFILL_3_BUFX2_insert941 gnd vdd FILL
XFILL_2__8251_ gnd vdd FILL
XFILL_3_BUFX2_insert952 gnd vdd FILL
XFILL_3_BUFX2_insert963 gnd vdd FILL
XFILL_4__9167_ gnd vdd FILL
XFILL_3_BUFX2_insert974 gnd vdd FILL
XSFILL98840x45050 gnd vdd FILL
X_10086_ _14245_/A _7411_/CLK _7411_/R vdd _10086_/D gnd vdd DFFSR
XFILL_2__7202_ gnd vdd FILL
X_14963_ _14963_/A _14962_/Y gnd _14964_/C vdd NOR2X1
XFILL_3_BUFX2_insert985 gnd vdd FILL
XFILL_2__8182_ gnd vdd FILL
XFILL_3_BUFX2_insert996 gnd vdd FILL
XFILL_2__10540_ gnd vdd FILL
XFILL_4__8118_ gnd vdd FILL
XFILL_1__9389_ gnd vdd FILL
XSFILL99480x11050 gnd vdd FILL
XFILL_4__9098_ gnd vdd FILL
XFILL_4__11100_ gnd vdd FILL
XFILL_5__9980_ gnd vdd FILL
X_13914_ _7697_/A gnd _15445_/D vdd INVX1
XFILL_5__10651_ gnd vdd FILL
XFILL_4__12080_ gnd vdd FILL
XFILL_3__11830_ gnd vdd FILL
X_14894_ _14892_/Y _14894_/B _14718_/C _14894_/D gnd _14898_/B vdd OAI22X1
XFILL_3_BUFX2_insert1002 gnd vdd FILL
XFILL_0__11650_ gnd vdd FILL
X_13845_ _9694_/Q gnd _13846_/C vdd INVX1
XFILL_3_BUFX2_insert1013 gnd vdd FILL
XFILL_5__13370_ gnd vdd FILL
XFILL_2__12210_ gnd vdd FILL
XFILL_4__11031_ gnd vdd FILL
XFILL_2__7064_ gnd vdd FILL
XFILL_3_BUFX2_insert1024 gnd vdd FILL
XFILL_3_BUFX2_insert1035 gnd vdd FILL
XFILL_3__11761_ gnd vdd FILL
XSFILL108840x30050 gnd vdd FILL
XFILL_3_BUFX2_insert1046 gnd vdd FILL
XFILL_3_BUFX2_insert1057 gnd vdd FILL
XFILL_5__12321_ gnd vdd FILL
XFILL_5__8862_ gnd vdd FILL
XFILL_0__11581_ gnd vdd FILL
XFILL_3__13500_ gnd vdd FILL
XSFILL13800x24050 gnd vdd FILL
X_13776_ _9352_/A gnd _13776_/Y vdd INVX1
XFILL_2__12141_ gnd vdd FILL
XFILL_3_BUFX2_insert1068 gnd vdd FILL
XFILL_0__13320_ gnd vdd FILL
XFILL_3__14480_ gnd vdd FILL
X_10988_ _12210_/Y _10988_/B gnd _10988_/Y vdd NOR2X1
XFILL_0__10532_ gnd vdd FILL
XFILL_1__12871_ gnd vdd FILL
XFILL_5__7813_ gnd vdd FILL
XFILL_3__11692_ gnd vdd FILL
XFILL112120x76050 gnd vdd FILL
XFILL_5__15040_ gnd vdd FILL
X_15515_ _10647_/A gnd _15517_/B vdd INVX1
X_12727_ _12727_/A _12721_/B _12726_/Y gnd _12727_/Y vdd OAI21X1
XFILL_5__12252_ gnd vdd FILL
XFILL_3__13431_ gnd vdd FILL
XFILL_4__15770_ gnd vdd FILL
XFILL_1__14610_ gnd vdd FILL
XFILL_2__12072_ gnd vdd FILL
XFILL_4__12982_ gnd vdd FILL
XFILL_3__10643_ gnd vdd FILL
XFILL_1__11822_ gnd vdd FILL
XFILL_0__13251_ gnd vdd FILL
XSFILL64040x61050 gnd vdd FILL
XFILL_5__7744_ gnd vdd FILL
XFILL_0_BUFX2_insert820 gnd vdd FILL
XFILL_1__15590_ gnd vdd FILL
XFILL_5__11203_ gnd vdd FILL
XFILL_4__14721_ gnd vdd FILL
XSFILL114440x28050 gnd vdd FILL
X_15446_ _15446_/A _15446_/B gnd _15454_/A vdd NOR2X1
X_12658_ vdd memoryOutData[30] gnd _12659_/C vdd NAND2X1
XFILL_2__15900_ gnd vdd FILL
XFILL_4__11933_ gnd vdd FILL
XFILL_0_BUFX2_insert831 gnd vdd FILL
XFILL_5__12183_ gnd vdd FILL
XFILL_2__11023_ gnd vdd FILL
XFILL_3__16150_ gnd vdd FILL
XFILL_3__13362_ gnd vdd FILL
XFILL_0__12202_ gnd vdd FILL
XFILL_0_BUFX2_insert842 gnd vdd FILL
XFILL_3__10574_ gnd vdd FILL
XFILL_0_BUFX2_insert853 gnd vdd FILL
XFILL_1__14541_ gnd vdd FILL
XFILL_2__7966_ gnd vdd FILL
XFILL_1__11753_ gnd vdd FILL
XFILL_0_BUFX2_insert864 gnd vdd FILL
XSFILL49080x1050 gnd vdd FILL
XFILL_0__10394_ gnd vdd FILL
X_11609_ _11587_/C _11597_/A _11596_/Y gnd _11609_/Y vdd NAND3X1
XFILL_5__11134_ gnd vdd FILL
XFILL_5__7675_ gnd vdd FILL
XFILL_3__15101_ gnd vdd FILL
X_15377_ _9310_/Q gnd _15378_/A vdd INVX1
XFILL_3__12313_ gnd vdd FILL
XFILL_0_BUFX2_insert875 gnd vdd FILL
XSFILL89240x6050 gnd vdd FILL
XFILL_4__14652_ gnd vdd FILL
X_12589_ vdd memoryOutData[7] gnd _12590_/C vdd NAND2X1
XFILL_0_BUFX2_insert886 gnd vdd FILL
XFILL_2__15831_ gnd vdd FILL
XFILL_0__6981_ gnd vdd FILL
XFILL_1_BUFX2_insert1050 gnd vdd FILL
XFILL_4__11864_ gnd vdd FILL
XFILL_2__6917_ gnd vdd FILL
XFILL_3__16081_ gnd vdd FILL
XFILL_1__10704_ gnd vdd FILL
XFILL_3__13293_ gnd vdd FILL
XFILL_1__14472_ gnd vdd FILL
XFILL_0_BUFX2_insert897 gnd vdd FILL
XFILL_5__9414_ gnd vdd FILL
XFILL_0__12133_ gnd vdd FILL
XFILL_1_BUFX2_insert1061 gnd vdd FILL
XFILL_3_BUFX2_insert13 gnd vdd FILL
XFILL_1__11684_ gnd vdd FILL
XFILL_1_BUFX2_insert1072 gnd vdd FILL
XFILL_0__8720_ gnd vdd FILL
XFILL_4__13603_ gnd vdd FILL
X_14328_ _10668_/A gnd _14330_/A vdd INVX1
XFILL_3_BUFX2_insert24 gnd vdd FILL
XFILL_4__10815_ gnd vdd FILL
XFILL_3__15032_ gnd vdd FILL
XFILL_5__15942_ gnd vdd FILL
XFILL_5__11065_ gnd vdd FILL
XFILL_3_BUFX2_insert35 gnd vdd FILL
XFILL_2__9636_ gnd vdd FILL
XFILL_4__14583_ gnd vdd FILL
XFILL_1__16211_ gnd vdd FILL
XFILL_1__13423_ gnd vdd FILL
XFILL_3__12244_ gnd vdd FILL
XFILL_1__10635_ gnd vdd FILL
XFILL_3_BUFX2_insert46 gnd vdd FILL
XFILL_2__6848_ gnd vdd FILL
XFILL_2__15762_ gnd vdd FILL
XFILL_4__11795_ gnd vdd FILL
XFILL_3_BUFX2_insert57 gnd vdd FILL
XFILL_5__9345_ gnd vdd FILL
XFILL_2__12974_ gnd vdd FILL
XFILL_0__12064_ gnd vdd FILL
XFILL_5__10016_ gnd vdd FILL
XFILL_4__16322_ gnd vdd FILL
XFILL_3_BUFX2_insert68 gnd vdd FILL
X_14259_ _14593_/C _14257_/Y _13850_/B _14258_/Y gnd _14260_/B vdd OAI22X1
XFILL_0__8651_ gnd vdd FILL
XFILL_3_BUFX2_insert79 gnd vdd FILL
XFILL_4__13534_ gnd vdd FILL
XFILL_2__14713_ gnd vdd FILL
XFILL_5__15873_ gnd vdd FILL
X_7190_ _7190_/A _7250_/B _7189_/Y gnd _7264_/D vdd OAI21X1
XFILL_4__10746_ gnd vdd FILL
XFILL_3__8360_ gnd vdd FILL
XFILL_1__13354_ gnd vdd FILL
XFILL_2__11925_ gnd vdd FILL
XFILL_3__12175_ gnd vdd FILL
XFILL_1__16142_ gnd vdd FILL
XFILL_0__11015_ gnd vdd FILL
XFILL_2__15693_ gnd vdd FILL
XFILL_1__10566_ gnd vdd FILL
XFILL_5__9276_ gnd vdd FILL
XSFILL59000x50050 gnd vdd FILL
XFILL_0__7602_ gnd vdd FILL
XFILL_5__14824_ gnd vdd FILL
XFILL_4__16253_ gnd vdd FILL
XFILL_3__7311_ gnd vdd FILL
XFILL_4__13465_ gnd vdd FILL
XFILL_2__8518_ gnd vdd FILL
XFILL_1__12305_ gnd vdd FILL
XFILL_3__11126_ gnd vdd FILL
XFILL_0__8582_ gnd vdd FILL
XFILL_4__10677_ gnd vdd FILL
XFILL_2__14644_ gnd vdd FILL
XFILL_1__16073_ gnd vdd FILL
XSFILL109400x17050 gnd vdd FILL
XFILL_1__13285_ gnd vdd FILL
XFILL_5__8227_ gnd vdd FILL
XFILL_2__9498_ gnd vdd FILL
XFILL_6_CLKBUF1_insert152 gnd vdd FILL
XFILL_0__15823_ gnd vdd FILL
XFILL_2__11856_ gnd vdd FILL
XFILL_1__10497_ gnd vdd FILL
XFILL_4__15204_ gnd vdd FILL
XFILL_4__12416_ gnd vdd FILL
XFILL_4__16184_ gnd vdd FILL
XFILL_5__11967_ gnd vdd FILL
XFILL_3__15934_ gnd vdd FILL
XFILL_1__15024_ gnd vdd FILL
XSFILL49080x38050 gnd vdd FILL
XFILL_3__11057_ gnd vdd FILL
XFILL_5__14755_ gnd vdd FILL
XFILL_2__10807_ gnd vdd FILL
XFILL_2__8449_ gnd vdd FILL
XFILL_3__7242_ gnd vdd FILL
XFILL112200x56050 gnd vdd FILL
XFILL_4__13396_ gnd vdd FILL
XFILL_1__12236_ gnd vdd FILL
XFILL_2__14575_ gnd vdd FILL
XFILL_2__11787_ gnd vdd FILL
XFILL_0__15754_ gnd vdd FILL
XFILL_0__12966_ gnd vdd FILL
XFILL_5__13706_ gnd vdd FILL
XFILL_4__15135_ gnd vdd FILL
X_9900_ _9960_/Q gnd _9900_/Y vdd INVX1
XFILL_0__7464_ gnd vdd FILL
XFILL_5__10918_ gnd vdd FILL
XFILL_4__12347_ gnd vdd FILL
XFILL_3__10008_ gnd vdd FILL
XFILL_2__16314_ gnd vdd FILL
XFILL_5__11898_ gnd vdd FILL
XFILL_5__14686_ gnd vdd FILL
XFILL_2__13526_ gnd vdd FILL
XFILL_3__15865_ gnd vdd FILL
XFILL_0__14705_ gnd vdd FILL
XFILL_5__7109_ gnd vdd FILL
XFILL_0__11917_ gnd vdd FILL
XFILL_1__12167_ gnd vdd FILL
XFILL_3__7173_ gnd vdd FILL
XFILL_0__15685_ gnd vdd FILL
XFILL_6__10119_ gnd vdd FILL
XFILL_0__12897_ gnd vdd FILL
XFILL_6__8971_ gnd vdd FILL
XFILL_5__8089_ gnd vdd FILL
XFILL_6__15976_ gnd vdd FILL
XFILL_5__13637_ gnd vdd FILL
XFILL_4__15066_ gnd vdd FILL
XFILL_3__14816_ gnd vdd FILL
X_9831_ _9831_/Q _7527_/CLK _8935_/R vdd _9831_/D gnd vdd DFFSR
XFILL_4__12278_ gnd vdd FILL
XFILL_1__11118_ gnd vdd FILL
XFILL_2__16245_ gnd vdd FILL
XFILL_0__14636_ gnd vdd FILL
XFILL_2__13457_ gnd vdd FILL
XFILL_3__15796_ gnd vdd FILL
XFILL_2__10669_ gnd vdd FILL
XFILL_1__12098_ gnd vdd FILL
XFILL_0__11848_ gnd vdd FILL
XFILL_4__14017_ gnd vdd FILL
XFILL_0__9134_ gnd vdd FILL
XFILL_6__14927_ gnd vdd FILL
XFILL_5__16356_ gnd vdd FILL
XFILL_5__13568_ gnd vdd FILL
XFILL_4__11229_ gnd vdd FILL
X_6974_ _6974_/A gnd _6974_/Y vdd INVX1
XFILL_2__12408_ gnd vdd FILL
X_9762_ _9760_/Y _9741_/B _9762_/C gnd _9828_/D vdd OAI21X1
XFILL_3__14747_ gnd vdd FILL
XSFILL18600x16050 gnd vdd FILL
XFILL_1__15926_ gnd vdd FILL
XFILL_3__11959_ gnd vdd FILL
XFILL_2__16176_ gnd vdd FILL
XFILL_1__11049_ gnd vdd FILL
XFILL_0__14567_ gnd vdd FILL
XFILL_2__13388_ gnd vdd FILL
XFILL_5__15307_ gnd vdd FILL
XFILL_0__11779_ gnd vdd FILL
XSFILL28760x60050 gnd vdd FILL
X_8713_ _8714_/B _9353_/B gnd _8713_/Y vdd NAND2X1
XFILL_5__12519_ gnd vdd FILL
X_9693_ _9611_/A _9963_/CLK _9963_/R vdd _9693_/D gnd vdd DFFSR
XFILL_5__16287_ gnd vdd FILL
XFILL_2__15127_ gnd vdd FILL
XFILL_5__13499_ gnd vdd FILL
XFILL_2__12339_ gnd vdd FILL
XFILL_0__16306_ gnd vdd FILL
XFILL_3__14678_ gnd vdd FILL
XFILL_0__13518_ gnd vdd FILL
XFILL_6_BUFX2_insert336 gnd vdd FILL
XFILL_1__15857_ gnd vdd FILL
XFILL_0__14498_ gnd vdd FILL
XFILL_6_BUFX2_insert347 gnd vdd FILL
XSFILL64200x3050 gnd vdd FILL
XFILL_0__8016_ gnd vdd FILL
XFILL_5__15238_ gnd vdd FILL
X_8644_ _8688_/Q gnd _8646_/A vdd INVX1
XFILL_3__13629_ gnd vdd FILL
XFILL_6__14789_ gnd vdd FILL
XFILL_0__16237_ gnd vdd FILL
XFILL_1__14808_ gnd vdd FILL
XSFILL8680x58050 gnd vdd FILL
XFILL_2__15058_ gnd vdd FILL
XFILL_4__15968_ gnd vdd FILL
XFILL_0__13449_ gnd vdd FILL
XFILL_1__15788_ gnd vdd FILL
X_8575_ _8665_/Q gnd _8575_/Y vdd INVX1
XFILL_5__15169_ gnd vdd FILL
XFILL_2__14009_ gnd vdd FILL
XFILL_3__16348_ gnd vdd FILL
XFILL_4__14919_ gnd vdd FILL
XFILL_3__9745_ gnd vdd FILL
XFILL_4__15899_ gnd vdd FILL
XFILL_0__16168_ gnd vdd FILL
XFILL_1__14739_ gnd vdd FILL
XFILL_3__6957_ gnd vdd FILL
X_7526_ _7526_/Q _8306_/CLK _7533_/R vdd _7464_/Y gnd vdd DFFSR
XFILL_1__8760_ gnd vdd FILL
XSFILL48920x73050 gnd vdd FILL
XFILL_0__15119_ gnd vdd FILL
XFILL_3__16279_ gnd vdd FILL
XFILL_3__9676_ gnd vdd FILL
XSFILL64200x21050 gnd vdd FILL
XFILL_0__16099_ gnd vdd FILL
XFILL_3__6888_ gnd vdd FILL
XFILL_1__7711_ gnd vdd FILL
X_7457_ _7457_/A _7329_/B gnd _7458_/C vdd NAND2X1
XFILL_1__16409_ gnd vdd FILL
XFILL_4__7420_ gnd vdd FILL
XFILL_3__8627_ gnd vdd FILL
XFILL_0__9898_ gnd vdd FILL
XSFILL27960x12050 gnd vdd FILL
XFILL_0__8849_ gnd vdd FILL
X_7388_ _7388_/Q _7406_/CLK _8430_/R vdd _7388_/D gnd vdd DFFSR
XFILL_4__7351_ gnd vdd FILL
XFILL_6__8267_ gnd vdd FILL
X_9127_ _9164_/B _7079_/B gnd _9128_/C vdd NAND2X1
XFILL_3__7509_ gnd vdd FILL
XFILL_1__7573_ gnd vdd FILL
XSFILL28840x40050 gnd vdd FILL
XFILL_3_BUFX2_insert226 gnd vdd FILL
XFILL_3__8489_ gnd vdd FILL
XFILL_6__7218_ gnd vdd FILL
XFILL_3_BUFX2_insert237 gnd vdd FILL
XSFILL54120x73050 gnd vdd FILL
XFILL_3_BUFX2_insert248 gnd vdd FILL
X_9058_ _8986_/A _7382_/CLK _8674_/R vdd _9058_/D gnd vdd DFFSR
XFILL_4__9021_ gnd vdd FILL
XFILL_3_BUFX2_insert259 gnd vdd FILL
X_8009_ _8009_/A _7997_/B _8008_/Y gnd _8049_/D vdd OAI21X1
XFILL_1__9243_ gnd vdd FILL
XFILL_2_BUFX2_insert904 gnd vdd FILL
XSFILL53880x2050 gnd vdd FILL
XFILL_2_BUFX2_insert915 gnd vdd FILL
XFILL_2_BUFX2_insert926 gnd vdd FILL
XSFILL33960x31050 gnd vdd FILL
X_11960_ _11975_/A _12083_/B gnd _11961_/C vdd NAND2X1
XFILL_2_BUFX2_insert937 gnd vdd FILL
XFILL_2_BUFX2_insert948 gnd vdd FILL
XFILL_2_BUFX2_insert959 gnd vdd FILL
X_10911_ _10911_/A _10898_/Y _10911_/C gnd _10911_/Y vdd OAI21X1
XFILL_1__8125_ gnd vdd FILL
X_11891_ _11969_/A _11991_/B gnd _11891_/Y vdd NAND2X1
XFILL_4__9923_ gnd vdd FILL
X_13630_ _13628_/Y _13630_/B _14456_/C _13629_/Y gnd _13634_/A vdd OAI22X1
X_10842_ _15237_/A _9818_/CLK _8688_/R vdd _10842_/D gnd vdd DFFSR
XFILL_1__8056_ gnd vdd FILL
XSFILL13720x39050 gnd vdd FILL
XFILL_4__9854_ gnd vdd FILL
XSFILL99240x1050 gnd vdd FILL
X_13561_ _10364_/A gnd _15149_/A vdd INVX1
XSFILL23880x83050 gnd vdd FILL
XBUFX2_insert903 _10913_/Y gnd _12777_/A vdd BUFX2
X_10773_ _10773_/A _7061_/B gnd _10774_/C vdd NAND2X1
XBUFX2_insert914 _12360_/Y gnd _9094_/B vdd BUFX2
XFILL_0_BUFX2_insert105 gnd vdd FILL
X_15300_ _15300_/A gnd _15301_/A vdd INVX1
X_12512_ vdd _12512_/B gnd _12513_/C vdd NAND2X1
XSFILL13320x41050 gnd vdd FILL
XFILL_4__9785_ gnd vdd FILL
XBUFX2_insert925 _12351_/Y gnd _7293_/B vdd BUFX2
XBUFX2_insert936 _13423_/Y gnd _13857_/B vdd BUFX2
XFILL_4__6997_ gnd vdd FILL
XSFILL94200x37050 gnd vdd FILL
X_16280_ _16280_/A _16280_/B gnd _16281_/B vdd NOR2X1
XFILL_2__7820_ gnd vdd FILL
XBUFX2_insert947 _11987_/Y gnd _12073_/B vdd BUFX2
X_13492_ _13491_/Y _14744_/B gnd _13493_/C vdd NOR2X1
XBUFX2_insert958 _13361_/Y gnd _10426_/B vdd BUFX2
XBUFX2_insert969 _12417_/Y gnd _7743_/B vdd BUFX2
XFILL_4__8736_ gnd vdd FILL
X_15231_ _9818_/Q _15390_/B gnd _15241_/A vdd NAND2X1
XSFILL54200x53050 gnd vdd FILL
X_12443_ vdd _11993_/A gnd _12443_/Y vdd NAND2X1
XFILL_1__8958_ gnd vdd FILL
XFILL_2__7751_ gnd vdd FILL
XFILL_5__7460_ gnd vdd FILL
XSFILL13640x5050 gnd vdd FILL
X_15162_ _15449_/C _15162_/B _13577_/B _16314_/A gnd _15162_/Y vdd OAI22X1
X_12374_ _12419_/A _12673_/Q gnd _12375_/C vdd NAND2X1
XFILL_3__10290_ gnd vdd FILL
XFILL_2__7682_ gnd vdd FILL
XFILL_1__8889_ gnd vdd FILL
XFILL_4__7618_ gnd vdd FILL
X_14113_ _9699_/Q gnd _14115_/A vdd INVX1
X_11325_ _11324_/Y _11325_/B gnd _11325_/Y vdd NOR2X1
XFILL_4__8598_ gnd vdd FILL
XFILL_2__9421_ gnd vdd FILL
X_15093_ _13485_/A _15357_/B _16294_/C _13497_/A gnd _15093_/Y vdd AOI22X1
XFILL_4__11580_ gnd vdd FILL
XFILL_1__10420_ gnd vdd FILL
XFILL_5__9130_ gnd vdd FILL
XSFILL18840x72050 gnd vdd FILL
XFILL_4__7549_ gnd vdd FILL
X_14044_ _7194_/A gnd _14044_/Y vdd INVX1
X_11256_ _11247_/Y _11253_/Y _11256_/C gnd _11256_/Y vdd OAI21X1
XFILL_4__10531_ gnd vdd FILL
XFILL_5__12870_ gnd vdd FILL
XFILL_2__9352_ gnd vdd FILL
XFILL_2__11710_ gnd vdd FILL
XSFILL108840x25050 gnd vdd FILL
XSFILL99320x70050 gnd vdd FILL
X_10207_ _13892_/A _7647_/CLK _9823_/R vdd _10207_/D gnd vdd DFFSR
XFILL_5__11821_ gnd vdd FILL
XFILL_4__13250_ gnd vdd FILL
X_11187_ _12318_/Y gnd _11188_/B vdd INVX1
XSFILL59000x4050 gnd vdd FILL
XFILL_4__9219_ gnd vdd FILL
XFILL_5__8012_ gnd vdd FILL
XFILL_3__13980_ gnd vdd FILL
XFILL_2__11641_ gnd vdd FILL
XFILL_2__9283_ gnd vdd FILL
XFILL_1__10282_ gnd vdd FILL
X_10138_ _10138_/A gnd _10140_/A vdd INVX1
XFILL_3_BUFX2_insert760 gnd vdd FILL
XSFILL23160x44050 gnd vdd FILL
XFILL_4__12201_ gnd vdd FILL
XFILL_5__14540_ gnd vdd FILL
XFILL_3_BUFX2_insert771 gnd vdd FILL
XFILL_5__11752_ gnd vdd FILL
X_15995_ _8891_/A _16037_/B _15995_/C gnd _15995_/Y vdd NAND3X1
XFILL_1__12021_ gnd vdd FILL
XSFILL109720x53050 gnd vdd FILL
XFILL_3_BUFX2_insert782 gnd vdd FILL
XFILL_2__8234_ gnd vdd FILL
XFILL_4__10393_ gnd vdd FILL
XFILL_2__14360_ gnd vdd FILL
XFILL112280x30050 gnd vdd FILL
XFILL_3_BUFX2_insert793 gnd vdd FILL
XFILL_2__11572_ gnd vdd FILL
XFILL_0__12751_ gnd vdd FILL
XSFILL64840x75050 gnd vdd FILL
XSFILL64040x56050 gnd vdd FILL
XFILL_5__10703_ gnd vdd FILL
XFILL_5__14471_ gnd vdd FILL
X_10069_ _10067_/Y _9993_/A _10069_/C gnd _10101_/D vdd OAI21X1
X_14946_ _14946_/A _14946_/B _14945_/Y _13879_/B gnd _14946_/Y vdd OAI22X1
XFILL_4__12132_ gnd vdd FILL
XFILL_2__13311_ gnd vdd FILL
XFILL_3__15650_ gnd vdd FILL
XFILL_2__10523_ gnd vdd FILL
XFILL_5__11683_ gnd vdd FILL
XFILL_0__11702_ gnd vdd FILL
XFILL_3__12862_ gnd vdd FILL
XFILL_2__14291_ gnd vdd FILL
XFILL_0__15470_ gnd vdd FILL
XFILL_5__16210_ gnd vdd FILL
XFILL_5__13422_ gnd vdd FILL
XFILL_0__7180_ gnd vdd FILL
XFILL_3__14601_ gnd vdd FILL
XFILL_5__10634_ gnd vdd FILL
XFILL_6__15761_ gnd vdd FILL
XFILL_2__7116_ gnd vdd FILL
X_14877_ _14557_/C _8269_/A _10867_/Q _14877_/D gnd _14877_/Y vdd AOI22X1
XFILL_2__16030_ gnd vdd FILL
XFILL_4__12063_ gnd vdd FILL
XFILL_3__11813_ gnd vdd FILL
XFILL_2__13242_ gnd vdd FILL
XFILL_0__14421_ gnd vdd FILL
XFILL_3__15581_ gnd vdd FILL
XSFILL43880x14050 gnd vdd FILL
XSFILL3480x63050 gnd vdd FILL
XFILL_2__8096_ gnd vdd FILL
XFILL_0__11633_ gnd vdd FILL
XFILL_5__8914_ gnd vdd FILL
XFILL_1__13972_ gnd vdd FILL
X_13828_ _7947_/A gnd _13828_/Y vdd INVX1
XFILL_5__13353_ gnd vdd FILL
XFILL_5__9894_ gnd vdd FILL
XFILL_4__11014_ gnd vdd FILL
XFILL_5__16141_ gnd vdd FILL
XFILL_3__14532_ gnd vdd FILL
XFILL_5__10565_ gnd vdd FILL
XFILL_1__15711_ gnd vdd FILL
XFILL_2__13173_ gnd vdd FILL
XFILL_2__7047_ gnd vdd FILL
XFILL_3__11744_ gnd vdd FILL
XFILL_0__14352_ gnd vdd FILL
XFILL_2__10385_ gnd vdd FILL
XFILL_5__8845_ gnd vdd FILL
XFILL_5__12304_ gnd vdd FILL
XFILL_0__11564_ gnd vdd FILL
XSFILL84200x69050 gnd vdd FILL
XFILL_5__16072_ gnd vdd FILL
XFILL_5__13284_ gnd vdd FILL
X_13759_ _13759_/A _13758_/Y gnd _13759_/Y vdd NOR2X1
XFILL_4__15822_ gnd vdd FILL
XFILL_6__11855_ gnd vdd FILL
XFILL_5__10496_ gnd vdd FILL
XFILL_0__13303_ gnd vdd FILL
XFILL_3__14463_ gnd vdd FILL
XFILL_2__12124_ gnd vdd FILL
XFILL_1__15642_ gnd vdd FILL
XFILL_3__11675_ gnd vdd FILL
XFILL_0__10515_ gnd vdd FILL
XFILL_3__7860_ gnd vdd FILL
XFILL_1__12854_ gnd vdd FILL
XFILL_0__14283_ gnd vdd FILL
XFILL_6__10806_ gnd vdd FILL
XFILL_3__16202_ gnd vdd FILL
XFILL_5__15023_ gnd vdd FILL
XSFILL59000x45050 gnd vdd FILL
XFILL_5__12235_ gnd vdd FILL
XFILL_0__11495_ gnd vdd FILL
XFILL_5__8776_ gnd vdd FILL
XFILL_6__14574_ gnd vdd FILL
XFILL_3__13414_ gnd vdd FILL
XFILL_0__16022_ gnd vdd FILL
XFILL_3__10626_ gnd vdd FILL
XFILL_4__12965_ gnd vdd FILL
XFILL_2__12055_ gnd vdd FILL
XFILL_4__15753_ gnd vdd FILL
XFILL_0__13234_ gnd vdd FILL
XSFILL99400x50050 gnd vdd FILL
XFILL_3__14394_ gnd vdd FILL
XFILL_1__11805_ gnd vdd FILL
XFILL_1__12785_ gnd vdd FILL
XFILL_0__10446_ gnd vdd FILL
XFILL_2__8998_ gnd vdd FILL
XFILL_1__15573_ gnd vdd FILL
XFILL_5__7727_ gnd vdd FILL
XFILL_0_BUFX2_insert650 gnd vdd FILL
X_15429_ _15841_/C _13924_/D _15429_/C _15813_/C gnd _15432_/B vdd OAI22X1
X_8360_ _8360_/A _8360_/B _8359_/Y gnd _8422_/D vdd OAI21X1
XFILL_4__11916_ gnd vdd FILL
XFILL_4__14704_ gnd vdd FILL
XFILL_0_BUFX2_insert661 gnd vdd FILL
XFILL_5__12166_ gnd vdd FILL
XFILL_2__11006_ gnd vdd FILL
XFILL_3__16133_ gnd vdd FILL
XFILL_3__13345_ gnd vdd FILL
XFILL_4__15684_ gnd vdd FILL
XFILL_0_BUFX2_insert672 gnd vdd FILL
XFILL111720x44050 gnd vdd FILL
XFILL_3__9530_ gnd vdd FILL
XFILL_2__7949_ gnd vdd FILL
XFILL_4__12896_ gnd vdd FILL
XFILL_3__10557_ gnd vdd FILL
XFILL_1__14524_ gnd vdd FILL
XFILL_0_BUFX2_insert683 gnd vdd FILL
XFILL_0__13165_ gnd vdd FILL
XFILL_0_BUFX2_insert694 gnd vdd FILL
XFILL_1__11736_ gnd vdd FILL
X_7311_ _7297_/B _8719_/B gnd _7311_/Y vdd NAND2X1
XFILL_0__10377_ gnd vdd FILL
XSFILL89480x38050 gnd vdd FILL
XFILL_5__11117_ gnd vdd FILL
XFILL_0__9752_ gnd vdd FILL
XFILL112360x10050 gnd vdd FILL
XFILL_4__14635_ gnd vdd FILL
XFILL_5__12097_ gnd vdd FILL
XSFILL64120x36050 gnd vdd FILL
XFILL_2__15814_ gnd vdd FILL
X_8291_ _8221_/A _7651_/CLK _9711_/R vdd _8223_/Y gnd vdd DFFSR
XFILL_0__6964_ gnd vdd FILL
XFILL_3__16064_ gnd vdd FILL
XFILL_4__11847_ gnd vdd FILL
XFILL_3__13276_ gnd vdd FILL
XFILL_0__12116_ gnd vdd FILL
XFILL_1__14455_ gnd vdd FILL
XFILL_3__10488_ gnd vdd FILL
XFILL_1__11667_ gnd vdd FILL
XFILL_0__8703_ gnd vdd FILL
XFILL_0__13096_ gnd vdd FILL
X_7242_ _7282_/Q gnd _7242_/Y vdd INVX1
XFILL_5__15925_ gnd vdd FILL
XFILL_5__7589_ gnd vdd FILL
XFILL_3__15015_ gnd vdd FILL
XFILL_5__11048_ gnd vdd FILL
XFILL_4__14566_ gnd vdd FILL
XFILL_0__9683_ gnd vdd FILL
XFILL_3__12227_ gnd vdd FILL
XFILL_2__9619_ gnd vdd FILL
XFILL_1__13406_ gnd vdd FILL
XFILL_1__10618_ gnd vdd FILL
XFILL_0__6895_ gnd vdd FILL
XFILL_4__11778_ gnd vdd FILL
XFILL_2__15745_ gnd vdd FILL
XFILL_0__12047_ gnd vdd FILL
XFILL_3__9392_ gnd vdd FILL
XFILL_1__14386_ gnd vdd FILL
XFILL_2__12957_ gnd vdd FILL
XFILL_1__11598_ gnd vdd FILL
XFILL_0__8634_ gnd vdd FILL
XFILL_4__16305_ gnd vdd FILL
XFILL_4__13517_ gnd vdd FILL
XSFILL3560x43050 gnd vdd FILL
XFILL_5__15856_ gnd vdd FILL
X_7173_ _7173_/A gnd _7173_/Y vdd INVX1
XFILL_4__14497_ gnd vdd FILL
XFILL_2__11908_ gnd vdd FILL
XFILL_3__12158_ gnd vdd FILL
XFILL_3__8343_ gnd vdd FILL
XFILL_1__16125_ gnd vdd FILL
XFILL_1__13337_ gnd vdd FILL
XFILL_1__10549_ gnd vdd FILL
XFILL_2__15676_ gnd vdd FILL
XFILL_2__12888_ gnd vdd FILL
XFILL_5__9259_ gnd vdd FILL
XFILL_5__14807_ gnd vdd FILL
XFILL_4__16236_ gnd vdd FILL
XSFILL28760x55050 gnd vdd FILL
XFILL_4__13448_ gnd vdd FILL
XFILL_3__11109_ gnd vdd FILL
XFILL_2__14627_ gnd vdd FILL
XFILL_5__15787_ gnd vdd FILL
XFILL_1__13268_ gnd vdd FILL
XFILL_3__12089_ gnd vdd FILL
XFILL_5__12999_ gnd vdd FILL
XFILL_0__15806_ gnd vdd FILL
XFILL_1__16056_ gnd vdd FILL
XFILL_3__8274_ gnd vdd FILL
XFILL_2__11839_ gnd vdd FILL
XFILL_0__13998_ gnd vdd FILL
XFILL_4__16167_ gnd vdd FILL
XFILL_5__14738_ gnd vdd FILL
XFILL_3__15917_ gnd vdd FILL
XFILL_1__15007_ gnd vdd FILL
XFILL_3__7225_ gnd vdd FILL
XFILL_4__13379_ gnd vdd FILL
XFILL_0__8496_ gnd vdd FILL
XFILL_1__12219_ gnd vdd FILL
XFILL_2__14558_ gnd vdd FILL
XFILL_0__15737_ gnd vdd FILL
XFILL_4__15118_ gnd vdd FILL
XFILL_0__7447_ gnd vdd FILL
XSFILL33880x46050 gnd vdd FILL
XFILL_4__16098_ gnd vdd FILL
XFILL_5__14669_ gnd vdd FILL
XFILL_2__13509_ gnd vdd FILL
XFILL_3__15848_ gnd vdd FILL
XFILL_2__14489_ gnd vdd FILL
XFILL_5__16408_ gnd vdd FILL
XFILL_0__15668_ gnd vdd FILL
X_9814_ _9718_/A _8022_/CLK _7644_/R vdd _9814_/D gnd vdd DFFSR
XFILL_4__15049_ gnd vdd FILL
XFILL_2__16228_ gnd vdd FILL
XFILL_0__7378_ gnd vdd FILL
XFILL_3__15779_ gnd vdd FILL
XFILL_0__14619_ gnd vdd FILL
XFILL_3__7087_ gnd vdd FILL
XFILL_0__9117_ gnd vdd FILL
XFILL_5__16339_ gnd vdd FILL
XFILL_0__15599_ gnd vdd FILL
X_6957_ _6948_/A _6957_/B gnd _6958_/C vdd NAND2X1
X_9745_ _9745_/A gnd _9745_/Y vdd INVX1
XFILL_1__15909_ gnd vdd FILL
XFILL_4__6920_ gnd vdd FILL
XFILL_2__16159_ gnd vdd FILL
XFILL_1__9930_ gnd vdd FILL
X_9676_ _9676_/A _9675_/A _9676_/C gnd _9676_/Y vdd OAI21X1
X_6888_ _6888_/A gnd memoryWriteData[18] vdd BUFX2
XSFILL89400x82050 gnd vdd FILL
XFILL_4__6851_ gnd vdd FILL
XSFILL3640x23050 gnd vdd FILL
XFILL_5_BUFX2_insert800 gnd vdd FILL
XSFILL93640x45050 gnd vdd FILL
XFILL_1__9861_ gnd vdd FILL
X_8627_ _8657_/A _8243_/B gnd _8628_/C vdd NAND2X1
XFILL_5_BUFX2_insert811 gnd vdd FILL
XFILL_3__7989_ gnd vdd FILL
XSFILL28840x35050 gnd vdd FILL
XFILL_5_BUFX2_insert822 gnd vdd FILL
XFILL_5_BUFX2_insert833 gnd vdd FILL
XSFILL94280x11050 gnd vdd FILL
XSFILL54120x68050 gnd vdd FILL
XFILL_5_BUFX2_insert844 gnd vdd FILL
XFILL_1__9792_ gnd vdd FILL
XFILL_3__9728_ gnd vdd FILL
X_8558_ _8558_/Q _7406_/CLK _8430_/R vdd _8512_/Y gnd vdd DFFSR
XFILL_4__8521_ gnd vdd FILL
XFILL_5_BUFX2_insert855 gnd vdd FILL
XBUFX2_insert1030 _13333_/Y gnd _9282_/A vdd BUFX2
XFILL_5_BUFX2_insert866 gnd vdd FILL
XFILL_5_BUFX2_insert877 gnd vdd FILL
XBUFX2_insert1041 _13297_/Y gnd _7672_/B vdd BUFX2
XFILL_1__8743_ gnd vdd FILL
X_7509_ _7507_/Y _7416_/B _7508_/Y gnd _7509_/Y vdd OAI21X1
XBUFX2_insert1052 _12806_/Q gnd _12297_/D vdd BUFX2
XFILL_5_BUFX2_insert888 gnd vdd FILL
XFILL_5_BUFX2_insert899 gnd vdd FILL
X_8489_ _8551_/Q gnd _8489_/Y vdd INVX1
XBUFX2_insert1063 _14992_/Y gnd _15802_/A vdd BUFX2
XFILL_3__9659_ gnd vdd FILL
XFILL_4__8452_ gnd vdd FILL
XBUFX2_insert1085 rst gnd BUFX2_insert559/A vdd BUFX2
XSFILL33960x26050 gnd vdd FILL
X_11110_ _11108_/Y _11109_/Y gnd _11110_/Y vdd NOR2X1
XFILL_4__8383_ gnd vdd FILL
X_12090_ _12090_/A _12090_/B _12089_/Y gnd _13155_/B vdd NAND3X1
XFILL_1__7625_ gnd vdd FILL
XFILL_4__7334_ gnd vdd FILL
X_11041_ _11041_/A _11021_/Y _11041_/C gnd _11041_/Y vdd OAI21X1
XFILL_1__7556_ gnd vdd FILL
XSFILL23880x78050 gnd vdd FILL
XSFILL23080x59050 gnd vdd FILL
XFILL_4__9004_ gnd vdd FILL
XFILL_1__7487_ gnd vdd FILL
XFILL_2_BUFX2_insert701 gnd vdd FILL
XSFILL109640x68050 gnd vdd FILL
X_14800_ _14796_/Y _14799_/Y gnd _14800_/Y vdd NOR2X1
XFILL_2_BUFX2_insert712 gnd vdd FILL
XFILL_4__7196_ gnd vdd FILL
XFILL_1__9226_ gnd vdd FILL
XFILL_2_BUFX2_insert723 gnd vdd FILL
X_15780_ _16225_/C _14349_/Y _15558_/D _14346_/Y gnd _15784_/B vdd OAI22X1
XFILL_2_BUFX2_insert734 gnd vdd FILL
X_12992_ _12990_/Y vdd _12992_/C gnd _13060_/D vdd OAI21X1
XFILL_2_BUFX2_insert745 gnd vdd FILL
XSFILL28920x15050 gnd vdd FILL
X_14731_ _16105_/A gnd _14731_/Y vdd INVX1
XFILL_2_BUFX2_insert756 gnd vdd FILL
XFILL_2_BUFX2_insert767 gnd vdd FILL
X_11943_ _11941_/Y _11895_/B _11943_/C gnd _6856_/A vdd OAI21X1
XFILL_2_BUFX2_insert778 gnd vdd FILL
XFILL_1__9157_ gnd vdd FILL
XFILL_2_BUFX2_insert789 gnd vdd FILL
XSFILL79160x52050 gnd vdd FILL
XFILL_5__6960_ gnd vdd FILL
XFILL_1__8108_ gnd vdd FILL
X_14662_ _16079_/A _14901_/B _14894_/B _14662_/D gnd _14666_/B vdd OAI22X1
X_11874_ _11874_/A _11874_/B _11873_/Y gnd _13305_/A vdd OAI21X1
XFILL_1__9088_ gnd vdd FILL
X_16401_ _16401_/A gnd _16401_/C gnd _16443_/D vdd OAI21X1
XFILL_4__9906_ gnd vdd FILL
X_13613_ _8409_/Q gnd _13613_/Y vdd INVX1
XFILL_5__6891_ gnd vdd FILL
X_10825_ _10823_/Y _10797_/A _10825_/C gnd _10865_/D vdd OAI21X1
XSFILL83640x77050 gnd vdd FILL
X_14593_ _14592_/Y _13614_/C _14593_/C _14591_/Y gnd _14594_/A vdd OAI22X1
XFILL_2__10170_ gnd vdd FILL
XFILL_5__8630_ gnd vdd FILL
XBUFX2_insert700 _12420_/Y gnd _6978_/B vdd BUFX2
XSFILL18840x67050 gnd vdd FILL
X_16332_ _16332_/A gnd _16332_/C gnd _16332_/Y vdd OAI21X1
XBUFX2_insert711 _12816_/Q gnd _14986_/A vdd BUFX2
XSFILL84280x43050 gnd vdd FILL
XFILL_6__11640_ gnd vdd FILL
XBUFX2_insert722 _13352_/Y gnd _10106_/A vdd BUFX2
X_13544_ _13544_/A _13544_/B _13540_/Y gnd _13560_/B vdd NAND3X1
X_10756_ _10756_/A _10792_/B _10756_/C gnd _10842_/D vdd OAI21X1
XFILL_5__10281_ gnd vdd FILL
XBUFX2_insert733 _15020_/Y gnd _15631_/B vdd BUFX2
XFILL_0__10300_ gnd vdd FILL
XFILL_2__8852_ gnd vdd FILL
XFILL_3__11460_ gnd vdd FILL
XBUFX2_insert744 _15055_/Y gnd _15378_/B vdd BUFX2
XFILL_4__9768_ gnd vdd FILL
XFILL_5__12020_ gnd vdd FILL
XBUFX2_insert755 _12213_/Y gnd _12224_/C vdd BUFX2
XFILL_0__11280_ gnd vdd FILL
XBUFX2_insert766 _12393_/Y gnd _9383_/B vdd BUFX2
X_16263_ _16263_/A _14983_/A _15715_/C gnd _16266_/A vdd NOR3X1
XFILL_4__12750_ gnd vdd FILL
XSFILL99320x65050 gnd vdd FILL
XBUFX2_insert777 _10911_/Y gnd _12137_/A vdd BUFX2
X_13475_ _13475_/A _13451_/Y gnd _13476_/B vdd NOR2X1
XFILL_3__10411_ gnd vdd FILL
XFILL_2__7803_ gnd vdd FILL
X_10687_ _10661_/B _7743_/B gnd _10688_/C vdd NAND2X1
XBUFX2_insert788 _13486_/Y gnd _13853_/C vdd BUFX2
XFILL_4__8719_ gnd vdd FILL
XFILL_1__12570_ gnd vdd FILL
XFILL_2__8783_ gnd vdd FILL
XFILL_0__10231_ gnd vdd FILL
XFILL_3__11391_ gnd vdd FILL
XBUFX2_insert799 _13334_/Y gnd _9359_/A vdd BUFX2
X_15214_ _13653_/Y _16002_/A gnd _15215_/C vdd NOR2X1
XSFILL23960x58050 gnd vdd FILL
XFILL_6__10522_ gnd vdd FILL
X_12426_ _12424_/Y _12395_/A _12426_/C gnd _12426_/Y vdd OAI21X1
XFILL_5__8492_ gnd vdd FILL
XFILL_4__11701_ gnd vdd FILL
X_16194_ _15972_/C _16194_/B _16194_/C gnd _16194_/Y vdd OAI21X1
XFILL_3__13130_ gnd vdd FILL
XFILL_2__7734_ gnd vdd FILL
XFILL_1__11521_ gnd vdd FILL
XFILL_2__13860_ gnd vdd FILL
XFILL112280x25050 gnd vdd FILL
XFILL_0__10162_ gnd vdd FILL
XFILL_5__7443_ gnd vdd FILL
XFILL_4__14420_ gnd vdd FILL
X_15145_ _16141_/A _15145_/B _16141_/C gnd _15166_/B vdd NOR3X1
XFILL_1_CLKBUF1_insert160 gnd vdd FILL
X_12357_ _12355_/Y _12371_/A _12357_/C gnd _12357_/Y vdd OAI21X1
XFILL_4__11632_ gnd vdd FILL
XFILL_1__14240_ gnd vdd FILL
XFILL_5__13971_ gnd vdd FILL
XSFILL24040x67050 gnd vdd FILL
XFILL_3__10273_ gnd vdd FILL
XFILL_1_CLKBUF1_insert171 gnd vdd FILL
XFILL_1__11452_ gnd vdd FILL
XFILL_2__13791_ gnd vdd FILL
XFILL_1_CLKBUF1_insert182 gnd vdd FILL
XFILL_1_CLKBUF1_insert193 gnd vdd FILL
XFILL_5__15710_ gnd vdd FILL
XFILL_5__7374_ gnd vdd FILL
XFILL_0__14970_ gnd vdd FILL
X_11308_ _11297_/Y _11597_/A _11308_/C gnd _11550_/C vdd OAI21X1
XFILL_2__9404_ gnd vdd FILL
X_15076_ _15076_/A _15075_/Y _15076_/C gnd _15077_/B vdd NOR3X1
XFILL_3__12012_ gnd vdd FILL
XFILL_4__14351_ gnd vdd FILL
XFILL_1__10403_ gnd vdd FILL
XFILL_2__15530_ gnd vdd FILL
XFILL_2_BUFX2_insert3 gnd vdd FILL
X_12288_ _12224_/A _12308_/B _12224_/C gnd _12290_/B vdd NAND3X1
XFILL_4__11563_ gnd vdd FILL
XFILL_2__12742_ gnd vdd FILL
XFILL_1__14171_ gnd vdd FILL
XFILL_5__9113_ gnd vdd FILL
XSFILL79240x32050 gnd vdd FILL
XSFILL3480x58050 gnd vdd FILL
XFILL_2__7596_ gnd vdd FILL
XFILL_0__13921_ gnd vdd FILL
XFILL_1__11383_ gnd vdd FILL
XFILL_4__13302_ gnd vdd FILL
X_14027_ _14025_/Y _13630_/B _14640_/C _14026_/Y gnd _14027_/Y vdd OAI22X1
XFILL_5__15641_ gnd vdd FILL
XFILL_4__10514_ gnd vdd FILL
X_11239_ _12218_/Y _12117_/Y gnd _11239_/Y vdd NAND2X1
XFILL_2__9335_ gnd vdd FILL
XFILL_1__13122_ gnd vdd FILL
XFILL_5__12853_ gnd vdd FILL
XFILL_4__14282_ gnd vdd FILL
XSFILL69160x5050 gnd vdd FILL
XFILL_4__11494_ gnd vdd FILL
XFILL_2__15461_ gnd vdd FILL
XFILL_0__13852_ gnd vdd FILL
XFILL_5__9044_ gnd vdd FILL
XFILL_4__16021_ gnd vdd FILL
XSFILL114440x41050 gnd vdd FILL
XFILL_4__13233_ gnd vdd FILL
XFILL_0__8350_ gnd vdd FILL
XFILL_5__11804_ gnd vdd FILL
XFILL_4__10445_ gnd vdd FILL
XFILL_5__15572_ gnd vdd FILL
XFILL_2__14412_ gnd vdd FILL
XFILL_5__12784_ gnd vdd FILL
XFILL_2__9266_ gnd vdd FILL
XFILL_2__11624_ gnd vdd FILL
XFILL_3__13963_ gnd vdd FILL
XFILL_2__15392_ gnd vdd FILL
XFILL_1__10265_ gnd vdd FILL
XSFILL84360x23050 gnd vdd FILL
XFILL_0__13783_ gnd vdd FILL
XFILL_3_BUFX2_insert590 gnd vdd FILL
XFILL_0__7301_ gnd vdd FILL
XFILL_5__14523_ gnd vdd FILL
XFILL_0__10995_ gnd vdd FILL
X_15978_ _8379_/A _15978_/B _15978_/C _8507_/A gnd _15978_/Y vdd AOI22X1
XFILL_3__15702_ gnd vdd FILL
XFILL_4__13164_ gnd vdd FILL
XFILL_1__12004_ gnd vdd FILL
XFILL_2__8217_ gnd vdd FILL
XFILL_3__12914_ gnd vdd FILL
XFILL_5__11735_ gnd vdd FILL
XFILL_4__10376_ gnd vdd FILL
XFILL_2__14343_ gnd vdd FILL
XFILL_0__12734_ gnd vdd FILL
XFILL_0__15522_ gnd vdd FILL
XFILL_3__13894_ gnd vdd FILL
XFILL_2__11555_ gnd vdd FILL
XFILL_1__10196_ gnd vdd FILL
XFILL_0__7232_ gnd vdd FILL
XFILL_4__12115_ gnd vdd FILL
X_14929_ _14929_/A _14929_/B _14402_/C gnd _13042_/B vdd AOI21X1
XFILL_5__14454_ gnd vdd FILL
XFILL_3__15633_ gnd vdd FILL
XFILL_5__11666_ gnd vdd FILL
X_7860_ _7860_/A _7878_/B _7860_/C gnd _7914_/D vdd OAI21X1
XFILL_3__12845_ gnd vdd FILL
XFILL_2__10506_ gnd vdd FILL
XFILL_4__13095_ gnd vdd FILL
XFILL_2__8148_ gnd vdd FILL
XFILL_2__14274_ gnd vdd FILL
XFILL_2__11486_ gnd vdd FILL
XFILL_0__15453_ gnd vdd FILL
XFILL_5__13405_ gnd vdd FILL
XSFILL109800x28050 gnd vdd FILL
XFILL_5__10617_ gnd vdd FILL
XFILL_0__7163_ gnd vdd FILL
XFILL_2__16013_ gnd vdd FILL
XFILL_4__12046_ gnd vdd FILL
XFILL_2__13225_ gnd vdd FILL
XFILL_3__15564_ gnd vdd FILL
XFILL_5__14385_ gnd vdd FILL
X_7791_ _7791_/Q _7791_/CLK _9711_/R vdd _7791_/D gnd vdd DFFSR
XFILL_5__11597_ gnd vdd FILL
XFILL_3__8961_ gnd vdd FILL
XFILL_2__8079_ gnd vdd FILL
XFILL_3__12776_ gnd vdd FILL
XFILL_2__10437_ gnd vdd FILL
XFILL_6_BUFX2_insert50 gnd vdd FILL
XFILL_0__11616_ gnd vdd FILL
XFILL_0__14404_ gnd vdd FILL
XFILL_0__15384_ gnd vdd FILL
XFILL_1__13955_ gnd vdd FILL
XSFILL74280x75050 gnd vdd FILL
XFILL_0__12596_ gnd vdd FILL
XFILL_5__16124_ gnd vdd FILL
XFILL_5__13336_ gnd vdd FILL
XFILL_0__7094_ gnd vdd FILL
XFILL_3__14515_ gnd vdd FILL
X_9530_ _9530_/A _9529_/A _9530_/C gnd _9530_/Y vdd OAI21X1
XFILL_5__9877_ gnd vdd FILL
XFILL_5__10548_ gnd vdd FILL
XFILL_6__12887_ gnd vdd FILL
XFILL_3__11727_ gnd vdd FILL
XFILL_2__10368_ gnd vdd FILL
XFILL_2__13156_ gnd vdd FILL
XFILL_0__14335_ gnd vdd FILL
XFILL_1__12906_ gnd vdd FILL
XFILL_3__15495_ gnd vdd FILL
XFILL_3__8892_ gnd vdd FILL
XFILL_6__7621_ gnd vdd FILL
XFILL_0__11547_ gnd vdd FILL
XFILL_1__13886_ gnd vdd FILL
XFILL_6__14626_ gnd vdd FILL
XFILL_5__8828_ gnd vdd FILL
XSFILL79320x12050 gnd vdd FILL
XFILL_5__13267_ gnd vdd FILL
X_9461_ _9461_/Q _7010_/CLK _7413_/R vdd _9429_/Y gnd vdd DFFSR
XFILL_4__15805_ gnd vdd FILL
XFILL_5__16055_ gnd vdd FILL
XFILL_2__12107_ gnd vdd FILL
XSFILL3560x38050 gnd vdd FILL
XFILL_3__14446_ gnd vdd FILL
XFILL_3__7843_ gnd vdd FILL
XFILL_1__15625_ gnd vdd FILL
XFILL_5_BUFX2_insert107 gnd vdd FILL
XFILL_3__11658_ gnd vdd FILL
XFILL_2__10299_ gnd vdd FILL
XFILL_1__12837_ gnd vdd FILL
XFILL_2__13087_ gnd vdd FILL
XFILL_4__13997_ gnd vdd FILL
XFILL_0__14266_ gnd vdd FILL
XFILL_5__8759_ gnd vdd FILL
XFILL_5__15006_ gnd vdd FILL
XFILL_5__12218_ gnd vdd FILL
XFILL_0__11478_ gnd vdd FILL
X_8412_ _8328_/A _7534_/CLK _8430_/R vdd _8412_/D gnd vdd DFFSR
X_9392_ _9401_/A _8496_/B gnd _9393_/C vdd NAND2X1
XFILL_4__15736_ gnd vdd FILL
XFILL_0__13217_ gnd vdd FILL
XFILL_0__16005_ gnd vdd FILL
XFILL_2__12038_ gnd vdd FILL
XFILL_3__14377_ gnd vdd FILL
XFILL_0__10429_ gnd vdd FILL
XFILL_1__15556_ gnd vdd FILL
XFILL_3__11589_ gnd vdd FILL
XFILL_1__12768_ gnd vdd FILL
XFILL_0__14197_ gnd vdd FILL
XFILL_0__9804_ gnd vdd FILL
XFILL_0_BUFX2_insert480 gnd vdd FILL
XFILL_3__16116_ gnd vdd FILL
X_8343_ _8343_/A gnd _8343_/Y vdd INVX1
XFILL_5__12149_ gnd vdd FILL
XFILL_0_BUFX2_insert491 gnd vdd FILL
XFILL_3__13328_ gnd vdd FILL
XFILL_3__9513_ gnd vdd FILL
XFILL_4__15667_ gnd vdd FILL
XFILL_0__7996_ gnd vdd FILL
XFILL_1__14507_ gnd vdd FILL
XFILL_4_BUFX2_insert807 gnd vdd FILL
XFILL_4__12879_ gnd vdd FILL
XFILL_0__13148_ gnd vdd FILL
XFILL_1__11719_ gnd vdd FILL
XFILL_6__16227_ gnd vdd FILL
XFILL_4_BUFX2_insert818 gnd vdd FILL
XFILL_1__15487_ gnd vdd FILL
XFILL_1__12699_ gnd vdd FILL
XFILL_4_BUFX2_insert829 gnd vdd FILL
XFILL_6__13439_ gnd vdd FILL
XFILL_0__9735_ gnd vdd FILL
XFILL_4__14618_ gnd vdd FILL
XFILL_0__6947_ gnd vdd FILL
XSFILL3560x7050 gnd vdd FILL
XFILL_3__16047_ gnd vdd FILL
X_8274_ _8274_/A _8216_/A _8273_/Y gnd _8274_/Y vdd OAI21X1
XFILL_3__13259_ gnd vdd FILL
XSFILL69240x64050 gnd vdd FILL
XFILL_4__15598_ gnd vdd FILL
XFILL_1__14438_ gnd vdd FILL
XFILL_0__13079_ gnd vdd FILL
XFILL_2__13989_ gnd vdd FILL
XFILL_5__15908_ gnd vdd FILL
X_7225_ _7202_/B _9017_/B gnd _7225_/Y vdd NAND2X1
XFILL_0__9666_ gnd vdd FILL
XFILL_2__15728_ gnd vdd FILL
XFILL_4__14549_ gnd vdd FILL
XFILL_0__6878_ gnd vdd FILL
XFILL_3__9375_ gnd vdd FILL
XSFILL104440x73050 gnd vdd FILL
XFILL_1__14369_ gnd vdd FILL
XFILL_0__8617_ gnd vdd FILL
XFILL_6__16089_ gnd vdd FILL
XFILL_5__15839_ gnd vdd FILL
X_7156_ _7156_/Q _7156_/CLK _7775_/R vdd _7156_/D gnd vdd DFFSR
XSFILL8680x71050 gnd vdd FILL
XFILL_1__8390_ gnd vdd FILL
XFILL_1__16108_ gnd vdd FILL
XFILL_0__9597_ gnd vdd FILL
XFILL_3__8326_ gnd vdd FILL
XSFILL23720x20050 gnd vdd FILL
XFILL_2__15659_ gnd vdd FILL
XCLKBUF1_insert170 CLKBUF1_insert150/A gnd _7537_/CLK vdd CLKBUF1
XCLKBUF1_insert181 CLKBUF1_insert187/A gnd _12809_/CLK vdd CLKBUF1
XFILL_4__16219_ gnd vdd FILL
XFILL_1__7341_ gnd vdd FILL
XCLKBUF1_insert192 CLKBUF1_insert192/A gnd _7790_/CLK vdd CLKBUF1
X_7087_ _7145_/Q gnd _7087_/Y vdd INVX1
XFILL_1__16039_ gnd vdd FILL
XFILL_4__7050_ gnd vdd FILL
XFILL_3__8257_ gnd vdd FILL
XSFILL3640x18050 gnd vdd FILL
XFILL_3__7208_ gnd vdd FILL
XFILL_0__8479_ gnd vdd FILL
XFILL_3__8188_ gnd vdd FILL
XFILL_1__9011_ gnd vdd FILL
XFILL_5_BUFX2_insert7 gnd vdd FILL
XSFILL13640x72050 gnd vdd FILL
XSFILL94520x68050 gnd vdd FILL
XFILL_1_BUFX2_insert708 gnd vdd FILL
XFILL_1_BUFX2_insert719 gnd vdd FILL
X_7989_ _7989_/A gnd _7989_/Y vdd INVX1
XFILL_4__7952_ gnd vdd FILL
X_9728_ _9764_/A _8576_/B gnd _9729_/C vdd NAND2X1
XFILL_4__6903_ gnd vdd FILL
XFILL_4__7883_ gnd vdd FILL
X_10610_ _16187_/A _9958_/CLK _8929_/R vdd _10610_/D gnd vdd DFFSR
XFILL_1__9913_ gnd vdd FILL
X_11590_ _11590_/A _11366_/B _11129_/Y _11574_/B gnd _11592_/B vdd OAI22X1
X_9659_ _9709_/Q gnd _9659_/Y vdd INVX1
XFILL_4__9622_ gnd vdd FILL
XSFILL8760x51050 gnd vdd FILL
X_10541_ _10505_/A _7853_/B gnd _10542_/C vdd NAND2X1
XSFILL33000x66050 gnd vdd FILL
XFILL_5_BUFX2_insert630 gnd vdd FILL
XFILL_5_BUFX2_insert641 gnd vdd FILL
XFILL_4__9553_ gnd vdd FILL
XFILL_5_BUFX2_insert652 gnd vdd FILL
X_13260_ _13295_/C _13260_/B gnd _13278_/B vdd NAND2X1
XFILL_5_BUFX2_insert663 gnd vdd FILL
XFILL_5_BUFX2_insert674 gnd vdd FILL
X_10472_ _10412_/A _7912_/CLK _7911_/R vdd _10472_/D gnd vdd DFFSR
XFILL_4__8504_ gnd vdd FILL
XFILL_1__9775_ gnd vdd FILL
XFILL_1__6987_ gnd vdd FILL
XFILL_5_BUFX2_insert685 gnd vdd FILL
XFILL_4__9484_ gnd vdd FILL
XFILL_5_BUFX2_insert696 gnd vdd FILL
X_12211_ _12216_/B gnd _12211_/Y vdd INVX8
X_13191_ _11935_/A _12537_/CLK _12536_/R vdd _13191_/D gnd vdd DFFSR
XFILL_1__8726_ gnd vdd FILL
X_12142_ _11914_/A gnd _12144_/A vdd INVX1
XSFILL63880x80050 gnd vdd FILL
XFILL_2__7450_ gnd vdd FILL
XFILL_1__8657_ gnd vdd FILL
XSFILL13720x52050 gnd vdd FILL
XFILL_2_CLKBUF1_insert200 gnd vdd FILL
XSFILL14200x59050 gnd vdd FILL
XFILL_2_CLKBUF1_insert211 gnd vdd FILL
XFILL_4__8366_ gnd vdd FILL
XFILL_2_CLKBUF1_insert222 gnd vdd FILL
XFILL_1__7608_ gnd vdd FILL
X_12073_ _12503_/B _12073_/B _12073_/C gnd gnd _12073_/Y vdd AOI22X1
XFILL_1__8588_ gnd vdd FILL
XFILL_2__7381_ gnd vdd FILL
XFILL_4__7317_ gnd vdd FILL
X_15901_ _15901_/A _15901_/B gnd _15902_/B vdd NOR2X1
XFILL_5__7090_ gnd vdd FILL
X_11024_ _11025_/A _12129_/Y gnd _11026_/C vdd AND2X2
XFILL_2__9120_ gnd vdd FILL
XSFILL28920x2050 gnd vdd FILL
XFILL_4__7248_ gnd vdd FILL
X_15832_ _16106_/A _15830_/Y _15832_/C _15948_/D gnd _15833_/B vdd OAI22X1
XFILL_4__10230_ gnd vdd FILL
XSFILL84280x38050 gnd vdd FILL
XFILL_2_BUFX2_insert520 gnd vdd FILL
XFILL_3__10960_ gnd vdd FILL
XFILL_1__10050_ gnd vdd FILL
XSFILL8840x31050 gnd vdd FILL
XFILL_2_BUFX2_insert531 gnd vdd FILL
XFILL_4__7179_ gnd vdd FILL
XFILL_0__10780_ gnd vdd FILL
XFILL_2_BUFX2_insert542 gnd vdd FILL
XFILL_5__11520_ gnd vdd FILL
XFILL_2_BUFX2_insert553 gnd vdd FILL
X_15763_ _9257_/A gnd _15765_/A vdd INVX1
XFILL_2__8002_ gnd vdd FILL
XFILL_1__9209_ gnd vdd FILL
X_12975_ _6878_/A gnd _12977_/A vdd INVX1
XFILL_4__10161_ gnd vdd FILL
XSFILL59080x14050 gnd vdd FILL
XFILL_2_BUFX2_insert564 gnd vdd FILL
XFILL_2__11340_ gnd vdd FILL
XFILL_2_BUFX2_insert575 gnd vdd FILL
XFILL_3__10891_ gnd vdd FILL
XFILL_5__9800_ gnd vdd FILL
X_14714_ _14714_/A _14712_/Y _14714_/C gnd _14715_/A vdd NAND3X1
XFILL_2_BUFX2_insert586 gnd vdd FILL
XFILL_5__7992_ gnd vdd FILL
X_11926_ _13188_/Q gnd _11926_/Y vdd INVX1
XFILL_5__11451_ gnd vdd FILL
XFILL_2_BUFX2_insert597 gnd vdd FILL
XFILL_3__12630_ gnd vdd FILL
X_15694_ _15694_/A _15693_/Y gnd _15694_/Y vdd NOR2X1
XFILL_2__11271_ gnd vdd FILL
XFILL_0__12450_ gnd vdd FILL
XFILL_5__9731_ gnd vdd FILL
XFILL_5__10402_ gnd vdd FILL
XFILL_5__6943_ gnd vdd FILL
X_14645_ _14645_/A _14645_/B gnd _14645_/Y vdd NAND2X1
XFILL_5__14170_ gnd vdd FILL
XFILL_2__13010_ gnd vdd FILL
XFILL_4__13920_ gnd vdd FILL
X_11857_ _11856_/Y _11857_/B _11675_/A gnd _11857_/Y vdd NAND3X1
XFILL_5__11382_ gnd vdd FILL
XFILL_0__11401_ gnd vdd FILL
XFILL_1__13740_ gnd vdd FILL
XFILL_1__10952_ gnd vdd FILL
XFILL_5__9662_ gnd vdd FILL
XFILL_0__12381_ gnd vdd FILL
XFILL_5__13121_ gnd vdd FILL
XSFILL38360x15050 gnd vdd FILL
XFILL_5__6874_ gnd vdd FILL
X_10808_ _14522_/A gnd _10810_/A vdd INVX1
XFILL_3__14300_ gnd vdd FILL
X_14576_ _7355_/A gnd _15986_/A vdd INVX1
XFILL_2__8904_ gnd vdd FILL
XSFILL13800x32050 gnd vdd FILL
XFILL_3__11512_ gnd vdd FILL
XFILL_4__13851_ gnd vdd FILL
XFILL_2__10153_ gnd vdd FILL
XFILL_0__14120_ gnd vdd FILL
XFILL_3__15280_ gnd vdd FILL
X_11788_ _11025_/A _11032_/Y _11786_/Y gnd _11789_/B vdd OAI21X1
XFILL_5__8613_ gnd vdd FILL
XFILL_2__9884_ gnd vdd FILL
XBUFX2_insert530 BUFX2_insert556/A gnd _7649_/R vdd BUFX2
XFILL_3__12492_ gnd vdd FILL
XFILL_0__11332_ gnd vdd FILL
XFILL_1__13671_ gnd vdd FILL
XFILL_1__10883_ gnd vdd FILL
X_16315_ _14942_/A gnd _16316_/A vdd INVX1
XFILL_6__14411_ gnd vdd FILL
XBUFX2_insert541 BUFX2_insert494/A gnd _8431_/R vdd BUFX2
X_13527_ _13879_/B gnd _13527_/Y vdd INVX8
XFILL_5__9593_ gnd vdd FILL
XBUFX2_insert552 BUFX2_insert524/A gnd _8433_/R vdd BUFX2
X_10739_ _10739_/Q _7661_/CLK _7789_/R vdd _10739_/D gnd vdd DFFSR
XFILL_3__14231_ gnd vdd FILL
XFILL_5__10264_ gnd vdd FILL
XBUFX2_insert563 BUFX2_insert559/A gnd _9054_/R vdd BUFX2
XFILL_1__15410_ gnd vdd FILL
XFILL_2__8835_ gnd vdd FILL
XFILL_4__13782_ gnd vdd FILL
XFILL_3__11443_ gnd vdd FILL
XFILL_1__12622_ gnd vdd FILL
XFILL_0__14051_ gnd vdd FILL
XFILL_2__14961_ gnd vdd FILL
XBUFX2_insert574 BUFX2_insert607/A gnd _8165_/R vdd BUFX2
XFILL_4__10994_ gnd vdd FILL
XFILL_1__16390_ gnd vdd FILL
XFILL_5__12003_ gnd vdd FILL
XBUFX2_insert585 BUFX2_insert496/A gnd _8034_/R vdd BUFX2
XFILL_0__11263_ gnd vdd FILL
XBUFX2_insert596 BUFX2_insert600/A gnd _8676_/R vdd BUFX2
XSFILL114440x36050 gnd vdd FILL
X_16246_ _16246_/A gnd _16246_/Y vdd INVX1
XFILL_4__12733_ gnd vdd FILL
X_13458_ _8022_/Q gnd _15048_/B vdd INVX1
XFILL_4__15521_ gnd vdd FILL
XFILL_0__7850_ gnd vdd FILL
XFILL_3__14162_ gnd vdd FILL
XFILL_5__10195_ gnd vdd FILL
XFILL_2__13912_ gnd vdd FILL
XFILL_0__13002_ gnd vdd FILL
XFILL_2__8766_ gnd vdd FILL
XFILL_1__15341_ gnd vdd FILL
XFILL_3__11374_ gnd vdd FILL
XFILL_2__14892_ gnd vdd FILL
X_12409_ _12409_/A gnd _12409_/Y vdd INVX1
XFILL_5__8475_ gnd vdd FILL
XFILL_0__11194_ gnd vdd FILL
X_16177_ _8394_/A _15978_/B _16212_/A _8690_/Q gnd _16178_/B vdd AOI22X1
XFILL_3__13113_ gnd vdd FILL
XFILL_6__14273_ gnd vdd FILL
XFILL_2__7717_ gnd vdd FILL
X_13389_ _13389_/A _13389_/B gnd _13390_/B vdd NOR2X1
XFILL_4__15452_ gnd vdd FILL
XFILL_3__10325_ gnd vdd FILL
XFILL_2__13843_ gnd vdd FILL
XFILL_3__14093_ gnd vdd FILL
XFILL_1__11504_ gnd vdd FILL
XFILL_6__16012_ gnd vdd FILL
XFILL_5__7426_ gnd vdd FILL
XFILL_1__12484_ gnd vdd FILL
XFILL_0__10145_ gnd vdd FILL
XFILL_3__7490_ gnd vdd FILL
XFILL_2__8697_ gnd vdd FILL
XFILL_1__15272_ gnd vdd FILL
XFILL_6__13224_ gnd vdd FILL
XFILL_0__9520_ gnd vdd FILL
X_15128_ _15569_/C gnd _15821_/B vdd INVX4
XFILL_4__11615_ gnd vdd FILL
XFILL_4__14403_ gnd vdd FILL
XFILL_4__15383_ gnd vdd FILL
XFILL_3__13044_ gnd vdd FILL
XFILL_5__13954_ gnd vdd FILL
XFILL_3__10256_ gnd vdd FILL
XFILL_4__12595_ gnd vdd FILL
XFILL_1__14223_ gnd vdd FILL
XFILL_1__11435_ gnd vdd FILL
XFILL_2__13774_ gnd vdd FILL
XSFILL84200x82050 gnd vdd FILL
XFILL_5__7357_ gnd vdd FILL
X_7010_ _6938_/A _7010_/CLK _8278_/R vdd _7010_/D gnd vdd DFFSR
XFILL_0__14953_ gnd vdd FILL
XFILL_6__10367_ gnd vdd FILL
X_15059_ _15036_/A _16037_/B _15212_/B gnd _15059_/Y vdd NAND3X1
XFILL_4__14334_ gnd vdd FILL
XFILL_5__12905_ gnd vdd FILL
XFILL_2__15513_ gnd vdd FILL
XFILL_4__11546_ gnd vdd FILL
XFILL_2__12725_ gnd vdd FILL
XFILL_5__13885_ gnd vdd FILL
XFILL_3__9160_ gnd vdd FILL
XFILL_3__10187_ gnd vdd FILL
XFILL_1__14154_ gnd vdd FILL
XFILL_2__7579_ gnd vdd FILL
XFILL_0__13904_ gnd vdd FILL
XFILL_1__11366_ gnd vdd FILL
XFILL_6__12106_ gnd vdd FILL
XFILL_0__8402_ gnd vdd FILL
XFILL_5__15624_ gnd vdd FILL
XFILL_5__7288_ gnd vdd FILL
XFILL_0__14884_ gnd vdd FILL
XFILL_0__9382_ gnd vdd FILL
XFILL_4__14265_ gnd vdd FILL
XFILL_5__12836_ gnd vdd FILL
XFILL_3__8111_ gnd vdd FILL
XFILL_1__10317_ gnd vdd FILL
XFILL_1__13105_ gnd vdd FILL
XFILL_4__11477_ gnd vdd FILL
XFILL_2__15444_ gnd vdd FILL
XFILL_2__12656_ gnd vdd FILL
XFILL_3__9091_ gnd vdd FILL
XFILL_3__14995_ gnd vdd FILL
XFILL_5__9027_ gnd vdd FILL
XFILL_1__14085_ gnd vdd FILL
XFILL_0__13835_ gnd vdd FILL
XFILL_1__11297_ gnd vdd FILL
XFILL_0__8333_ gnd vdd FILL
XFILL_4__13216_ gnd vdd FILL
XFILL_4__16004_ gnd vdd FILL
XFILL_4__10428_ gnd vdd FILL
XSFILL49080x46050 gnd vdd FILL
XFILL_5__15555_ gnd vdd FILL
X_8961_ _8961_/A _8961_/B _8960_/Y gnd _8961_/Y vdd OAI21X1
XFILL_5__12767_ gnd vdd FILL
XFILL112200x64050 gnd vdd FILL
XFILL_4__14196_ gnd vdd FILL
XFILL_2__9249_ gnd vdd FILL
XFILL_1__13036_ gnd vdd FILL
XFILL_2__11607_ gnd vdd FILL
XFILL_3__13946_ gnd vdd FILL
XFILL_1__10248_ gnd vdd FILL
XFILL_2__15375_ gnd vdd FILL
XFILL_2__12587_ gnd vdd FILL
XFILL_0__10978_ gnd vdd FILL
XFILL_0__13766_ gnd vdd FILL
XFILL_5__14506_ gnd vdd FILL
XFILL_4__13147_ gnd vdd FILL
X_7912_ _7852_/A _7912_/CLK _7911_/R vdd _7912_/D gnd vdd DFFSR
XFILL_5__11718_ gnd vdd FILL
XFILL_0__8264_ gnd vdd FILL
XFILL_4__10359_ gnd vdd FILL
XFILL_2__14326_ gnd vdd FILL
XFILL_5__15486_ gnd vdd FILL
XFILL_5__12698_ gnd vdd FILL
XFILL_3__13877_ gnd vdd FILL
X_8892_ _8893_/B _8764_/B gnd _8892_/Y vdd NAND2X1
XFILL_0__15505_ gnd vdd FILL
XFILL_2__11538_ gnd vdd FILL
XSFILL114520x16050 gnd vdd FILL
XFILL_0__12717_ gnd vdd FILL
XFILL_1__10179_ gnd vdd FILL
XFILL_0__7215_ gnd vdd FILL
XFILL_0__13697_ gnd vdd FILL
XFILL_5__14437_ gnd vdd FILL
X_7843_ _7909_/Q gnd _7843_/Y vdd INVX1
XFILL_0__8195_ gnd vdd FILL
XFILL_3__15616_ gnd vdd FILL
XFILL_5__11649_ gnd vdd FILL
XFILL_3__12828_ gnd vdd FILL
XFILL_2__14257_ gnd vdd FILL
XFILL_0__12648_ gnd vdd FILL
XFILL_3__9993_ gnd vdd FILL
XFILL_0__15436_ gnd vdd FILL
XFILL_2__11469_ gnd vdd FILL
XFILL_1__14987_ gnd vdd FILL
XFILL_5__9929_ gnd vdd FILL
XFILL_4__12029_ gnd vdd FILL
XFILL_2__13208_ gnd vdd FILL
XFILL_3__15547_ gnd vdd FILL
XFILL_5__14368_ gnd vdd FILL
X_7774_ _7694_/A _8942_/CLK _9561_/R vdd _7774_/D gnd vdd DFFSR
XFILL_3__12759_ gnd vdd FILL
XFILL_0_CLKBUF1_insert119 gnd vdd FILL
XFILL_2__14188_ gnd vdd FILL
XFILL_1__13938_ gnd vdd FILL
XFILL_0__12579_ gnd vdd FILL
XFILL_0__15367_ gnd vdd FILL
XFILL_5__16107_ gnd vdd FILL
XFILL_5__13319_ gnd vdd FILL
X_9513_ _9575_/Q gnd _9515_/A vdd INVX1
XFILL_0__7077_ gnd vdd FILL
XFILL_2__13139_ gnd vdd FILL
XFILL_5__14299_ gnd vdd FILL
XFILL_3__15478_ gnd vdd FILL
XFILL_0__14318_ gnd vdd FILL
XFILL_3__8875_ gnd vdd FILL
XFILL_1__13869_ gnd vdd FILL
XSFILL104440x68050 gnd vdd FILL
XFILL_0__15298_ gnd vdd FILL
XFILL_5__16038_ gnd vdd FILL
XFILL_1__6910_ gnd vdd FILL
X_9444_ _9376_/A _7642_/CLK _7258_/R vdd _9444_/D gnd vdd DFFSR
XFILL_3__14429_ gnd vdd FILL
XFILL_1__15608_ gnd vdd FILL
XFILL_3__7826_ gnd vdd FILL
XFILL_1__7890_ gnd vdd FILL
XFILL_0__14249_ gnd vdd FILL
XSFILL23720x15050 gnd vdd FILL
XFILL_1__6841_ gnd vdd FILL
XFILL_4__15719_ gnd vdd FILL
X_9375_ _9373_/Y _9339_/B _9375_/C gnd _9375_/Y vdd OAI21X1
XFILL_3__7757_ gnd vdd FILL
XFILL_1__15539_ gnd vdd FILL
XFILL_4_BUFX2_insert604 gnd vdd FILL
XSFILL74760x71050 gnd vdd FILL
XFILL_4_BUFX2_insert615 gnd vdd FILL
XFILL_4_BUFX2_insert626 gnd vdd FILL
XSFILL24600x43050 gnd vdd FILL
X_8326_ _8315_/B _9478_/B gnd _8327_/C vdd NAND2X1
XSFILL48920x81050 gnd vdd FILL
XFILL_0__7979_ gnd vdd FILL
XFILL_4_BUFX2_insert637 gnd vdd FILL
XFILL_3__7688_ gnd vdd FILL
XFILL_4_BUFX2_insert648 gnd vdd FILL
XFILL_1__8511_ gnd vdd FILL
XFILL_0__9718_ gnd vdd FILL
XFILL_4_BUFX2_insert659 gnd vdd FILL
XSFILL94440x8050 gnd vdd FILL
X_8257_ _8303_/Q gnd _8257_/Y vdd INVX1
XFILL_4__8220_ gnd vdd FILL
XFILL_3__9427_ gnd vdd FILL
XSFILL43720x4050 gnd vdd FILL
XFILL_1__9491_ gnd vdd FILL
XFILL_6__9136_ gnd vdd FILL
XSFILL13640x67050 gnd vdd FILL
X_7208_ _7208_/A _7207_/A _7208_/C gnd _7208_/Y vdd OAI21X1
XFILL_0__9649_ gnd vdd FILL
XFILL_1__8442_ gnd vdd FILL
X_8188_ _8280_/Q gnd _8190_/A vdd INVX1
XFILL_3__9358_ gnd vdd FILL
XFILL_2_BUFX2_insert70 gnd vdd FILL
XFILL_2_BUFX2_insert81 gnd vdd FILL
XFILL_2_BUFX2_insert92 gnd vdd FILL
X_7139_ _7139_/Q _7651_/CLK _9711_/R vdd _7139_/D gnd vdd DFFSR
XFILL_1__8373_ gnd vdd FILL
XFILL_4__7102_ gnd vdd FILL
XSFILL79480x83050 gnd vdd FILL
XFILL_3__9289_ gnd vdd FILL
XFILL_4__8082_ gnd vdd FILL
XSFILL54120x81050 gnd vdd FILL
XFILL_1__7324_ gnd vdd FILL
XSFILL104520x48050 gnd vdd FILL
XFILL_4__7033_ gnd vdd FILL
XSFILL8760x46050 gnd vdd FILL
X_12760_ _12758_/Y _12721_/B _12760_/C gnd _12812_/D vdd OAI21X1
XFILL_1_BUFX2_insert505 gnd vdd FILL
XFILL_1_BUFX2_insert516 gnd vdd FILL
XFILL_1__7186_ gnd vdd FILL
XSFILL74040x32050 gnd vdd FILL
XFILL_1_BUFX2_insert527 gnd vdd FILL
XFILL_4__8984_ gnd vdd FILL
XFILL_1_BUFX2_insert538 gnd vdd FILL
X_11711_ _11073_/Y gnd _11713_/A vdd INVX1
XFILL_1_BUFX2_insert549 gnd vdd FILL
X_12691_ _12428_/B _12809_/CLK _12685_/R vdd _12691_/D gnd vdd DFFSR
XFILL_4__7935_ gnd vdd FILL
X_14430_ _14429_/Y _14430_/B gnd _14430_/Y vdd NOR2X1
X_11642_ _11092_/Y _11641_/Y gnd _11642_/Y vdd NOR2X1
XFILL_2__6950_ gnd vdd FILL
XSFILL13720x47050 gnd vdd FILL
XFILL_4__7866_ gnd vdd FILL
XSFILL78680x35050 gnd vdd FILL
X_14361_ _7401_/Q gnd _14361_/Y vdd INVX1
X_11573_ _11115_/Y _11509_/B _11573_/C _11116_/Y gnd _11574_/C vdd AOI22X1
XSFILL109640x81050 gnd vdd FILL
XSFILL38680x51050 gnd vdd FILL
X_16100_ _16100_/A _16100_/B gnd _16100_/Y vdd NOR2X1
XFILL_2__6881_ gnd vdd FILL
XFILL_4__9605_ gnd vdd FILL
X_13312_ _13312_/A _13311_/Y _13295_/C gnd _13312_/Y vdd OAI21X1
X_10524_ _10522_/Y _10505_/A _10524_/C gnd _10594_/D vdd OAI21X1
XSFILL113880x44050 gnd vdd FILL
XFILL_2__8620_ gnd vdd FILL
X_14292_ _9831_/Q gnd _14292_/Y vdd INVX1
XFILL_5_BUFX2_insert460 gnd vdd FILL
XFILL_5_BUFX2_insert471 gnd vdd FILL
XFILL_4__9536_ gnd vdd FILL
X_16031_ _15392_/C _14599_/Y _15677_/D _14634_/Y gnd _16032_/B vdd OAI22X1
XFILL_5_BUFX2_insert482 gnd vdd FILL
X_13243_ _13295_/C _13302_/C gnd _13244_/B vdd NAND2X1
XFILL_5_BUFX2_insert493 gnd vdd FILL
X_10455_ _13528_/A _7515_/CLK _7000_/R vdd _10363_/Y gnd vdd DFFSR
XFILL_1__9758_ gnd vdd FILL
XFILL_5__8260_ gnd vdd FILL
XFILL_4__9467_ gnd vdd FILL
XSFILL8840x26050 gnd vdd FILL
XFILL_2__7502_ gnd vdd FILL
X_13174_ _13174_/A _13173_/A _13174_/C gnd _13206_/D vdd OAI21X1
XFILL_3__10110_ gnd vdd FILL
XFILL_1__8709_ gnd vdd FILL
X_10386_ _10450_/B _7954_/B gnd _10386_/Y vdd NAND2X1
XFILL_2__8482_ gnd vdd FILL
XFILL_3__11090_ gnd vdd FILL
XFILL_5__7211_ gnd vdd FILL
XFILL_5__8191_ gnd vdd FILL
XFILL_4__9398_ gnd vdd FILL
X_12125_ _12137_/A _12125_/B gnd _12126_/C vdd NAND2X1
XFILL_4__11400_ gnd vdd FILL
XSFILL99480x14050 gnd vdd FILL
XFILL_5__10951_ gnd vdd FILL
XFILL_4__12380_ gnd vdd FILL
XFILL_2__7433_ gnd vdd FILL
XFILL_3__10041_ gnd vdd FILL
XFILL_1__11220_ gnd vdd FILL
XSFILL74120x12050 gnd vdd FILL
XFILL_0__11950_ gnd vdd FILL
XFILL_2__10771_ gnd vdd FILL
XFILL_4__8349_ gnd vdd FILL
X_12056_ _11988_/B _11885_/B _12096_/C gnd _12056_/Y vdd NAND3X1
XFILL_4__11331_ gnd vdd FILL
XFILL_5__13670_ gnd vdd FILL
XFILL_2__12510_ gnd vdd FILL
XFILL_5__10882_ gnd vdd FILL
XFILL_0__10901_ gnd vdd FILL
XFILL_2__7364_ gnd vdd FILL
XFILL_1__11151_ gnd vdd FILL
XFILL_2__13490_ gnd vdd FILL
XFILL_0__11881_ gnd vdd FILL
XFILL_5__7073_ gnd vdd FILL
X_11007_ _12120_/Y gnd _11007_/Y vdd INVX1
XFILL_5__12621_ gnd vdd FILL
XFILL_2__9103_ gnd vdd FILL
XFILL_3__13800_ gnd vdd FILL
XSFILL63960x55050 gnd vdd FILL
XFILL_4__14050_ gnd vdd FILL
XFILL_1__10102_ gnd vdd FILL
XFILL_4__11262_ gnd vdd FILL
XFILL_2__12441_ gnd vdd FILL
XFILL_3__14780_ gnd vdd FILL
XFILL_2__7295_ gnd vdd FILL
XFILL_0__13620_ gnd vdd FILL
XFILL_3__11992_ gnd vdd FILL
XFILL_1__11082_ gnd vdd FILL
XFILL_0__10832_ gnd vdd FILL
XFILL_4__13001_ gnd vdd FILL
XFILL_5__15340_ gnd vdd FILL
X_15815_ _16225_/C _15815_/B _15726_/A _15815_/D gnd _15816_/B vdd OAI22X1
XFILL_2__9034_ gnd vdd FILL
XFILL_3__13731_ gnd vdd FILL
XFILL_3__10943_ gnd vdd FILL
XFILL_1__10033_ gnd vdd FILL
XFILL_2_BUFX2_insert350 gnd vdd FILL
XFILL_2__15160_ gnd vdd FILL
XFILL_1__14910_ gnd vdd FILL
XFILL_4__11193_ gnd vdd FILL
XSFILL64040x64050 gnd vdd FILL
XFILL_2__12372_ gnd vdd FILL
XFILL_2_BUFX2_insert361 gnd vdd FILL
XFILL_0__13551_ gnd vdd FILL
XFILL_2_BUFX2_insert372 gnd vdd FILL
XFILL_0__10763_ gnd vdd FILL
XFILL_1__15890_ gnd vdd FILL
X_15746_ _15745_/Y _15746_/B _15736_/Y gnd _15770_/A vdd NOR3X1
XFILL_5__11503_ gnd vdd FILL
XFILL_2_BUFX2_insert383 gnd vdd FILL
XFILL_3__16450_ gnd vdd FILL
XFILL_4__10144_ gnd vdd FILL
XFILL_5__12483_ gnd vdd FILL
XFILL_2_BUFX2_insert394 gnd vdd FILL
XFILL_2__14111_ gnd vdd FILL
XFILL_5__15271_ gnd vdd FILL
X_12958_ vdd _13584_/Y gnd _12958_/Y vdd NAND2X1
XFILL_0__12502_ gnd vdd FILL
XFILL_3__13662_ gnd vdd FILL
XFILL_2__11323_ gnd vdd FILL
XFILL_1__14841_ gnd vdd FILL
XFILL_3__10874_ gnd vdd FILL
XFILL_2__15091_ gnd vdd FILL
XSFILL49080x4050 gnd vdd FILL
XFILL_0__13482_ gnd vdd FILL
XFILL_0__16270_ gnd vdd FILL
XFILL_5__7975_ gnd vdd FILL
XFILL_5__14222_ gnd vdd FILL
XFILL_3__15401_ gnd vdd FILL
X_11909_ _11909_/A _12364_/A gnd _11910_/C vdd NAND2X1
XFILL_0__10694_ gnd vdd FILL
XFILL_5__11434_ gnd vdd FILL
X_15677_ _15677_/A _15676_/Y _14187_/Y _15677_/D gnd _15678_/C vdd OAI22X1
XFILL_3__12613_ gnd vdd FILL
X_12889_ _12889_/A gnd _12889_/Y vdd INVX1
XFILL_2__14042_ gnd vdd FILL
XFILL_4__14952_ gnd vdd FILL
XFILL_3__16381_ gnd vdd FILL
XSFILL43880x22050 gnd vdd FILL
XSFILL3480x71050 gnd vdd FILL
XFILL_3__13593_ gnd vdd FILL
XFILL_0__15221_ gnd vdd FILL
XFILL_0__12433_ gnd vdd FILL
XFILL_2__11254_ gnd vdd FILL
XFILL_3__6990_ gnd vdd FILL
XFILL_5__6926_ gnd vdd FILL
XFILL_1__14772_ gnd vdd FILL
X_14628_ _14628_/A _14203_/B gnd _14629_/C vdd NOR2X1
XFILL_1__11984_ gnd vdd FILL
XFILL_3__15332_ gnd vdd FILL
XFILL_5__14153_ gnd vdd FILL
XFILL_4__13903_ gnd vdd FILL
XFILL_5__11365_ gnd vdd FILL
XFILL_1__13723_ gnd vdd FILL
XFILL_2__11185_ gnd vdd FILL
XFILL_0__15152_ gnd vdd FILL
XFILL_2__9936_ gnd vdd FILL
XFILL_4__14883_ gnd vdd FILL
XFILL_1__10935_ gnd vdd FILL
XFILL_0__12364_ gnd vdd FILL
XFILL_5__10316_ gnd vdd FILL
XFILL_5__13104_ gnd vdd FILL
XFILL_5__6857_ gnd vdd FILL
XFILL_5__9645_ gnd vdd FILL
XFILL_6__12655_ gnd vdd FILL
X_14559_ _14559_/A _14558_/Y _14559_/C gnd _14570_/B vdd NAND3X1
XFILL_0__8951_ gnd vdd FILL
XFILL_5__14084_ gnd vdd FILL
XFILL_4__13834_ gnd vdd FILL
XFILL_2__10136_ gnd vdd FILL
XFILL_0__14103_ gnd vdd FILL
XFILL_5__11296_ gnd vdd FILL
X_7490_ _7430_/A _7490_/B gnd _7490_/Y vdd NAND2X1
XFILL_3__15263_ gnd vdd FILL
XFILL_2__9867_ gnd vdd FILL
XFILL_3__12475_ gnd vdd FILL
XFILL_0__11315_ gnd vdd FILL
XBUFX2_insert360 _11352_/Y gnd _11360_/C vdd BUFX2
XFILL_3__8660_ gnd vdd FILL
XFILL_2__15993_ gnd vdd FILL
XFILL_1__13654_ gnd vdd FILL
XFILL_0__15083_ gnd vdd FILL
XBUFX2_insert371 _13338_/Y gnd _9554_/B vdd BUFX2
XFILL_0__12295_ gnd vdd FILL
XFILL_3__14214_ gnd vdd FILL
XSFILL59000x53050 gnd vdd FILL
XFILL_5__13035_ gnd vdd FILL
XFILL_5__10247_ gnd vdd FILL
XBUFX2_insert382 _13331_/Y gnd _9170_/B vdd BUFX2
XFILL_3__7611_ gnd vdd FILL
XBUFX2_insert393 _12387_/Y gnd _9889_/B vdd BUFX2
XFILL_0__8882_ gnd vdd FILL
XFILL_3__11426_ gnd vdd FILL
XFILL_1__12605_ gnd vdd FILL
XFILL_4__10977_ gnd vdd FILL
XFILL_3__15194_ gnd vdd FILL
XFILL_4__13765_ gnd vdd FILL
XFILL_0__14034_ gnd vdd FILL
XFILL_2__10067_ gnd vdd FILL
XFILL_2__14944_ gnd vdd FILL
XFILL_3__8591_ gnd vdd FILL
XFILL_5__8527_ gnd vdd FILL
XFILL_2__9798_ gnd vdd FILL
XFILL_0__11246_ gnd vdd FILL
XFILL_1__16373_ gnd vdd FILL
XFILL_1__13585_ gnd vdd FILL
X_16229_ _16002_/C _14870_/Y _14849_/A _15170_/D gnd _16230_/B vdd OAI22X1
XFILL_1__10797_ gnd vdd FILL
XFILL_0__7833_ gnd vdd FILL
XFILL_4__15504_ gnd vdd FILL
X_9160_ _9086_/B _7240_/B gnd _9161_/C vdd NAND2X1
XFILL_4__12716_ gnd vdd FILL
XFILL_3__14145_ gnd vdd FILL
XFILL_5__10178_ gnd vdd FILL
XFILL112200x59050 gnd vdd FILL
XFILL_1__15324_ gnd vdd FILL
XFILL_3__7542_ gnd vdd FILL
XFILL_2__8749_ gnd vdd FILL
XSFILL23240x32050 gnd vdd FILL
XFILL_4__13696_ gnd vdd FILL
XFILL_3__11357_ gnd vdd FILL
XFILL_2__14875_ gnd vdd FILL
XFILL_5__8458_ gnd vdd FILL
X_8111_ _8169_/Q gnd _8111_/Y vdd INVX1
XSFILL38840x11050 gnd vdd FILL
XFILL_0__11177_ gnd vdd FILL
XSFILL109000x22050 gnd vdd FILL
X_9091_ _9101_/B _9475_/B gnd _9092_/C vdd NAND2X1
XSFILL64120x44050 gnd vdd FILL
XFILL_3__10308_ gnd vdd FILL
XFILL_0__7764_ gnd vdd FILL
XFILL_4__15435_ gnd vdd FILL
XFILL_4__12647_ gnd vdd FILL
XFILL_2__13826_ gnd vdd FILL
XFILL_5__14986_ gnd vdd FILL
XFILL_3__14076_ gnd vdd FILL
XFILL_0__10128_ gnd vdd FILL
XFILL_1__15255_ gnd vdd FILL
XFILL_3__7473_ gnd vdd FILL
XFILL_3__11288_ gnd vdd FILL
XFILL_1__12467_ gnd vdd FILL
XFILL_0__9503_ gnd vdd FILL
XFILL_0__15985_ gnd vdd FILL
XFILL_5__8389_ gnd vdd FILL
XFILL_6__10419_ gnd vdd FILL
X_8042_ _8042_/Q _8169_/CLK _8937_/R vdd _8042_/D gnd vdd DFFSR
XFILL_3__13027_ gnd vdd FILL
XFILL_5__13937_ gnd vdd FILL
XFILL_3__9212_ gnd vdd FILL
XFILL_0__7695_ gnd vdd FILL
XFILL_4__12578_ gnd vdd FILL
XFILL_3__10239_ gnd vdd FILL
XFILL_4__15366_ gnd vdd FILL
XFILL_1__14206_ gnd vdd FILL
XFILL_2__13757_ gnd vdd FILL
XFILL_1__11418_ gnd vdd FILL
XFILL_2__10969_ gnd vdd FILL
XFILL_1__12398_ gnd vdd FILL
XFILL_1__15186_ gnd vdd FILL
XFILL_0__10059_ gnd vdd FILL
XFILL_0__14936_ gnd vdd FILL
XSFILL3560x51050 gnd vdd FILL
XFILL_4__14317_ gnd vdd FILL
XFILL_4__11529_ gnd vdd FILL
XFILL_3__9143_ gnd vdd FILL
XFILL_2__12708_ gnd vdd FILL
XFILL_5__13868_ gnd vdd FILL
XFILL_4__15297_ gnd vdd FILL
XFILL_1__14137_ gnd vdd FILL
XFILL_2__13688_ gnd vdd FILL
XFILL_1__11349_ gnd vdd FILL
XFILL_0__14867_ gnd vdd FILL
XFILL_5__15607_ gnd vdd FILL
XSFILL28760x63050 gnd vdd FILL
XFILL_0__9365_ gnd vdd FILL
XFILL_4__14248_ gnd vdd FILL
XFILL_2__15427_ gnd vdd FILL
XFILL_5__13799_ gnd vdd FILL
XFILL_2__12639_ gnd vdd FILL
X_9993_ _9993_/A _9993_/B gnd _9994_/C vdd NAND2X1
XSFILL44040x11050 gnd vdd FILL
XFILL_0__13818_ gnd vdd FILL
XFILL_1__14068_ gnd vdd FILL
XFILL_3__14978_ gnd vdd FILL
XFILL_0__8316_ gnd vdd FILL
XFILL_0__14798_ gnd vdd FILL
XFILL_5__15538_ gnd vdd FILL
XFILL_4__14179_ gnd vdd FILL
X_8944_ _8900_/A _9328_/CLK _7408_/R vdd _8902_/Y gnd vdd DFFSR
XFILL_0__9296_ gnd vdd FILL
XFILL_2__15358_ gnd vdd FILL
XFILL_1__13019_ gnd vdd FILL
XFILL_3__13929_ gnd vdd FILL
XFILL_0__13749_ gnd vdd FILL
XFILL_1__7040_ gnd vdd FILL
XFILL_0__8247_ gnd vdd FILL
XSFILL33880x54050 gnd vdd FILL
XFILL_2__14309_ gnd vdd FILL
XFILL_5__15469_ gnd vdd FILL
X_8875_ _8875_/A _8859_/A _8874_/Y gnd _8935_/D vdd OAI21X1
XFILL_2__15289_ gnd vdd FILL
X_7826_ _7878_/B _8466_/B gnd _7827_/C vdd NAND2X1
XSFILL89560x26050 gnd vdd FILL
XFILL_0__15419_ gnd vdd FILL
XFILL_3__9976_ gnd vdd FILL
XSFILL64200x24050 gnd vdd FILL
XFILL_0__16399_ gnd vdd FILL
X_7757_ _7757_/A gnd _7759_/A vdd INVX1
XFILL_4__7720_ gnd vdd FILL
XFILL_1__8991_ gnd vdd FILL
XFILL_1__7942_ gnd vdd FILL
X_7688_ _7688_/A gnd _7688_/Y vdd INVX1
XFILL_3__8858_ gnd vdd FILL
XSFILL3640x31050 gnd vdd FILL
X_9427_ _9461_/Q gnd _9427_/Y vdd INVX1
XFILL_1__7873_ gnd vdd FILL
XFILL_3__7809_ gnd vdd FILL
XFILL_4__7582_ gnd vdd FILL
XFILL_3__8789_ gnd vdd FILL
XFILL_1__9612_ gnd vdd FILL
XFILL_4_BUFX2_insert401 gnd vdd FILL
X_9358_ _9438_/Q gnd _9358_/Y vdd INVX1
XFILL_4_BUFX2_insert412 gnd vdd FILL
XFILL_4_BUFX2_insert423 gnd vdd FILL
XFILL_4_BUFX2_insert434 gnd vdd FILL
X_10240_ _10318_/A _9600_/B gnd _10241_/C vdd NAND2X1
XFILL_4_BUFX2_insert445 gnd vdd FILL
XSFILL79080x80050 gnd vdd FILL
XFILL_1__9543_ gnd vdd FILL
X_8309_ _8275_/A _9589_/CLK _7285_/R vdd _8309_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert456 gnd vdd FILL
XFILL_4__9252_ gnd vdd FILL
XFILL_4_BUFX2_insert467 gnd vdd FILL
X_9289_ _9287_/Y _9301_/B _9289_/C gnd _9289_/Y vdd OAI21X1
XFILL_4_BUFX2_insert478 gnd vdd FILL
X_10171_ _10171_/A gnd _10171_/Y vdd INVX1
XFILL_4_BUFX2_insert489 gnd vdd FILL
XSFILL33960x34050 gnd vdd FILL
XFILL_1__9474_ gnd vdd FILL
XSFILL58760x79050 gnd vdd FILL
XFILL_4__8203_ gnd vdd FILL
XFILL_4__8134_ gnd vdd FILL
X_13930_ _13930_/A _13930_/B _14402_/C gnd _12979_/B vdd AOI21X1
XFILL_1__8356_ gnd vdd FILL
XFILL_4__8065_ gnd vdd FILL
XFILL_3_CLKBUF1_insert114 gnd vdd FILL
X_13861_ _13860_/Y _13857_/Y gnd _13862_/C vdd NOR2X1
XFILL_1__7307_ gnd vdd FILL
XFILL_3_CLKBUF1_insert125 gnd vdd FILL
XFILL_5_CLKBUF1_insert1074 gnd vdd FILL
XFILL_3_CLKBUF1_insert136 gnd vdd FILL
XFILL_2__7080_ gnd vdd FILL
XFILL_3_CLKBUF1_insert147 gnd vdd FILL
XSFILL3720x11050 gnd vdd FILL
XFILL_3_CLKBUF1_insert158 gnd vdd FILL
X_15600_ _7139_/Q gnd _15601_/B vdd INVX1
X_12812_ _12812_/Q _7005_/CLK _12799_/R vdd _12812_/D gnd vdd DFFSR
XFILL_3_CLKBUF1_insert169 gnd vdd FILL
X_13792_ _13792_/A _14496_/A _13791_/Y gnd _13792_/Y vdd OAI21X1
XFILL_1__7238_ gnd vdd FILL
XFILL_1_BUFX2_insert302 gnd vdd FILL
XSFILL113880x39050 gnd vdd FILL
XSFILL28920x23050 gnd vdd FILL
XFILL_1_BUFX2_insert313 gnd vdd FILL
X_15531_ _7575_/A gnd _15531_/Y vdd INVX1
XFILL_1_BUFX2_insert324 gnd vdd FILL
X_12743_ _12807_/Q gnd _12745_/A vdd INVX1
XFILL_1_BUFX2_insert335 gnd vdd FILL
XFILL_1_BUFX2_insert346 gnd vdd FILL
XFILL_1__7169_ gnd vdd FILL
XFILL_1_BUFX2_insert357 gnd vdd FILL
XFILL_1_BUFX2_insert368 gnd vdd FILL
XSFILL13640x8050 gnd vdd FILL
XFILL_5__7760_ gnd vdd FILL
XFILL_1_BUFX2_insert379 gnd vdd FILL
XFILL_4__8967_ gnd vdd FILL
X_15462_ _15458_/Y _15462_/B _15461_/Y gnd _15466_/C vdd NOR3X1
X_12674_ _12600_/A _12685_/CLK _12685_/R vdd _12674_/D gnd vdd DFFSR
XFILL_6__10770_ gnd vdd FILL
XSFILL48840x50 gnd vdd FILL
XFILL_2__7982_ gnd vdd FILL
XSFILL104200x25050 gnd vdd FILL
X_14413_ _14413_/A _8242_/A _15863_/B _13621_/B gnd _14413_/Y vdd AOI22X1
XFILL_5__7691_ gnd vdd FILL
XFILL_4__10900_ gnd vdd FILL
XFILL_4__8898_ gnd vdd FILL
XFILL_5__11150_ gnd vdd FILL
X_11625_ _11614_/A _11625_/B gnd _11627_/A vdd NOR2X1
X_15393_ _10462_/Q gnd _15394_/A vdd INVX1
XFILL_2__9721_ gnd vdd FILL
XFILL_4__11880_ gnd vdd FILL
XFILL_2__6933_ gnd vdd FILL
XSFILL18840x75050 gnd vdd FILL
XSFILL84280x51050 gnd vdd FILL
X_14344_ _15787_/A _14344_/B _14344_/C _7084_/A gnd _14344_/Y vdd AOI22X1
XFILL_4__7849_ gnd vdd FILL
XFILL_4__10831_ gnd vdd FILL
XFILL_5__11081_ gnd vdd FILL
X_11556_ _11110_/Y _11509_/B _11555_/Y gnd _11556_/Y vdd AOI21X1
XSFILL58440x61050 gnd vdd FILL
XFILL_3__12260_ gnd vdd FILL
XFILL_0__11100_ gnd vdd FILL
XFILL_2__9652_ gnd vdd FILL
XFILL_2__6864_ gnd vdd FILL
XFILL_1__10651_ gnd vdd FILL
XFILL_0__12080_ gnd vdd FILL
XFILL_5__9361_ gnd vdd FILL
XFILL_2__12990_ gnd vdd FILL
X_10507_ _10589_/Q gnd _10509_/A vdd INVX1
XFILL_5__10032_ gnd vdd FILL
XSFILL99320x73050 gnd vdd FILL
XFILL_2__8603_ gnd vdd FILL
XFILL_4__13550_ gnd vdd FILL
XFILL_3__11211_ gnd vdd FILL
X_14275_ _14275_/A _14275_/B _14275_/C gnd _14288_/A vdd NAND3X1
XFILL_4__10762_ gnd vdd FILL
XFILL_5_BUFX2_insert290 gnd vdd FILL
X_11487_ _11360_/C _11473_/C _11487_/C gnd _11487_/Y vdd NAND3X1
XFILL_5__8312_ gnd vdd FILL
XFILL_2__11941_ gnd vdd FILL
XSFILL59000x7050 gnd vdd FILL
XFILL_3__12191_ gnd vdd FILL
XFILL_0__11031_ gnd vdd FILL
X_16014_ _7230_/A _15177_/B _16014_/C _8254_/A gnd _16020_/B vdd AOI22X1
XFILL_1__13370_ gnd vdd FILL
XFILL_4__9519_ gnd vdd FILL
X_13226_ _13225_/Y _13226_/B gnd _13335_/A vdd NOR2X1
XFILL_5__9292_ gnd vdd FILL
XFILL_5__14840_ gnd vdd FILL
XFILL_4__12501_ gnd vdd FILL
X_10438_ _10438_/A _10372_/B _10437_/Y gnd _10438_/Y vdd OAI21X1
XFILL_3__11142_ gnd vdd FILL
XFILL_4__13481_ gnd vdd FILL
XFILL_4__10693_ gnd vdd FILL
XFILL112280x33050 gnd vdd FILL
XFILL_1__12321_ gnd vdd FILL
XFILL_2__14660_ gnd vdd FILL
XFILL_2__11872_ gnd vdd FILL
XFILL_5__8243_ gnd vdd FILL
XFILL_4__12432_ gnd vdd FILL
X_13157_ _13157_/A gnd _13157_/Y vdd INVX1
XFILL_4__15220_ gnd vdd FILL
X_10369_ _10367_/Y _10443_/A _10369_/C gnd _10457_/D vdd OAI21X1
XFILL_2__13611_ gnd vdd FILL
XFILL_4_BUFX2_insert990 gnd vdd FILL
XFILL_5__14771_ gnd vdd FILL
XFILL_5__11983_ gnd vdd FILL
XFILL_1__15040_ gnd vdd FILL
XFILL_3__15950_ gnd vdd FILL
XFILL_1__12252_ gnd vdd FILL
XFILL_3__11073_ gnd vdd FILL
XFILL_2__8465_ gnd vdd FILL
XFILL_2__10823_ gnd vdd FILL
XFILL_2__14591_ gnd vdd FILL
X_12108_ _11988_/B _12108_/B _12096_/C gnd _12110_/B vdd NAND3X1
XFILL_0__15770_ gnd vdd FILL
XSFILL74200x1050 gnd vdd FILL
XFILL_0__12982_ gnd vdd FILL
XFILL_4__15151_ gnd vdd FILL
XFILL_5__13722_ gnd vdd FILL
XFILL_5__10934_ gnd vdd FILL
XFILL_4__12363_ gnd vdd FILL
XFILL_2__16330_ gnd vdd FILL
X_13088_ _11896_/A gnd _13090_/A vdd INVX1
XFILL_3__10024_ gnd vdd FILL
XFILL_2__7416_ gnd vdd FILL
XFILL_0__7480_ gnd vdd FILL
XFILL_3__14901_ gnd vdd FILL
XSFILL79240x40050 gnd vdd FILL
XSFILL43880x17050 gnd vdd FILL
XFILL_2__13542_ gnd vdd FILL
XFILL_1__11203_ gnd vdd FILL
XFILL_2__8396_ gnd vdd FILL
XFILL_2__10754_ gnd vdd FILL
XFILL_5__7125_ gnd vdd FILL
XFILL_0__14721_ gnd vdd FILL
XFILL_1__12183_ gnd vdd FILL
XFILL_3__15881_ gnd vdd FILL
XFILL_0__11933_ gnd vdd FILL
XFILL_6__10135_ gnd vdd FILL
X_12039_ _12031_/A _12382_/A _12031_/C gnd _12042_/A vdd NAND3X1
XFILL_4__14102_ gnd vdd FILL
XFILL_4__11314_ gnd vdd FILL
XFILL_5__13653_ gnd vdd FILL
XFILL_6__15992_ gnd vdd FILL
XFILL_4__15082_ gnd vdd FILL
XFILL_3__14832_ gnd vdd FILL
XFILL_4__12294_ gnd vdd FILL
XFILL_1__11134_ gnd vdd FILL
XFILL_2__16261_ gnd vdd FILL
XFILL_2__7347_ gnd vdd FILL
XFILL_2__13473_ gnd vdd FILL
XFILL_2__10685_ gnd vdd FILL
XFILL_5__7056_ gnd vdd FILL
XFILL_0__11864_ gnd vdd FILL
XFILL_0__14652_ gnd vdd FILL
XFILL_5__12604_ gnd vdd FILL
XFILL_0__9150_ gnd vdd FILL
XFILL_4__14033_ gnd vdd FILL
XFILL_6__14943_ gnd vdd FILL
XFILL_2__15212_ gnd vdd FILL
XFILL_5__16372_ gnd vdd FILL
XFILL_4__11245_ gnd vdd FILL
XFILL_2__12424_ gnd vdd FILL
XFILL_5__13584_ gnd vdd FILL
XFILL_3__14763_ gnd vdd FILL
X_6990_ _6951_/A _8910_/B gnd _6991_/C vdd NAND2X1
XFILL_0__13603_ gnd vdd FILL
XFILL_3__11975_ gnd vdd FILL
XFILL_2__16192_ gnd vdd FILL
XFILL_1__15942_ gnd vdd FILL
XFILL_5__10796_ gnd vdd FILL
XSFILL84360x31050 gnd vdd FILL
XFILL_1__11065_ gnd vdd FILL
XFILL_0__10815_ gnd vdd FILL
XFILL_0__8101_ gnd vdd FILL
XFILL_0__14583_ gnd vdd FILL
XFILL_5__15323_ gnd vdd FILL
XFILL_0__11795_ gnd vdd FILL
XSFILL59000x48050 gnd vdd FILL
XFILL_2__9017_ gnd vdd FILL
XFILL_0__9081_ gnd vdd FILL
XFILL_3__10926_ gnd vdd FILL
XFILL_1__10016_ gnd vdd FILL
XFILL_2__15143_ gnd vdd FILL
XFILL_4__11176_ gnd vdd FILL
XFILL_3__13714_ gnd vdd FILL
XFILL_0__16322_ gnd vdd FILL
XFILL_2__12355_ gnd vdd FILL
XFILL_3__14694_ gnd vdd FILL
XSFILL99400x53050 gnd vdd FILL
XFILL_1__15873_ gnd vdd FILL
XFILL_0__10746_ gnd vdd FILL
XFILL_0__13534_ gnd vdd FILL
XFILL_4__10127_ gnd vdd FILL
X_15729_ _15729_/A _15729_/B gnd _15730_/B vdd NOR2X1
XFILL_5__15254_ gnd vdd FILL
XFILL_3__13645_ gnd vdd FILL
XFILL_5__12466_ gnd vdd FILL
XFILL_2__11306_ gnd vdd FILL
X_8660_ _8607_/B _9172_/B gnd _8660_/Y vdd NAND2X1
XFILL_4__15984_ gnd vdd FILL
XFILL_1__14824_ gnd vdd FILL
XFILL_2__15074_ gnd vdd FILL
XFILL_0__13465_ gnd vdd FILL
XFILL_0__16253_ gnd vdd FILL
XFILL_2__12286_ gnd vdd FILL
XFILL_0__10677_ gnd vdd FILL
XFILL_5__14205_ gnd vdd FILL
X_7611_ _7611_/A gnd _7613_/A vdd INVX1
XFILL_6__13756_ gnd vdd FILL
XFILL_5__7958_ gnd vdd FILL
XFILL112360x13050 gnd vdd FILL
XFILL_5__11417_ gnd vdd FILL
XFILL_5__15185_ gnd vdd FILL
XFILL_4__10058_ gnd vdd FILL
XFILL_2__14025_ gnd vdd FILL
XSFILL64120x39050 gnd vdd FILL
XFILL_4__14935_ gnd vdd FILL
XFILL_1_BUFX2_insert880 gnd vdd FILL
X_8591_ _8577_/B _8207_/B gnd _8592_/C vdd NAND2X1
XFILL_1_BUFX2_insert891 gnd vdd FILL
XFILL_0__15204_ gnd vdd FILL
XFILL_3__9761_ gnd vdd FILL
XFILL_3__16364_ gnd vdd FILL
XFILL_5__12397_ gnd vdd FILL
XFILL_3__13576_ gnd vdd FILL
XFILL_2__11237_ gnd vdd FILL
XFILL_3__6973_ gnd vdd FILL
XFILL_3__10788_ gnd vdd FILL
XFILL_0__12416_ gnd vdd FILL
XFILL_1__14755_ gnd vdd FILL
XFILL_6__12707_ gnd vdd FILL
XFILL_0__16184_ gnd vdd FILL
XFILL_1__11967_ gnd vdd FILL
XFILL_0__13396_ gnd vdd FILL
XFILL_5__6909_ gnd vdd FILL
XFILL_5__14136_ gnd vdd FILL
XFILL_0__9983_ gnd vdd FILL
XFILL_3__8712_ gnd vdd FILL
XFILL_3__15315_ gnd vdd FILL
XFILL_3__12527_ gnd vdd FILL
X_7542_ _7638_/Q gnd _7542_/Y vdd INVX1
XFILL_5__7889_ gnd vdd FILL
XFILL_5__11348_ gnd vdd FILL
XFILL_4__14866_ gnd vdd FILL
XFILL_2__9919_ gnd vdd FILL
XFILL_3__16295_ gnd vdd FILL
XFILL_1__13706_ gnd vdd FILL
XFILL_1__10918_ gnd vdd FILL
XFILL_0__12347_ gnd vdd FILL
XFILL_0__15135_ gnd vdd FILL
XFILL_2__11168_ gnd vdd FILL
XFILL_5__9628_ gnd vdd FILL
XFILL_1__14686_ gnd vdd FILL
XFILL_1__11898_ gnd vdd FILL
XSFILL79320x20050 gnd vdd FILL
XFILL_4__13817_ gnd vdd FILL
XFILL_3__15246_ gnd vdd FILL
XFILL_5__14067_ gnd vdd FILL
X_7473_ _7473_/A _7472_/A _7473_/C gnd _7473_/Y vdd OAI21X1
XFILL_5__11279_ gnd vdd FILL
XFILL_3__12458_ gnd vdd FILL
XSFILL3560x46050 gnd vdd FILL
XFILL_3__8643_ gnd vdd FILL
XFILL_2__10119_ gnd vdd FILL
XFILL_1__13637_ gnd vdd FILL
XFILL_4__14797_ gnd vdd FILL
XSFILL13160x79050 gnd vdd FILL
XFILL_2__15976_ gnd vdd FILL
XFILL_0__15066_ gnd vdd FILL
XFILL_0__12278_ gnd vdd FILL
XFILL_2__11099_ gnd vdd FILL
XFILL_6__15357_ gnd vdd FILL
XFILL_5__13018_ gnd vdd FILL
X_9212_ _9304_/Q gnd _9212_/Y vdd INVX1
XFILL_0__8865_ gnd vdd FILL
XFILL_3__11409_ gnd vdd FILL
XFILL_3__15177_ gnd vdd FILL
XFILL_4__13748_ gnd vdd FILL
XFILL_3__12389_ gnd vdd FILL
XFILL_0__14017_ gnd vdd FILL
XFILL_1__16356_ gnd vdd FILL
XFILL_3__8574_ gnd vdd FILL
XFILL_0__11229_ gnd vdd FILL
XFILL_2__14927_ gnd vdd FILL
XFILL_6__14308_ gnd vdd FILL
XFILL_1__13568_ gnd vdd FILL
XFILL_0__7816_ gnd vdd FILL
X_9143_ _9141_/Y _9101_/B _9143_/C gnd _9143_/Y vdd OAI21X1
XFILL_3__14128_ gnd vdd FILL
XFILL_1__15307_ gnd vdd FILL
XFILL_2__14858_ gnd vdd FILL
XFILL_4__13679_ gnd vdd FILL
XFILL_1__12519_ gnd vdd FILL
XFILL_1__16287_ gnd vdd FILL
XFILL_6__7234_ gnd vdd FILL
XFILL_1__13499_ gnd vdd FILL
X_9074_ _9034_/A _8306_/CLK _7533_/R vdd _9036_/Y gnd vdd DFFSR
XFILL_0__7747_ gnd vdd FILL
XFILL_4__15418_ gnd vdd FILL
XFILL_3_BUFX2_insert408 gnd vdd FILL
XFILL_2__13809_ gnd vdd FILL
XSFILL33880x49050 gnd vdd FILL
XFILL_3__14059_ gnd vdd FILL
XFILL_5__14969_ gnd vdd FILL
XFILL_1__15238_ gnd vdd FILL
XFILL_3__7456_ gnd vdd FILL
XFILL_3_BUFX2_insert419 gnd vdd FILL
XFILL_4__16398_ gnd vdd FILL
XFILL_2__14789_ gnd vdd FILL
XFILL_0__15968_ gnd vdd FILL
XFILL111800x27050 gnd vdd FILL
X_8025_ _8025_/Q _8025_/CLK _8025_/R vdd _8025_/D gnd vdd DFFSR
XFILL_4__15349_ gnd vdd FILL
XFILL_0__7678_ gnd vdd FILL
XSFILL104440x81050 gnd vdd FILL
XFILL_1__15169_ gnd vdd FILL
XFILL_0__14919_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1080 gnd vdd FILL
XFILL_0__9417_ gnd vdd FILL
XFILL_1__8210_ gnd vdd FILL
XSFILL64200x19050 gnd vdd FILL
XFILL_0__15899_ gnd vdd FILL
XFILL_3__9126_ gnd vdd FILL
XFILL_1__8141_ gnd vdd FILL
XFILL_0__9348_ gnd vdd FILL
X_9976_ _9974_/Y _9975_/B _9976_/C gnd _9976_/Y vdd OAI21X1
XFILL_0__9279_ gnd vdd FILL
XFILL_1__8072_ gnd vdd FILL
X_8927_ _8927_/Q _7007_/CLK _8047_/R vdd _8927_/D gnd vdd DFFSR
XFILL_3__8008_ gnd vdd FILL
XFILL_4__9870_ gnd vdd FILL
XSFILL94280x14050 gnd vdd FILL
XFILL112120x7050 gnd vdd FILL
XFILL_4_CLKBUF1_insert209 gnd vdd FILL
X_8858_ _8930_/Q gnd _8860_/A vdd INVX1
X_7809_ _7807_/Y _7872_/B _7809_/C gnd _7897_/D vdd OAI21X1
XFILL_0_BUFX2_insert309 gnd vdd FILL
X_8789_ _8789_/A _8788_/A _8789_/C gnd _8821_/D vdd OAI21X1
XFILL_4__8752_ gnd vdd FILL
XSFILL33960x29050 gnd vdd FILL
XFILL_6__9668_ gnd vdd FILL
XFILL_1__8974_ gnd vdd FILL
XFILL_4__7703_ gnd vdd FILL
X_11410_ _11185_/C gnd _11411_/C vdd INVX1
XFILL_6__8619_ gnd vdd FILL
X_12390_ _12390_/A _12422_/A _12390_/C gnd _12390_/Y vdd OAI21X1
XFILL_4__7634_ gnd vdd FILL
X_11341_ _10991_/Y _11341_/B _11340_/Y gnd _11341_/Y vdd OAI21X1
XFILL_1__7856_ gnd vdd FILL
XFILL_4__7565_ gnd vdd FILL
X_14060_ _8986_/A gnd _14060_/Y vdd INVX1
X_11272_ _12262_/Y gnd _11274_/A vdd INVX1
XFILL_4_BUFX2_insert231 gnd vdd FILL
XFILL_4_BUFX2_insert242 gnd vdd FILL
XFILL_4_BUFX2_insert253 gnd vdd FILL
XFILL_4_BUFX2_insert264 gnd vdd FILL
X_13011_ _6890_/A gnd _13011_/Y vdd INVX1
XFILL_4__7496_ gnd vdd FILL
XFILL_4_BUFX2_insert275 gnd vdd FILL
X_10223_ _10177_/A _7647_/CLK _9056_/R vdd _10223_/D gnd vdd DFFSR
XFILL_1__9526_ gnd vdd FILL
XFILL_4_BUFX2_insert286 gnd vdd FILL
XFILL_4__9235_ gnd vdd FILL
XFILL_4_BUFX2_insert297 gnd vdd FILL
XSFILL28920x18050 gnd vdd FILL
XFILL_3_BUFX2_insert920 gnd vdd FILL
X_10154_ _10140_/B _8874_/B gnd _10155_/C vdd NAND2X1
XFILL_3_BUFX2_insert931 gnd vdd FILL
XFILL_2__8250_ gnd vdd FILL
XFILL_3_BUFX2_insert942 gnd vdd FILL
XSFILL13720x60050 gnd vdd FILL
XFILL_4__9166_ gnd vdd FILL
XFILL_3_BUFX2_insert953 gnd vdd FILL
XSFILL79160x55050 gnd vdd FILL
XFILL_3_BUFX2_insert964 gnd vdd FILL
XSFILL28520x20050 gnd vdd FILL
XFILL_2__7201_ gnd vdd FILL
XFILL_3_BUFX2_insert975 gnd vdd FILL
X_14962_ _14960_/Y _14697_/C _14640_/C _14961_/Y gnd _14962_/Y vdd OAI22X1
XFILL_3_BUFX2_insert986 gnd vdd FILL
X_10085_ _10019_/A _7269_/CLK _9061_/R vdd _10085_/D gnd vdd DFFSR
XFILL_4__8117_ gnd vdd FILL
XFILL_3_BUFX2_insert997 gnd vdd FILL
XFILL_1__9388_ gnd vdd FILL
XFILL_4__9097_ gnd vdd FILL
X_13913_ _13911_/Y _14506_/C _14718_/B _13912_/Y gnd _13917_/B vdd OAI22X1
XFILL_5__10650_ gnd vdd FILL
XFILL_1__8339_ gnd vdd FILL
X_14893_ _9424_/A gnd _14894_/D vdd INVX1
XFILL_3_BUFX2_insert1003 gnd vdd FILL
X_13844_ _10206_/Q gnd _13844_/Y vdd INVX1
XFILL_4__11030_ gnd vdd FILL
XFILL_3_BUFX2_insert1014 gnd vdd FILL
XFILL_5__10581_ gnd vdd FILL
XFILL_3_BUFX2_insert1025 gnd vdd FILL
XFILL_2__7063_ gnd vdd FILL
XFILL_3__11760_ gnd vdd FILL
XFILL_3_BUFX2_insert1036 gnd vdd FILL
XFILL_1_BUFX2_insert110 gnd vdd FILL
XFILL_0__11580_ gnd vdd FILL
XFILL_3_BUFX2_insert1047 gnd vdd FILL
XFILL_5__12320_ gnd vdd FILL
XFILL_5__8861_ gnd vdd FILL
XSFILL99320x68050 gnd vdd FILL
X_13775_ _13773_/Y _13775_/B _13882_/B _13774_/Y gnd _13779_/A vdd OAI22X1
XFILL_6__11871_ gnd vdd FILL
XFILL_3_BUFX2_insert1058 gnd vdd FILL
XSFILL59080x22050 gnd vdd FILL
X_10987_ _10987_/Q _12692_/CLK _12692_/R vdd _10983_/Y gnd vdd DFFSR
XFILL_2__12140_ gnd vdd FILL
XFILL_3_BUFX2_insert1069 gnd vdd FILL
XFILL_0__10531_ gnd vdd FILL
XFILL_3__11691_ gnd vdd FILL
XFILL_5__7812_ gnd vdd FILL
XFILL_1__12870_ gnd vdd FILL
X_12726_ _12768_/A memoryOutData[10] gnd _12726_/Y vdd NAND2X1
X_15514_ _15632_/A _15514_/B _15514_/C gnd _15518_/A vdd OAI21X1
XFILL_6__10822_ gnd vdd FILL
XFILL_6__14590_ gnd vdd FILL
XFILL_3__13430_ gnd vdd FILL
XFILL_5__12251_ gnd vdd FILL
XFILL_4__9999_ gnd vdd FILL
XFILL_3__10642_ gnd vdd FILL
XFILL_0__13250_ gnd vdd FILL
XFILL_2__12071_ gnd vdd FILL
XFILL112280x28050 gnd vdd FILL
XFILL_4__12981_ gnd vdd FILL
XFILL_1__11821_ gnd vdd FILL
XFILL_5__7743_ gnd vdd FILL
XFILL_6__13541_ gnd vdd FILL
XFILL_0_BUFX2_insert810 gnd vdd FILL
X_15445_ _13901_/Y _15958_/B _15010_/A _15445_/D gnd _15446_/A vdd OAI22X1
XFILL_5__11202_ gnd vdd FILL
X_12657_ _12693_/Q gnd _12657_/Y vdd INVX1
XFILL_4__14720_ gnd vdd FILL
XFILL_5__12182_ gnd vdd FILL
XFILL_0_BUFX2_insert821 gnd vdd FILL
XFILL_3__13361_ gnd vdd FILL
XFILL_4__11932_ gnd vdd FILL
XFILL_0_BUFX2_insert832 gnd vdd FILL
XFILL_0__12201_ gnd vdd FILL
XFILL_2__11022_ gnd vdd FILL
XFILL_3__10573_ gnd vdd FILL
XFILL_1__14540_ gnd vdd FILL
XFILL_2__7965_ gnd vdd FILL
XFILL_0_BUFX2_insert843 gnd vdd FILL
XFILL_1__11752_ gnd vdd FILL
XFILL_0_BUFX2_insert854 gnd vdd FILL
XFILL_3__15100_ gnd vdd FILL
XFILL_0__10393_ gnd vdd FILL
X_11608_ _11608_/A _11608_/B gnd _11608_/Y vdd NOR2X1
XFILL_5__7674_ gnd vdd FILL
XFILL_5__11133_ gnd vdd FILL
X_15376_ _13866_/Y _15376_/B gnd _15379_/C vdd NOR2X1
XSFILL13800x40050 gnd vdd FILL
XFILL_3__12312_ gnd vdd FILL
XFILL_0_BUFX2_insert865 gnd vdd FILL
X_12588_ _12588_/A gnd _12590_/A vdd INVX1
XFILL_2__6916_ gnd vdd FILL
XFILL_0_BUFX2_insert876 gnd vdd FILL
XFILL_0__6980_ gnd vdd FILL
XFILL_4__14651_ gnd vdd FILL
XFILL_3__16080_ gnd vdd FILL
XFILL_1_BUFX2_insert1040 gnd vdd FILL
XFILL_3__13292_ gnd vdd FILL
XFILL_1__10703_ gnd vdd FILL
XFILL_0_BUFX2_insert887 gnd vdd FILL
XFILL_2__15830_ gnd vdd FILL
XFILL_4__11863_ gnd vdd FILL
XFILL_0__12132_ gnd vdd FILL
XFILL_1__14471_ gnd vdd FILL
XFILL_5__9413_ gnd vdd FILL
XFILL_1_BUFX2_insert1051 gnd vdd FILL
XFILL_0_BUFX2_insert898 gnd vdd FILL
XFILL_6__12423_ gnd vdd FILL
XFILL_1_BUFX2_insert1062 gnd vdd FILL
X_14327_ _13879_/B _14325_/Y _14640_/C _15790_/B gnd _14327_/Y vdd OAI22X1
XFILL_1__11683_ gnd vdd FILL
XFILL_4__13602_ gnd vdd FILL
XFILL_1_BUFX2_insert1073 gnd vdd FILL
XFILL_6__16191_ gnd vdd FILL
XFILL_3__15031_ gnd vdd FILL
XFILL_5__15941_ gnd vdd FILL
XFILL_3_BUFX2_insert14 gnd vdd FILL
X_11539_ _11538_/Y _11544_/A _11107_/B gnd _11539_/Y vdd OAI21X1
XFILL_5__11064_ gnd vdd FILL
XFILL_4__10814_ gnd vdd FILL
XFILL_1_BUFX2_insert1084 gnd vdd FILL
XFILL_1__16210_ gnd vdd FILL
XFILL_3__12243_ gnd vdd FILL
XFILL_3_BUFX2_insert25 gnd vdd FILL
XFILL_4__14582_ gnd vdd FILL
XFILL_2__9635_ gnd vdd FILL
XFILL_3_BUFX2_insert36 gnd vdd FILL
XFILL_1__13422_ gnd vdd FILL
XFILL_2__6847_ gnd vdd FILL
XFILL_4__11794_ gnd vdd FILL
XFILL_2__15761_ gnd vdd FILL
XFILL_2__12973_ gnd vdd FILL
XFILL_1__10634_ gnd vdd FILL
XFILL_0__12063_ gnd vdd FILL
XFILL_3_BUFX2_insert47 gnd vdd FILL
XSFILL69160x8050 gnd vdd FILL
XFILL_5__9344_ gnd vdd FILL
XFILL_5__10015_ gnd vdd FILL
XFILL_6__15142_ gnd vdd FILL
X_14258_ _7526_/Q gnd _14258_/Y vdd INVX1
XFILL_0__8650_ gnd vdd FILL
XFILL_4__16321_ gnd vdd FILL
XFILL_3_BUFX2_insert58 gnd vdd FILL
XFILL_3_BUFX2_insert69 gnd vdd FILL
XFILL_2__14712_ gnd vdd FILL
XFILL_5__15872_ gnd vdd FILL
XFILL_4__10745_ gnd vdd FILL
XFILL_4__13533_ gnd vdd FILL
XFILL_2__11924_ gnd vdd FILL
XFILL_3__12174_ gnd vdd FILL
XFILL_0__11014_ gnd vdd FILL
XFILL_1__16141_ gnd vdd FILL
XFILL_1__13353_ gnd vdd FILL
XFILL_2__15692_ gnd vdd FILL
XSFILL84360x26050 gnd vdd FILL
X_13209_ _13220_/A _13209_/B gnd _13209_/Y vdd NOR2X1
XFILL_5__9275_ gnd vdd FILL
XFILL_1__10565_ gnd vdd FILL
XFILL_0__7601_ gnd vdd FILL
XFILL_5__14823_ gnd vdd FILL
XFILL_3__7310_ gnd vdd FILL
X_14189_ _14187_/Y _14636_/C _14555_/C _14188_/Y gnd _14193_/B vdd OAI22X1
XFILL_2__8517_ gnd vdd FILL
XFILL_3__11125_ gnd vdd FILL
XFILL_0__8581_ gnd vdd FILL
XFILL_4__16252_ gnd vdd FILL
XFILL_6__12285_ gnd vdd FILL
XFILL_2__14643_ gnd vdd FILL
XFILL_4__13464_ gnd vdd FILL
XFILL_1__12304_ gnd vdd FILL
XFILL_4__10676_ gnd vdd FILL
XFILL_6_CLKBUF1_insert142 gnd vdd FILL
XFILL_2__9497_ gnd vdd FILL
XFILL_5__8226_ gnd vdd FILL
XFILL_0__15822_ gnd vdd FILL
XFILL_1__16072_ gnd vdd FILL
XFILL_2__11855_ gnd vdd FILL
XFILL_1__13284_ gnd vdd FILL
XFILL_1__10496_ gnd vdd FILL
XSFILL18520x52050 gnd vdd FILL
XSFILL99400x48050 gnd vdd FILL
XFILL_4__15203_ gnd vdd FILL
XSFILL84360x2050 gnd vdd FILL
XFILL_6__11236_ gnd vdd FILL
XFILL_4__12415_ gnd vdd FILL
XFILL_5__14754_ gnd vdd FILL
XFILL_2__10806_ gnd vdd FILL
XFILL_2__8448_ gnd vdd FILL
XFILL_4__16183_ gnd vdd FILL
XFILL_5__11966_ gnd vdd FILL
XFILL_3__15933_ gnd vdd FILL
XFILL_1__15023_ gnd vdd FILL
XFILL_4__13395_ gnd vdd FILL
XFILL_3__11056_ gnd vdd FILL
XFILL_3__7241_ gnd vdd FILL
XFILL_2__14574_ gnd vdd FILL
XFILL_1__12235_ gnd vdd FILL
XFILL_2__11786_ gnd vdd FILL
XFILL_0__15753_ gnd vdd FILL
XFILL_0__12965_ gnd vdd FILL
XFILL_5__13705_ gnd vdd FILL
XFILL_0__7463_ gnd vdd FILL
XFILL_5__10917_ gnd vdd FILL
XFILL_3__10007_ gnd vdd FILL
XFILL_4__12346_ gnd vdd FILL
XFILL_2__16313_ gnd vdd FILL
XFILL_4__15134_ gnd vdd FILL
XFILL_5__14685_ gnd vdd FILL
XFILL_2__13525_ gnd vdd FILL
XFILL_2__8379_ gnd vdd FILL
XFILL_5__11897_ gnd vdd FILL
XFILL_3__7172_ gnd vdd FILL
XFILL_0__14704_ gnd vdd FILL
XFILL_5__7108_ gnd vdd FILL
XFILL_3__15864_ gnd vdd FILL
XFILL_0__11916_ gnd vdd FILL
XFILL_1__12166_ gnd vdd FILL
XFILL_0__15684_ gnd vdd FILL
XFILL_5__8088_ gnd vdd FILL
X_9830_ _9766_/A _8038_/CLK _8038_/R vdd _9768_/Y gnd vdd DFFSR
XFILL_5__13636_ gnd vdd FILL
XFILL_0__12896_ gnd vdd FILL
XSFILL44680x3050 gnd vdd FILL
XFILL_2__16244_ gnd vdd FILL
XFILL_3__14815_ gnd vdd FILL
XFILL_4__15065_ gnd vdd FILL
XFILL_4__12277_ gnd vdd FILL
XFILL_6__11098_ gnd vdd FILL
XFILL_2__13456_ gnd vdd FILL
XFILL_1__11117_ gnd vdd FILL
XFILL_5__7039_ gnd vdd FILL
XFILL_0__14635_ gnd vdd FILL
XFILL_1__12097_ gnd vdd FILL
XFILL_3__15795_ gnd vdd FILL
XFILL_2__10668_ gnd vdd FILL
XFILL_0__9133_ gnd vdd FILL
XFILL_0__11847_ gnd vdd FILL
XSFILL49080x54050 gnd vdd FILL
XFILL_5__16355_ gnd vdd FILL
XFILL_4__14016_ gnd vdd FILL
XFILL_4__11228_ gnd vdd FILL
XFILL_2__12407_ gnd vdd FILL
X_9761_ _9741_/B _9633_/B gnd _9762_/C vdd NAND2X1
XFILL_5__13567_ gnd vdd FILL
X_6973_ _6971_/Y _6951_/A _6972_/Y gnd _7021_/D vdd OAI21X1
XFILL_1__15925_ gnd vdd FILL
XFILL_2__16175_ gnd vdd FILL
XFILL_3__11958_ gnd vdd FILL
XFILL_5__10779_ gnd vdd FILL
XFILL_1__11048_ gnd vdd FILL
XFILL_3__14746_ gnd vdd FILL
XFILL_2__13387_ gnd vdd FILL
XFILL_0__14566_ gnd vdd FILL
XFILL_5__15306_ gnd vdd FILL
X_8712_ _8796_/Q gnd _8714_/A vdd INVX1
XFILL_5__12518_ gnd vdd FILL
XFILL_0__11778_ gnd vdd FILL
XFILL_3__10909_ gnd vdd FILL
XFILL_5__16286_ gnd vdd FILL
XFILL_4__11159_ gnd vdd FILL
XFILL_2__15126_ gnd vdd FILL
X_9692_ _9608_/A _8046_/CLK _9692_/R vdd _9692_/D gnd vdd DFFSR
XFILL_0__16305_ gnd vdd FILL
XFILL_2__12338_ gnd vdd FILL
XFILL_5__13498_ gnd vdd FILL
XSFILL114520x24050 gnd vdd FILL
XFILL_6_BUFX2_insert326 gnd vdd FILL
XFILL_3__11889_ gnd vdd FILL
XFILL_1__15856_ gnd vdd FILL
XFILL_3__14677_ gnd vdd FILL
XFILL_0__13517_ gnd vdd FILL
XFILL_0__8015_ gnd vdd FILL
XFILL_0__14497_ gnd vdd FILL
XFILL_5__15237_ gnd vdd FILL
XFILL_5__12449_ gnd vdd FILL
XFILL_3__16416_ gnd vdd FILL
X_8643_ _8641_/Y _8607_/B _8643_/C gnd _8643_/Y vdd OAI21X1
XFILL_3__13628_ gnd vdd FILL
XFILL_1__14807_ gnd vdd FILL
XFILL_2__15057_ gnd vdd FILL
XFILL_4__15967_ gnd vdd FILL
XFILL_3__9813_ gnd vdd FILL
XFILL_0__16236_ gnd vdd FILL
XFILL_2__12269_ gnd vdd FILL
XFILL_0__13448_ gnd vdd FILL
XFILL_1__15787_ gnd vdd FILL
XFILL_1__12999_ gnd vdd FILL
XFILL_5__15168_ gnd vdd FILL
XFILL_2__14008_ gnd vdd FILL
XFILL_4__14918_ gnd vdd FILL
XFILL_3__16347_ gnd vdd FILL
XSFILL69240x67050 gnd vdd FILL
XFILL_3__13559_ gnd vdd FILL
X_8574_ _8574_/A _8619_/B _8574_/C gnd _8664_/D vdd OAI21X1
XFILL_3__9744_ gnd vdd FILL
XFILL_4__15898_ gnd vdd FILL
XFILL_3__6956_ gnd vdd FILL
XFILL_1__14738_ gnd vdd FILL
XFILL_0__16167_ gnd vdd FILL
XFILL_0__13379_ gnd vdd FILL
XFILL_5__14119_ gnd vdd FILL
X_7525_ _7459_/A _8165_/CLK _8165_/R vdd _7525_/D gnd vdd DFFSR
XFILL_4__14849_ gnd vdd FILL
XFILL_5__15099_ gnd vdd FILL
XFILL_0__15118_ gnd vdd FILL
XFILL_3__16278_ gnd vdd FILL
XFILL_3__9675_ gnd vdd FILL
XFILL_1__14669_ gnd vdd FILL
XFILL_3__6887_ gnd vdd FILL
XSFILL104440x76050 gnd vdd FILL
XFILL_0__16098_ gnd vdd FILL
XFILL_1__7710_ gnd vdd FILL
XFILL_6__9384_ gnd vdd FILL
XFILL_0__8917_ gnd vdd FILL
XFILL_1__16408_ gnd vdd FILL
XFILL_3__15229_ gnd vdd FILL
X_7456_ _7456_/A gnd _7456_/Y vdd INVX1
XFILL_0__9897_ gnd vdd FILL
XSFILL8680x74050 gnd vdd FILL
XFILL_3__8626_ gnd vdd FILL
XSFILL23720x23050 gnd vdd FILL
XFILL_0__15049_ gnd vdd FILL
XFILL_2__15959_ gnd vdd FILL
XFILL_6__8335_ gnd vdd FILL
XFILL_0__8848_ gnd vdd FILL
XFILL_4__7350_ gnd vdd FILL
XFILL_1__16339_ gnd vdd FILL
X_7387_ _7301_/A _9447_/CLK _9447_/R vdd _7387_/D gnd vdd DFFSR
X_9126_ _9190_/Q gnd _9126_/Y vdd INVX1
XFILL_0__8779_ gnd vdd FILL
XFILL_3__7508_ gnd vdd FILL
XFILL_1__7572_ gnd vdd FILL
XFILL_3__8488_ gnd vdd FILL
XFILL_3_BUFX2_insert227 gnd vdd FILL
XFILL_4__9020_ gnd vdd FILL
X_9057_ _9057_/Q _9453_/CLK _9453_/R vdd _8985_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert238 gnd vdd FILL
XFILL_3__7439_ gnd vdd FILL
XFILL_3_BUFX2_insert249 gnd vdd FILL
XSFILL13640x75050 gnd vdd FILL
XFILL_1__9242_ gnd vdd FILL
X_8008_ _7997_/B _8008_/B gnd _8008_/Y vdd NAND2X1
XFILL_2_BUFX2_insert905 gnd vdd FILL
XFILL_2_BUFX2_insert916 gnd vdd FILL
XFILL_6__7079_ gnd vdd FILL
XFILL_2_BUFX2_insert927 gnd vdd FILL
XFILL_2_BUFX2_insert938 gnd vdd FILL
XFILL_3__9109_ gnd vdd FILL
XFILL_1__9173_ gnd vdd FILL
XFILL_2_BUFX2_insert949 gnd vdd FILL
X_10910_ _10897_/Y _10910_/B _10944_/A gnd _10911_/C vdd OAI21X1
XFILL_1__8124_ gnd vdd FILL
X_11890_ _11890_/A gnd _11892_/A vdd INVX1
X_9959_ _9897_/A _8551_/CLK _9959_/R vdd _9959_/D gnd vdd DFFSR
XSFILL104520x56050 gnd vdd FILL
XFILL_4__9922_ gnd vdd FILL
X_10841_ _10751_/A _9817_/CLK _8942_/R vdd _10841_/D gnd vdd DFFSR
XSFILL73960x31050 gnd vdd FILL
XSFILL8760x54050 gnd vdd FILL
XFILL_1__8055_ gnd vdd FILL
XSFILL73400x74050 gnd vdd FILL
XFILL_4__9853_ gnd vdd FILL
X_13560_ _13559_/Y _13560_/B gnd _13584_/A vdd NOR2X1
X_10772_ _10848_/Q gnd _10772_/Y vdd INVX1
XBUFX2_insert904 _10913_/Y gnd _12768_/A vdd BUFX2
X_12511_ _12083_/B gnd _12511_/Y vdd INVX1
XFILL_0_BUFX2_insert106 gnd vdd FILL
XBUFX2_insert915 _12360_/Y gnd _6918_/B vdd BUFX2
XFILL_4__6996_ gnd vdd FILL
XFILL_4__9784_ gnd vdd FILL
XBUFX2_insert926 _12351_/Y gnd _9597_/B vdd BUFX2
XBUFX2_insert937 _13423_/Y gnd _14320_/C vdd BUFX2
X_13491_ _7511_/Q gnd _13491_/Y vdd INVX1
XBUFX2_insert948 _11987_/Y gnd _12105_/B vdd BUFX2
X_15230_ _15229_/Y _15230_/B gnd _15259_/B vdd NOR2X1
XBUFX2_insert959 _13361_/Y gnd _10450_/B vdd BUFX2
XFILL_4__8735_ gnd vdd FILL
X_12442_ _11991_/B gnd _12442_/Y vdd INVX1
XSFILL68600x4050 gnd vdd FILL
XSFILL63880x83050 gnd vdd FILL
XFILL_2__7750_ gnd vdd FILL
XSFILL13720x55050 gnd vdd FILL
XFILL_1__8957_ gnd vdd FILL
X_15161_ _8280_/Q gnd _15162_/B vdd INVX1
X_12373_ _12027_/B gnd _12373_/Y vdd INVX1
XFILL_2__7681_ gnd vdd FILL
XFILL_1__8888_ gnd vdd FILL
XFILL_4__7617_ gnd vdd FILL
X_14112_ _9373_/A _13883_/B _14112_/C gnd _14112_/Y vdd AOI21X1
XFILL_4__8597_ gnd vdd FILL
X_11324_ _11494_/A _11498_/A gnd _11324_/Y vdd NAND2X1
XFILL_2__9420_ gnd vdd FILL
X_15092_ _15239_/B gnd _15357_/B vdd INVX4
XFILL_1__7839_ gnd vdd FILL
XSFILL28920x5050 gnd vdd FILL
XFILL_4__7548_ gnd vdd FILL
X_14043_ _14043_/A gnd _14045_/D vdd INVX1
XFILL_4__10530_ gnd vdd FILL
X_11255_ _11019_/Y _11254_/Y _11383_/A gnd _11256_/C vdd AOI21X1
XFILL_2__9351_ gnd vdd FILL
XSFILL8840x34050 gnd vdd FILL
X_10206_ _10206_/Q _8025_/CLK _7262_/R vdd _10206_/D gnd vdd DFFSR
XFILL_4__7479_ gnd vdd FILL
XFILL_6__12070_ gnd vdd FILL
XFILL_5__11820_ gnd vdd FILL
XFILL_1__9509_ gnd vdd FILL
XSFILL7800x70050 gnd vdd FILL
X_11186_ _12189_/Y _11180_/Y gnd _11186_/Y vdd NAND2X1
XSFILL59080x17050 gnd vdd FILL
XFILL_5__8011_ gnd vdd FILL
XFILL_2__11640_ gnd vdd FILL
XFILL_2__9282_ gnd vdd FILL
XFILL_4__9218_ gnd vdd FILL
XFILL_1__10281_ gnd vdd FILL
XFILL_3_BUFX2_insert750 gnd vdd FILL
XFILL_4__12200_ gnd vdd FILL
XSFILL99480x22050 gnd vdd FILL
XFILL_6__11021_ gnd vdd FILL
X_10137_ _10137_/A _10169_/A _10137_/C gnd _10209_/D vdd OAI21X1
XFILL_3_BUFX2_insert761 gnd vdd FILL
XFILL_5__11751_ gnd vdd FILL
XSFILL74120x20050 gnd vdd FILL
XFILL_2__8233_ gnd vdd FILL
X_15994_ _15994_/A _15993_/Y gnd _16005_/C vdd NAND2X1
XFILL_1__12020_ gnd vdd FILL
XFILL_4__10392_ gnd vdd FILL
XFILL_3_BUFX2_insert772 gnd vdd FILL
XFILL_4__9149_ gnd vdd FILL
XFILL_3_BUFX2_insert783 gnd vdd FILL
XFILL_2__11571_ gnd vdd FILL
XFILL_0__12750_ gnd vdd FILL
XFILL_3_BUFX2_insert794 gnd vdd FILL
XFILL_5__10702_ gnd vdd FILL
XFILL_4__12131_ gnd vdd FILL
XFILL_2__13310_ gnd vdd FILL
XFILL_5__14470_ gnd vdd FILL
X_10068_ _9993_/A _9556_/B gnd _10069_/C vdd NAND2X1
X_14945_ _9811_/A gnd _14945_/Y vdd INVX1
XFILL_2__10522_ gnd vdd FILL
XFILL_3__12861_ gnd vdd FILL
XFILL_5__11682_ gnd vdd FILL
XFILL_2__14290_ gnd vdd FILL
XFILL_0__11701_ gnd vdd FILL
XFILL_5__13421_ gnd vdd FILL
XFILL_2__7115_ gnd vdd FILL
XFILL_3__14600_ gnd vdd FILL
XFILL_5__10633_ gnd vdd FILL
XFILL_4__12062_ gnd vdd FILL
XSFILL13800x35050 gnd vdd FILL
XFILL_3__11812_ gnd vdd FILL
XFILL_2__13241_ gnd vdd FILL
X_14876_ _14876_/A _14876_/B gnd _14879_/C vdd NOR2X1
XFILL_2__10453_ gnd vdd FILL
XFILL_0__14420_ gnd vdd FILL
XFILL_2__8095_ gnd vdd FILL
XFILL_3__15580_ gnd vdd FILL
XFILL_0__11632_ gnd vdd FILL
XFILL_1__13971_ gnd vdd FILL
XFILL_5__8913_ gnd vdd FILL
XFILL_4__11013_ gnd vdd FILL
XFILL_5__16140_ gnd vdd FILL
XFILL_5__13352_ gnd vdd FILL
XFILL_5__9893_ gnd vdd FILL
X_13827_ _14868_/A _10717_/Q _10763_/A _14877_/D gnd _13838_/A vdd AOI22X1
XFILL_1__15710_ gnd vdd FILL
XFILL_3__14531_ gnd vdd FILL
XFILL_5__10564_ gnd vdd FILL
XFILL_2__7046_ gnd vdd FILL
XFILL_3__11743_ gnd vdd FILL
XSFILL64040x72050 gnd vdd FILL
XFILL_2__13172_ gnd vdd FILL
XFILL_2__10384_ gnd vdd FILL
XFILL_0__14351_ gnd vdd FILL
XFILL_0__11563_ gnd vdd FILL
XFILL_5__8844_ gnd vdd FILL
XFILL_5__12303_ gnd vdd FILL
X_13758_ _13871_/A _13758_/B _13850_/B _13758_/D gnd _13758_/Y vdd OAI22X1
XFILL_4__15821_ gnd vdd FILL
XFILL_5__16071_ gnd vdd FILL
XFILL_5__13283_ gnd vdd FILL
XFILL_5__10495_ gnd vdd FILL
XFILL_3__14462_ gnd vdd FILL
XFILL_2__12123_ gnd vdd FILL
XFILL_0__13302_ gnd vdd FILL
XFILL_1__15641_ gnd vdd FILL
XFILL_3__11674_ gnd vdd FILL
XFILL_0__10514_ gnd vdd FILL
XFILL_1__12853_ gnd vdd FILL
X_12709_ _12709_/A _10944_/C _12709_/C gnd _12795_/D vdd OAI21X1
XFILL_5__15022_ gnd vdd FILL
XFILL_0__11494_ gnd vdd FILL
XFILL_0__14282_ gnd vdd FILL
XFILL_3__16201_ gnd vdd FILL
XFILL_3__13413_ gnd vdd FILL
XFILL_5__12234_ gnd vdd FILL
XFILL_5__8775_ gnd vdd FILL
XFILL_3__10625_ gnd vdd FILL
XSFILL43880x30050 gnd vdd FILL
X_13689_ _13689_/A _14320_/C gnd _13690_/C vdd NOR2X1
XFILL_4__15752_ gnd vdd FILL
XFILL_0__16021_ gnd vdd FILL
XFILL_4__12964_ gnd vdd FILL
XFILL_2__12054_ gnd vdd FILL
XFILL_3__14393_ gnd vdd FILL
XFILL_1__11804_ gnd vdd FILL
XFILL_0__13233_ gnd vdd FILL
XFILL_0__10445_ gnd vdd FILL
XFILL_1__15572_ gnd vdd FILL
XFILL_1__12784_ gnd vdd FILL
XFILL_2__8997_ gnd vdd FILL
XFILL_5__7726_ gnd vdd FILL
XFILL_0_BUFX2_insert640 gnd vdd FILL
XFILL_0_BUFX2_insert651 gnd vdd FILL
XFILL_4__14703_ gnd vdd FILL
X_15428_ _15225_/A _7647_/Q _7441_/A _15383_/D gnd _15433_/B vdd AOI22X1
XFILL_3__13344_ gnd vdd FILL
XFILL_4__11915_ gnd vdd FILL
XFILL_5__12165_ gnd vdd FILL
XFILL_0_BUFX2_insert662 gnd vdd FILL
XFILL_2__11005_ gnd vdd FILL
XFILL_3__16132_ gnd vdd FILL
XFILL_4__15683_ gnd vdd FILL
XFILL_3__10556_ gnd vdd FILL
XFILL_1__14523_ gnd vdd FILL
XFILL_2__7948_ gnd vdd FILL
XFILL_4__12895_ gnd vdd FILL
XFILL_0__13164_ gnd vdd FILL
XFILL_0_BUFX2_insert673 gnd vdd FILL
XFILL_1__11735_ gnd vdd FILL
XFILL_0__10376_ gnd vdd FILL
XFILL_0_BUFX2_insert684 gnd vdd FILL
XFILL_0_BUFX2_insert695 gnd vdd FILL
X_7310_ _7390_/Q gnd _7312_/A vdd INVX1
X_15359_ _16002_/C _15358_/Y _13808_/Y _15912_/D gnd _15359_/Y vdd OAI22X1
XFILL_0__9751_ gnd vdd FILL
XFILL_5__11116_ gnd vdd FILL
XFILL_4__14634_ gnd vdd FILL
XSFILL99000x45050 gnd vdd FILL
XFILL_5__12096_ gnd vdd FILL
XFILL_6__10667_ gnd vdd FILL
XFILL_0__6963_ gnd vdd FILL
XFILL_3__16063_ gnd vdd FILL
XFILL_3__13275_ gnd vdd FILL
XFILL_0__12115_ gnd vdd FILL
X_8290_ _8290_/Q _7010_/CLK _7413_/R vdd _8290_/D gnd vdd DFFSR
XFILL_2__15813_ gnd vdd FILL
XFILL_4__11846_ gnd vdd FILL
XFILL_1__14454_ gnd vdd FILL
XFILL_3__10487_ gnd vdd FILL
XFILL_2__7879_ gnd vdd FILL
XFILL_0__13095_ gnd vdd FILL
XFILL_0__8702_ gnd vdd FILL
XFILL_1__11666_ gnd vdd FILL
XFILL_5__15924_ gnd vdd FILL
XFILL_5__7588_ gnd vdd FILL
XFILL_3__15014_ gnd vdd FILL
XSFILL23640x38050 gnd vdd FILL
XFILL_5__11047_ gnd vdd FILL
XFILL_3__12226_ gnd vdd FILL
XFILL_0__9682_ gnd vdd FILL
X_7241_ _7241_/A _7210_/A _7240_/Y gnd _7281_/D vdd OAI21X1
XFILL_4__14565_ gnd vdd FILL
XFILL_1__13405_ gnd vdd FILL
XFILL_0__6894_ gnd vdd FILL
XFILL_2__9618_ gnd vdd FILL
XFILL_0__12046_ gnd vdd FILL
XFILL_3__9391_ gnd vdd FILL
XFILL_1__10617_ gnd vdd FILL
XFILL_2__12956_ gnd vdd FILL
XFILL_4__11777_ gnd vdd FILL
XFILL_2__15744_ gnd vdd FILL
XFILL_1__14385_ gnd vdd FILL
XFILL_0__8633_ gnd vdd FILL
XFILL_4__16304_ gnd vdd FILL
XFILL_1__11597_ gnd vdd FILL
X_7172_ _7172_/A _7181_/B _7172_/C gnd _7172_/Y vdd OAI21X1
XFILL_5__15855_ gnd vdd FILL
XFILL_4__13516_ gnd vdd FILL
XFILL112200x67050 gnd vdd FILL
XFILL_2__11907_ gnd vdd FILL
XFILL_3__12157_ gnd vdd FILL
XFILL_1__16124_ gnd vdd FILL
XFILL_3__8342_ gnd vdd FILL
XFILL_2__9549_ gnd vdd FILL
XFILL_1__13336_ gnd vdd FILL
XFILL_2__15675_ gnd vdd FILL
XFILL_4__14496_ gnd vdd FILL
XFILL_2__12887_ gnd vdd FILL
XFILL_1__10548_ gnd vdd FILL
XFILL_5__14806_ gnd vdd FILL
XFILL_5__9258_ gnd vdd FILL
XFILL_4__16235_ gnd vdd FILL
XSFILL64120x52050 gnd vdd FILL
XFILL_3__11108_ gnd vdd FILL
XFILL_4__10659_ gnd vdd FILL
XFILL_2__14626_ gnd vdd FILL
XFILL_4__13447_ gnd vdd FILL
XFILL_5__15786_ gnd vdd FILL
XSFILL49480x70050 gnd vdd FILL
XFILL_5__12998_ gnd vdd FILL
XFILL_3__12088_ gnd vdd FILL
XFILL_0__15805_ gnd vdd FILL
XFILL_1__16055_ gnd vdd FILL
XFILL_3__8273_ gnd vdd FILL
XFILL_2__11838_ gnd vdd FILL
XFILL_1__13267_ gnd vdd FILL
XFILL_6__14007_ gnd vdd FILL
XFILL_5__8209_ gnd vdd FILL
XFILL_0__13997_ gnd vdd FILL
XFILL_5__14737_ gnd vdd FILL
XFILL_3__15916_ gnd vdd FILL
XFILL_4__16166_ gnd vdd FILL
XFILL_5__11949_ gnd vdd FILL
XFILL_3__7224_ gnd vdd FILL
XFILL_1__15006_ gnd vdd FILL
XFILL_0__8495_ gnd vdd FILL
XFILL_3__11039_ gnd vdd FILL
XFILL_2__14557_ gnd vdd FILL
XFILL_4__13378_ gnd vdd FILL
XFILL_1__12218_ gnd vdd FILL
XFILL_2__11769_ gnd vdd FILL
XFILL_0__15736_ gnd vdd FILL
XSFILL43960x10050 gnd vdd FILL
XFILL_0__7446_ gnd vdd FILL
XFILL_4__15117_ gnd vdd FILL
XFILL_4__12329_ gnd vdd FILL
XFILL_5__14668_ gnd vdd FILL
XFILL_2__13508_ gnd vdd FILL
XFILL_4__16097_ gnd vdd FILL
XFILL_3__15847_ gnd vdd FILL
XSFILL18600x27050 gnd vdd FILL
XFILL_2__14488_ gnd vdd FILL
XFILL_1__12149_ gnd vdd FILL
XFILL_0__15667_ gnd vdd FILL
XFILL_5__16407_ gnd vdd FILL
XSFILL28760x71050 gnd vdd FILL
XFILL_5__13619_ gnd vdd FILL
XFILL_0__12879_ gnd vdd FILL
X_9813_ _9811_/Y _9813_/B _9812_/Y gnd _9845_/D vdd OAI21X1
XFILL_4__15048_ gnd vdd FILL
XFILL_0__7377_ gnd vdd FILL
XFILL_5__14599_ gnd vdd FILL
XFILL_2__16227_ gnd vdd FILL
XFILL_2__13439_ gnd vdd FILL
XFILL_0__14618_ gnd vdd FILL
XFILL_3__15778_ gnd vdd FILL
XFILL_3__7086_ gnd vdd FILL
XFILL_0__9116_ gnd vdd FILL
XFILL_5__16338_ gnd vdd FILL
XFILL_0__15598_ gnd vdd FILL
X_9744_ _9742_/Y _9764_/A _9744_/C gnd _9822_/D vdd OAI21X1
XFILL_6_BUFX2_insert101 gnd vdd FILL
XFILL_3__14729_ gnd vdd FILL
X_6956_ _6956_/A gnd _6956_/Y vdd INVX1
XFILL_2__16158_ gnd vdd FILL
XFILL_6__15889_ gnd vdd FILL
XSFILL8680x69050 gnd vdd FILL
XFILL_1__15908_ gnd vdd FILL
XSFILL23720x18050 gnd vdd FILL
XFILL_0__14549_ gnd vdd FILL
XSFILL33880x62050 gnd vdd FILL
XFILL_2__15109_ gnd vdd FILL
XFILL_5__16269_ gnd vdd FILL
X_9675_ _9675_/A _9803_/B gnd _9676_/C vdd NAND2X1
XFILL_4__6850_ gnd vdd FILL
XFILL_2__16089_ gnd vdd FILL
XFILL_1__15839_ gnd vdd FILL
X_6887_ _6887_/A gnd memoryWriteData[17] vdd BUFX2
XFILL_1__9860_ gnd vdd FILL
X_8626_ _8626_/A gnd _8626_/Y vdd INVX1
XFILL_0__16219_ gnd vdd FILL
XFILL_5_BUFX2_insert801 gnd vdd FILL
XFILL_5_BUFX2_insert812 gnd vdd FILL
XFILL_5_BUFX2_insert823 gnd vdd FILL
XFILL_3__7988_ gnd vdd FILL
XFILL_1__9791_ gnd vdd FILL
X_8557_ _8507_/A _8306_/CLK _7533_/R vdd _8557_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert834 gnd vdd FILL
XFILL_3__9727_ gnd vdd FILL
XFILL_4__8520_ gnd vdd FILL
XFILL_5_BUFX2_insert845 gnd vdd FILL
XFILL_5_BUFX2_insert856 gnd vdd FILL
XBUFX2_insert1020 _13340_/Y gnd _9613_/B vdd BUFX2
XFILL_3__6939_ gnd vdd FILL
XBUFX2_insert1031 _13333_/Y gnd _9301_/B vdd BUFX2
XFILL_5_BUFX2_insert867 gnd vdd FILL
XBUFX2_insert1042 _13297_/Y gnd _7690_/B vdd BUFX2
XFILL_1__8742_ gnd vdd FILL
XFILL_5_BUFX2_insert878 gnd vdd FILL
X_7508_ _7416_/B _7508_/B gnd _7508_/Y vdd NAND2X1
XBUFX2_insert1053 _13527_/Y gnd _14213_/A vdd BUFX2
X_8488_ _8488_/A _8508_/A _8488_/C gnd _8488_/Y vdd OAI21X1
XFILL_4__8451_ gnd vdd FILL
XFILL_5_BUFX2_insert889 gnd vdd FILL
XBUFX2_insert1064 _14992_/Y gnd _15204_/A vdd BUFX2
XFILL_3__9658_ gnd vdd FILL
XBUFX2_insert1086 rst gnd BUFX2_insert518/A vdd BUFX2
X_7439_ _7425_/B _7439_/B gnd _7439_/Y vdd NAND2X1
XFILL_3__8609_ gnd vdd FILL
XFILL_4__8382_ gnd vdd FILL
XSFILL28840x51050 gnd vdd FILL
XFILL_1__7624_ gnd vdd FILL
XSFILL99320x50 gnd vdd FILL
XFILL_4__7333_ gnd vdd FILL
X_11040_ _11037_/Y _11035_/Y _11040_/C gnd _11041_/C vdd AOI21X1
X_9109_ _9170_/B _6933_/B gnd _9110_/C vdd NAND2X1
XFILL_1__7555_ gnd vdd FILL
XSFILL8760x49050 gnd vdd FILL
XFILL_4__9003_ gnd vdd FILL
XFILL_1__7486_ gnd vdd FILL
XFILL_2_BUFX2_insert702 gnd vdd FILL
XFILL_4__7195_ gnd vdd FILL
XFILL_1__9225_ gnd vdd FILL
XFILL_2_BUFX2_insert713 gnd vdd FILL
X_12991_ vdd _12991_/B gnd _12992_/C vdd NAND2X1
XFILL_2_BUFX2_insert724 gnd vdd FILL
XFILL_2_BUFX2_insert735 gnd vdd FILL
XFILL_2_BUFX2_insert746 gnd vdd FILL
X_11942_ _11955_/B _12553_/Q gnd _11943_/C vdd NAND2X1
X_14730_ _14730_/A _14730_/B gnd _14741_/A vdd NAND2X1
XFILL_2_BUFX2_insert757 gnd vdd FILL
XFILL_2_BUFX2_insert768 gnd vdd FILL
XFILL_1__9156_ gnd vdd FILL
XFILL_2_BUFX2_insert779 gnd vdd FILL
X_14661_ _7919_/Q gnd _16079_/A vdd INVX1
XFILL_1__8107_ gnd vdd FILL
X_11873_ _12802_/Q _11874_/B gnd _11873_/Y vdd NAND2X1
XFILL_1__9087_ gnd vdd FILL
XFILL_4__9905_ gnd vdd FILL
X_13612_ _8665_/Q gnd _13612_/Y vdd INVX1
X_16400_ gnd gnd gnd _16401_/C vdd NAND2X1
X_10824_ _10797_/A _8008_/B gnd _10825_/C vdd NAND2X1
XFILL_5__6890_ gnd vdd FILL
X_14592_ _8685_/Q gnd _14592_/Y vdd INVX1
XSFILL113880x47050 gnd vdd FILL
XSFILL28920x31050 gnd vdd FILL
XBUFX2_insert701 _12420_/Y gnd _9282_/B vdd BUFX2
X_16331_ gnd gnd gnd _16332_/C vdd NAND2X1
X_13543_ _7256_/Q _13434_/B _14323_/B _8280_/Q gnd _13544_/B vdd AOI22X1
XFILL_5__10280_ gnd vdd FILL
XBUFX2_insert712 _15023_/Y gnd _15924_/B vdd BUFX2
X_10755_ _10792_/B _7555_/B gnd _10756_/C vdd NAND2X1
XBUFX2_insert723 _13352_/Y gnd _10169_/A vdd BUFX2
XBUFX2_insert734 _15020_/Y gnd _16232_/B vdd BUFX2
XFILL_2__8851_ gnd vdd FILL
XBUFX2_insert745 _15055_/Y gnd _15795_/B vdd BUFX2
XFILL_4__9767_ gnd vdd FILL
XBUFX2_insert756 _12213_/Y gnd _12248_/C vdd BUFX2
X_16262_ _9844_/Q _15390_/B _16262_/C gnd _16267_/C vdd AOI21X1
X_13474_ _13474_/A _13473_/Y gnd _13475_/A vdd NAND2X1
XFILL_3__10410_ gnd vdd FILL
XFILL_4__6979_ gnd vdd FILL
X_10686_ _14598_/A gnd _10688_/A vdd INVX1
XBUFX2_insert767 _12393_/Y gnd _9895_/B vdd BUFX2
XFILL_2__7802_ gnd vdd FILL
XFILL_2__8782_ gnd vdd FILL
XBUFX2_insert778 _10911_/Y gnd _12179_/A vdd BUFX2
XFILL_0__10230_ gnd vdd FILL
XFILL_3__11390_ gnd vdd FILL
XFILL_4__8718_ gnd vdd FILL
X_15213_ _15213_/A _15656_/B _15656_/C gnd _15215_/B vdd NOR3X1
XBUFX2_insert789 _15052_/Y gnd _15899_/C vdd BUFX2
XFILL_1__9989_ gnd vdd FILL
X_12425_ _12359_/A _12648_/A gnd _12426_/C vdd NAND2X1
XFILL_5__8491_ gnd vdd FILL
XSFILL99480x17050 gnd vdd FILL
X_16193_ _9970_/Q _16035_/B _16037_/C gnd _16194_/C vdd NAND3X1
XFILL_4__11700_ gnd vdd FILL
XFILL_2__7733_ gnd vdd FILL
XFILL_1__11520_ gnd vdd FILL
XSFILL18840x83050 gnd vdd FILL
XFILL_0__10161_ gnd vdd FILL
XFILL_5__7442_ gnd vdd FILL
X_15144_ _15144_/A _15144_/B gnd _15167_/A vdd NOR2X1
XFILL_4__8649_ gnd vdd FILL
X_12356_ _12422_/A _12667_/Q gnd _12357_/C vdd NAND2X1
XSFILL34120x31050 gnd vdd FILL
XFILL_1_CLKBUF1_insert150 gnd vdd FILL
XFILL_4__11631_ gnd vdd FILL
XFILL_5__13970_ gnd vdd FILL
XFILL_3__10272_ gnd vdd FILL
XFILL_1_CLKBUF1_insert161 gnd vdd FILL
XFILL_2__13790_ gnd vdd FILL
XFILL_1_CLKBUF1_insert172 gnd vdd FILL
XFILL_1__11451_ gnd vdd FILL
XFILL_5__7373_ gnd vdd FILL
XFILL_1_CLKBUF1_insert183 gnd vdd FILL
X_11307_ _11307_/A gnd _11308_/C vdd INVX1
XSFILL99320x81050 gnd vdd FILL
XFILL_3__12011_ gnd vdd FILL
X_15075_ _15075_/A _15074_/Y gnd _15075_/Y vdd NAND2X1
XFILL_6__13171_ gnd vdd FILL
XFILL_1_CLKBUF1_insert194 gnd vdd FILL
XFILL_6__10383_ gnd vdd FILL
XFILL_2__9403_ gnd vdd FILL
XFILL_4__14350_ gnd vdd FILL
X_12287_ _12216_/A gnd _12311_/C gnd _12287_/Y vdd NAND3X1
XFILL_4__11562_ gnd vdd FILL
XFILL_2__12741_ gnd vdd FILL
XFILL_1__10402_ gnd vdd FILL
XFILL_1__14170_ gnd vdd FILL
XFILL_2_BUFX2_insert4 gnd vdd FILL
XFILL_5__9112_ gnd vdd FILL
XFILL_2__7595_ gnd vdd FILL
XFILL_0__13920_ gnd vdd FILL
X_14026_ _7522_/Q gnd _14026_/Y vdd INVX1
XFILL_1__11382_ gnd vdd FILL
XFILL_4__13301_ gnd vdd FILL
XFILL_5__15640_ gnd vdd FILL
XFILL_4__10513_ gnd vdd FILL
X_11238_ _12222_/Y _12120_/Y gnd _11238_/Y vdd NOR2X1
XFILL_2__9334_ gnd vdd FILL
XFILL_5__12852_ gnd vdd FILL
XFILL_1__13121_ gnd vdd FILL
XFILL112280x41050 gnd vdd FILL
XFILL_4__11493_ gnd vdd FILL
XFILL_2__15460_ gnd vdd FILL
XFILL_4__14281_ gnd vdd FILL
XSFILL64040x67050 gnd vdd FILL
XFILL_5__9043_ gnd vdd FILL
XFILL_0__13851_ gnd vdd FILL
XSFILL38200x77050 gnd vdd FILL
XFILL_4__16020_ gnd vdd FILL
XFILL_5__11803_ gnd vdd FILL
XFILL_4__13232_ gnd vdd FILL
XFILL_4__10444_ gnd vdd FILL
XFILL_5__15571_ gnd vdd FILL
XFILL_2__14411_ gnd vdd FILL
X_11169_ _11166_/Y _11477_/B gnd _11480_/A vdd NOR2X1
XFILL_5__12783_ gnd vdd FILL
XFILL_2__9265_ gnd vdd FILL
XFILL_2__11623_ gnd vdd FILL
XFILL_2__15391_ gnd vdd FILL
XFILL_1__10264_ gnd vdd FILL
XFILL_3__13962_ gnd vdd FILL
XFILL_0__7300_ gnd vdd FILL
XFILL_3_BUFX2_insert580 gnd vdd FILL
XFILL_0__13782_ gnd vdd FILL
XFILL_3_BUFX2_insert591 gnd vdd FILL
XFILL_5__14522_ gnd vdd FILL
XSFILL49080x7050 gnd vdd FILL
XFILL_3__15701_ gnd vdd FILL
XFILL_4__13163_ gnd vdd FILL
XFILL_2__8216_ gnd vdd FILL
XFILL_5__11734_ gnd vdd FILL
XFILL_0__10994_ gnd vdd FILL
X_15977_ _7277_/Q _15177_/B gnd _15983_/A vdd NAND2X1
XFILL_1__12003_ gnd vdd FILL
XFILL_2__14342_ gnd vdd FILL
XFILL_3__12913_ gnd vdd FILL
XFILL_4__10375_ gnd vdd FILL
XFILL_0__15521_ gnd vdd FILL
XFILL_2__11554_ gnd vdd FILL
XFILL_0__12733_ gnd vdd FILL
XFILL_1__10195_ gnd vdd FILL
XFILL_3__13893_ gnd vdd FILL
XFILL_0__7231_ gnd vdd FILL
XFILL_6__15812_ gnd vdd FILL
XFILL_5__14453_ gnd vdd FILL
XFILL_4__12114_ gnd vdd FILL
X_14928_ _14917_/Y _14928_/B gnd _14929_/A vdd NOR2X1
XFILL_2__10505_ gnd vdd FILL
XFILL_3__15632_ gnd vdd FILL
XFILL_4__13094_ gnd vdd FILL
XFILL_2__8147_ gnd vdd FILL
XFILL_5__11665_ gnd vdd FILL
XFILL_3__12844_ gnd vdd FILL
XFILL_2__14273_ gnd vdd FILL
XSFILL8520x11050 gnd vdd FILL
XFILL_0__15452_ gnd vdd FILL
XFILL_2__11485_ gnd vdd FILL
XFILL_5__13404_ gnd vdd FILL
XFILL_2__16012_ gnd vdd FILL
XFILL_5__10616_ gnd vdd FILL
XFILL_4__12045_ gnd vdd FILL
XFILL_6__12955_ gnd vdd FILL
XFILL_0__7162_ gnd vdd FILL
XFILL_2__13224_ gnd vdd FILL
X_14859_ _14859_/A _14859_/B gnd _14881_/A vdd NOR2X1
XSFILL18920x63050 gnd vdd FILL
XFILL_5__14384_ gnd vdd FILL
X_7790_ _7790_/Q _7790_/CLK _9561_/R vdd _7790_/D gnd vdd DFFSR
XFILL_2__8078_ gnd vdd FILL
XFILL_3__12775_ gnd vdd FILL
XFILL_6_BUFX2_insert40 gnd vdd FILL
XFILL_2__10436_ gnd vdd FILL
XFILL_3__15563_ gnd vdd FILL
XFILL_5__11596_ gnd vdd FILL
XFILL_0__14403_ gnd vdd FILL
XFILL_3__8960_ gnd vdd FILL
XFILL_1__13954_ gnd vdd FILL
XFILL_0__11615_ gnd vdd FILL
XFILL_0__15383_ gnd vdd FILL
XFILL_6__11906_ gnd vdd FILL
XFILL_5__16123_ gnd vdd FILL
XFILL_5__13335_ gnd vdd FILL
XFILL_6__15674_ gnd vdd FILL
XFILL_0__12595_ gnd vdd FILL
XSFILL59000x56050 gnd vdd FILL
XFILL_5__9876_ gnd vdd FILL
XFILL_0__7093_ gnd vdd FILL
XFILL_3__14514_ gnd vdd FILL
XFILL_5__10547_ gnd vdd FILL
XFILL_2__13155_ gnd vdd FILL
XFILL_3__11726_ gnd vdd FILL
XFILL_1__12905_ gnd vdd FILL
XFILL_2__10367_ gnd vdd FILL
XFILL_0__14334_ gnd vdd FILL
XFILL_3__15494_ gnd vdd FILL
XFILL_1__13885_ gnd vdd FILL
XFILL_3__8891_ gnd vdd FILL
XFILL_0__11546_ gnd vdd FILL
XFILL_5__8827_ gnd vdd FILL
XFILL_4__15804_ gnd vdd FILL
XFILL_5__16054_ gnd vdd FILL
XFILL_5__13266_ gnd vdd FILL
XFILL_2__12106_ gnd vdd FILL
X_9460_ _9424_/A _9578_/CLK _9460_/R vdd _9426_/Y gnd vdd DFFSR
XFILL_1__15624_ gnd vdd FILL
XFILL_3__11657_ gnd vdd FILL
XFILL_3__14445_ gnd vdd FILL
XFILL_1__12836_ gnd vdd FILL
XFILL_3__7842_ gnd vdd FILL
XFILL_2__13086_ gnd vdd FILL
XFILL_4__13996_ gnd vdd FILL
XFILL_5_BUFX2_insert108 gnd vdd FILL
XFILL_0__14265_ gnd vdd FILL
XSFILL109800x44050 gnd vdd FILL
XFILL_5__15005_ gnd vdd FILL
XFILL_2__10298_ gnd vdd FILL
XSFILL38840x14050 gnd vdd FILL
XFILL_0__11477_ gnd vdd FILL
XSFILL109000x25050 gnd vdd FILL
XFILL_5__8758_ gnd vdd FILL
XFILL_5__12217_ gnd vdd FILL
X_8411_ _8411_/Q _8151_/CLK _9048_/R vdd _8411_/D gnd vdd DFFSR
XFILL112360x21050 gnd vdd FILL
XSFILL64120x47050 gnd vdd FILL
XFILL_6__11768_ gnd vdd FILL
XFILL_4__15735_ gnd vdd FILL
XFILL_0__16004_ gnd vdd FILL
XFILL_2__12037_ gnd vdd FILL
XFILL_3__14376_ gnd vdd FILL
X_9391_ _9449_/Q gnd _9393_/A vdd INVX1
XFILL_0__13216_ gnd vdd FILL
XFILL_1__15555_ gnd vdd FILL
XFILL_3__11588_ gnd vdd FILL
XFILL_0__10428_ gnd vdd FILL
XFILL_1__12767_ gnd vdd FILL
XFILL_0_BUFX2_insert470 gnd vdd FILL
XFILL_5__7709_ gnd vdd FILL
XFILL_0__14196_ gnd vdd FILL
XSFILL24120x63050 gnd vdd FILL
XFILL_0__9803_ gnd vdd FILL
XFILL_6__7482_ gnd vdd FILL
XFILL_0_BUFX2_insert481 gnd vdd FILL
XFILL_6__14487_ gnd vdd FILL
XFILL_5__12148_ gnd vdd FILL
XFILL_3__16115_ gnd vdd FILL
X_8342_ _8342_/A _8372_/B _8341_/Y gnd _8342_/Y vdd OAI21X1
XFILL_3__13327_ gnd vdd FILL
XFILL_4__15666_ gnd vdd FILL
XFILL_0__7995_ gnd vdd FILL
XFILL_3__9512_ gnd vdd FILL
XFILL_3__10539_ gnd vdd FILL
XFILL_1__14506_ gnd vdd FILL
XFILL_0_BUFX2_insert492 gnd vdd FILL
XFILL_4__12878_ gnd vdd FILL
XFILL_1__11718_ gnd vdd FILL
XSFILL65000x75050 gnd vdd FILL
XFILL_0__10359_ gnd vdd FILL
XFILL_0__13147_ gnd vdd FILL
XFILL_4_BUFX2_insert808 gnd vdd FILL
XFILL_1__15486_ gnd vdd FILL
XFILL_1__12698_ gnd vdd FILL
XFILL_4_BUFX2_insert819 gnd vdd FILL
XFILL_4__14617_ gnd vdd FILL
XFILL_0__6946_ gnd vdd FILL
XFILL_0__9734_ gnd vdd FILL
XFILL_3__13258_ gnd vdd FILL
XFILL_3__16046_ gnd vdd FILL
XFILL_5__12079_ gnd vdd FILL
XSFILL3560x54050 gnd vdd FILL
XFILL_4__11829_ gnd vdd FILL
X_8273_ _8216_/A _8273_/B gnd _8273_/Y vdd NAND2X1
XFILL_4__15597_ gnd vdd FILL
XFILL_1__14437_ gnd vdd FILL
XFILL_2__13988_ gnd vdd FILL
XFILL_1__11649_ gnd vdd FILL
XSFILL84840x17050 gnd vdd FILL
XSFILL28760x66050 gnd vdd FILL
XFILL_5__15907_ gnd vdd FILL
X_7224_ _7276_/Q gnd _7226_/A vdd INVX1
XFILL_3__12209_ gnd vdd FILL
XFILL_0__9665_ gnd vdd FILL
XSFILL109560x1050 gnd vdd FILL
XFILL_0__6877_ gnd vdd FILL
XFILL_4__14548_ gnd vdd FILL
XFILL_2__15727_ gnd vdd FILL
XFILL_3__9374_ gnd vdd FILL
XFILL_0__12029_ gnd vdd FILL
XFILL_1__14368_ gnd vdd FILL
XFILL_0__8616_ gnd vdd FILL
X_7155_ _7155_/Q _8038_/CLK _7789_/R vdd _7155_/D gnd vdd DFFSR
XFILL_5__15838_ gnd vdd FILL
XFILL_1__16107_ gnd vdd FILL
XFILL_0__9596_ gnd vdd FILL
XFILL_3__8325_ gnd vdd FILL
XFILL_1__13319_ gnd vdd FILL
XFILL_4__14479_ gnd vdd FILL
XFILL_2__15658_ gnd vdd FILL
XCLKBUF1_insert160 CLKBUF1_insert192/A gnd _7282_/CLK vdd CLKBUF1
XFILL_1__14299_ gnd vdd FILL
XFILL_4__16218_ gnd vdd FILL
XFILL_1__7340_ gnd vdd FILL
X_7086_ _7084_/Y _7067_/A _7086_/C gnd _7144_/D vdd OAI21X1
XFILL_5__15769_ gnd vdd FILL
XCLKBUF1_insert171 CLKBUF1_insert182/A gnd _7530_/CLK vdd CLKBUF1
XFILL_3__8256_ gnd vdd FILL
XFILL_2__14609_ gnd vdd FILL
XFILL_1__16038_ gnd vdd FILL
XCLKBUF1_insert182 CLKBUF1_insert182/A gnd _7535_/CLK vdd CLKBUF1
XCLKBUF1_insert193 CLKBUF1_insert193/A gnd _8679_/CLK vdd CLKBUF1
XFILL_2__15589_ gnd vdd FILL
XFILL_3__7207_ gnd vdd FILL
XFILL_4__16149_ gnd vdd FILL
XFILL_0__8478_ gnd vdd FILL
XSFILL48920x79050 gnd vdd FILL
XSFILL89560x29050 gnd vdd FILL
XFILL_0__15719_ gnd vdd FILL
XFILL_3__8187_ gnd vdd FILL
XSFILL64200x27050 gnd vdd FILL
XFILL_1__9010_ gnd vdd FILL
XFILL_0__7429_ gnd vdd FILL
XFILL_5_BUFX2_insert8 gnd vdd FILL
XFILL_1_BUFX2_insert709 gnd vdd FILL
XFILL_3__7069_ gnd vdd FILL
X_7988_ _7988_/A _8006_/B _7988_/C gnd _8042_/D vdd OAI21X1
XFILL_4__7951_ gnd vdd FILL
XSFILL3640x34050 gnd vdd FILL
X_9727_ _9817_/Q gnd _9727_/Y vdd INVX1
XFILL_6__8867_ gnd vdd FILL
X_6939_ _6948_/A _9371_/B gnd _6939_/Y vdd NAND2X1
XFILL_4__6902_ gnd vdd FILL
XSFILL28840x46050 gnd vdd FILL
XSFILL53640x72050 gnd vdd FILL
XFILL_4__7882_ gnd vdd FILL
XFILL_6__7818_ gnd vdd FILL
XSFILL94280x22050 gnd vdd FILL
XFILL_1__9912_ gnd vdd FILL
X_9658_ _9658_/A _9625_/B _9658_/C gnd _9708_/D vdd OAI21X1
XFILL_4__9621_ gnd vdd FILL
X_10540_ _15806_/A gnd _10540_/Y vdd INVX1
X_8609_ _8609_/A _7713_/B gnd _8610_/C vdd NAND2X1
XFILL_5_BUFX2_insert620 gnd vdd FILL
X_9589_ _9555_/A _9589_/CLK _7911_/R vdd _9589_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert631 gnd vdd FILL
XFILL_5_BUFX2_insert642 gnd vdd FILL
XFILL_4__9552_ gnd vdd FILL
XSFILL33960x37050 gnd vdd FILL
XFILL_5_BUFX2_insert653 gnd vdd FILL
X_10471_ _10409_/A _7016_/CLK _9064_/R vdd _10471_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert664 gnd vdd FILL
XFILL_4__8503_ gnd vdd FILL
XFILL_1__6986_ gnd vdd FILL
XFILL_5_BUFX2_insert675 gnd vdd FILL
XFILL_1__9774_ gnd vdd FILL
XFILL_5_BUFX2_insert686 gnd vdd FILL
X_12210_ _12210_/A _12201_/B _12210_/C gnd _12210_/Y vdd OAI21X1
XFILL_4__9483_ gnd vdd FILL
XFILL_5_BUFX2_insert697 gnd vdd FILL
X_13190_ _13190_/Q _12669_/CLK _9050_/R vdd _13190_/D gnd vdd DFFSR
XFILL_1__8725_ gnd vdd FILL
X_12141_ _12139_/Y _12137_/A _12141_/C gnd _12141_/Y vdd OAI21X1
XFILL_1__8656_ gnd vdd FILL
XSFILL89240x11050 gnd vdd FILL
XFILL_4__8365_ gnd vdd FILL
XSFILL59080x2050 gnd vdd FILL
XFILL_2_CLKBUF1_insert201 gnd vdd FILL
XFILL_1__7607_ gnd vdd FILL
XFILL_2_CLKBUF1_insert212 gnd vdd FILL
X_12072_ _12072_/A _11881_/A _12072_/C gnd _12072_/Y vdd NAND3X1
XFILL_2_CLKBUF1_insert223 gnd vdd FILL
XFILL_1__8587_ gnd vdd FILL
XFILL_2__7380_ gnd vdd FILL
XFILL_4__7316_ gnd vdd FILL
X_15900_ _15204_/A _14492_/Y _14491_/Y _15980_/C gnd _15901_/B vdd OAI22X1
XSFILL110120x67050 gnd vdd FILL
X_11023_ _12238_/Y _11030_/A gnd _11026_/B vdd NOR2X1
XSFILL28920x26050 gnd vdd FILL
XFILL_4__7247_ gnd vdd FILL
X_15831_ _6959_/A gnd _15832_/C vdd INVX1
XFILL_2_BUFX2_insert510 gnd vdd FILL
XFILL_1__7469_ gnd vdd FILL
XFILL_2_BUFX2_insert521 gnd vdd FILL
XFILL_2_BUFX2_insert532 gnd vdd FILL
XFILL_4__7178_ gnd vdd FILL
XSFILL79160x63050 gnd vdd FILL
XFILL_2_BUFX2_insert543 gnd vdd FILL
XFILL_2__8001_ gnd vdd FILL
X_12974_ _12972_/Y vdd _12974_/C gnd _13054_/D vdd OAI21X1
XFILL_1__9208_ gnd vdd FILL
XFILL_4__10160_ gnd vdd FILL
X_15762_ _15762_/A _15761_/Y gnd _15762_/Y vdd NOR2X1
XFILL_2_BUFX2_insert554 gnd vdd FILL
XFILL_2_BUFX2_insert565 gnd vdd FILL
XFILL_3__10890_ gnd vdd FILL
XFILL_2_BUFX2_insert576 gnd vdd FILL
X_14713_ _14713_/A _14344_/B _13645_/C _9924_/A gnd _14714_/A vdd AOI22X1
XFILL_2_BUFX2_insert587 gnd vdd FILL
XFILL_5__7991_ gnd vdd FILL
X_11925_ _11925_/A _11921_/A _11925_/C gnd _6850_/A vdd OAI21X1
XFILL_5__11450_ gnd vdd FILL
XFILL_1__9139_ gnd vdd FILL
XFILL_2_BUFX2_insert598 gnd vdd FILL
X_15693_ _16002_/A _14237_/A _15321_/C _14237_/D gnd _15693_/Y vdd OAI22X1
XFILL_2__11270_ gnd vdd FILL
XFILL_5__9730_ gnd vdd FILL
XFILL_5__10401_ gnd vdd FILL
XFILL_5__6942_ gnd vdd FILL
X_14644_ _14644_/A _14644_/B gnd _14645_/B vdd NOR2X1
X_11856_ _11856_/A _11856_/B gnd _11856_/Y vdd OR2X2
XFILL_5__11381_ gnd vdd FILL
XFILL_0__11400_ gnd vdd FILL
XFILL_1__10951_ gnd vdd FILL
XFILL_0__12380_ gnd vdd FILL
XFILL_6_BUFX2_insert1073 gnd vdd FILL
XFILL_5__9661_ gnd vdd FILL
X_10807_ _10805_/Y _10831_/B _10806_/Y gnd _10859_/D vdd OAI21X1
XFILL_5__13120_ gnd vdd FILL
XFILL_5__6873_ gnd vdd FILL
X_14575_ _14573_/Y _14203_/B _14575_/C _14574_/Y gnd _14575_/Y vdd OAI22X1
XSFILL59080x30050 gnd vdd FILL
XFILL_3__11511_ gnd vdd FILL
XFILL_4__13850_ gnd vdd FILL
XFILL_2__8903_ gnd vdd FILL
X_11787_ _11787_/A _11786_/Y _11787_/C gnd _11790_/B vdd AOI21X1
XFILL_2__10152_ gnd vdd FILL
XFILL_3__12491_ gnd vdd FILL
XBUFX2_insert520 BUFX2_insert520/A gnd _7920_/R vdd BUFX2
XFILL_0__11331_ gnd vdd FILL
XFILL_1__13670_ gnd vdd FILL
XFILL_5__8612_ gnd vdd FILL
XFILL_2__9883_ gnd vdd FILL
XFILL_1__10882_ gnd vdd FILL
X_16314_ _16314_/A _16314_/B _16313_/Y _16314_/D gnd _16314_/Y vdd OAI22X1
XBUFX2_insert531 BUFX2_insert496/A gnd _8935_/R vdd BUFX2
XFILL_3__14230_ gnd vdd FILL
X_10738_ _10738_/Q _8537_/CLK _8166_/R vdd _10700_/Y gnd vdd DFFSR
XBUFX2_insert542 BUFX2_insert600/A gnd _12536_/R vdd BUFX2
XFILL_5__9592_ gnd vdd FILL
X_13526_ _13525_/Y _13526_/B gnd _13531_/C vdd NOR2X1
XBUFX2_insert553 BUFX2_insert559/A gnd _8942_/R vdd BUFX2
XFILL_5__10263_ gnd vdd FILL
XFILL_3__11442_ gnd vdd FILL
XFILL_1__12621_ gnd vdd FILL
XFILL_2__8834_ gnd vdd FILL
XFILL_4__13781_ gnd vdd FILL
XBUFX2_insert564 BUFX2_insert494/A gnd _8682_/R vdd BUFX2
XBUFX2_insert575 BUFX2_insert518/A gnd _9453_/R vdd BUFX2
XFILL_0__14050_ gnd vdd FILL
XFILL112280x36050 gnd vdd FILL
XFILL_2__14960_ gnd vdd FILL
XFILL_4__10993_ gnd vdd FILL
XFILL_0__11262_ gnd vdd FILL
XFILL_5__12002_ gnd vdd FILL
X_13457_ _9078_/A gnd _13457_/Y vdd INVX1
XFILL_4__15520_ gnd vdd FILL
XBUFX2_insert586 BUFX2_insert524/A gnd _7537_/R vdd BUFX2
XFILL_6__11553_ gnd vdd FILL
X_16245_ _14885_/A _15863_/A gnd _16245_/Y vdd NAND2X1
XFILL_4__12732_ gnd vdd FILL
XFILL_3__14161_ gnd vdd FILL
X_10669_ _10615_/B _9005_/B gnd _10670_/C vdd NAND2X1
XBUFX2_insert597 BUFX2_insert496/A gnd _9704_/R vdd BUFX2
XFILL_5__10194_ gnd vdd FILL
XFILL_1__15340_ gnd vdd FILL
XFILL_0__13001_ gnd vdd FILL
XFILL_2__13911_ gnd vdd FILL
XFILL_3__11373_ gnd vdd FILL
XFILL_2__8765_ gnd vdd FILL
XFILL_2__14891_ gnd vdd FILL
X_12408_ _12406_/Y _12407_/A _12408_/C gnd _12408_/Y vdd OAI21X1
XSFILL74200x4050 gnd vdd FILL
XFILL_0__11193_ gnd vdd FILL
XFILL_5__8474_ gnd vdd FILL
XFILL_3__13112_ gnd vdd FILL
XSFILL113800x4050 gnd vdd FILL
X_16176_ _15175_/B _10442_/A _14793_/C _15357_/B gnd _16178_/A vdd AOI22X1
X_13388_ _12808_/Q _12807_/Q gnd _13389_/B vdd NAND2X1
XFILL_4__15451_ gnd vdd FILL
XFILL_3__10324_ gnd vdd FILL
XFILL_2__13842_ gnd vdd FILL
XFILL_2__7716_ gnd vdd FILL
XSFILL79240x43050 gnd vdd FILL
XFILL_3__14092_ gnd vdd FILL
XFILL_1__11503_ gnd vdd FILL
XFILL_0__10144_ gnd vdd FILL
XFILL_2__8696_ gnd vdd FILL
XFILL_1__15271_ gnd vdd FILL
XFILL_5__7425_ gnd vdd FILL
XFILL_1__12483_ gnd vdd FILL
X_12339_ _12327_/A gnd _12319_/C gnd _12342_/A vdd NAND3X1
XFILL_4__14402_ gnd vdd FILL
X_15127_ _15127_/A _15127_/B _15812_/C gnd _15127_/Y vdd AOI21X1
XFILL_5__13953_ gnd vdd FILL
XFILL_4__11614_ gnd vdd FILL
XFILL_3__13043_ gnd vdd FILL
XFILL_1__14222_ gnd vdd FILL
XFILL_3__10255_ gnd vdd FILL
XFILL_4__15382_ gnd vdd FILL
XFILL_2__13773_ gnd vdd FILL
XFILL_4__12594_ gnd vdd FILL
XFILL_1__11434_ gnd vdd FILL
XFILL_0__14952_ gnd vdd FILL
XFILL_5__7356_ gnd vdd FILL
XSFILL114440x52050 gnd vdd FILL
X_15058_ _15057_/Y _15058_/B gnd _15076_/C vdd NAND2X1
XFILL_5__12904_ gnd vdd FILL
XFILL_4__14333_ gnd vdd FILL
XFILL_5__13884_ gnd vdd FILL
XFILL_2__12724_ gnd vdd FILL
XFILL_2__15512_ gnd vdd FILL
XFILL_4__11545_ gnd vdd FILL
XFILL_3__10186_ gnd vdd FILL
XFILL_1__14153_ gnd vdd FILL
XFILL_2__7578_ gnd vdd FILL
XFILL_0__13903_ gnd vdd FILL
X_14009_ _9313_/Q gnd _14010_/A vdd INVX1
XFILL_1__11365_ gnd vdd FILL
XFILL_0__8401_ gnd vdd FILL
XFILL_5__15623_ gnd vdd FILL
XFILL_5__7287_ gnd vdd FILL
XFILL_0__14883_ gnd vdd FILL
XFILL_0__9381_ gnd vdd FILL
XFILL_5__12835_ gnd vdd FILL
XFILL_3__8110_ gnd vdd FILL
XFILL_4__14264_ gnd vdd FILL
XFILL_1__13104_ gnd vdd FILL
XFILL_2__12655_ gnd vdd FILL
XFILL_3__9090_ gnd vdd FILL
XFILL_1__10316_ gnd vdd FILL
XFILL_4__11476_ gnd vdd FILL
XFILL_2__15443_ gnd vdd FILL
XFILL_0__13834_ gnd vdd FILL
XSFILL99400x56050 gnd vdd FILL
XFILL_3__14994_ gnd vdd FILL
XFILL_5__9026_ gnd vdd FILL
XSFILL59160x10050 gnd vdd FILL
XFILL_1__14084_ gnd vdd FILL
XFILL_0__8332_ gnd vdd FILL
XFILL_4__16003_ gnd vdd FILL
XFILL_1__11296_ gnd vdd FILL
XFILL_4__13215_ gnd vdd FILL
XFILL_5__15554_ gnd vdd FILL
X_8960_ _8961_/B _8832_/B gnd _8960_/Y vdd NAND2X1
XFILL_5__12766_ gnd vdd FILL
XFILL_4__10427_ gnd vdd FILL
XFILL_2__11606_ gnd vdd FILL
XSFILL59400x72050 gnd vdd FILL
XFILL_2__15374_ gnd vdd FILL
XFILL_4__14195_ gnd vdd FILL
XFILL_2__9248_ gnd vdd FILL
XFILL_1__13035_ gnd vdd FILL
XFILL_3__13945_ gnd vdd FILL
XFILL_2__12586_ gnd vdd FILL
XFILL_1__10247_ gnd vdd FILL
XFILL_0__13765_ gnd vdd FILL
XFILL_5__14505_ gnd vdd FILL
XFILL_0__10977_ gnd vdd FILL
X_7911_ _7911_/Q _7912_/CLK _7911_/R vdd _7851_/Y gnd vdd DFFSR
XFILL_5__11717_ gnd vdd FILL
XFILL_0__8263_ gnd vdd FILL
XFILL_4__10358_ gnd vdd FILL
XFILL_4__13146_ gnd vdd FILL
XFILL_2__14325_ gnd vdd FILL
XFILL_5__15485_ gnd vdd FILL
XFILL112360x16050 gnd vdd FILL
XFILL_5__12697_ gnd vdd FILL
X_8891_ _8891_/A gnd _8893_/A vdd INVX1
XFILL_0__15504_ gnd vdd FILL
XFILL_2__11537_ gnd vdd FILL
XFILL_0__12716_ gnd vdd FILL
XFILL_3__13876_ gnd vdd FILL
XSFILL23640x51050 gnd vdd FILL
XFILL_0__7214_ gnd vdd FILL
XFILL_1__10178_ gnd vdd FILL
XFILL_0__13696_ gnd vdd FILL
XFILL_5__14436_ gnd vdd FILL
XFILL_0__8194_ gnd vdd FILL
XFILL_3__15615_ gnd vdd FILL
X_7842_ _7842_/A _7821_/B _7842_/C gnd _7842_/Y vdd OAI21X1
XFILL_5__11648_ gnd vdd FILL
XFILL_2__14256_ gnd vdd FILL
XFILL_4__10289_ gnd vdd FILL
XFILL_3__12827_ gnd vdd FILL
XFILL_0__15435_ gnd vdd FILL
XFILL_2__11468_ gnd vdd FILL
XFILL_0__12647_ gnd vdd FILL
XFILL_3__9992_ gnd vdd FILL
XFILL_1__14986_ gnd vdd FILL
XFILL_5__9928_ gnd vdd FILL
XSFILL49080x62050 gnd vdd FILL
XSFILL79320x23050 gnd vdd FILL
XFILL112200x80050 gnd vdd FILL
XFILL_2__13207_ gnd vdd FILL
XFILL_4__12028_ gnd vdd FILL
XFILL_5__14367_ gnd vdd FILL
X_7773_ _7773_/Q _7261_/CLK _8669_/R vdd _7773_/D gnd vdd DFFSR
XSFILL3560x49050 gnd vdd FILL
XFILL_3__15546_ gnd vdd FILL
XFILL_2__10419_ gnd vdd FILL
XFILL_5__11579_ gnd vdd FILL
XFILL_3__12758_ gnd vdd FILL
XFILL_2__14187_ gnd vdd FILL
XFILL_1__13937_ gnd vdd FILL
XFILL_0__15366_ gnd vdd FILL
XFILL_5__16106_ gnd vdd FILL
XFILL_2__11399_ gnd vdd FILL
XFILL_5__13318_ gnd vdd FILL
XFILL_0__12578_ gnd vdd FILL
XFILL_5__9859_ gnd vdd FILL
X_9512_ _9512_/A _9533_/B _9512_/C gnd _9512_/Y vdd OAI21X1
XFILL_0__7076_ gnd vdd FILL
XFILL_2__13138_ gnd vdd FILL
XFILL_5__14298_ gnd vdd FILL
XFILL_3__11709_ gnd vdd FILL
XFILL_0__14317_ gnd vdd FILL
XSFILL114520x32050 gnd vdd FILL
XFILL_3__15477_ gnd vdd FILL
XFILL_1__13868_ gnd vdd FILL
XFILL_0__11529_ gnd vdd FILL
XFILL_3__8874_ gnd vdd FILL
XFILL_5__16037_ gnd vdd FILL
XFILL_0__15297_ gnd vdd FILL
XFILL_5__13249_ gnd vdd FILL
X_9443_ _9373_/A _7515_/CLK _7011_/R vdd _9375_/Y gnd vdd DFFSR
XFILL_6__8583_ gnd vdd FILL
XFILL_3__14428_ gnd vdd FILL
XFILL_4__13979_ gnd vdd FILL
XFILL_1__15607_ gnd vdd FILL
XFILL_3__7825_ gnd vdd FILL
XFILL_0__14248_ gnd vdd FILL
XFILL_1__13799_ gnd vdd FILL
XFILL_4__15718_ gnd vdd FILL
XFILL_1__6840_ gnd vdd FILL
XFILL_6__14539_ gnd vdd FILL
XSFILL69240x75050 gnd vdd FILL
X_9374_ _9339_/B _9374_/B gnd _9375_/C vdd NAND2X1
XFILL_1__15538_ gnd vdd FILL
XFILL_3__14359_ gnd vdd FILL
XFILL_3__7756_ gnd vdd FILL
XFILL_0__14179_ gnd vdd FILL
XFILL_4_BUFX2_insert605 gnd vdd FILL
X_8325_ _8411_/Q gnd _8325_/Y vdd INVX1
XFILL_4__15649_ gnd vdd FILL
XFILL_4_BUFX2_insert616 gnd vdd FILL
XFILL_0__7978_ gnd vdd FILL
XFILL_4_BUFX2_insert627 gnd vdd FILL
XFILL_4_BUFX2_insert638 gnd vdd FILL
XFILL_1__15469_ gnd vdd FILL
XFILL_3__7687_ gnd vdd FILL
XFILL_1__8510_ gnd vdd FILL
XFILL_4_BUFX2_insert649 gnd vdd FILL
X_8256_ _8254_/Y _8208_/B _8256_/C gnd _8302_/D vdd OAI21X1
XFILL_3__16029_ gnd vdd FILL
XFILL_0__6929_ gnd vdd FILL
XFILL_1__9490_ gnd vdd FILL
XSFILL8680x82050 gnd vdd FILL
XFILL_3__9426_ gnd vdd FILL
X_7207_ _7207_/A _7079_/B gnd _7208_/C vdd NAND2X1
XFILL_1__8441_ gnd vdd FILL
XFILL_0__9648_ gnd vdd FILL
XFILL_2_BUFX2_insert60 gnd vdd FILL
X_8187_ _8185_/Y _8187_/B _8187_/C gnd _8279_/D vdd OAI21X1
XFILL_3__9357_ gnd vdd FILL
XSFILL49160x42050 gnd vdd FILL
XFILL_2_BUFX2_insert71 gnd vdd FILL
XFILL_2_BUFX2_insert82 gnd vdd FILL
XSFILL3640x29050 gnd vdd FILL
XFILL_4__7101_ gnd vdd FILL
XFILL_2_BUFX2_insert93 gnd vdd FILL
X_7138_ _7138_/Q _7778_/CLK _8424_/R vdd _7138_/D gnd vdd DFFSR
XFILL_1__8372_ gnd vdd FILL
XFILL_4__8081_ gnd vdd FILL
XFILL_3__9288_ gnd vdd FILL
XFILL_1__7323_ gnd vdd FILL
XSFILL94280x17050 gnd vdd FILL
XFILL_4__7032_ gnd vdd FILL
X_7069_ _7139_/Q gnd _7069_/Y vdd INVX1
XFILL_3__8239_ gnd vdd FILL
XSFILL13640x83050 gnd vdd FILL
XSFILL28440x43050 gnd vdd FILL
XSFILL69320x55050 gnd vdd FILL
XFILL_1_BUFX2_insert506 gnd vdd FILL
XFILL_1__7185_ gnd vdd FILL
XFILL_1_BUFX2_insert517 gnd vdd FILL
XFILL_1_BUFX2_insert528 gnd vdd FILL
X_11710_ _11708_/Y _11710_/B gnd _11710_/Y vdd AND2X2
XFILL_1_BUFX2_insert539 gnd vdd FILL
XFILL_4__8983_ gnd vdd FILL
X_12690_ _12648_/A _12809_/CLK _12809_/R vdd _12690_/D gnd vdd DFFSR
XSFILL104520x64050 gnd vdd FILL
XFILL_4__7934_ gnd vdd FILL
X_11641_ _11663_/C _11687_/C _11641_/C gnd _11641_/Y vdd AOI21X1
XSFILL8760x62050 gnd vdd FILL
XSFILL23800x11050 gnd vdd FILL
XFILL_4__7865_ gnd vdd FILL
X_14360_ _9647_/A gnd _14360_/Y vdd INVX1
X_11572_ _11117_/Y _11570_/Y _11572_/C gnd _11579_/B vdd AOI21X1
XFILL_4__9604_ gnd vdd FILL
XFILL_2__6880_ gnd vdd FILL
X_13311_ _13311_/A gnd _13311_/Y vdd INVX1
X_10523_ _10505_/A _7579_/B gnd _10524_/C vdd NAND2X1
X_14291_ _10409_/A gnd _14293_/A vdd INVX1
XFILL_5_BUFX2_insert450 gnd vdd FILL
XFILL_5_BUFX2_insert461 gnd vdd FILL
XFILL_4__9535_ gnd vdd FILL
XFILL_5_BUFX2_insert472 gnd vdd FILL
X_13242_ _13295_/C _13242_/B _13241_/Y gnd _13245_/B vdd AOI21X1
X_16030_ _16030_/A _15378_/B _16029_/Y gnd _16032_/A vdd OAI21X1
X_10454_ _10358_/A _9436_/CLK _9454_/R vdd _10454_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert483 gnd vdd FILL
XFILL_5_BUFX2_insert494 gnd vdd FILL
XSFILL13720x63050 gnd vdd FILL
XSFILL94600x59050 gnd vdd FILL
XFILL_1__9757_ gnd vdd FILL
XFILL_1__6969_ gnd vdd FILL
XFILL_4__9466_ gnd vdd FILL
XFILL_2__7501_ gnd vdd FILL
XSFILL79160x58050 gnd vdd FILL
X_13173_ _13173_/A _13173_/B gnd _13174_/C vdd NAND2X1
XFILL_1__8708_ gnd vdd FILL
X_10385_ _15437_/A gnd _10387_/A vdd INVX1
XFILL_2__8481_ gnd vdd FILL
XFILL_5__7210_ gnd vdd FILL
XSFILL94200x61050 gnd vdd FILL
X_12124_ _11896_/A gnd _12126_/A vdd INVX1
XFILL_5__8190_ gnd vdd FILL
XFILL_4__9397_ gnd vdd FILL
XFILL_5__10950_ gnd vdd FILL
XFILL_2__7432_ gnd vdd FILL
XFILL_3__10040_ gnd vdd FILL
XFILL_1__8639_ gnd vdd FILL
XSFILL114360x67050 gnd vdd FILL
XFILL_2__10770_ gnd vdd FILL
XFILL_4__8348_ gnd vdd FILL
X_12055_ _12111_/A _12055_/B _12111_/C gnd _12055_/Y vdd NAND3X1
XFILL_4__11330_ gnd vdd FILL
XFILL_5__10881_ gnd vdd FILL
XFILL_2__7363_ gnd vdd FILL
XFILL_0__10900_ gnd vdd FILL
XFILL_1__11150_ gnd vdd FILL
XFILL_5__7072_ gnd vdd FILL
X_11006_ _11006_/A _11005_/Y _11006_/C gnd _11006_/Y vdd AOI21X1
XFILL_5__12620_ gnd vdd FILL
XFILL_0__11880_ gnd vdd FILL
XFILL_2__9102_ gnd vdd FILL
XFILL_4__11261_ gnd vdd FILL
XSFILL59080x25050 gnd vdd FILL
XFILL_2__12440_ gnd vdd FILL
XFILL_3__11991_ gnd vdd FILL
XFILL_2__7294_ gnd vdd FILL
XFILL_0__10831_ gnd vdd FILL
XSFILL99480x30050 gnd vdd FILL
XFILL_1__11081_ gnd vdd FILL
XFILL_4__13000_ gnd vdd FILL
X_15814_ _14359_/D gnd _15815_/B vdd INVX1
XFILL_2__9033_ gnd vdd FILL
XFILL_2_BUFX2_insert340 gnd vdd FILL
XFILL_3__13730_ gnd vdd FILL
XFILL_4__11192_ gnd vdd FILL
XFILL_3__10942_ gnd vdd FILL
XFILL_2__12371_ gnd vdd FILL
XFILL_1__10032_ gnd vdd FILL
XFILL_2_BUFX2_insert351 gnd vdd FILL
XFILL_2_BUFX2_insert362 gnd vdd FILL
XFILL_0__13550_ gnd vdd FILL
XFILL_0__10762_ gnd vdd FILL
XFILL_5__11502_ gnd vdd FILL
XFILL_2_BUFX2_insert373 gnd vdd FILL
XFILL_2__14110_ gnd vdd FILL
XFILL_4__10143_ gnd vdd FILL
XFILL_5__15270_ gnd vdd FILL
X_15745_ _15742_/Y _15744_/Y _15745_/C gnd _15745_/Y vdd NAND3X1
XFILL_5__12482_ gnd vdd FILL
XFILL_2_BUFX2_insert384 gnd vdd FILL
XFILL_2__11322_ gnd vdd FILL
X_12957_ _6872_/A gnd _12957_/Y vdd INVX1
XFILL_1__14840_ gnd vdd FILL
XFILL_3__13661_ gnd vdd FILL
XFILL_0__12501_ gnd vdd FILL
XFILL_2__15090_ gnd vdd FILL
XFILL_3__10873_ gnd vdd FILL
XFILL_2_BUFX2_insert395 gnd vdd FILL
XSFILL63960x71050 gnd vdd FILL
XFILL_5__14221_ gnd vdd FILL
XFILL_0__13481_ gnd vdd FILL
XFILL_5__7974_ gnd vdd FILL
XFILL_3__15400_ gnd vdd FILL
X_11908_ _13182_/Q gnd _11910_/A vdd INVX1
XFILL_0__10693_ gnd vdd FILL
XFILL_5__11433_ gnd vdd FILL
X_15676_ _10019_/A gnd _15676_/Y vdd INVX1
XFILL_3__12612_ gnd vdd FILL
XFILL_2__14041_ gnd vdd FILL
XFILL_4__14951_ gnd vdd FILL
X_12888_ _12888_/A vdd _12888_/C gnd _12940_/D vdd OAI21X1
XFILL_0__15220_ gnd vdd FILL
XSFILL79240x38050 gnd vdd FILL
XFILL_3__16380_ gnd vdd FILL
XFILL_2__11253_ gnd vdd FILL
XFILL_0__12432_ gnd vdd FILL
XFILL_3__13592_ gnd vdd FILL
XFILL_1__14771_ gnd vdd FILL
XFILL_5__6925_ gnd vdd FILL
XFILL_1__11983_ gnd vdd FILL
XFILL_6__15511_ gnd vdd FILL
X_14627_ _9710_/Q gnd _14628_/A vdd INVX1
XFILL_5__14152_ gnd vdd FILL
XFILL_4__13902_ gnd vdd FILL
XFILL_3__15331_ gnd vdd FILL
XFILL_5__11364_ gnd vdd FILL
X_11839_ _11839_/A _11838_/Y gnd _11839_/Y vdd NAND2X1
XSFILL64040x80050 gnd vdd FILL
XFILL_2__9935_ gnd vdd FILL
XFILL_1__13722_ gnd vdd FILL
XFILL_4__14882_ gnd vdd FILL
XFILL_1__10934_ gnd vdd FILL
XFILL_2__11184_ gnd vdd FILL
XFILL_0__15151_ gnd vdd FILL
XFILL_0__12363_ gnd vdd FILL
XFILL_5__13103_ gnd vdd FILL
XFILL_5__9644_ gnd vdd FILL
XFILL_5__10315_ gnd vdd FILL
XFILL_5__6856_ gnd vdd FILL
XFILL_0__8950_ gnd vdd FILL
X_14558_ _8891_/A _14482_/B _13854_/B _9325_/Q gnd _14558_/Y vdd AOI22X1
XFILL_4__13833_ gnd vdd FILL
XFILL_5__14083_ gnd vdd FILL
XFILL_3__12474_ gnd vdd FILL
XFILL_2__10135_ gnd vdd FILL
XFILL_0__14102_ gnd vdd FILL
XFILL_5__11295_ gnd vdd FILL
XFILL_3__15262_ gnd vdd FILL
XFILL_1__13653_ gnd vdd FILL
XFILL_2__9866_ gnd vdd FILL
XBUFX2_insert350 _10927_/Y gnd _12239_/A vdd BUFX2
XFILL_0__11314_ gnd vdd FILL
XFILL_2__15992_ gnd vdd FILL
XSFILL84360x29050 gnd vdd FILL
XBUFX2_insert361 _11352_/Y gnd _11553_/C vdd BUFX2
XFILL_0__15082_ gnd vdd FILL
XBUFX2_insert372 _13338_/Y gnd _9551_/B vdd BUFX2
XFILL_0__12294_ gnd vdd FILL
XFILL_5__13034_ gnd vdd FILL
X_13509_ _9175_/Q gnd _13509_/Y vdd INVX1
XFILL_3__14213_ gnd vdd FILL
XFILL_5__10246_ gnd vdd FILL
XFILL_3__11425_ gnd vdd FILL
XBUFX2_insert383 _13331_/Y gnd _9086_/B vdd BUFX2
XFILL_0__8881_ gnd vdd FILL
XFILL_3__7610_ gnd vdd FILL
XFILL_1__12604_ gnd vdd FILL
X_14489_ _14488_/Y _14567_/D _14489_/C _15895_/A gnd _14489_/Y vdd OAI22X1
XFILL_4__13764_ gnd vdd FILL
XBUFX2_insert394 _13293_/Y gnd _7624_/A vdd BUFX2
XFILL_3__8590_ gnd vdd FILL
XFILL_4__10976_ gnd vdd FILL
XFILL_3__15193_ gnd vdd FILL
XSFILL98920x44050 gnd vdd FILL
XFILL_0__14033_ gnd vdd FILL
XFILL_2__14943_ gnd vdd FILL
XFILL_1__16372_ gnd vdd FILL
XFILL_2__10066_ gnd vdd FILL
XFILL_5__8526_ gnd vdd FILL
XFILL_2__9797_ gnd vdd FILL
XFILL_6__14324_ gnd vdd FILL
XFILL_1__13584_ gnd vdd FILL
XFILL_0__11245_ gnd vdd FILL
X_16228_ _14842_/Y _16228_/B _15726_/A _16227_/Y gnd _16230_/A vdd OAI22X1
XFILL_0__7832_ gnd vdd FILL
XFILL_4__15503_ gnd vdd FILL
XFILL_1__10796_ gnd vdd FILL
XSFILL84360x5050 gnd vdd FILL
XFILL_4__12715_ gnd vdd FILL
XFILL_3__14144_ gnd vdd FILL
XFILL_1__15323_ gnd vdd FILL
XFILL_3__11356_ gnd vdd FILL
XFILL_5__10177_ gnd vdd FILL
XFILL_2__8748_ gnd vdd FILL
XFILL_4__13695_ gnd vdd FILL
XFILL_2__14874_ gnd vdd FILL
XFILL_0__11176_ gnd vdd FILL
XFILL_5__8457_ gnd vdd FILL
X_8110_ _8108_/Y _8100_/A _8110_/C gnd _8168_/D vdd OAI21X1
XFILL_0__7763_ gnd vdd FILL
XFILL_3__10307_ gnd vdd FILL
XFILL_4__15434_ gnd vdd FILL
X_16159_ _14763_/B gnd _16160_/B vdd INVX1
X_9090_ _9090_/A gnd _9090_/Y vdd INVX1
XFILL_4__12646_ gnd vdd FILL
XFILL_5__14985_ gnd vdd FILL
XFILL_3__14075_ gnd vdd FILL
XFILL_0__10127_ gnd vdd FILL
XFILL_2__13825_ gnd vdd FILL
XFILL_1__15254_ gnd vdd FILL
XFILL_3__7472_ gnd vdd FILL
XFILL_3__11287_ gnd vdd FILL
XFILL_1__12466_ gnd vdd FILL
XFILL_0__15984_ gnd vdd FILL
XSFILL23640x46050 gnd vdd FILL
XFILL_0__9502_ gnd vdd FILL
XFILL_6__14186_ gnd vdd FILL
XFILL_5__8388_ gnd vdd FILL
X_8041_ _8041_/Q _9328_/CLK _7408_/R vdd _8041_/D gnd vdd DFFSR
XFILL_3__13026_ gnd vdd FILL
XFILL_5__13936_ gnd vdd FILL
XFILL_0__7694_ gnd vdd FILL
XFILL_4__15365_ gnd vdd FILL
XFILL_1__14205_ gnd vdd FILL
XFILL_3__10238_ gnd vdd FILL
XFILL_3__9211_ gnd vdd FILL
XFILL_4__12577_ gnd vdd FILL
XFILL_1__11417_ gnd vdd FILL
XFILL_2__10968_ gnd vdd FILL
XFILL_1__15185_ gnd vdd FILL
XFILL_0__10058_ gnd vdd FILL
XFILL_2__13756_ gnd vdd FILL
XFILL_0__14935_ gnd vdd FILL
XFILL_1__12397_ gnd vdd FILL
XFILL_5__7339_ gnd vdd FILL
XFILL_4__14316_ gnd vdd FILL
XFILL_5__13867_ gnd vdd FILL
XSFILL49080x57050 gnd vdd FILL
XFILL_4__11528_ gnd vdd FILL
XFILL_3__9142_ gnd vdd FILL
XFILL112200x75050 gnd vdd FILL
XFILL_2__12707_ gnd vdd FILL
XFILL_1__14136_ gnd vdd FILL
XFILL_3__10169_ gnd vdd FILL
XFILL_4__15296_ gnd vdd FILL
XFILL_2__13687_ gnd vdd FILL
XFILL_1__11348_ gnd vdd FILL
XFILL_0__14866_ gnd vdd FILL
XFILL_2__10899_ gnd vdd FILL
XFILL_0__9364_ gnd vdd FILL
XFILL_5__15606_ gnd vdd FILL
XFILL_4__14247_ gnd vdd FILL
XFILL_2__12638_ gnd vdd FILL
XFILL_5__13798_ gnd vdd FILL
X_9992_ _9992_/A gnd _9994_/A vdd INVX1
XFILL_4__11459_ gnd vdd FILL
XFILL_2__15426_ gnd vdd FILL
XFILL_0__13817_ gnd vdd FILL
XFILL_1__14067_ gnd vdd FILL
XFILL_5__9009_ gnd vdd FILL
XFILL_3__14977_ gnd vdd FILL
XSFILL114520x27050 gnd vdd FILL
XFILL_6__12019_ gnd vdd FILL
XFILL_1__11279_ gnd vdd FILL
XFILL_0__8315_ gnd vdd FILL
XFILL_0__14797_ gnd vdd FILL
XFILL_5__15537_ gnd vdd FILL
XFILL_5__12749_ gnd vdd FILL
XFILL_0__9295_ gnd vdd FILL
X_8943_ _8943_/Q _9823_/CLK _9056_/R vdd _8943_/D gnd vdd DFFSR
XFILL_4__14178_ gnd vdd FILL
XFILL_1__13018_ gnd vdd FILL
XFILL_3__13928_ gnd vdd FILL
XFILL_2__12569_ gnd vdd FILL
XFILL_2__15357_ gnd vdd FILL
XFILL_0__13748_ gnd vdd FILL
XFILL_0__8246_ gnd vdd FILL
XFILL_4__13129_ gnd vdd FILL
XFILL_5__15468_ gnd vdd FILL
XFILL_2__14308_ gnd vdd FILL
X_8874_ _8859_/A _8874_/B gnd _8874_/Y vdd NAND2X1
XFILL_3__13859_ gnd vdd FILL
XFILL_2__15288_ gnd vdd FILL
XFILL_0__13679_ gnd vdd FILL
XFILL_5__14419_ gnd vdd FILL
XFILL_6__6965_ gnd vdd FILL
X_7825_ _7903_/Q gnd _7827_/A vdd INVX1
XFILL_5__15399_ gnd vdd FILL
XFILL_2__14239_ gnd vdd FILL
XFILL_0__15418_ gnd vdd FILL
XFILL_3__9975_ gnd vdd FILL
XFILL_1__14969_ gnd vdd FILL
XFILL_0__16398_ gnd vdd FILL
XFILL_6__9684_ gnd vdd FILL
X_7756_ _7754_/Y _7690_/B _7756_/C gnd _7756_/Y vdd OAI21X1
XFILL_3__15529_ gnd vdd FILL
XSFILL8680x77050 gnd vdd FILL
XFILL_1__8990_ gnd vdd FILL
XFILL_0__15349_ gnd vdd FILL
XFILL_6__8635_ gnd vdd FILL
XFILL_0__7059_ gnd vdd FILL
XSFILL33880x70050 gnd vdd FILL
XFILL_1__7941_ gnd vdd FILL
X_7687_ _7685_/Y _7723_/B _7687_/C gnd _7771_/D vdd OAI21X1
XFILL_3__8857_ gnd vdd FILL
X_9426_ _9424_/Y _9425_/A _9426_/C gnd _9426_/Y vdd OAI21X1
XFILL_1__7872_ gnd vdd FILL
XSFILL90040x30050 gnd vdd FILL
XFILL_3__7808_ gnd vdd FILL
XSFILL64200x40050 gnd vdd FILL
XFILL_4__7581_ gnd vdd FILL
XFILL_3__8788_ gnd vdd FILL
XFILL_1__9611_ gnd vdd FILL
XFILL_4_BUFX2_insert402 gnd vdd FILL
X_9357_ _9355_/Y _9356_/A _9357_/C gnd _9357_/Y vdd OAI21X1
XFILL_4_BUFX2_insert413 gnd vdd FILL
XFILL_3__7739_ gnd vdd FILL
XFILL_4_BUFX2_insert424 gnd vdd FILL
XSFILL54280x28050 gnd vdd FILL
X_8308_ _8272_/A _8297_/CLK _7796_/R vdd _8274_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert435 gnd vdd FILL
XFILL_4_BUFX2_insert446 gnd vdd FILL
XFILL_1__9542_ gnd vdd FILL
XFILL_4_BUFX2_insert457 gnd vdd FILL
X_9288_ _9301_/B _7496_/B gnd _9289_/C vdd NAND2X1
XFILL_4_BUFX2_insert468 gnd vdd FILL
XFILL_4__9251_ gnd vdd FILL
X_10170_ _10170_/A _10169_/A _10169_/Y gnd _10170_/Y vdd OAI21X1
XFILL_4_BUFX2_insert479 gnd vdd FILL
XFILL_1__9473_ gnd vdd FILL
X_8239_ _8297_/Q gnd _8241_/A vdd INVX1
XFILL_4__8202_ gnd vdd FILL
XFILL_3__9409_ gnd vdd FILL
XSFILL104520x59050 gnd vdd FILL
XFILL_4__8133_ gnd vdd FILL
XFILL_1__8355_ gnd vdd FILL
XFILL_4__8064_ gnd vdd FILL
XFILL_1__7306_ gnd vdd FILL
XFILL_3_CLKBUF1_insert115 gnd vdd FILL
X_13860_ _13859_/Y _13860_/B _14203_/C _13860_/D gnd _13860_/Y vdd OAI22X1
XFILL_3_CLKBUF1_insert126 gnd vdd FILL
XFILL_5_CLKBUF1_insert1075 gnd vdd FILL
XSFILL74040x43050 gnd vdd FILL
XFILL_3_CLKBUF1_insert137 gnd vdd FILL
XFILL_3_CLKBUF1_insert148 gnd vdd FILL
X_12811_ _12811_/Q _8171_/CLK _8171_/R vdd _12757_/Y gnd vdd DFFSR
XFILL_3_CLKBUF1_insert159 gnd vdd FILL
XFILL_1__7237_ gnd vdd FILL
X_13791_ _16342_/A _14344_/B gnd _13791_/Y vdd NAND2X1
XFILL_1_BUFX2_insert303 gnd vdd FILL
XFILL_1_BUFX2_insert314 gnd vdd FILL
X_15530_ _15646_/D _14002_/Y _15530_/C _15070_/C gnd _15533_/A vdd OAI22X1
X_12742_ _12740_/Y _12718_/B _12742_/C gnd _12742_/Y vdd OAI21X1
XFILL_1_BUFX2_insert325 gnd vdd FILL
XFILL_1__7168_ gnd vdd FILL
XFILL_1_BUFX2_insert336 gnd vdd FILL
XFILL_1_BUFX2_insert347 gnd vdd FILL
XSFILL13720x58050 gnd vdd FILL
XFILL_1_BUFX2_insert358 gnd vdd FILL
XFILL_4__8966_ gnd vdd FILL
X_12673_ _12673_/Q _9060_/CLK _9060_/R vdd _12673_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert369 gnd vdd FILL
X_15461_ _15461_/A _15848_/A gnd _15461_/Y vdd NOR2X1
XFILL_1__7099_ gnd vdd FILL
XFILL_2__7981_ gnd vdd FILL
X_11624_ _11617_/A _12282_/Y _11624_/C gnd _11625_/B vdd OAI21X1
X_14412_ _14403_/Y _14404_/Y _14412_/C gnd _14412_/Y vdd NAND3X1
XFILL_5__7690_ gnd vdd FILL
XFILL_4__8897_ gnd vdd FILL
X_15392_ _15391_/Y _15392_/B _15392_/C _13877_/Y gnd _15395_/A vdd OAI22X1
XFILL_2__9720_ gnd vdd FILL
XFILL_2__6932_ gnd vdd FILL
XSFILL28920x8050 gnd vdd FILL
XFILL_4__7848_ gnd vdd FILL
X_14343_ _8808_/Q _13853_/B _14343_/C gnd _14345_/A vdd AOI21X1
X_11555_ _11111_/Y _11423_/B gnd _11555_/Y vdd NOR2X1
XFILL_4__10830_ gnd vdd FILL
XFILL_5__11080_ gnd vdd FILL
XFILL_2__9651_ gnd vdd FILL
XFILL_2__6863_ gnd vdd FILL
XFILL_1__10650_ gnd vdd FILL
XFILL_5__9360_ gnd vdd FILL
X_10506_ _10504_/Y _10505_/A _10506_/C gnd _10506_/Y vdd OAI21X1
XSFILL8840x37050 gnd vdd FILL
XFILL_5__10031_ gnd vdd FILL
XFILL_3__11210_ gnd vdd FILL
X_14274_ _7271_/Q _13434_/B _14323_/B _8233_/A gnd _14275_/B vdd AOI22X1
XFILL_5_BUFX2_insert280 gnd vdd FILL
XFILL_2__8602_ gnd vdd FILL
X_11486_ _11174_/C _11327_/Y _11486_/C gnd _11487_/C vdd NAND3X1
XFILL_1__9809_ gnd vdd FILL
XFILL_4__10761_ gnd vdd FILL
XFILL_2__11940_ gnd vdd FILL
XFILL_5_BUFX2_insert291 gnd vdd FILL
XFILL_0__11030_ gnd vdd FILL
XFILL_3__12190_ gnd vdd FILL
XFILL_5__8311_ gnd vdd FILL
XFILL_4__9518_ gnd vdd FILL
X_13225_ _13209_/Y _13359_/A _13244_/A _13225_/D gnd _13225_/Y vdd OAI22X1
X_16013_ _7790_/Q _15969_/C gnd _16013_/Y vdd NAND2X1
XFILL_1__10581_ gnd vdd FILL
XFILL_4__12500_ gnd vdd FILL
XFILL_5__9291_ gnd vdd FILL
X_10437_ _10372_/B _9413_/B gnd _10437_/Y vdd NAND2X1
XSFILL99480x25050 gnd vdd FILL
XFILL_3__11141_ gnd vdd FILL
XSFILL74120x23050 gnd vdd FILL
XFILL_2__8533_ gnd vdd FILL
XFILL_1__12320_ gnd vdd FILL
XFILL_4__13480_ gnd vdd FILL
XFILL_4__10692_ gnd vdd FILL
XFILL_2__11871_ gnd vdd FILL
XFILL_5__8242_ gnd vdd FILL
X_13156_ _13154_/Y _13155_/A _13156_/C gnd _13200_/D vdd OAI21X1
X_10368_ _10443_/A _7424_/B gnd _10369_/C vdd NAND2X1
XFILL_4__12431_ gnd vdd FILL
XFILL_5__14770_ gnd vdd FILL
XFILL_2__13610_ gnd vdd FILL
XFILL_5__11982_ gnd vdd FILL
XFILL_4_BUFX2_insert980 gnd vdd FILL
XFILL_2__10822_ gnd vdd FILL
XFILL_3__11072_ gnd vdd FILL
XFILL_4_BUFX2_insert991 gnd vdd FILL
XFILL_2__8464_ gnd vdd FILL
XFILL_2__14590_ gnd vdd FILL
XFILL_1__12251_ gnd vdd FILL
X_12107_ _12111_/A _12107_/B _12111_/C gnd _12110_/A vdd NAND3X1
XFILL_0__12981_ gnd vdd FILL
XFILL_5__13721_ gnd vdd FILL
XFILL_5__10933_ gnd vdd FILL
XFILL_3__10023_ gnd vdd FILL
X_13087_ _13087_/A _13134_/A _13087_/C gnd _13087_/Y vdd OAI21X1
XSFILL13800x38050 gnd vdd FILL
XFILL_3__14900_ gnd vdd FILL
XFILL_4__15150_ gnd vdd FILL
X_10299_ _10349_/Q gnd _10299_/Y vdd INVX1
XFILL_4__12362_ gnd vdd FILL
XFILL_2__7415_ gnd vdd FILL
XFILL_2__13541_ gnd vdd FILL
XFILL_1__11202_ gnd vdd FILL
XFILL_2__10753_ gnd vdd FILL
XFILL_2__8395_ gnd vdd FILL
XFILL_0__14720_ gnd vdd FILL
XSFILL109480x10050 gnd vdd FILL
XFILL_3__15880_ gnd vdd FILL
XFILL_0__11932_ gnd vdd FILL
XFILL_5__7124_ gnd vdd FILL
XFILL_1__12182_ gnd vdd FILL
XSFILL23960x82050 gnd vdd FILL
X_12038_ _12038_/A _12036_/Y _12037_/Y gnd _13116_/B vdd NAND3X1
XFILL_4__14101_ gnd vdd FILL
XFILL_5__13652_ gnd vdd FILL
XFILL_4__11313_ gnd vdd FILL
XFILL_3__14831_ gnd vdd FILL
XFILL_4__15081_ gnd vdd FILL
XFILL_2__7346_ gnd vdd FILL
XFILL_2__13472_ gnd vdd FILL
XFILL_4__12293_ gnd vdd FILL
XFILL_1__11133_ gnd vdd FILL
XFILL_2__16260_ gnd vdd FILL
XFILL_2__10684_ gnd vdd FILL
XFILL_5__7055_ gnd vdd FILL
XFILL_0__14651_ gnd vdd FILL
XFILL_5__12603_ gnd vdd FILL
XFILL_0__11863_ gnd vdd FILL
XFILL_5__16371_ gnd vdd FILL
XFILL_4__14032_ gnd vdd FILL
XFILL_2__15211_ gnd vdd FILL
XFILL_2__12423_ gnd vdd FILL
XFILL_5__13583_ gnd vdd FILL
XFILL_4__11244_ gnd vdd FILL
XFILL_0__13602_ gnd vdd FILL
XFILL_2__16191_ gnd vdd FILL
XFILL_5__10795_ gnd vdd FILL
XFILL_3__14762_ gnd vdd FILL
XFILL_0__8100_ gnd vdd FILL
XFILL_0__10814_ gnd vdd FILL
XFILL_3__11974_ gnd vdd FILL
XFILL_1__15941_ gnd vdd FILL
XFILL_1__11064_ gnd vdd FILL
XFILL_0__14582_ gnd vdd FILL
XFILL_5__15322_ gnd vdd FILL
XFILL_0__9080_ gnd vdd FILL
XFILL_5__12534_ gnd vdd FILL
XFILL_0__11794_ gnd vdd FILL
XFILL_2__9016_ gnd vdd FILL
XFILL_3__13713_ gnd vdd FILL
XFILL_2__15142_ gnd vdd FILL
XFILL_4__11175_ gnd vdd FILL
XFILL_2__12354_ gnd vdd FILL
XFILL_3__10925_ gnd vdd FILL
XFILL_0__16321_ gnd vdd FILL
X_13989_ _7191_/A _14458_/C _14481_/C _6935_/A gnd _13997_/B vdd AOI22X1
XFILL_1__10015_ gnd vdd FILL
XFILL_3__14693_ gnd vdd FILL
XFILL_0__13533_ gnd vdd FILL
XFILL_1__15872_ gnd vdd FILL
XFILL_0__10745_ gnd vdd FILL
X_15728_ _15180_/C _15728_/B _15170_/D _14229_/Y gnd _15729_/A vdd OAI22X1
XFILL_5__15253_ gnd vdd FILL
XFILL_4__10126_ gnd vdd FILL
XFILL_5__12465_ gnd vdd FILL
XFILL_2__11305_ gnd vdd FILL
XFILL_4__15983_ gnd vdd FILL
XFILL_3__13644_ gnd vdd FILL
XFILL_2__15073_ gnd vdd FILL
XFILL_1__14823_ gnd vdd FILL
XFILL_0__16252_ gnd vdd FILL
XFILL_2__12285_ gnd vdd FILL
XFILL_5__14204_ gnd vdd FILL
XFILL_0__13464_ gnd vdd FILL
XSFILL68280x80050 gnd vdd FILL
X_7610_ _7610_/A _7592_/B _7609_/Y gnd _7660_/D vdd OAI21X1
XFILL_5__7957_ gnd vdd FILL
XFILL_0__10676_ gnd vdd FILL
XFILL_5__11416_ gnd vdd FILL
XFILL_5__15184_ gnd vdd FILL
X_15659_ _9317_/Q _15892_/B _15380_/C _9957_/Q gnd _15659_/Y vdd AOI22X1
XFILL_2__14024_ gnd vdd FILL
XFILL_4__14934_ gnd vdd FILL
XFILL_4__10057_ gnd vdd FILL
X_8590_ _8670_/Q gnd _8590_/Y vdd INVX1
XFILL_0__15203_ gnd vdd FILL
XFILL_3__16363_ gnd vdd FILL
XFILL_5__12396_ gnd vdd FILL
XFILL_1_BUFX2_insert870 gnd vdd FILL
XFILL_2__11236_ gnd vdd FILL
XFILL_3__10787_ gnd vdd FILL
XFILL_0__12415_ gnd vdd FILL
XFILL_3__9760_ gnd vdd FILL
XFILL_1_BUFX2_insert881 gnd vdd FILL
XFILL_3__13575_ gnd vdd FILL
XFILL_1__14754_ gnd vdd FILL
XFILL_3__6972_ gnd vdd FILL
XFILL_1_BUFX2_insert892 gnd vdd FILL
XFILL_0__16183_ gnd vdd FILL
XFILL_1__11966_ gnd vdd FILL
XFILL_5__6908_ gnd vdd FILL
XSFILL59000x64050 gnd vdd FILL
XFILL_5__14135_ gnd vdd FILL
XFILL_0__13395_ gnd vdd FILL
XFILL_3__15314_ gnd vdd FILL
X_7541_ _7541_/Q _7010_/CLK _8278_/R vdd _7509_/Y gnd vdd DFFSR
XFILL_5__7888_ gnd vdd FILL
XFILL_5__11347_ gnd vdd FILL
XFILL_4__14865_ gnd vdd FILL
XFILL_2__9918_ gnd vdd FILL
XFILL_3__12526_ gnd vdd FILL
XFILL_3__8711_ gnd vdd FILL
XFILL_0__9982_ gnd vdd FILL
XFILL_1__13705_ gnd vdd FILL
XFILL_1__10917_ gnd vdd FILL
XFILL_0__15134_ gnd vdd FILL
XFILL_2__11167_ gnd vdd FILL
XFILL_3__16294_ gnd vdd FILL
XFILL_5__9627_ gnd vdd FILL
XFILL_0__12346_ gnd vdd FILL
XFILL_1__14685_ gnd vdd FILL
XFILL_1__11897_ gnd vdd FILL
XFILL_5__6839_ gnd vdd FILL
XFILL_4__13816_ gnd vdd FILL
XFILL_5__14066_ gnd vdd FILL
XFILL_3__15245_ gnd vdd FILL
X_7472_ _7472_/A _8496_/B gnd _7473_/C vdd NAND2X1
XFILL_2__10118_ gnd vdd FILL
XFILL_5__11278_ gnd vdd FILL
XFILL_1__13636_ gnd vdd FILL
XFILL_3__12457_ gnd vdd FILL
XFILL_4__14796_ gnd vdd FILL
XFILL_2__9849_ gnd vdd FILL
XFILL_3__8642_ gnd vdd FILL
XFILL_2__15975_ gnd vdd FILL
XFILL_0__15065_ gnd vdd FILL
XFILL_2__11098_ gnd vdd FILL
XSFILL38840x22050 gnd vdd FILL
XFILL_5__13017_ gnd vdd FILL
XFILL_0__12277_ gnd vdd FILL
XSFILL109000x33050 gnd vdd FILL
XFILL_6__8351_ gnd vdd FILL
X_9211_ _9211_/A _9238_/B _9210_/Y gnd _9211_/Y vdd OAI21X1
XFILL_6__12568_ gnd vdd FILL
XFILL_4__13747_ gnd vdd FILL
XFILL_0__8864_ gnd vdd FILL
XSFILL64120x55050 gnd vdd FILL
XFILL_3__11408_ gnd vdd FILL
XFILL_4__10959_ gnd vdd FILL
XFILL_3__15176_ gnd vdd FILL
XFILL_3__12388_ gnd vdd FILL
XFILL_1__16355_ gnd vdd FILL
XFILL_0__14016_ gnd vdd FILL
XFILL_2__10049_ gnd vdd FILL
XFILL_2__14926_ gnd vdd FILL
XFILL_5__8509_ gnd vdd FILL
XFILL_3__8573_ gnd vdd FILL
XFILL_1__13567_ gnd vdd FILL
XFILL_0__11228_ gnd vdd FILL
XFILL_6__7302_ gnd vdd FILL
XFILL_1__10779_ gnd vdd FILL
X_9142_ _9101_/B _9782_/B gnd _9143_/C vdd NAND2X1
XFILL_0__7815_ gnd vdd FILL
XFILL_5__9489_ gnd vdd FILL
XFILL_3__14127_ gnd vdd FILL
XFILL_1__15306_ gnd vdd FILL
XFILL_4__13678_ gnd vdd FILL
XFILL_1__12518_ gnd vdd FILL
XFILL_3__11339_ gnd vdd FILL
XFILL_2__14857_ gnd vdd FILL
XFILL_1__16286_ gnd vdd FILL
XSFILL43960x13050 gnd vdd FILL
XFILL_1__13498_ gnd vdd FILL
XFILL_0__11159_ gnd vdd FILL
XFILL_4__15417_ gnd vdd FILL
XFILL_4__12629_ gnd vdd FILL
XFILL_0__7746_ gnd vdd FILL
X_9073_ _9031_/A _8433_/CLK _7921_/R vdd _9073_/D gnd vdd DFFSR
XFILL_2__13808_ gnd vdd FILL
XFILL_3_BUFX2_insert409 gnd vdd FILL
XFILL_1__15237_ gnd vdd FILL
XFILL_3__14058_ gnd vdd FILL
XFILL_5__14968_ gnd vdd FILL
XFILL_4__16397_ gnd vdd FILL
XFILL_1__12449_ gnd vdd FILL
XFILL_3__7455_ gnd vdd FILL
XFILL_0__15967_ gnd vdd FILL
XFILL_2__14788_ gnd vdd FILL
X_8024_ _8024_/Q _8152_/CLK _9944_/R vdd _8024_/D gnd vdd DFFSR
XSFILL28760x74050 gnd vdd FILL
XFILL_4__15348_ gnd vdd FILL
XFILL_3__13009_ gnd vdd FILL
XFILL_0__7677_ gnd vdd FILL
XFILL_5__13919_ gnd vdd FILL
XFILL_5__14899_ gnd vdd FILL
XSFILL44040x22050 gnd vdd FILL
XFILL_1__15168_ gnd vdd FILL
XFILL_2__13739_ gnd vdd FILL
XFILL_0__14918_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1081 gnd vdd FILL
XFILL_0__15898_ gnd vdd FILL
XFILL_0__9416_ gnd vdd FILL
XFILL_3__9125_ gnd vdd FILL
XFILL_1__14119_ gnd vdd FILL
XFILL_4__15279_ gnd vdd FILL
XFILL_0__14849_ gnd vdd FILL
XFILL_1__15099_ gnd vdd FILL
XFILL_1__8140_ gnd vdd FILL
XFILL_0__9347_ gnd vdd FILL
XFILL_2__15409_ gnd vdd FILL
XSFILL33880x65050 gnd vdd FILL
X_9975_ _8567_/A _9975_/B gnd _9976_/C vdd NAND2X1
XFILL_2__16389_ gnd vdd FILL
X_8926_ _8926_/Q _8926_/CLK _7262_/R vdd _8848_/Y gnd vdd DFFSR
XFILL_0__9278_ gnd vdd FILL
XFILL_1__8071_ gnd vdd FILL
XFILL_3__8007_ gnd vdd FILL
XFILL_0__8229_ gnd vdd FILL
X_8857_ _8855_/Y _8893_/B _8857_/C gnd _8929_/D vdd OAI21X1
XFILL_6__9736_ gnd vdd FILL
XSFILL39000x11050 gnd vdd FILL
X_7808_ _7872_/B _8832_/B gnd _7809_/C vdd NAND2X1
X_8788_ _8788_/A _9940_/B gnd _8789_/C vdd NAND2X1
XFILL_4__8751_ gnd vdd FILL
XSFILL3640x42050 gnd vdd FILL
X_7739_ _7739_/A gnd _7741_/A vdd INVX1
XFILL_3__8909_ gnd vdd FILL
XFILL_1__8973_ gnd vdd FILL
XFILL_4__7702_ gnd vdd FILL
XFILL_3__9889_ gnd vdd FILL
XSFILL28840x54050 gnd vdd FILL
XFILL_4__7633_ gnd vdd FILL
X_11340_ _10991_/Y _11341_/B _11835_/C gnd _11340_/Y vdd AOI21X1
X_9409_ _9455_/Q gnd _9411_/A vdd INVX1
XFILL_1__7855_ gnd vdd FILL
XFILL_4__7564_ gnd vdd FILL
XSFILL33960x45050 gnd vdd FILL
X_11271_ _11268_/Y _11270_/Y _11732_/A gnd _11271_/Y vdd AOI21X1
XFILL_4_BUFX2_insert232 gnd vdd FILL
XFILL_4_BUFX2_insert243 gnd vdd FILL
X_13010_ _13008_/Y vdd _13010_/C gnd _13066_/D vdd OAI21X1
X_10222_ _10222_/Q _8046_/CLK _9692_/R vdd _10222_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert254 gnd vdd FILL
XFILL_4_BUFX2_insert265 gnd vdd FILL
XFILL_4__7495_ gnd vdd FILL
XFILL_1__9525_ gnd vdd FILL
XFILL_4_BUFX2_insert276 gnd vdd FILL
XFILL_4_BUFX2_insert287 gnd vdd FILL
XFILL_4__9234_ gnd vdd FILL
XFILL_3_BUFX2_insert910 gnd vdd FILL
XFILL_4_BUFX2_insert298 gnd vdd FILL
X_10153_ _10215_/Q gnd _10153_/Y vdd INVX1
XFILL_3_BUFX2_insert921 gnd vdd FILL
XFILL_3_BUFX2_insert932 gnd vdd FILL
XFILL_3_BUFX2_insert943 gnd vdd FILL
XFILL_3_BUFX2_insert954 gnd vdd FILL
XFILL_4__9165_ gnd vdd FILL
XFILL_3_BUFX2_insert965 gnd vdd FILL
XFILL_2__7200_ gnd vdd FILL
X_10084_ _10016_/A _8541_/CLK _7258_/R vdd _10084_/D gnd vdd DFFSR
X_14961_ _7541_/Q gnd _14961_/Y vdd INVX1
XFILL_3_BUFX2_insert976 gnd vdd FILL
XFILL_4__8116_ gnd vdd FILL
XFILL_1__9387_ gnd vdd FILL
XFILL_3_BUFX2_insert987 gnd vdd FILL
XSFILL3720x22050 gnd vdd FILL
XFILL_3_BUFX2_insert998 gnd vdd FILL
XFILL_4__9096_ gnd vdd FILL
X_13912_ _9567_/Q gnd _13912_/Y vdd INVX1
XSFILL28920x34050 gnd vdd FILL
XFILL_1__8338_ gnd vdd FILL
X_14892_ _10100_/Q gnd _14892_/Y vdd INVX1
XSFILL94360x10050 gnd vdd FILL
X_13843_ _13842_/Y _14045_/A _13843_/C _13843_/D gnd _13847_/A vdd OAI22X1
XFILL_1__8269_ gnd vdd FILL
XFILL_3_BUFX2_insert1004 gnd vdd FILL
XFILL_2__7062_ gnd vdd FILL
XFILL_5__10580_ gnd vdd FILL
XFILL_3_BUFX2_insert1015 gnd vdd FILL
XFILL_3_BUFX2_insert1026 gnd vdd FILL
XSFILL79160x71050 gnd vdd FILL
XFILL_3_BUFX2_insert1037 gnd vdd FILL
XFILL_1_BUFX2_insert100 gnd vdd FILL
XFILL_5__8860_ gnd vdd FILL
XFILL_3_BUFX2_insert1048 gnd vdd FILL
X_13774_ _7944_/A gnd _13774_/Y vdd INVX1
X_10986_ _10906_/A _12667_/CLK _12689_/R vdd _10986_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert1059 gnd vdd FILL
XFILL_3__11690_ gnd vdd FILL
XFILL_5__7811_ gnd vdd FILL
XFILL_0__10530_ gnd vdd FILL
X_15513_ _7319_/A _15631_/B _15636_/B gnd _15514_/C vdd NAND3X1
X_12725_ _12801_/Q gnd _12727_/A vdd INVX1
XFILL_4__9998_ gnd vdd FILL
XFILL_5__12250_ gnd vdd FILL
XFILL_3__10641_ gnd vdd FILL
XFILL_2__12070_ gnd vdd FILL
XFILL_4__12980_ gnd vdd FILL
XFILL_1__11820_ gnd vdd FILL
XSFILL74120x18050 gnd vdd FILL
XFILL_5__7742_ gnd vdd FILL
XFILL_0_BUFX2_insert800 gnd vdd FILL
XFILL_5__11201_ gnd vdd FILL
XSFILL84280x62050 gnd vdd FILL
XFILL_0_BUFX2_insert811 gnd vdd FILL
X_15444_ _15444_/A _15527_/A _14999_/A _15442_/Y gnd _15446_/B vdd OAI22X1
X_12656_ _12656_/A vdd _12655_/Y gnd _12692_/D vdd OAI21X1
XFILL_4__11931_ gnd vdd FILL
XFILL_5__12181_ gnd vdd FILL
XFILL_2__11021_ gnd vdd FILL
XFILL_3__13360_ gnd vdd FILL
XFILL_3__10572_ gnd vdd FILL
XFILL_0__12200_ gnd vdd FILL
XFILL_0_BUFX2_insert822 gnd vdd FILL
XFILL_2__7964_ gnd vdd FILL
XFILL_0_BUFX2_insert833 gnd vdd FILL
XFILL_1__11751_ gnd vdd FILL
XFILL_0__10392_ gnd vdd FILL
XFILL_0_BUFX2_insert844 gnd vdd FILL
XFILL_0_BUFX2_insert855 gnd vdd FILL
X_11607_ _11121_/Y _11484_/B _11621_/C _11120_/Y gnd _11608_/A vdd OAI22X1
XFILL_5__11132_ gnd vdd FILL
XFILL_5__7673_ gnd vdd FILL
X_12587_ _12587_/A vdd _12587_/C gnd _12669_/D vdd OAI21X1
X_15375_ _13875_/Y _15169_/D gnd _15379_/A vdd NOR2X1
XFILL_3__12311_ gnd vdd FILL
XFILL_4__14650_ gnd vdd FILL
XFILL_3__13291_ gnd vdd FILL
XFILL_1__10702_ gnd vdd FILL
XFILL_2__6915_ gnd vdd FILL
XFILL_0_BUFX2_insert866 gnd vdd FILL
XFILL_1_BUFX2_insert1030 gnd vdd FILL
XFILL_4__11862_ gnd vdd FILL
XFILL_1__14470_ gnd vdd FILL
XFILL_5__9412_ gnd vdd FILL
XFILL_0_BUFX2_insert877 gnd vdd FILL
XFILL_1_BUFX2_insert1041 gnd vdd FILL
XFILL_0__12131_ gnd vdd FILL
XFILL_1_BUFX2_insert1052 gnd vdd FILL
XFILL_0_BUFX2_insert888 gnd vdd FILL
XFILL_1__11682_ gnd vdd FILL
XFILL_4__13601_ gnd vdd FILL
XFILL_0_BUFX2_insert899 gnd vdd FILL
X_14326_ _7468_/A gnd _15790_/B vdd INVX1
XFILL_4__10813_ gnd vdd FILL
XFILL_3_BUFX2_insert15 gnd vdd FILL
XFILL_3__15030_ gnd vdd FILL
XFILL_5__15940_ gnd vdd FILL
XFILL_3__12242_ gnd vdd FILL
X_11538_ _11437_/A _11537_/Y _11521_/C gnd _11538_/Y vdd AOI21X1
XFILL_5__11063_ gnd vdd FILL
XFILL_1_BUFX2_insert1063 gnd vdd FILL
XFILL_4__14581_ gnd vdd FILL
XFILL_2__9634_ gnd vdd FILL
XFILL_1__13421_ gnd vdd FILL
XFILL_3_BUFX2_insert26 gnd vdd FILL
XFILL_1_BUFX2_insert1085 gnd vdd FILL
XFILL_1__10633_ gnd vdd FILL
XFILL_2__6846_ gnd vdd FILL
XFILL112280x44050 gnd vdd FILL
XFILL_2__15760_ gnd vdd FILL
XFILL_4__11793_ gnd vdd FILL
XFILL_5__9343_ gnd vdd FILL
XFILL_2__12972_ gnd vdd FILL
XFILL_0__12062_ gnd vdd FILL
XFILL_3_BUFX2_insert37 gnd vdd FILL
XFILL_3_BUFX2_insert48 gnd vdd FILL
XFILL_4__16320_ gnd vdd FILL
XFILL_5__10014_ gnd vdd FILL
X_14257_ _9062_/Q gnd _14257_/Y vdd INVX1
XFILL_3_BUFX2_insert59 gnd vdd FILL
XSFILL79640x49050 gnd vdd FILL
X_11469_ _11226_/B _11195_/A _11423_/B gnd _11469_/Y vdd OAI21X1
XFILL_4__13532_ gnd vdd FILL
XFILL_4__10744_ gnd vdd FILL
XFILL_3__12173_ gnd vdd FILL
XFILL_2__14711_ gnd vdd FILL
XFILL_1__16140_ gnd vdd FILL
XFILL_5__15871_ gnd vdd FILL
XFILL_1__13352_ gnd vdd FILL
XFILL_2__11923_ gnd vdd FILL
XFILL_0__11013_ gnd vdd FILL
XFILL_2__15691_ gnd vdd FILL
XFILL_1__10564_ gnd vdd FILL
X_13208_ _13305_/A gnd _13209_/B vdd INVX2
XFILL_5__9274_ gnd vdd FILL
XFILL_0__7600_ gnd vdd FILL
XFILL_0__8580_ gnd vdd FILL
XFILL_5__14822_ gnd vdd FILL
XFILL_3__11124_ gnd vdd FILL
XFILL_4__16251_ gnd vdd FILL
X_14188_ _6947_/A gnd _14188_/Y vdd INVX1
XSFILL79240x51050 gnd vdd FILL
XFILL_2__8516_ gnd vdd FILL
XFILL_4__13463_ gnd vdd FILL
XFILL_1__12303_ gnd vdd FILL
XFILL_2__14642_ gnd vdd FILL
XSFILL114040x39050 gnd vdd FILL
XFILL_6_CLKBUF1_insert121 gnd vdd FILL
XFILL_0__15821_ gnd vdd FILL
XSFILL43880x28050 gnd vdd FILL
XFILL_1__16071_ gnd vdd FILL
XFILL_4__10675_ gnd vdd FILL
XFILL_2__11854_ gnd vdd FILL
XFILL_1__13283_ gnd vdd FILL
XFILL_2__9496_ gnd vdd FILL
XFILL_5__8225_ gnd vdd FILL
XFILL_6_CLKBUF1_insert132 gnd vdd FILL
XFILL_1__10495_ gnd vdd FILL
XFILL_4__15202_ gnd vdd FILL
XFILL_4__12414_ gnd vdd FILL
X_13139_ _11947_/A gnd _13139_/Y vdd INVX1
XFILL_5__14753_ gnd vdd FILL
XFILL_4__16182_ gnd vdd FILL
XFILL_5__11965_ gnd vdd FILL
XFILL_3__15932_ gnd vdd FILL
XFILL_1__15022_ gnd vdd FILL
XFILL_3__11055_ gnd vdd FILL
XFILL_3__7240_ gnd vdd FILL
XFILL_2__10805_ gnd vdd FILL
XFILL_2__8447_ gnd vdd FILL
XFILL_4__13394_ gnd vdd FILL
XFILL_1__12234_ gnd vdd FILL
XFILL_2__14573_ gnd vdd FILL
XFILL_2__11785_ gnd vdd FILL
XFILL_0__15752_ gnd vdd FILL
XSFILL114440x60050 gnd vdd FILL
XFILL_0__12964_ gnd vdd FILL
XSFILL8520x14050 gnd vdd FILL
XFILL_0__7462_ gnd vdd FILL
XFILL_5__10916_ gnd vdd FILL
XFILL_6_CLKBUF1_insert198 gnd vdd FILL
XFILL_3__10006_ gnd vdd FILL
XFILL_4__15133_ gnd vdd FILL
XFILL_5__13704_ gnd vdd FILL
XFILL_4__12345_ gnd vdd FILL
XFILL_2__16312_ gnd vdd FILL
XFILL_5__14684_ gnd vdd FILL
XFILL_3__7171_ gnd vdd FILL
XFILL_5__11896_ gnd vdd FILL
XFILL_0__14703_ gnd vdd FILL
XSFILL99640x2050 gnd vdd FILL
XFILL_2__13524_ gnd vdd FILL
XFILL_3__15863_ gnd vdd FILL
XFILL_2__8378_ gnd vdd FILL
XFILL_0__11915_ gnd vdd FILL
XFILL_1__12165_ gnd vdd FILL
XFILL_5__7107_ gnd vdd FILL
XFILL_0__15683_ gnd vdd FILL
XFILL_5__13635_ gnd vdd FILL
XFILL_0__12895_ gnd vdd FILL
XFILL_5__8087_ gnd vdd FILL
XSFILL59000x59050 gnd vdd FILL
XFILL_3__14814_ gnd vdd FILL
XFILL_4__15064_ gnd vdd FILL
XFILL_2__16243_ gnd vdd FILL
XFILL_2__7329_ gnd vdd FILL
XSFILL9400x42050 gnd vdd FILL
XFILL_4__12276_ gnd vdd FILL
XFILL_1__11116_ gnd vdd FILL
XFILL_0__14634_ gnd vdd FILL
XSFILL99400x64050 gnd vdd FILL
XFILL_2__13455_ gnd vdd FILL
XFILL_3__15794_ gnd vdd FILL
XFILL_2__10667_ gnd vdd FILL
XFILL_1__12096_ gnd vdd FILL
XFILL_0__9132_ gnd vdd FILL
XFILL_5__7038_ gnd vdd FILL
XFILL_0__11846_ gnd vdd FILL
XFILL_4__14015_ gnd vdd FILL
X_9760_ _9760_/A gnd _9760_/Y vdd INVX1
XFILL_5__16354_ gnd vdd FILL
XFILL_5__13566_ gnd vdd FILL
XFILL_4__11227_ gnd vdd FILL
X_6972_ _6951_/A _7868_/B gnd _6972_/Y vdd NAND2X1
XFILL_2__12406_ gnd vdd FILL
XFILL_5__10778_ gnd vdd FILL
XFILL_3__14745_ gnd vdd FILL
XFILL_1__15924_ gnd vdd FILL
XFILL_2__16174_ gnd vdd FILL
XFILL_3__11957_ gnd vdd FILL
XFILL_2__13386_ gnd vdd FILL
XFILL_1__11047_ gnd vdd FILL
XFILL_0__14565_ gnd vdd FILL
XFILL_5__15305_ gnd vdd FILL
XFILL_5__12517_ gnd vdd FILL
X_8711_ _8711_/A _8698_/A _8710_/Y gnd _8795_/D vdd OAI21X1
XFILL_0__11777_ gnd vdd FILL
XFILL_6__14856_ gnd vdd FILL
XFILL_5__16285_ gnd vdd FILL
XFILL_3__10908_ gnd vdd FILL
XFILL_0__16304_ gnd vdd FILL
X_9691_ _9691_/Q _8151_/CLK _9048_/R vdd _9691_/D gnd vdd DFFSR
XFILL_5__13497_ gnd vdd FILL
XFILL_4__11158_ gnd vdd FILL
XFILL_2__15125_ gnd vdd FILL
XFILL_2__12337_ gnd vdd FILL
XFILL_3__14676_ gnd vdd FILL
XFILL_0__13516_ gnd vdd FILL
XFILL_0__8014_ gnd vdd FILL
XSFILL49480x68050 gnd vdd FILL
XFILL_3__11888_ gnd vdd FILL
XFILL_6_BUFX2_insert316 gnd vdd FILL
XFILL_1__15855_ gnd vdd FILL
XFILL_0__14496_ gnd vdd FILL
XFILL_6__13807_ gnd vdd FILL
XFILL_5__15236_ gnd vdd FILL
XFILL_5__12448_ gnd vdd FILL
XFILL_3__16415_ gnd vdd FILL
X_8642_ _8607_/B _8642_/B gnd _8643_/C vdd NAND2X1
XFILL_5__8989_ gnd vdd FILL
XFILL_4__10109_ gnd vdd FILL
XFILL_3__13627_ gnd vdd FILL
XFILL_3__9812_ gnd vdd FILL
XFILL_0__16235_ gnd vdd FILL
XFILL_1__14806_ gnd vdd FILL
XFILL_2__15056_ gnd vdd FILL
XFILL_4__15966_ gnd vdd FILL
XFILL_2__12268_ gnd vdd FILL
XFILL_4__11089_ gnd vdd FILL
XFILL_0__13447_ gnd vdd FILL
XFILL_0__10659_ gnd vdd FILL
XFILL_1__12998_ gnd vdd FILL
XFILL_1__15786_ gnd vdd FILL
XSFILL79320x31050 gnd vdd FILL
XFILL_5__15167_ gnd vdd FILL
XFILL_3__16346_ gnd vdd FILL
XFILL_2__14007_ gnd vdd FILL
XFILL_5__12379_ gnd vdd FILL
X_8573_ _8619_/B _9981_/B gnd _8574_/C vdd NAND2X1
XFILL_4__14917_ gnd vdd FILL
XFILL_2__11219_ gnd vdd FILL
XFILL_3__9743_ gnd vdd FILL
XFILL_4__15897_ gnd vdd FILL
XFILL_3__13558_ gnd vdd FILL
XFILL_0__16166_ gnd vdd FILL
XFILL_1__11949_ gnd vdd FILL
XFILL_1__14737_ gnd vdd FILL
XFILL_2__12199_ gnd vdd FILL
XFILL_3__6955_ gnd vdd FILL
XFILL_0__13378_ gnd vdd FILL
XFILL_5__14118_ gnd vdd FILL
X_7524_ _7456_/A _8161_/CLK _7140_/R vdd _7524_/D gnd vdd DFFSR
XFILL_4__14848_ gnd vdd FILL
XSFILL28760x69050 gnd vdd FILL
XFILL_6__13669_ gnd vdd FILL
XFILL_3__12509_ gnd vdd FILL
XFILL_5__15098_ gnd vdd FILL
XFILL_0__15117_ gnd vdd FILL
XFILL_3__16277_ gnd vdd FILL
XFILL_3__9674_ gnd vdd FILL
XFILL_0__12329_ gnd vdd FILL
XFILL_3__13489_ gnd vdd FILL
XSFILL44040x17050 gnd vdd FILL
XFILL_6__15408_ gnd vdd FILL
XFILL_3__6886_ gnd vdd FILL
XFILL_0__16097_ gnd vdd FILL
XFILL_1__14668_ gnd vdd FILL
XFILL_5__14049_ gnd vdd FILL
XFILL_0__8916_ gnd vdd FILL
XFILL_3__15228_ gnd vdd FILL
X_7455_ _7455_/A _7430_/A _7454_/Y gnd _7455_/Y vdd OAI21X1
XFILL_0__9896_ gnd vdd FILL
XFILL_1__16407_ gnd vdd FILL
XFILL_3__8625_ gnd vdd FILL
XFILL_4__14779_ gnd vdd FILL
XFILL_1__13619_ gnd vdd FILL
XFILL_0__15048_ gnd vdd FILL
XFILL_2__15958_ gnd vdd FILL
XFILL_1__14599_ gnd vdd FILL
XFILL_0__8847_ gnd vdd FILL
XSFILL69240x83050 gnd vdd FILL
X_7386_ _7298_/A _8541_/CLK _7258_/R vdd _7386_/D gnd vdd DFFSR
XFILL_3__15159_ gnd vdd FILL
XFILL_2__14909_ gnd vdd FILL
XFILL_1__16338_ gnd vdd FILL
XFILL_2__15889_ gnd vdd FILL
X_9125_ _9125_/A _9163_/A _9125_/C gnd _9189_/D vdd OAI21X1
XFILL111800x38050 gnd vdd FILL
XFILL_4__16449_ gnd vdd FILL
XFILL_1__7571_ gnd vdd FILL
XFILL_0__8778_ gnd vdd FILL
XFILL_3__7507_ gnd vdd FILL
XFILL_3__8487_ gnd vdd FILL
XFILL_1__16269_ gnd vdd FILL
XFILL_3_BUFX2_insert228 gnd vdd FILL
XFILL_6__8196_ gnd vdd FILL
XFILL_0__7729_ gnd vdd FILL
X_9056_ _8980_/A _7647_/CLK _9056_/R vdd _8982_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert239 gnd vdd FILL
XFILL_3__7438_ gnd vdd FILL
X_8007_ _8049_/Q gnd _8009_/A vdd INVX1
XFILL_1__9241_ gnd vdd FILL
XFILL_2_BUFX2_insert906 gnd vdd FILL
XSFILL49160x50050 gnd vdd FILL
XFILL_3__7369_ gnd vdd FILL
XFILL_2_BUFX2_insert917 gnd vdd FILL
XSFILL3640x37050 gnd vdd FILL
XFILL_1__9172_ gnd vdd FILL
XFILL_3__9108_ gnd vdd FILL
XFILL_2_BUFX2_insert928 gnd vdd FILL
XFILL_2_BUFX2_insert939 gnd vdd FILL
XFILL_1__8123_ gnd vdd FILL
XSFILL28840x49050 gnd vdd FILL
XSFILL114600x20050 gnd vdd FILL
XSFILL94280x25050 gnd vdd FILL
XFILL_3__9039_ gnd vdd FILL
X_9958_ _9958_/Q _9958_/CLK _7270_/R vdd _9958_/D gnd vdd DFFSR
XFILL_4__9921_ gnd vdd FILL
X_10840_ _13568_/C _7640_/CLK _7515_/R vdd _10750_/Y gnd vdd DFFSR
XFILL_1__8054_ gnd vdd FILL
X_8909_ _8909_/A gnd _8909_/Y vdd INVX1
X_9889_ _9868_/A _9889_/B gnd _9890_/C vdd NAND2X1
XFILL_4__9852_ gnd vdd FILL
X_10771_ _10769_/Y _10773_/A _10771_/C gnd _10847_/D vdd OAI21X1
XBUFX2_insert905 _10913_/Y gnd _12762_/A vdd BUFX2
XFILL_4__9783_ gnd vdd FILL
X_12510_ _12508_/Y vdd _12509_/Y gnd _12510_/Y vdd OAI21X1
XBUFX2_insert916 _15069_/Y gnd _16002_/A vdd BUFX2
X_13490_ _13587_/C gnd _13490_/Y vdd INVX8
XFILL_0_BUFX2_insert107 gnd vdd FILL
XFILL_4__6995_ gnd vdd FILL
XBUFX2_insert927 _12351_/Y gnd _7037_/B vdd BUFX2
XBUFX2_insert938 _13423_/Y gnd _13978_/B vdd BUFX2
XFILL_6_BUFX2_insert894 gnd vdd FILL
XBUFX2_insert949 _11987_/Y gnd _12093_/B vdd BUFX2
XFILL_4__8734_ gnd vdd FILL
X_12441_ _12441_/A vdd _12440_/Y gnd _12535_/D vdd OAI21X1
XSFILL74440x54050 gnd vdd FILL
XFILL_1__8956_ gnd vdd FILL
XSFILL89240x14050 gnd vdd FILL
X_12372_ _12370_/Y _12419_/A _12372_/C gnd _12372_/Y vdd OAI21X1
X_15160_ _15160_/A _15157_/Y gnd _15165_/B vdd NOR2X1
XFILL_2__7680_ gnd vdd FILL
XFILL_1__8887_ gnd vdd FILL
XFILL_4__7616_ gnd vdd FILL
XSFILL3720x17050 gnd vdd FILL
X_11323_ _11182_/Y _11181_/Y gnd _11498_/A vdd NOR2X1
X_14111_ _14111_/A _14752_/C gnd _14112_/C vdd NOR2X1
XFILL_4__8596_ gnd vdd FILL
X_15091_ _16225_/C gnd _15091_/Y vdd INVX8
XFILL_1__7838_ gnd vdd FILL
XFILL_4__7547_ gnd vdd FILL
X_14042_ _14041_/Y _13843_/C gnd _14046_/A vdd NOR2X1
X_11254_ _11018_/Y gnd _11254_/Y vdd INVX1
XFILL_2__9350_ gnd vdd FILL
XSFILL13720x71050 gnd vdd FILL
XSFILL14200x78050 gnd vdd FILL
X_10205_ _10205_/Q _7261_/CLK _7531_/R vdd _10125_/Y gnd vdd DFFSR
XFILL_4__7478_ gnd vdd FILL
XSFILL79160x66050 gnd vdd FILL
XFILL_1__9508_ gnd vdd FILL
XSFILL29000x38050 gnd vdd FILL
X_11185_ _11185_/A _11185_/B _11185_/C gnd _11207_/B vdd OAI21X1
XFILL_4__9217_ gnd vdd FILL
XFILL_5__8010_ gnd vdd FILL
XFILL_2__9281_ gnd vdd FILL
XFILL_1__10280_ gnd vdd FILL
XFILL_3_BUFX2_insert740 gnd vdd FILL
X_10136_ _10169_/A _8088_/B gnd _10137_/C vdd NAND2X1
XFILL_3_BUFX2_insert751 gnd vdd FILL
XFILL_5__11750_ gnd vdd FILL
XSFILL114360x75050 gnd vdd FILL
X_15993_ _15991_/Y _15993_/B gnd _15993_/Y vdd NOR2X1
XFILL_2__8232_ gnd vdd FILL
XFILL_4__10391_ gnd vdd FILL
XFILL_3_BUFX2_insert762 gnd vdd FILL
XSFILL8440x29050 gnd vdd FILL
XFILL_3_BUFX2_insert773 gnd vdd FILL
XFILL_2__11570_ gnd vdd FILL
XFILL_4__9148_ gnd vdd FILL
XFILL_3_BUFX2_insert784 gnd vdd FILL
XFILL_5__10701_ gnd vdd FILL
XSFILL33640x22050 gnd vdd FILL
XSFILL84280x57050 gnd vdd FILL
XFILL_3_BUFX2_insert795 gnd vdd FILL
X_10067_ _10067_/A gnd _10067_/Y vdd INVX1
X_14944_ _10741_/Q gnd _14946_/B vdd INVX1
XFILL_4__12130_ gnd vdd FILL
XFILL_2__10521_ gnd vdd FILL
XFILL_5__11681_ gnd vdd FILL
XFILL_3__12860_ gnd vdd FILL
XFILL_0__11700_ gnd vdd FILL
XSFILL98840x72050 gnd vdd FILL
XSFILL9320x57050 gnd vdd FILL
XFILL_4__9079_ gnd vdd FILL
XFILL_5__13420_ gnd vdd FILL
XFILL_5__10632_ gnd vdd FILL
XFILL_2__13240_ gnd vdd FILL
XFILL_2__7114_ gnd vdd FILL
X_14875_ _14873_/Y _13871_/D _13467_/A _14875_/D gnd _14876_/A vdd OAI22X1
XFILL_4__12061_ gnd vdd FILL
XFILL_6__12971_ gnd vdd FILL
XSFILL59080x33050 gnd vdd FILL
XFILL_3__11811_ gnd vdd FILL
XFILL_2__10452_ gnd vdd FILL
XFILL_2__8094_ gnd vdd FILL
XFILL_0__11631_ gnd vdd FILL
XFILL_1__13970_ gnd vdd FILL
XFILL_5__8912_ gnd vdd FILL
XFILL_5__13351_ gnd vdd FILL
XFILL_5__9892_ gnd vdd FILL
X_13826_ _13826_/A _13826_/B _13825_/Y gnd _13839_/A vdd NAND3X1
XFILL_6__11922_ gnd vdd FILL
XFILL_4__11012_ gnd vdd FILL
XFILL_6__15690_ gnd vdd FILL
XFILL_3__14530_ gnd vdd FILL
XFILL_2__7045_ gnd vdd FILL
XFILL_5__10563_ gnd vdd FILL
XFILL_2__13171_ gnd vdd FILL
XFILL_3__11742_ gnd vdd FILL
XFILL_2__10383_ gnd vdd FILL
XFILL_0__14350_ gnd vdd FILL
XFILL_5__8843_ gnd vdd FILL
XFILL_5__12302_ gnd vdd FILL
XFILL_0__11562_ gnd vdd FILL
XFILL_6__14641_ gnd vdd FILL
XFILL_5__16070_ gnd vdd FILL
XFILL_5__13282_ gnd vdd FILL
X_13757_ _7432_/A gnd _13758_/D vdd INVX1
XFILL_4__15820_ gnd vdd FILL
XFILL_2__12122_ gnd vdd FILL
XFILL_0__13301_ gnd vdd FILL
X_10969_ _10935_/A _10934_/Y _10969_/C _10969_/D gnd _10970_/A vdd OAI22X1
XFILL_3__14461_ gnd vdd FILL
XFILL_5__10494_ gnd vdd FILL
XFILL_1__15640_ gnd vdd FILL
XFILL_3__11673_ gnd vdd FILL
XFILL_1__12852_ gnd vdd FILL
XFILL_0__10513_ gnd vdd FILL
XFILL_5__15021_ gnd vdd FILL
XFILL_0__14281_ gnd vdd FILL
X_12708_ _10944_/C memoryOutData[4] gnd _12709_/C vdd NAND2X1
XFILL_3__16200_ gnd vdd FILL
XSFILL13800x51050 gnd vdd FILL
XFILL_5__8774_ gnd vdd FILL
XFILL_5__12233_ gnd vdd FILL
XSFILL74200x7050 gnd vdd FILL
XFILL_0__11493_ gnd vdd FILL
XFILL_3__13412_ gnd vdd FILL
XFILL_4__15751_ gnd vdd FILL
XFILL_6__11784_ gnd vdd FILL
XFILL_3__10624_ gnd vdd FILL
XFILL_0__16020_ gnd vdd FILL
XFILL_4__12963_ gnd vdd FILL
XFILL_2__12053_ gnd vdd FILL
X_13688_ _8069_/A gnd _13689_/A vdd INVX1
XFILL_1__11803_ gnd vdd FILL
XFILL_0__13232_ gnd vdd FILL
XSFILL79240x46050 gnd vdd FILL
XFILL_1__15571_ gnd vdd FILL
XFILL_3__14392_ gnd vdd FILL
XFILL_1__12783_ gnd vdd FILL
XFILL_0__10444_ gnd vdd FILL
XFILL_2__8996_ gnd vdd FILL
XFILL_0_BUFX2_insert630 gnd vdd FILL
XFILL_5__7725_ gnd vdd FILL
XFILL_4__14702_ gnd vdd FILL
X_15427_ _7007_/Q _15382_/B _16096_/C _7391_/Q gnd _15433_/A vdd AOI22X1
X_12639_ _12639_/A gnd _12639_/Y vdd INVX1
XFILL_4__11914_ gnd vdd FILL
XFILL_5__12164_ gnd vdd FILL
XFILL_3__16131_ gnd vdd FILL
XFILL_2__11004_ gnd vdd FILL
XFILL_0_BUFX2_insert641 gnd vdd FILL
XFILL_3__13343_ gnd vdd FILL
XFILL_4__15682_ gnd vdd FILL
XFILL_0_BUFX2_insert652 gnd vdd FILL
XFILL_2__7947_ gnd vdd FILL
XFILL_4__12894_ gnd vdd FILL
XFILL_3__10555_ gnd vdd FILL
XFILL_1__14522_ gnd vdd FILL
XFILL_1__11734_ gnd vdd FILL
XFILL_0_BUFX2_insert663 gnd vdd FILL
XFILL_0__13163_ gnd vdd FILL
XFILL_0_BUFX2_insert674 gnd vdd FILL
XFILL_6__16242_ gnd vdd FILL
XFILL_0__10375_ gnd vdd FILL
XFILL_5__11115_ gnd vdd FILL
XSFILL43480x25050 gnd vdd FILL
X_15358_ _9995_/A gnd _15358_/Y vdd INVX1
XFILL_4__14633_ gnd vdd FILL
XFILL_6__13454_ gnd vdd FILL
XFILL_0_BUFX2_insert685 gnd vdd FILL
XFILL_0__9750_ gnd vdd FILL
XFILL_0_BUFX2_insert696 gnd vdd FILL
XFILL_5__12095_ gnd vdd FILL
XFILL_2__15812_ gnd vdd FILL
XFILL_0__6962_ gnd vdd FILL
XFILL_3__16062_ gnd vdd FILL
XFILL_4__11845_ gnd vdd FILL
XFILL_3__13274_ gnd vdd FILL
XFILL_1__14453_ gnd vdd FILL
XFILL_3__10486_ gnd vdd FILL
XFILL_0__12114_ gnd vdd FILL
XSFILL84360x37050 gnd vdd FILL
XFILL_2__7878_ gnd vdd FILL
XFILL_1__11665_ gnd vdd FILL
XFILL_0__13094_ gnd vdd FILL
X_14309_ _7911_/Q _13865_/B _14309_/C gnd _14310_/B vdd AOI21X1
XFILL_0__8701_ gnd vdd FILL
XFILL_5__15923_ gnd vdd FILL
XFILL_5__7587_ gnd vdd FILL
XFILL_3__15013_ gnd vdd FILL
XFILL_5__11046_ gnd vdd FILL
X_7240_ _7210_/A _7240_/B gnd _7240_/Y vdd NAND2X1
XFILL_0__6893_ gnd vdd FILL
XFILL_4__14564_ gnd vdd FILL
XFILL_1__13404_ gnd vdd FILL
XFILL_3__12225_ gnd vdd FILL
X_15289_ _15289_/A _15286_/Y gnd _15294_/B vdd NOR2X1
XFILL_2__9617_ gnd vdd FILL
XFILL_0__9681_ gnd vdd FILL
XFILL_1__10616_ gnd vdd FILL
XFILL_4__11776_ gnd vdd FILL
XFILL_2__15743_ gnd vdd FILL
XFILL_0__12045_ gnd vdd FILL
XFILL_3__9390_ gnd vdd FILL
XFILL_1__14384_ gnd vdd FILL
XFILL_2__12955_ gnd vdd FILL
XSFILL99400x59050 gnd vdd FILL
XFILL_4__16303_ gnd vdd FILL
XFILL_6__12336_ gnd vdd FILL
XFILL_1__11596_ gnd vdd FILL
XSFILL59160x13050 gnd vdd FILL
XFILL_0__8632_ gnd vdd FILL
XFILL_4__13515_ gnd vdd FILL
X_7171_ _7181_/B _9347_/B gnd _7172_/C vdd NAND2X1
XFILL_5__15854_ gnd vdd FILL
XFILL_1__13335_ gnd vdd FILL
XFILL_2__9548_ gnd vdd FILL
XFILL_4__14495_ gnd vdd FILL
XFILL_2__11906_ gnd vdd FILL
XFILL_1__16123_ gnd vdd FILL
XFILL_3__8341_ gnd vdd FILL
XFILL_3__12156_ gnd vdd FILL
XFILL_2__15674_ gnd vdd FILL
XFILL_1__10547_ gnd vdd FILL
XFILL_2__12886_ gnd vdd FILL
XFILL_5__9257_ gnd vdd FILL
XFILL_5__14805_ gnd vdd FILL
XFILL_4__16234_ gnd vdd FILL
XFILL_6__15055_ gnd vdd FILL
XFILL111880x12050 gnd vdd FILL
XFILL_4__13446_ gnd vdd FILL
XFILL_3__11107_ gnd vdd FILL
XFILL112360x19050 gnd vdd FILL
XFILL_5__12997_ gnd vdd FILL
XFILL_2__14625_ gnd vdd FILL
XFILL_4__10658_ gnd vdd FILL
XFILL_3__12087_ gnd vdd FILL
XFILL_5__15785_ gnd vdd FILL
XFILL_1__16054_ gnd vdd FILL
XFILL_5__8208_ gnd vdd FILL
XFILL_1__13266_ gnd vdd FILL
XFILL_0__15804_ gnd vdd FILL
XFILL_2__9479_ gnd vdd FILL
XFILL_3__8272_ gnd vdd FILL
XFILL_2__11837_ gnd vdd FILL
XFILL_0__13996_ gnd vdd FILL
XFILL_3__15915_ gnd vdd FILL
XFILL_4__16165_ gnd vdd FILL
XFILL_5__11948_ gnd vdd FILL
XFILL_1__15005_ gnd vdd FILL
XFILL_5__14736_ gnd vdd FILL
XFILL_6__12198_ gnd vdd FILL
XFILL_0__8494_ gnd vdd FILL
XFILL_3__11038_ gnd vdd FILL
XFILL_3__7223_ gnd vdd FILL
XFILL_4__13377_ gnd vdd FILL
XFILL_1__12217_ gnd vdd FILL
XFILL_2__14556_ gnd vdd FILL
XFILL_5__8139_ gnd vdd FILL
XFILL_2__11768_ gnd vdd FILL
XFILL_0__15735_ gnd vdd FILL
XFILL_0__7445_ gnd vdd FILL
XFILL_6__11149_ gnd vdd FILL
XFILL_4__15116_ gnd vdd FILL
XSFILL49080x65050 gnd vdd FILL
XFILL_4__12328_ gnd vdd FILL
XSFILL79320x26050 gnd vdd FILL
XFILL112200x83050 gnd vdd FILL
XFILL_5__11879_ gnd vdd FILL
XFILL_4__16096_ gnd vdd FILL
XFILL_3__15846_ gnd vdd FILL
XSFILL63880x6050 gnd vdd FILL
XFILL_5__14667_ gnd vdd FILL
XFILL_2__13507_ gnd vdd FILL
XFILL_1__12148_ gnd vdd FILL
XFILL_0__15666_ gnd vdd FILL
XFILL_2__14487_ gnd vdd FILL
XFILL_2__11699_ gnd vdd FILL
XFILL_5__16406_ gnd vdd FILL
XFILL_0__12878_ gnd vdd FILL
XFILL_5__13618_ gnd vdd FILL
XFILL_4__15047_ gnd vdd FILL
X_9812_ _9813_/B _9940_/B gnd _9812_/Y vdd NAND2X1
XFILL_0__7376_ gnd vdd FILL
XFILL_5__14598_ gnd vdd FILL
XFILL_2__16226_ gnd vdd FILL
XFILL_4__12259_ gnd vdd FILL
XFILL_0__14617_ gnd vdd FILL
XSFILL114520x35050 gnd vdd FILL
XFILL_3__15777_ gnd vdd FILL
XFILL_3__7085_ gnd vdd FILL
XFILL_2__13438_ gnd vdd FILL
XFILL_1__12079_ gnd vdd FILL
XFILL_3__12989_ gnd vdd FILL
XFILL_0__11829_ gnd vdd FILL
XFILL_0__9115_ gnd vdd FILL
XSFILL83960x10050 gnd vdd FILL
XFILL_0__15597_ gnd vdd FILL
XFILL_5__13549_ gnd vdd FILL
XFILL_6__8883_ gnd vdd FILL
XFILL_5__16337_ gnd vdd FILL
X_9743_ _9764_/A _9487_/B gnd _9744_/C vdd NAND2X1
XFILL_3__14728_ gnd vdd FILL
X_6955_ _6955_/A _6955_/B _6954_/Y gnd _7015_/D vdd OAI21X1
XFILL_1__15907_ gnd vdd FILL
XFILL_2__16157_ gnd vdd FILL
XFILL_2__13369_ gnd vdd FILL
XFILL_0__14548_ gnd vdd FILL
XFILL_6__7834_ gnd vdd FILL
XSFILL44440x33050 gnd vdd FILL
X_9674_ _9674_/A gnd _9676_/A vdd INVX1
XFILL_5__16268_ gnd vdd FILL
XFILL_2__15108_ gnd vdd FILL
X_6886_ _6886_/A gnd memoryWriteData[16] vdd BUFX2
XFILL_3__14659_ gnd vdd FILL
XFILL_2__16088_ gnd vdd FILL
XFILL_1__15838_ gnd vdd FILL
XFILL_0__14479_ gnd vdd FILL
XFILL_5__15219_ gnd vdd FILL
X_8625_ _8623_/Y _8609_/A _8624_/Y gnd _8681_/D vdd OAI21X1
XFILL_5__16199_ gnd vdd FILL
XFILL_0__16218_ gnd vdd FILL
XFILL_2__15039_ gnd vdd FILL
XFILL_4__15949_ gnd vdd FILL
XFILL_5_BUFX2_insert802 gnd vdd FILL
XFILL_1__15769_ gnd vdd FILL
XFILL_3__7987_ gnd vdd FILL
XFILL_5_BUFX2_insert813 gnd vdd FILL
X_8556_ _8556_/Q _9453_/CLK _9453_/R vdd _8506_/Y gnd vdd DFFSR
XFILL_3__16329_ gnd vdd FILL
XFILL_5_BUFX2_insert824 gnd vdd FILL
XFILL_1__9790_ gnd vdd FILL
XFILL_5_BUFX2_insert835 gnd vdd FILL
XFILL_3__9726_ gnd vdd FILL
XBUFX2_insert1010 _13569_/Y gnd _13645_/C vdd BUFX2
XFILL_3__6938_ gnd vdd FILL
XFILL_0__16149_ gnd vdd FILL
XFILL_5_BUFX2_insert846 gnd vdd FILL
XBUFX2_insert1021 _13340_/Y gnd _9652_/B vdd BUFX2
X_7507_ _7541_/Q gnd _7507_/Y vdd INVX1
XFILL_5_BUFX2_insert857 gnd vdd FILL
XFILL_1__8741_ gnd vdd FILL
XBUFX2_insert1032 _13333_/Y gnd _9277_/B vdd BUFX2
XFILL_5_BUFX2_insert868 gnd vdd FILL
XBUFX2_insert1043 _13297_/Y gnd _7759_/B vdd BUFX2
X_8487_ _8508_/A _9383_/B gnd _8488_/C vdd NAND2X1
XFILL_5_BUFX2_insert879 gnd vdd FILL
XSFILL18840x2050 gnd vdd FILL
XBUFX2_insert1054 _13527_/Y gnd _14470_/B vdd BUFX2
XFILL_4__8450_ gnd vdd FILL
XFILL_3__9657_ gnd vdd FILL
XFILL_3__6869_ gnd vdd FILL
XBUFX2_insert1065 _14992_/Y gnd _16261_/A vdd BUFX2
X_7438_ _7518_/Q gnd _7440_/A vdd INVX1
XBUFX2_insert1087 rst gnd BUFX2_insert607/A vdd BUFX2
XFILL_3__8608_ gnd vdd FILL
XFILL_0__9879_ gnd vdd FILL
XFILL_4__8381_ gnd vdd FILL
XFILL_1__7623_ gnd vdd FILL
X_7369_ _7367_/Y _7369_/B _7369_/C gnd _7409_/D vdd OAI21X1
XFILL_4__7332_ gnd vdd FILL
X_9108_ _9184_/Q gnd _9108_/Y vdd INVX1
XFILL_1__7554_ gnd vdd FILL
XSFILL4120x62050 gnd vdd FILL
X_9039_ _9037_/Y _8961_/B _9039_/C gnd _9075_/D vdd OAI21X1
XSFILL69320x58050 gnd vdd FILL
XFILL_1__7485_ gnd vdd FILL
XSFILL108600x8050 gnd vdd FILL
XFILL_4__9002_ gnd vdd FILL
XFILL_4__7194_ gnd vdd FILL
XFILL_1__9224_ gnd vdd FILL
XFILL_2_BUFX2_insert703 gnd vdd FILL
XFILL_2_BUFX2_insert714 gnd vdd FILL
X_12990_ _6883_/A gnd _12990_/Y vdd INVX1
XSFILL104520x67050 gnd vdd FILL
XFILL_2_BUFX2_insert725 gnd vdd FILL
XFILL_2_BUFX2_insert736 gnd vdd FILL
X_11941_ _13133_/A gnd _11941_/Y vdd INVX1
XFILL_2_BUFX2_insert747 gnd vdd FILL
XFILL_2_BUFX2_insert758 gnd vdd FILL
XFILL_1__9155_ gnd vdd FILL
XFILL_2_BUFX2_insert769 gnd vdd FILL
XSFILL84200x2050 gnd vdd FILL
X_14660_ _14660_/A gnd _14662_/D vdd INVX1
XFILL_1__8106_ gnd vdd FILL
X_11872_ _12807_/Q gnd _11874_/A vdd INVX1
XFILL_4__9904_ gnd vdd FILL
XFILL_1__9086_ gnd vdd FILL
XSFILL74040x51050 gnd vdd FILL
X_13611_ _13611_/A _13611_/B gnd _13637_/A vdd NOR2X1
X_10823_ _14774_/D gnd _10823_/Y vdd INVX1
X_14591_ _9069_/Q gnd _14591_/Y vdd INVX1
X_16330_ _13594_/A gnd _16332_/A vdd INVX1
XSFILL44520x3050 gnd vdd FILL
XBUFX2_insert702 _11985_/Y gnd _11996_/C vdd BUFX2
X_13542_ _7292_/A _14353_/A _14273_/C _8536_/Q gnd _13544_/A vdd AOI22X1
X_10754_ _15237_/A gnd _10756_/A vdd INVX1
XBUFX2_insert713 _15023_/Y gnd _15527_/C vdd BUFX2
XBUFX2_insert724 _13352_/Y gnd _10166_/A vdd BUFX2
XFILL_2__8850_ gnd vdd FILL
XSFILL13720x66050 gnd vdd FILL
XFILL_4__9766_ gnd vdd FILL
XBUFX2_insert735 _15020_/Y gnd _15114_/B vdd BUFX2
XBUFX2_insert746 _15055_/Y gnd _15203_/B vdd BUFX2
XFILL_4__6978_ gnd vdd FILL
X_16261_ _16261_/A _14911_/Y _14910_/Y _16261_/D gnd _16262_/C vdd OAI22X1
X_10685_ _10685_/A _10678_/A _10685_/C gnd _10733_/D vdd OAI21X1
X_13473_ _13473_/A _13467_/Y gnd _13473_/Y vdd NOR2X1
XBUFX2_insert757 _12213_/Y gnd _12272_/C vdd BUFX2
XFILL_2__7801_ gnd vdd FILL
XBUFX2_insert768 _12393_/Y gnd _7975_/B vdd BUFX2
XFILL_2__8781_ gnd vdd FILL
XFILL_4__8717_ gnd vdd FILL
XFILL_1__9988_ gnd vdd FILL
XBUFX2_insert779 _10911_/Y gnd _12201_/B vdd BUFX2
X_15212_ _15064_/A _15212_/B gnd _15656_/C vdd NAND2X1
X_12424_ _11969_/B gnd _12424_/Y vdd INVX1
XFILL_5__8490_ gnd vdd FILL
X_16192_ _15170_/D _14830_/D _16191_/Y gnd _16195_/A vdd OAI21X1
XFILL_2__7732_ gnd vdd FILL
XFILL_0__10160_ gnd vdd FILL
XFILL_5__7441_ gnd vdd FILL
XFILL_4__8648_ gnd vdd FILL
X_15143_ _15143_/A _15143_/B _15142_/Y gnd _15144_/A vdd NAND3X1
XFILL_1_CLKBUF1_insert140 gnd vdd FILL
X_12355_ _12355_/A gnd _12355_/Y vdd INVX1
XFILL_4__11630_ gnd vdd FILL
XFILL_3__10271_ gnd vdd FILL
XFILL_1_CLKBUF1_insert151 gnd vdd FILL
XFILL_1__11450_ gnd vdd FILL
XFILL_1_CLKBUF1_insert162 gnd vdd FILL
XFILL_5__7372_ gnd vdd FILL
XFILL_1_CLKBUF1_insert173 gnd vdd FILL
XFILL_4__8579_ gnd vdd FILL
X_11306_ _11591_/A _11121_/Y _11591_/C gnd _11307_/A vdd OAI21X1
X_15074_ _15073_/Y _15074_/B gnd _15074_/Y vdd NOR2X1
XFILL_1_CLKBUF1_insert184 gnd vdd FILL
XFILL_3__12010_ gnd vdd FILL
XFILL_2__9402_ gnd vdd FILL
X_12286_ _12283_/Y _12286_/B _12286_/C gnd _11150_/B vdd NAND3X1
XFILL_1_CLKBUF1_insert195 gnd vdd FILL
XFILL_1__10401_ gnd vdd FILL
XSFILL59080x28050 gnd vdd FILL
XFILL_4__11561_ gnd vdd FILL
XFILL_2__12740_ gnd vdd FILL
XFILL_5__9111_ gnd vdd FILL
XFILL_6__12121_ gnd vdd FILL
XFILL_2_BUFX2_insert5 gnd vdd FILL
XFILL_2__7594_ gnd vdd FILL
XFILL_1__11381_ gnd vdd FILL
XFILL_4__13300_ gnd vdd FILL
X_14025_ _10778_/A gnd _14025_/Y vdd INVX1
XSFILL99480x33050 gnd vdd FILL
X_11237_ _11236_/Y _11235_/Y gnd _11241_/C vdd NOR2X1
XFILL_4__10512_ gnd vdd FILL
XFILL_5__12851_ gnd vdd FILL
XFILL_1__13120_ gnd vdd FILL
XFILL_4__14280_ gnd vdd FILL
XFILL_4__11492_ gnd vdd FILL
XFILL_0__13850_ gnd vdd FILL
XFILL_5__9042_ gnd vdd FILL
XFILL_5__11802_ gnd vdd FILL
XFILL_4__13231_ gnd vdd FILL
X_11168_ _11167_/Y gnd _11477_/B vdd INVX1
XFILL_5__12782_ gnd vdd FILL
XFILL_4__10443_ gnd vdd FILL
XFILL_5__15570_ gnd vdd FILL
XFILL_2__14410_ gnd vdd FILL
XFILL_2__9264_ gnd vdd FILL
XFILL_2__11622_ gnd vdd FILL
XFILL_3__13961_ gnd vdd FILL
XFILL_2__15390_ gnd vdd FILL
XSFILL108840x52050 gnd vdd FILL
XFILL_1__10263_ gnd vdd FILL
XFILL_3_BUFX2_insert570 gnd vdd FILL
XFILL_0__13781_ gnd vdd FILL
X_10119_ _10117_/Y _10106_/A _10119_/C gnd _10203_/D vdd OAI21X1
XFILL_3_BUFX2_insert581 gnd vdd FILL
XFILL_3__15700_ gnd vdd FILL
XFILL_5__14521_ gnd vdd FILL
XFILL_0__10993_ gnd vdd FILL
XFILL_5__11733_ gnd vdd FILL
XFILL_3_BUFX2_insert592 gnd vdd FILL
X_15976_ _15969_/Y _15976_/B _15975_/Y gnd _15984_/B vdd NAND3X1
XFILL_3__12912_ gnd vdd FILL
XFILL_1__12002_ gnd vdd FILL
XSFILL13800x46050 gnd vdd FILL
XFILL_2__8215_ gnd vdd FILL
XFILL_4__13162_ gnd vdd FILL
X_11099_ _12183_/Y _12306_/Y gnd _11099_/Y vdd NAND2X1
XFILL_0__15520_ gnd vdd FILL
XFILL_2__14341_ gnd vdd FILL
XFILL_4__10374_ gnd vdd FILL
XFILL_2__11553_ gnd vdd FILL
XFILL_0__12732_ gnd vdd FILL
XFILL_3__13892_ gnd vdd FILL
XFILL_0__7230_ gnd vdd FILL
XFILL_1__10194_ gnd vdd FILL
XFILL_5__14452_ gnd vdd FILL
XFILL_4__12113_ gnd vdd FILL
X_14927_ _14925_/Y _14927_/B _14924_/Y gnd _14928_/B vdd NAND3X1
XFILL_2__10504_ gnd vdd FILL
XFILL_3__15631_ gnd vdd FILL
XFILL_5__11664_ gnd vdd FILL
XFILL_3__12843_ gnd vdd FILL
XFILL_4__13093_ gnd vdd FILL
XFILL_2__8146_ gnd vdd FILL
XFILL_0__15451_ gnd vdd FILL
XFILL_2__11484_ gnd vdd FILL
XFILL_2__14272_ gnd vdd FILL
XFILL_5__13403_ gnd vdd FILL
XSFILL80120x50050 gnd vdd FILL
XFILL_5__10615_ gnd vdd FILL
XFILL_0__7161_ gnd vdd FILL
X_14858_ _14858_/A _14850_/Y _14858_/C gnd _14859_/A vdd NAND3X1
XFILL_2__16011_ gnd vdd FILL
XFILL_4__12044_ gnd vdd FILL
XFILL_5__14383_ gnd vdd FILL
XFILL_2__13223_ gnd vdd FILL
XFILL_3__15562_ gnd vdd FILL
XFILL_0__14402_ gnd vdd FILL
XFILL_2__10435_ gnd vdd FILL
XFILL_5__11595_ gnd vdd FILL
XFILL_3__12774_ gnd vdd FILL
XFILL_2__8077_ gnd vdd FILL
XFILL_0__11614_ gnd vdd FILL
XFILL_0__15382_ gnd vdd FILL
XFILL_1__13953_ gnd vdd FILL
XFILL_5__13334_ gnd vdd FILL
X_13809_ _7005_/Q gnd _13809_/Y vdd INVX1
XFILL_0__12594_ gnd vdd FILL
XFILL_5__16122_ gnd vdd FILL
XFILL_5__9875_ gnd vdd FILL
XFILL_3__14513_ gnd vdd FILL
XFILL_0__7092_ gnd vdd FILL
XFILL_5__10546_ gnd vdd FILL
XFILL_2__13154_ gnd vdd FILL
XSFILL43880x41050 gnd vdd FILL
XFILL_3__11725_ gnd vdd FILL
X_14789_ _14783_/Y _14789_/B _14789_/C gnd _14789_/Y vdd NAND3X1
XFILL_0__14333_ gnd vdd FILL
XFILL_1__12904_ gnd vdd FILL
XFILL_2__10366_ gnd vdd FILL
XFILL_3__15493_ gnd vdd FILL
XFILL_3__8890_ gnd vdd FILL
XFILL_5__8826_ gnd vdd FILL
XFILL_0__11545_ gnd vdd FILL
XFILL_1__13884_ gnd vdd FILL
XFILL_6_BUFX2_insert96 gnd vdd FILL
XFILL_5__16053_ gnd vdd FILL
XFILL_5__13265_ gnd vdd FILL
XFILL_2__12105_ gnd vdd FILL
XFILL_4__15803_ gnd vdd FILL
XFILL_3__14444_ gnd vdd FILL
XFILL_1__15623_ gnd vdd FILL
XFILL_3__7841_ gnd vdd FILL
XFILL_2__13085_ gnd vdd FILL
XFILL_4__13995_ gnd vdd FILL
XFILL_3__11656_ gnd vdd FILL
XFILL_0__14264_ gnd vdd FILL
XFILL_1__12835_ gnd vdd FILL
XFILL_2__10297_ gnd vdd FILL
XSFILL74200x11050 gnd vdd FILL
XFILL_5__15004_ gnd vdd FILL
XFILL_5__8757_ gnd vdd FILL
X_8410_ _8410_/Q _9306_/CLK _9306_/R vdd _8410_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert109 gnd vdd FILL
XFILL_5__12216_ gnd vdd FILL
XFILL_6__7550_ gnd vdd FILL
XFILL_0__11476_ gnd vdd FILL
XFILL_0__16003_ gnd vdd FILL
XFILL_2__12036_ gnd vdd FILL
X_9390_ _9388_/Y _9372_/B _9389_/Y gnd _9390_/Y vdd OAI21X1
XFILL_4__15734_ gnd vdd FILL
XFILL_0__13215_ gnd vdd FILL
XFILL_3__14375_ gnd vdd FILL
XFILL_1__12766_ gnd vdd FILL
XFILL_0__10427_ gnd vdd FILL
XFILL_5__7708_ gnd vdd FILL
XFILL_1__15554_ gnd vdd FILL
XFILL_3__11587_ gnd vdd FILL
XFILL_2__8979_ gnd vdd FILL
XFILL_0__14195_ gnd vdd FILL
XFILL_0__9802_ gnd vdd FILL
XFILL_0_BUFX2_insert460 gnd vdd FILL
XFILL_0_BUFX2_insert471 gnd vdd FILL
XFILL_3__16114_ gnd vdd FILL
X_8341_ _8372_/B _8853_/B gnd _8341_/Y vdd NAND2X1
XFILL_5__12147_ gnd vdd FILL
XFILL_3__13326_ gnd vdd FILL
XFILL_4__15665_ gnd vdd FILL
XFILL_3__9511_ gnd vdd FILL
XFILL_0_BUFX2_insert482 gnd vdd FILL
XFILL_0_BUFX2_insert493 gnd vdd FILL
XFILL_0__7994_ gnd vdd FILL
XSFILL109400x39050 gnd vdd FILL
XFILL_1__14505_ gnd vdd FILL
XFILL_4__12877_ gnd vdd FILL
XFILL_1__11717_ gnd vdd FILL
XFILL_3__10538_ gnd vdd FILL
XFILL_0__13146_ gnd vdd FILL
XFILL_1__12697_ gnd vdd FILL
XFILL_0__10358_ gnd vdd FILL
XFILL_1__15485_ gnd vdd FILL
XFILL_4_BUFX2_insert809 gnd vdd FILL
XFILL_4__14616_ gnd vdd FILL
XFILL_0__9733_ gnd vdd FILL
XFILL_3__16045_ gnd vdd FILL
XFILL_0__6945_ gnd vdd FILL
XFILL_5__12078_ gnd vdd FILL
XFILL_4__11828_ gnd vdd FILL
X_8272_ _8272_/A gnd _8274_/A vdd INVX1
XFILL_3__13257_ gnd vdd FILL
XFILL112200x78050 gnd vdd FILL
XFILL_4__15596_ gnd vdd FILL
XSFILL38840x30050 gnd vdd FILL
XFILL_1__11648_ gnd vdd FILL
XFILL_1__14436_ gnd vdd FILL
XFILL_6__9151_ gnd vdd FILL
XFILL_2__13987_ gnd vdd FILL
X_7223_ _7223_/A _7181_/B _7222_/Y gnd _7223_/Y vdd OAI21X1
XFILL_5__15906_ gnd vdd FILL
XFILL_0__10289_ gnd vdd FILL
XFILL_5__11029_ gnd vdd FILL
XFILL_0__9664_ gnd vdd FILL
XSFILL64120x63050 gnd vdd FILL
XFILL_4__14547_ gnd vdd FILL
XFILL_3__12208_ gnd vdd FILL
XFILL_2__15726_ gnd vdd FILL
XFILL_0__6876_ gnd vdd FILL
XFILL_4__11759_ gnd vdd FILL
XFILL_6__8102_ gnd vdd FILL
XFILL_0__12028_ gnd vdd FILL
XFILL_1__14367_ gnd vdd FILL
XFILL_3__9373_ gnd vdd FILL
XFILL_1__11579_ gnd vdd FILL
XFILL_0__8615_ gnd vdd FILL
X_7154_ _7114_/A _7902_/CLK _7150_/R vdd _7154_/D gnd vdd DFFSR
XFILL_5__15837_ gnd vdd FILL
XFILL_4__14478_ gnd vdd FILL
XFILL_1__13318_ gnd vdd FILL
XFILL_3__8324_ gnd vdd FILL
XFILL_3__12139_ gnd vdd FILL
XFILL_1__16106_ gnd vdd FILL
XFILL_0__9595_ gnd vdd FILL
XFILL_2__15657_ gnd vdd FILL
XFILL_2__12869_ gnd vdd FILL
XFILL_1__14298_ gnd vdd FILL
XCLKBUF1_insert150 CLKBUF1_insert150/A gnd _9958_/CLK vdd CLKBUF1
XSFILL43960x21050 gnd vdd FILL
XSFILL3560x70050 gnd vdd FILL
XFILL_4__16217_ gnd vdd FILL
XFILL_4__13429_ gnd vdd FILL
XCLKBUF1_insert161 CLKBUF1_insert182/A gnd _7651_/CLK vdd CLKBUF1
XFILL_2__14608_ gnd vdd FILL
X_7085_ _7067_/A _9005_/B gnd _7086_/C vdd NAND2X1
XFILL_5__15768_ gnd vdd FILL
XCLKBUF1_insert172 CLKBUF1_insert193/A gnd _7640_/CLK vdd CLKBUF1
XFILL_1__13249_ gnd vdd FILL
XFILL_3__8255_ gnd vdd FILL
XFILL_1__16037_ gnd vdd FILL
XCLKBUF1_insert183 CLKBUF1_insert150/A gnd _9705_/CLK vdd CLKBUF1
XFILL_2__15588_ gnd vdd FILL
XCLKBUF1_insert194 CLKBUF1_insert187/A gnd _12692_/CLK vdd CLKBUF1
XFILL_0__13979_ gnd vdd FILL
XSFILL28760x82050 gnd vdd FILL
XFILL_5__14719_ gnd vdd FILL
XFILL_4__16148_ gnd vdd FILL
XFILL_3__7206_ gnd vdd FILL
XFILL_0__8477_ gnd vdd FILL
XFILL_5__15699_ gnd vdd FILL
XFILL_2__14539_ gnd vdd FILL
XSFILL44040x30050 gnd vdd FILL
XFILL_0__15718_ gnd vdd FILL
XFILL_3__8186_ gnd vdd FILL
XFILL_6__9984_ gnd vdd FILL
XFILL_0__7428_ gnd vdd FILL
XFILL_4__16079_ gnd vdd FILL
XFILL_3__15829_ gnd vdd FILL
XFILL_5_BUFX2_insert9 gnd vdd FILL
XFILL_0__15649_ gnd vdd FILL
XSFILL33880x73050 gnd vdd FILL
XFILL_2__16209_ gnd vdd FILL
XFILL_0__7359_ gnd vdd FILL
X_7987_ _8006_/B _9267_/B gnd _7988_/C vdd NAND2X1
XFILL_4__7950_ gnd vdd FILL
XFILL_3__7068_ gnd vdd FILL
XFILL111800x51050 gnd vdd FILL
X_6938_ _6938_/A gnd _6940_/A vdd INVX1
X_9726_ _9726_/A _9813_/B _9725_/Y gnd _9816_/D vdd OAI21X1
XFILL_4__6901_ gnd vdd FILL
XFILL_4__7881_ gnd vdd FILL
XFILL_1__9911_ gnd vdd FILL
XFILL_0__9029_ gnd vdd FILL
X_6869_ _6869_/A gnd memoryAddress[31] vdd BUFX2
X_9657_ _9625_/B _9657_/B gnd _9658_/C vdd NAND2X1
XFILL_4__9620_ gnd vdd FILL
XFILL_5_BUFX2_insert610 gnd vdd FILL
X_8608_ _8608_/A gnd _8610_/A vdd INVX1
XFILL_5_BUFX2_insert621 gnd vdd FILL
X_9588_ _9552_/A _9194_/CLK _7914_/R vdd _9588_/D gnd vdd DFFSR
XFILL_4__9551_ gnd vdd FILL
XFILL_5_BUFX2_insert632 gnd vdd FILL
XSFILL3640x50050 gnd vdd FILL
X_10470_ _10406_/A _8038_/CLK _8038_/R vdd _10408_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert643 gnd vdd FILL
XFILL_6__7679_ gnd vdd FILL
XFILL_5_BUFX2_insert654 gnd vdd FILL
X_8539_ _8453_/A _7143_/CLK _7131_/R vdd _8539_/D gnd vdd DFFSR
XFILL_4__8502_ gnd vdd FILL
XFILL_1__9773_ gnd vdd FILL
XFILL_5_BUFX2_insert665 gnd vdd FILL
XFILL_1__6985_ gnd vdd FILL
XFILL_4__9482_ gnd vdd FILL
XFILL_5_BUFX2_insert676 gnd vdd FILL
XFILL_5_BUFX2_insert687 gnd vdd FILL
XFILL_1__8724_ gnd vdd FILL
XFILL_5_BUFX2_insert698 gnd vdd FILL
X_12140_ _12137_/A _12847_/A gnd _12141_/C vdd NAND2X1
XSFILL85000x22050 gnd vdd FILL
XFILL_1__8655_ gnd vdd FILL
XFILL_4__8364_ gnd vdd FILL
X_12071_ _11999_/A _12406_/A _11999_/C gnd _12074_/A vdd NAND3X1
XSFILL33960x53050 gnd vdd FILL
XFILL_2_CLKBUF1_insert202 gnd vdd FILL
XSFILL79160x50 gnd vdd FILL
XFILL_1__7606_ gnd vdd FILL
XFILL_2_CLKBUF1_insert213 gnd vdd FILL
XFILL_2_CLKBUF1_insert224 gnd vdd FILL
XFILL_1__8586_ gnd vdd FILL
XFILL_4__7315_ gnd vdd FILL
X_11022_ _12238_/Y _11030_/A gnd _11026_/A vdd AND2X2
XSFILL79160x9050 gnd vdd FILL
XFILL_4__7246_ gnd vdd FILL
X_15830_ _10671_/A gnd _15830_/Y vdd INVX1
XFILL_2_BUFX2_insert500 gnd vdd FILL
XFILL_2_BUFX2_insert511 gnd vdd FILL
XFILL_1__7468_ gnd vdd FILL
XFILL_4__7177_ gnd vdd FILL
XFILL_2_BUFX2_insert522 gnd vdd FILL
XFILL_2__8000_ gnd vdd FILL
XFILL_2_BUFX2_insert533 gnd vdd FILL
XFILL_1__9207_ gnd vdd FILL
X_15761_ _16301_/A _14294_/Y _15761_/C _15761_/D gnd _15761_/Y vdd OAI22X1
X_12973_ vdd _12973_/B gnd _12974_/C vdd NAND2X1
XFILL_2_BUFX2_insert544 gnd vdd FILL
XSFILL3720x30050 gnd vdd FILL
XFILL_2_BUFX2_insert555 gnd vdd FILL
XFILL_2_BUFX2_insert566 gnd vdd FILL
X_14712_ _9796_/A _14712_/B _14711_/Y gnd _14712_/Y vdd AOI21X1
XSFILL94360x3050 gnd vdd FILL
XFILL_5__7990_ gnd vdd FILL
XFILL_2_BUFX2_insert577 gnd vdd FILL
X_11924_ _11921_/A _12035_/B gnd _11925_/C vdd NAND2X1
X_15692_ _15692_/A _15203_/B _16225_/C _14223_/D gnd _15694_/A vdd OAI22X1
XFILL_2_BUFX2_insert588 gnd vdd FILL
XFILL_1__9138_ gnd vdd FILL
XFILL_2_BUFX2_insert599 gnd vdd FILL
XFILL_5__10400_ gnd vdd FILL
XFILL_5__6941_ gnd vdd FILL
X_14643_ _14642_/Y _14643_/B _14643_/C _14641_/Y gnd _14644_/A vdd OAI22X1
XSFILL69000x35050 gnd vdd FILL
XFILL_5__11380_ gnd vdd FILL
X_11855_ _11700_/A _11855_/B _11629_/A gnd _11855_/Y vdd NAND3X1
XFILL_1__10950_ gnd vdd FILL
XFILL_5__9660_ gnd vdd FILL
XFILL_6_BUFX2_insert1063 gnd vdd FILL
X_10806_ _10831_/B _8630_/B gnd _10806_/Y vdd NAND2X1
XFILL_5__6872_ gnd vdd FILL
X_14574_ _9581_/Q gnd _14574_/Y vdd INVX1
XFILL_2__8902_ gnd vdd FILL
XFILL_3__11510_ gnd vdd FILL
XFILL_2__10151_ gnd vdd FILL
X_11786_ _11377_/Y _11379_/B _11444_/Y gnd _11786_/Y vdd OAI21X1
XBUFX2_insert510 BUFX2_insert570/A gnd _8171_/R vdd BUFX2
XFILL_2__9882_ gnd vdd FILL
XFILL_3__12490_ gnd vdd FILL
XFILL_5__8611_ gnd vdd FILL
XFILL_0__11330_ gnd vdd FILL
XSFILL33240x14050 gnd vdd FILL
XBUFX2_insert521 BUFX2_insert570/A gnd _12795_/R vdd BUFX2
XFILL_1__10881_ gnd vdd FILL
X_16313_ _9205_/Q gnd _16313_/Y vdd INVX1
XBUFX2_insert532 BUFX2_insert518/A gnd _8051_/R vdd BUFX2
XFILL_5__9591_ gnd vdd FILL
XSFILL99480x28050 gnd vdd FILL
X_13525_ _14211_/A _13524_/Y _13574_/C _13525_/D gnd _13525_/Y vdd OAI22X1
XBUFX2_insert543 BUFX2_insert494/A gnd _7914_/R vdd BUFX2
XFILL_5__10262_ gnd vdd FILL
X_10737_ _10737_/Q _9834_/CLK _7793_/R vdd _10697_/Y gnd vdd DFFSR
XFILL_2__8833_ gnd vdd FILL
XFILL_1__12620_ gnd vdd FILL
XFILL_4__13780_ gnd vdd FILL
XFILL_3__11441_ gnd vdd FILL
XSFILL74120x26050 gnd vdd FILL
XFILL_4__10992_ gnd vdd FILL
XBUFX2_insert554 BUFX2_insert524/A gnd _7285_/R vdd BUFX2
XBUFX2_insert565 BUFX2_insert607/A gnd _9454_/R vdd BUFX2
XFILL_5__12001_ gnd vdd FILL
XFILL_0__11261_ gnd vdd FILL
XFILL_4__9749_ gnd vdd FILL
XSFILL84280x70050 gnd vdd FILL
X_16244_ _16244_/A _16244_/B _14597_/C gnd _12911_/B vdd AOI21X1
XBUFX2_insert576 BUFX2_insert496/A gnd _9064_/R vdd BUFX2
XFILL_4__12731_ gnd vdd FILL
X_13456_ _13456_/A _15062_/A _13857_/C _13453_/Y gnd _13456_/Y vdd OAI22X1
XBUFX2_insert587 BUFX2_insert520/A gnd _8047_/R vdd BUFX2
XSFILL58440x80050 gnd vdd FILL
XBUFX2_insert598 BUFX2_insert556/A gnd _7411_/R vdd BUFX2
XFILL_0__13000_ gnd vdd FILL
XFILL_3__14160_ gnd vdd FILL
X_10668_ _10668_/A gnd _10670_/A vdd INVX1
XFILL_5__10193_ gnd vdd FILL
XFILL_2__13910_ gnd vdd FILL
XFILL_2__8764_ gnd vdd FILL
XFILL_3__11372_ gnd vdd FILL
XFILL_2__14890_ gnd vdd FILL
X_12407_ _12407_/A _12407_/B gnd _12408_/C vdd NAND2X1
XFILL_5__8473_ gnd vdd FILL
XFILL_0__11192_ gnd vdd FILL
X_16175_ _7794_/Q _15969_/C _16175_/C gnd _16178_/C vdd AOI21X1
XFILL_3__13111_ gnd vdd FILL
XFILL_4__15450_ gnd vdd FILL
XFILL_4__12662_ gnd vdd FILL
XFILL_2__7715_ gnd vdd FILL
X_13387_ _11881_/A _12809_/Q gnd _13389_/A vdd NAND2X1
XFILL_1__11502_ gnd vdd FILL
X_10599_ _14295_/A _7527_/CLK _8935_/R vdd _10599_/D gnd vdd DFFSR
XFILL_3__10323_ gnd vdd FILL
XFILL_2__13841_ gnd vdd FILL
XFILL_3__14091_ gnd vdd FILL
XSFILL109480x13050 gnd vdd FILL
XFILL_1__15270_ gnd vdd FILL
XFILL_5__7424_ gnd vdd FILL
XFILL_2__8695_ gnd vdd FILL
XFILL_1__12482_ gnd vdd FILL
XFILL_0__10143_ gnd vdd FILL
XFILL_4__14401_ gnd vdd FILL
XSFILL8760x4050 gnd vdd FILL
XFILL_6__10434_ gnd vdd FILL
X_15126_ _15126_/A _15104_/Y _15126_/C gnd _15127_/B vdd NOR3X1
XFILL_4__11613_ gnd vdd FILL
X_12338_ _12338_/A _12338_/B _12338_/C gnd _12338_/Y vdd NAND3X1
XFILL_3__10254_ gnd vdd FILL
XFILL_4__15381_ gnd vdd FILL
XFILL_1__14221_ gnd vdd FILL
XSFILL54120x6050 gnd vdd FILL
XFILL_5__13952_ gnd vdd FILL
XFILL_3__13042_ gnd vdd FILL
XFILL_4__12593_ gnd vdd FILL
XFILL112280x52050 gnd vdd FILL
XFILL_1__11433_ gnd vdd FILL
XSFILL64040x78050 gnd vdd FILL
XFILL_2__13772_ gnd vdd FILL
XFILL_5__7355_ gnd vdd FILL
XSFILL113960x38050 gnd vdd FILL
XFILL_0__14951_ gnd vdd FILL
X_15057_ _15057_/A _15057_/B gnd _15057_/Y vdd NOR2X1
XFILL_5__12903_ gnd vdd FILL
XFILL_4__14332_ gnd vdd FILL
XFILL_2__15511_ gnd vdd FILL
X_12269_ _6883_/A _12249_/B _12269_/C _12802_/Q gnd _12270_/C vdd AOI22X1
XFILL_4__11544_ gnd vdd FILL
XFILL_2__12723_ gnd vdd FILL
XFILL_5__13883_ gnd vdd FILL
XFILL_1__14152_ gnd vdd FILL
XFILL_3__10185_ gnd vdd FILL
XFILL_2__7577_ gnd vdd FILL
XFILL_0__13902_ gnd vdd FILL
XFILL_1__11364_ gnd vdd FILL
X_14008_ _9569_/Q gnd _14008_/Y vdd INVX1
XFILL_0__14882_ gnd vdd FILL
XFILL_0__8400_ gnd vdd FILL
XFILL_5__7286_ gnd vdd FILL
XFILL_5__15622_ gnd vdd FILL
XFILL_6__13084_ gnd vdd FILL
XFILL_0__9380_ gnd vdd FILL
XFILL_4__14263_ gnd vdd FILL
XFILL_5__12834_ gnd vdd FILL
XFILL_1__13103_ gnd vdd FILL
XFILL_1__10315_ gnd vdd FILL
XSFILL43880x36050 gnd vdd FILL
XFILL_4__11475_ gnd vdd FILL
XFILL_2__15442_ gnd vdd FILL
XFILL_2__12654_ gnd vdd FILL
XFILL_0__13833_ gnd vdd FILL
XFILL_3__14993_ gnd vdd FILL
XFILL_5__9025_ gnd vdd FILL
XFILL_1__14083_ gnd vdd FILL
XFILL_4__16002_ gnd vdd FILL
XFILL_1__11295_ gnd vdd FILL
XFILL_0__8331_ gnd vdd FILL
XFILL_4__13214_ gnd vdd FILL
XFILL_5__12765_ gnd vdd FILL
XFILL_5__15553_ gnd vdd FILL
XFILL_4__10426_ gnd vdd FILL
XFILL_4__14194_ gnd vdd FILL
XFILL_1__13034_ gnd vdd FILL
XFILL_2__9247_ gnd vdd FILL
XFILL_2__11605_ gnd vdd FILL
XFILL_3__13944_ gnd vdd FILL
XFILL_2__15373_ gnd vdd FILL
XFILL_1__10246_ gnd vdd FILL
XSFILL18680x12050 gnd vdd FILL
XFILL_2__12585_ gnd vdd FILL
XFILL_0__13764_ gnd vdd FILL
XFILL_0__10976_ gnd vdd FILL
XFILL_5__14504_ gnd vdd FILL
X_7910_ _7910_/Q _8921_/CLK _9049_/R vdd _7848_/Y gnd vdd DFFSR
XFILL_4__13145_ gnd vdd FILL
X_15959_ _15959_/A _15956_/Y gnd _15959_/Y vdd NOR2X1
XFILL_0__8262_ gnd vdd FILL
XFILL_5__11716_ gnd vdd FILL
XFILL_5__12696_ gnd vdd FILL
X_8890_ _8888_/Y _8893_/B _8889_/Y gnd _8940_/D vdd OAI21X1
XFILL_2__14324_ gnd vdd FILL
XFILL_5__15484_ gnd vdd FILL
XFILL_0__12715_ gnd vdd FILL
XFILL_3__13875_ gnd vdd FILL
XSFILL84360x50050 gnd vdd FILL
XFILL_0__15503_ gnd vdd FILL
XFILL_2__11536_ gnd vdd FILL
XFILL_1__10177_ gnd vdd FILL
XFILL_0__7213_ gnd vdd FILL
XFILL_0__13695_ gnd vdd FILL
XFILL_0__8193_ gnd vdd FILL
XSFILL59000x67050 gnd vdd FILL
XFILL_3__15614_ gnd vdd FILL
X_7841_ _7821_/B _7329_/B gnd _7842_/C vdd NAND2X1
XFILL_6__6981_ gnd vdd FILL
XFILL_5__14435_ gnd vdd FILL
XFILL_5__11647_ gnd vdd FILL
XFILL_6__13986_ gnd vdd FILL
XFILL_2__8129_ gnd vdd FILL
XFILL_3__12826_ gnd vdd FILL
XFILL_2__14255_ gnd vdd FILL
XFILL_4__10288_ gnd vdd FILL
XFILL_0__15434_ gnd vdd FILL
XFILL_2__11467_ gnd vdd FILL
XFILL_0__12646_ gnd vdd FILL
XFILL_3__9991_ gnd vdd FILL
XFILL_6__15725_ gnd vdd FILL
XFILL_1__14985_ gnd vdd FILL
XFILL_5__9927_ gnd vdd FILL
XFILL_4__12027_ gnd vdd FILL
X_7772_ _7688_/A _7781_/CLK _8670_/R vdd _7772_/D gnd vdd DFFSR
XFILL111720x66050 gnd vdd FILL
XFILL_3__15545_ gnd vdd FILL
XFILL_5__14366_ gnd vdd FILL
XFILL_5__11578_ gnd vdd FILL
XFILL_3__12757_ gnd vdd FILL
XFILL_2__10418_ gnd vdd FILL
XFILL_0__15365_ gnd vdd FILL
XFILL_2__14186_ gnd vdd FILL
XFILL_2__11398_ gnd vdd FILL
XFILL_1__13936_ gnd vdd FILL
XFILL_0__12577_ gnd vdd FILL
XFILL_5__9858_ gnd vdd FILL
XFILL_5__16105_ gnd vdd FILL
XSFILL38840x25050 gnd vdd FILL
XFILL_5__13317_ gnd vdd FILL
XFILL_0__7075_ gnd vdd FILL
X_9511_ _9533_/B _9895_/B gnd _9512_/C vdd NAND2X1
XFILL_5__10529_ gnd vdd FILL
XFILL112360x32050 gnd vdd FILL
XSFILL23800x50 gnd vdd FILL
XSFILL64120x58050 gnd vdd FILL
XFILL_3__11708_ gnd vdd FILL
XFILL_5__14297_ gnd vdd FILL
XFILL_2__13137_ gnd vdd FILL
XFILL_0__14316_ gnd vdd FILL
XFILL_3__15476_ gnd vdd FILL
XFILL_3__8873_ gnd vdd FILL
XFILL_0__11528_ gnd vdd FILL
XFILL_1__13867_ gnd vdd FILL
XFILL_0__15296_ gnd vdd FILL
XFILL_5__13248_ gnd vdd FILL
XFILL_5__9789_ gnd vdd FILL
XFILL_5__16036_ gnd vdd FILL
X_9442_ _9442_/Q _7010_/CLK _8278_/R vdd _9372_/Y gnd vdd DFFSR
XFILL_6__11819_ gnd vdd FILL
XFILL_6__15587_ gnd vdd FILL
XFILL_3__14427_ gnd vdd FILL
XFILL_3__7824_ gnd vdd FILL
XFILL_4_CLKBUF1_insert190 gnd vdd FILL
XFILL_3__11639_ gnd vdd FILL
XFILL_1__15606_ gnd vdd FILL
XFILL_0__14247_ gnd vdd FILL
XFILL_4__13978_ gnd vdd FILL
XFILL_0__11459_ gnd vdd FILL
XFILL_1__13798_ gnd vdd FILL
XSFILL114920x46050 gnd vdd FILL
XSFILL43960x16050 gnd vdd FILL
XSFILL3560x65050 gnd vdd FILL
XFILL_4__15717_ gnd vdd FILL
X_9373_ _9373_/A gnd _9373_/Y vdd INVX1
XFILL_2__12019_ gnd vdd FILL
XFILL_3__14358_ gnd vdd FILL
XFILL_3__7755_ gnd vdd FILL
XFILL_1__15537_ gnd vdd FILL
XFILL_1__12749_ gnd vdd FILL
XFILL_0__14178_ gnd vdd FILL
XFILL_0_BUFX2_insert290 gnd vdd FILL
X_8324_ _8322_/Y _8333_/B _8324_/C gnd _8410_/D vdd OAI21X1
XFILL_3__13309_ gnd vdd FILL
XSFILL28760x77050 gnd vdd FILL
XFILL_4_BUFX2_insert606 gnd vdd FILL
XFILL_4__15648_ gnd vdd FILL
XFILL_4_BUFX2_insert617 gnd vdd FILL
XFILL_0__7977_ gnd vdd FILL
XFILL_0__13129_ gnd vdd FILL
XFILL_3__14289_ gnd vdd FILL
XFILL_4_BUFX2_insert628 gnd vdd FILL
XFILL_1__15468_ gnd vdd FILL
XFILL_3__7686_ gnd vdd FILL
XFILL_4_BUFX2_insert639 gnd vdd FILL
X_8255_ _8208_/B _8255_/B gnd _8256_/C vdd NAND2X1
XFILL_0__6928_ gnd vdd FILL
XFILL_3__16028_ gnd vdd FILL
XFILL_3__9425_ gnd vdd FILL
XFILL_1__14419_ gnd vdd FILL
XFILL_4__15579_ gnd vdd FILL
XFILL_1__15399_ gnd vdd FILL
X_7206_ _7206_/A gnd _7208_/A vdd INVX1
XFILL_1__8440_ gnd vdd FILL
XFILL_0__9647_ gnd vdd FILL
XSFILL33880x68050 gnd vdd FILL
XFILL_2__15709_ gnd vdd FILL
XFILL_0__6859_ gnd vdd FILL
X_8186_ _8187_/B _9466_/B gnd _8187_/C vdd NAND2X1
XFILL_3__9356_ gnd vdd FILL
XFILL_2_BUFX2_insert50 gnd vdd FILL
XFILL_2_BUFX2_insert61 gnd vdd FILL
XFILL_2_BUFX2_insert72 gnd vdd FILL
XFILL111800x46050 gnd vdd FILL
XFILL_2_BUFX2_insert83 gnd vdd FILL
X_7137_ _7137_/Q _8560_/CLK _9313_/R vdd _7137_/D gnd vdd DFFSR
XSFILL23320x26050 gnd vdd FILL
XFILL_4__7100_ gnd vdd FILL
XSFILL49480x5050 gnd vdd FILL
XFILL_1__8371_ gnd vdd FILL
XFILL_2_BUFX2_insert94 gnd vdd FILL
XFILL_4__8080_ gnd vdd FILL
XFILL_3__9287_ gnd vdd FILL
XFILL112440x12050 gnd vdd FILL
XSFILL64200x38050 gnd vdd FILL
XFILL_1__7322_ gnd vdd FILL
XFILL_0__8529_ gnd vdd FILL
X_7068_ _7066_/Y _7068_/B _7067_/Y gnd _7138_/D vdd OAI21X1
XSFILL38920x6050 gnd vdd FILL
XFILL_4__7031_ gnd vdd FILL
XFILL_3__8238_ gnd vdd FILL
XFILL_1__7253_ gnd vdd FILL
XSFILL3640x45050 gnd vdd FILL
XFILL_1__7184_ gnd vdd FILL
XFILL_1_BUFX2_insert507 gnd vdd FILL
XFILL_1_BUFX2_insert518 gnd vdd FILL
XSFILL28840x57050 gnd vdd FILL
XFILL_4__8982_ gnd vdd FILL
XFILL_1_BUFX2_insert529 gnd vdd FILL
XSFILL94280x33050 gnd vdd FILL
XFILL_4__7933_ gnd vdd FILL
X_11640_ _11639_/Y _11086_/Y _11640_/C gnd _11687_/C vdd OAI21X1
X_9709_ _9709_/Q _7021_/CLK _9062_/R vdd _9709_/D gnd vdd DFFSR
XFILL_4__7864_ gnd vdd FILL
X_11571_ _11571_/A _11563_/C gnd _11572_/C vdd NAND2X1
XFILL_4__9603_ gnd vdd FILL
X_13310_ _13310_/A _13283_/A gnd _13312_/A vdd NOR2X1
X_10522_ _15545_/A gnd _10522_/Y vdd INVX1
XSFILL64120x1050 gnd vdd FILL
XSFILL103720x1050 gnd vdd FILL
X_14290_ _9257_/A _13854_/B _14290_/C _7593_/A gnd _14290_/Y vdd AOI22X1
XFILL_5_BUFX2_insert440 gnd vdd FILL
XFILL_5_BUFX2_insert451 gnd vdd FILL
XFILL_4__9534_ gnd vdd FILL
XSFILL34040x57050 gnd vdd FILL
XFILL_5_BUFX2_insert462 gnd vdd FILL
X_13241_ _13236_/B _13240_/Y gnd _13241_/Y vdd NOR2X1
XFILL_5_BUFX2_insert473 gnd vdd FILL
X_10453_ _10451_/Y _10395_/A _10452_/Y gnd _10485_/D vdd OAI21X1
XSFILL74440x62050 gnd vdd FILL
XFILL_5_BUFX2_insert484 gnd vdd FILL
XFILL_1__9756_ gnd vdd FILL
XFILL_1__6968_ gnd vdd FILL
XFILL_5_BUFX2_insert495 gnd vdd FILL
XSFILL89240x22050 gnd vdd FILL
XFILL_4__9465_ gnd vdd FILL
X_10384_ _10382_/Y _10443_/A _10384_/C gnd _10462_/D vdd OAI21X1
XFILL_2__7500_ gnd vdd FILL
XFILL_1__8707_ gnd vdd FILL
X_13172_ _13172_/A gnd _13174_/A vdd INVX1
XFILL_2__8480_ gnd vdd FILL
XSFILL3720x25050 gnd vdd FILL
XFILL_1__6899_ gnd vdd FILL
XFILL_4__9396_ gnd vdd FILL
X_12123_ _12123_/A _12123_/B _12122_/Y gnd _11013_/B vdd OAI21X1
XFILL_1__8638_ gnd vdd FILL
XFILL_2__7431_ gnd vdd FILL
XSFILL28920x37050 gnd vdd FILL
XFILL_4__8347_ gnd vdd FILL
XSFILL94360x13050 gnd vdd FILL
XFILL_6__10150_ gnd vdd FILL
X_12054_ _12051_/Y _12054_/B _12053_/Y gnd _12054_/Y vdd NAND3X1
XFILL_5__10880_ gnd vdd FILL
XFILL_2__7362_ gnd vdd FILL
XFILL_1__8569_ gnd vdd FILL
XSFILL79160x74050 gnd vdd FILL
XFILL_5__7071_ gnd vdd FILL
X_11005_ _11003_/Y _11015_/D gnd _11005_/Y vdd NAND2X1
XFILL_2__9101_ gnd vdd FILL
XFILL_4__11260_ gnd vdd FILL
XFILL_0__10830_ gnd vdd FILL
XFILL_4__7229_ gnd vdd FILL
XFILL_3__11990_ gnd vdd FILL
XFILL_1__11080_ gnd vdd FILL
XFILL_2__7293_ gnd vdd FILL
X_15813_ _15010_/A _14393_/B _15813_/C _14383_/A gnd _15813_/Y vdd OAI22X1
XSFILL114360x83050 gnd vdd FILL
XFILL_2_BUFX2_insert330 gnd vdd FILL
XFILL_2__9032_ gnd vdd FILL
XFILL_3__10941_ gnd vdd FILL
XFILL_2__12370_ gnd vdd FILL
XFILL_1__10031_ gnd vdd FILL
XFILL_4__11191_ gnd vdd FILL
XFILL_2_BUFX2_insert341 gnd vdd FILL
XFILL_0__10761_ gnd vdd FILL
XFILL_2_BUFX2_insert352 gnd vdd FILL
XFILL_5__11501_ gnd vdd FILL
XSFILL84280x65050 gnd vdd FILL
XSFILL33640x30050 gnd vdd FILL
XFILL_2_BUFX2_insert363 gnd vdd FILL
X_15744_ _7911_/Q _16204_/B _16014_/C _8233_/A gnd _15744_/Y vdd AOI22X1
XFILL_5__12481_ gnd vdd FILL
XFILL_4__10142_ gnd vdd FILL
XFILL_2__11321_ gnd vdd FILL
X_12956_ _12954_/Y vdd _12956_/C gnd _13048_/D vdd OAI21X1
XFILL_2_BUFX2_insert374 gnd vdd FILL
XFILL_2_BUFX2_insert385 gnd vdd FILL
XFILL_3__13660_ gnd vdd FILL
XFILL_0__12500_ gnd vdd FILL
XFILL_3__10872_ gnd vdd FILL
XFILL_2_BUFX2_insert396 gnd vdd FILL
XFILL_0__13480_ gnd vdd FILL
XFILL_5__14220_ gnd vdd FILL
XFILL_5__7973_ gnd vdd FILL
X_11907_ _11907_/A _11934_/B _11907_/C gnd _6844_/A vdd OAI21X1
XFILL_0__10692_ gnd vdd FILL
XFILL_5__11432_ gnd vdd FILL
X_15675_ _15675_/A _15672_/Y gnd _15675_/Y vdd NOR2X1
XFILL_3__12611_ gnd vdd FILL
XFILL_6__13771_ gnd vdd FILL
XSFILL59080x41050 gnd vdd FILL
X_12887_ vdd _12887_/B gnd _12888_/C vdd NAND2X1
XFILL_2__14040_ gnd vdd FILL
XFILL_4__14950_ gnd vdd FILL
XFILL_2__11252_ gnd vdd FILL
XFILL_0__12431_ gnd vdd FILL
XFILL_3__13591_ gnd vdd FILL
XFILL_5__6924_ gnd vdd FILL
XFILL_1__11982_ gnd vdd FILL
XFILL_1__14770_ gnd vdd FILL
X_14626_ _14626_/A _7406_/Q _7918_/Q _13865_/B gnd _14630_/A vdd AOI22X1
XFILL_6__12722_ gnd vdd FILL
XFILL_5__14151_ gnd vdd FILL
XFILL_3__15330_ gnd vdd FILL
XFILL_4__13901_ gnd vdd FILL
XFILL_5__11363_ gnd vdd FILL
X_11838_ _11837_/Y _11835_/A gnd _11838_/Y vdd NAND2X1
XFILL_2__9934_ gnd vdd FILL
XFILL_4__14881_ gnd vdd FILL
XFILL_1__10933_ gnd vdd FILL
XFILL112280x47050 gnd vdd FILL
XFILL_2__11183_ gnd vdd FILL
XFILL_0__15150_ gnd vdd FILL
XFILL_1__13721_ gnd vdd FILL
XFILL_0__12362_ gnd vdd FILL
XFILL_5__13102_ gnd vdd FILL
XFILL_5__9643_ gnd vdd FILL
XFILL_5__10314_ gnd vdd FILL
XFILL_5__6855_ gnd vdd FILL
X_14557_ _8379_/A _13848_/B _14557_/C _8301_/Q gnd _14559_/A vdd AOI22X1
XFILL_5__14082_ gnd vdd FILL
XFILL_4__13832_ gnd vdd FILL
XFILL_2__10134_ gnd vdd FILL
XFILL_5__11294_ gnd vdd FILL
XFILL_3__15261_ gnd vdd FILL
XFILL_0__14101_ gnd vdd FILL
X_11769_ _11769_/A _11020_/Y _11766_/Y gnd _11770_/B vdd OAI21X1
XFILL_2__9865_ gnd vdd FILL
XBUFX2_insert340 _12811_/Q gnd _13372_/A vdd BUFX2
XFILL_3__12473_ gnd vdd FILL
XFILL_0__11313_ gnd vdd FILL
XSFILL109320x72050 gnd vdd FILL
XFILL_1__13652_ gnd vdd FILL
XFILL_2__15991_ gnd vdd FILL
XFILL_0__15081_ gnd vdd FILL
XBUFX2_insert351 _10927_/Y gnd _12227_/A vdd BUFX2
XFILL_0__12293_ gnd vdd FILL
XFILL_6__11604_ gnd vdd FILL
XBUFX2_insert362 _11352_/Y gnd _11751_/C vdd BUFX2
X_13508_ _9849_/A gnd _13510_/D vdd INVX1
XFILL_5__13033_ gnd vdd FILL
XFILL_6__15372_ gnd vdd FILL
XFILL_3__14212_ gnd vdd FILL
XFILL_5__10245_ gnd vdd FILL
XBUFX2_insert373 _13338_/Y gnd _9533_/B vdd BUFX2
X_14488_ _8171_/Q gnd _14488_/Y vdd INVX1
XFILL_4__13763_ gnd vdd FILL
XFILL_0__8880_ gnd vdd FILL
XFILL_3__11424_ gnd vdd FILL
XFILL_1__12603_ gnd vdd FILL
XFILL_4__10975_ gnd vdd FILL
XFILL_3__15192_ gnd vdd FILL
XSFILL79240x54050 gnd vdd FILL
XFILL_0__14032_ gnd vdd FILL
XBUFX2_insert384 _13331_/Y gnd _9112_/A vdd BUFX2
XFILL_2__14942_ gnd vdd FILL
XFILL_2__10065_ gnd vdd FILL
XFILL_5__8525_ gnd vdd FILL
XFILL_1__16371_ gnd vdd FILL
XFILL_2__9796_ gnd vdd FILL
XFILL_1__13583_ gnd vdd FILL
XFILL_0__11244_ gnd vdd FILL
XBUFX2_insert395 _13293_/Y gnd _7598_/B vdd BUFX2
X_16227_ _7629_/A gnd _16227_/Y vdd INVX1
XFILL_1__10795_ gnd vdd FILL
XFILL_4__12714_ gnd vdd FILL
XFILL_0__7831_ gnd vdd FILL
X_13439_ _13865_/C _7766_/Q _8278_/Q _13592_/A gnd _13439_/Y vdd AOI22X1
XFILL_4__15502_ gnd vdd FILL
XFILL_5__10176_ gnd vdd FILL
XFILL_3__14143_ gnd vdd FILL
XFILL_1__15322_ gnd vdd FILL
XFILL_2__8747_ gnd vdd FILL
XFILL_4__13694_ gnd vdd FILL
XFILL_3__11355_ gnd vdd FILL
XFILL_2__14873_ gnd vdd FILL
XFILL_1__12534_ gnd vdd FILL
XSFILL83720x79050 gnd vdd FILL
XSFILL114440x63050 gnd vdd FILL
XFILL_5__8456_ gnd vdd FILL
XFILL_0__11175_ gnd vdd FILL
X_16158_ _16157_/Y _15581_/C _16314_/A _14756_/Y gnd _16161_/A vdd OAI22X1
XFILL_4__12645_ gnd vdd FILL
XFILL_3__10306_ gnd vdd FILL
XFILL_4__15433_ gnd vdd FILL
XFILL_6__11466_ gnd vdd FILL
XFILL_0__7762_ gnd vdd FILL
XFILL_2__13824_ gnd vdd FILL
XFILL_5__14984_ gnd vdd FILL
XFILL_3__14074_ gnd vdd FILL
XFILL_0__10126_ gnd vdd FILL
XFILL_1__15253_ gnd vdd FILL
XFILL_1__12465_ gnd vdd FILL
XSFILL84360x45050 gnd vdd FILL
XFILL_3__7471_ gnd vdd FILL
XFILL_3__11286_ gnd vdd FILL
XFILL_0__9501_ gnd vdd FILL
X_15109_ _15108_/Y _15109_/B gnd _15113_/A vdd NOR2X1
XFILL_0__15983_ gnd vdd FILL
X_8040_ _7980_/A _8680_/CLK _8034_/R vdd _8040_/D gnd vdd DFFSR
XFILL_5__8387_ gnd vdd FILL
XSFILL48920x1050 gnd vdd FILL
XFILL_4__15364_ gnd vdd FILL
XFILL_3__13025_ gnd vdd FILL
X_16089_ _14719_/Y _16089_/B gnd _16093_/A vdd NOR2X1
XFILL_5__13935_ gnd vdd FILL
XFILL_3__9210_ gnd vdd FILL
XFILL_4__12576_ gnd vdd FILL
XFILL_2__7629_ gnd vdd FILL
XFILL_0__7693_ gnd vdd FILL
XFILL_1__14204_ gnd vdd FILL
XFILL_3__10237_ gnd vdd FILL
XFILL_1__11416_ gnd vdd FILL
XFILL_1__15184_ gnd vdd FILL
XFILL_2__13755_ gnd vdd FILL
XFILL_2__10967_ gnd vdd FILL
XSFILL99400x67050 gnd vdd FILL
XFILL_1__12396_ gnd vdd FILL
XFILL_5__7338_ gnd vdd FILL
XFILL_0__14934_ gnd vdd FILL
XFILL_0__10057_ gnd vdd FILL
XSFILL59160x21050 gnd vdd FILL
XFILL_6__13136_ gnd vdd FILL
XFILL_4__14315_ gnd vdd FILL
XFILL_4__11527_ gnd vdd FILL
XFILL_3__9141_ gnd vdd FILL
XFILL_2__12706_ gnd vdd FILL
XFILL_5__13866_ gnd vdd FILL
XFILL_4__15295_ gnd vdd FILL
XFILL_1__14135_ gnd vdd FILL
XFILL_3__10168_ gnd vdd FILL
XFILL_1__11347_ gnd vdd FILL
XFILL_2__13686_ gnd vdd FILL
XFILL_2__10898_ gnd vdd FILL
XFILL_0__14865_ gnd vdd FILL
XSFILL59960x6050 gnd vdd FILL
XFILL_5__15605_ gnd vdd FILL
XFILL_4__14246_ gnd vdd FILL
XFILL_6__10279_ gnd vdd FILL
XFILL112360x27050 gnd vdd FILL
XFILL_0__9363_ gnd vdd FILL
XFILL_4__11458_ gnd vdd FILL
XFILL_2__15425_ gnd vdd FILL
XFILL_2__12637_ gnd vdd FILL
XFILL_5__13797_ gnd vdd FILL
XFILL_1__14066_ gnd vdd FILL
XFILL_5__9008_ gnd vdd FILL
XFILL_3__14976_ gnd vdd FILL
X_9991_ _9989_/Y _9979_/B _9990_/Y gnd _9991_/Y vdd OAI21X1
XFILL_0__13816_ gnd vdd FILL
XFILL_1__11278_ gnd vdd FILL
XFILL_0__14796_ gnd vdd FILL
XFILL_0__8314_ gnd vdd FILL
XFILL_5__15536_ gnd vdd FILL
XFILL_4__10409_ gnd vdd FILL
X_8942_ _8894_/A _8942_/CLK _8942_/R vdd _8942_/D gnd vdd DFFSR
XFILL_5__12748_ gnd vdd FILL
XFILL_0__9294_ gnd vdd FILL
XFILL_4__14177_ gnd vdd FILL
XFILL_1__13017_ gnd vdd FILL
XFILL_3__13927_ gnd vdd FILL
XFILL_2__15356_ gnd vdd FILL
XFILL_4__11389_ gnd vdd FILL
XFILL_2__12568_ gnd vdd FILL
XFILL_0__10959_ gnd vdd FILL
XFILL_0__13747_ gnd vdd FILL
XSFILL113640x15050 gnd vdd FILL
XSFILL49080x73050 gnd vdd FILL
XFILL_0__8245_ gnd vdd FILL
XFILL_4__13128_ gnd vdd FILL
XSFILL79320x34050 gnd vdd FILL
XFILL_2__14307_ gnd vdd FILL
XFILL_5__15467_ gnd vdd FILL
XFILL_3__13858_ gnd vdd FILL
X_8873_ _8873_/A gnd _8875_/A vdd INVX1
XFILL_2__11519_ gnd vdd FILL
XFILL_2__15287_ gnd vdd FILL
XFILL_0__13678_ gnd vdd FILL
XFILL_2__12499_ gnd vdd FILL
XFILL_5__14418_ gnd vdd FILL
X_7824_ _7822_/Y _7824_/B _7824_/C gnd _7824_/Y vdd OAI21X1
XSFILL109560x7050 gnd vdd FILL
XFILL_5__15398_ gnd vdd FILL
XFILL_2__14238_ gnd vdd FILL
XSFILL114520x43050 gnd vdd FILL
XFILL_0__12629_ gnd vdd FILL
XFILL_3__9974_ gnd vdd FILL
XFILL_3__13789_ gnd vdd FILL
XFILL_0__15417_ gnd vdd FILL
XFILL_1__14968_ gnd vdd FILL
XFILL_0__16397_ gnd vdd FILL
XFILL_3__15528_ gnd vdd FILL
XFILL_5__14349_ gnd vdd FILL
X_7755_ _7690_/B _7883_/B gnd _7756_/C vdd NAND2X1
XFILL_2__14169_ gnd vdd FILL
XFILL_1__13919_ gnd vdd FILL
XFILL_0__15348_ gnd vdd FILL
XFILL_6__15639_ gnd vdd FILL
XFILL_0__7058_ gnd vdd FILL
XFILL_1__14899_ gnd vdd FILL
XFILL_1__7940_ gnd vdd FILL
XFILL_3__15459_ gnd vdd FILL
X_7686_ _7723_/B _8582_/B gnd _7687_/C vdd NAND2X1
XFILL_3__8856_ gnd vdd FILL
XFILL_0__15279_ gnd vdd FILL
XFILL_5__16019_ gnd vdd FILL
X_9425_ _9425_/A _8529_/B gnd _9426_/C vdd NAND2X1
XFILL_1__7871_ gnd vdd FILL
XFILL_3__7807_ gnd vdd FILL
XFILL_4__7580_ gnd vdd FILL
XFILL_3__8787_ gnd vdd FILL
XFILL_1__9610_ gnd vdd FILL
X_9356_ _9356_/A _7564_/B gnd _9357_/C vdd NAND2X1
XFILL_4_BUFX2_insert403 gnd vdd FILL
XSFILL23720x42050 gnd vdd FILL
XFILL_3__7738_ gnd vdd FILL
XFILL_4_BUFX2_insert414 gnd vdd FILL
XFILL_4_BUFX2_insert425 gnd vdd FILL
X_8307_ _8269_/A _7661_/CLK _8819_/R vdd _8307_/D gnd vdd DFFSR
XFILL_1__9541_ gnd vdd FILL
XFILL_4_BUFX2_insert436 gnd vdd FILL
X_9287_ _9329_/Q gnd _9287_/Y vdd INVX1
XFILL_4__9250_ gnd vdd FILL
XFILL_4_BUFX2_insert447 gnd vdd FILL
XFILL_4_BUFX2_insert458 gnd vdd FILL
XSFILL49160x53050 gnd vdd FILL
XFILL_4_BUFX2_insert469 gnd vdd FILL
X_8238_ _8238_/A _8237_/A _8238_/C gnd _8238_/Y vdd OAI21X1
XFILL_6__7378_ gnd vdd FILL
XFILL_1__9472_ gnd vdd FILL
XFILL_3__9408_ gnd vdd FILL
XFILL_4__8201_ gnd vdd FILL
XSFILL94280x28050 gnd vdd FILL
XSFILL114600x23050 gnd vdd FILL
X_8169_ _8169_/Q _8169_/CLK _7408_/R vdd _8169_/D gnd vdd DFFSR
XFILL_4__8132_ gnd vdd FILL
XFILL_3__9339_ gnd vdd FILL
XFILL_1__8354_ gnd vdd FILL
XFILL_4__8063_ gnd vdd FILL
XFILL_1__7305_ gnd vdd FILL
XFILL_3_CLKBUF1_insert116 gnd vdd FILL
XFILL_3_CLKBUF1_insert127 gnd vdd FILL
XFILL_5_CLKBUF1_insert1076 gnd vdd FILL
XFILL_3_CLKBUF1_insert138 gnd vdd FILL
X_12810_ _11881_/A _12667_/CLK _12689_/R vdd _12810_/D gnd vdd DFFSR
XFILL_3_CLKBUF1_insert149 gnd vdd FILL
X_13790_ _10333_/Q gnd _13792_/A vdd INVX1
XFILL_1__7236_ gnd vdd FILL
XSFILL104520x75050 gnd vdd FILL
XFILL_1_BUFX2_insert304 gnd vdd FILL
XSFILL8760x73050 gnd vdd FILL
X_12741_ _12718_/B memoryOutData[15] gnd _12742_/C vdd NAND2X1
XFILL_1_BUFX2_insert315 gnd vdd FILL
XFILL_1_BUFX2_insert326 gnd vdd FILL
XSFILL23800x22050 gnd vdd FILL
XFILL_1__7167_ gnd vdd FILL
XSFILL59080x8050 gnd vdd FILL
XSFILL89240x17050 gnd vdd FILL
XFILL_1_BUFX2_insert337 gnd vdd FILL
XFILL_1_BUFX2_insert348 gnd vdd FILL
XFILL_4__8965_ gnd vdd FILL
X_15460_ _15459_/Y _15656_/B _15656_/C gnd _15462_/B vdd NOR3X1
XFILL_1_BUFX2_insert359 gnd vdd FILL
X_12672_ _12594_/A _8171_/CLK _8171_/R vdd _12672_/D gnd vdd DFFSR
XFILL_1__7098_ gnd vdd FILL
XFILL_2__7980_ gnd vdd FILL
X_14411_ _14411_/A _14411_/B gnd _14412_/C vdd NOR2X1
XFILL_4__8896_ gnd vdd FILL
X_11623_ _11623_/A _11623_/B _11138_/Y gnd _11624_/C vdd OAI21X1
X_15391_ _10846_/Q gnd _15391_/Y vdd INVX1
XFILL_2__6931_ gnd vdd FILL
XFILL_4__7847_ gnd vdd FILL
X_14342_ _14341_/Y _14342_/B gnd _14343_/C vdd NOR2X1
XSFILL113880x2050 gnd vdd FILL
XSFILL74280x2050 gnd vdd FILL
X_11554_ _11764_/A _11553_/B _11111_/Y _11495_/C gnd _11554_/Y vdd AOI22X1
XFILL_2__9650_ gnd vdd FILL
XSFILL13720x74050 gnd vdd FILL
XFILL_2__6862_ gnd vdd FILL
XSFILL79160x69050 gnd vdd FILL
X_10505_ _10505_/A _9737_/B gnd _10506_/C vdd NAND2X1
XFILL_5__10030_ gnd vdd FILL
XFILL_2__8601_ gnd vdd FILL
X_14273_ _7337_/A _14353_/A _14273_/C _8551_/Q gnd _14275_/A vdd AOI22X1
XFILL_1__9808_ gnd vdd FILL
XFILL_5_BUFX2_insert270 gnd vdd FILL
XFILL_4__10760_ gnd vdd FILL
X_11485_ _11485_/A _11483_/Y gnd _11485_/Y vdd NOR2X1
XFILL_5_BUFX2_insert281 gnd vdd FILL
XFILL_5__8310_ gnd vdd FILL
XFILL_4__9517_ gnd vdd FILL
XFILL_5_BUFX2_insert292 gnd vdd FILL
X_16012_ _16010_/Y _16012_/B _16009_/Y gnd _16012_/Y vdd NAND3X1
XFILL_1__10580_ gnd vdd FILL
X_13224_ _13289_/B _13302_/C gnd _13359_/A vdd NAND2X1
XFILL_5__9290_ gnd vdd FILL
X_10436_ _16105_/A gnd _10438_/A vdd INVX1
XFILL_1__9739_ gnd vdd FILL
XFILL_2__8532_ gnd vdd FILL
XFILL_3__11140_ gnd vdd FILL
XSFILL29400x62050 gnd vdd FILL
XFILL_4__10691_ gnd vdd FILL
XFILL_2__11870_ gnd vdd FILL
XFILL_5__8241_ gnd vdd FILL
XFILL_6__11251_ gnd vdd FILL
XFILL_4__12430_ gnd vdd FILL
X_13155_ _13155_/A _13155_/B gnd _13156_/C vdd NAND2X1
X_10367_ _10457_/Q gnd _10367_/Y vdd INVX1
XFILL_4_BUFX2_insert970 gnd vdd FILL
XFILL_2__8463_ gnd vdd FILL
XFILL_5__11981_ gnd vdd FILL
XFILL_1__12250_ gnd vdd FILL
XFILL_2__10821_ gnd vdd FILL
XFILL_4_BUFX2_insert981 gnd vdd FILL
XFILL_3__11071_ gnd vdd FILL
XSFILL44280x76050 gnd vdd FILL
XFILL_4__9379_ gnd vdd FILL
XFILL_4_BUFX2_insert992 gnd vdd FILL
X_12106_ _12103_/Y _12106_/B _12105_/Y gnd _13167_/B vdd NAND3X1
XFILL_0__12980_ gnd vdd FILL
XFILL_5__13720_ gnd vdd FILL
XFILL_5__10932_ gnd vdd FILL
XFILL_3__10022_ gnd vdd FILL
XFILL_4__12361_ gnd vdd FILL
XFILL_2__7414_ gnd vdd FILL
X_13086_ _13134_/A _13086_/B gnd _13087_/C vdd NAND2X1
X_10298_ _10298_/A _10280_/B _10297_/Y gnd _10298_/Y vdd OAI21X1
XSFILL59080x36050 gnd vdd FILL
XFILL_1__11201_ gnd vdd FILL
XSFILL104520x50 gnd vdd FILL
XFILL_2__13540_ gnd vdd FILL
XFILL_2__10752_ gnd vdd FILL
XFILL_2__8394_ gnd vdd FILL
XFILL_0__11931_ gnd vdd FILL
XFILL_1__12181_ gnd vdd FILL
XFILL_5__7123_ gnd vdd FILL
XSFILL99480x41050 gnd vdd FILL
XFILL_4__14100_ gnd vdd FILL
X_12037_ _12476_/B _12025_/B _12025_/C gnd gnd _12037_/Y vdd AOI22X1
XFILL_4__11312_ gnd vdd FILL
XFILL_5__13651_ gnd vdd FILL
XFILL_3__14830_ gnd vdd FILL
XFILL_4__15080_ gnd vdd FILL
XFILL_2__7345_ gnd vdd FILL
XFILL_4__12292_ gnd vdd FILL
XFILL_1__11132_ gnd vdd FILL
XFILL_2__13471_ gnd vdd FILL
XFILL_0__14650_ gnd vdd FILL
XFILL_2__10683_ gnd vdd FILL
XFILL_5__7054_ gnd vdd FILL
XFILL_0__11862_ gnd vdd FILL
XFILL_5__12602_ gnd vdd FILL
XFILL_4__14031_ gnd vdd FILL
XSFILL109880x24050 gnd vdd FILL
XFILL_2__15210_ gnd vdd FILL
XFILL_5__16370_ gnd vdd FILL
XFILL_4__11243_ gnd vdd FILL
XFILL_2__12422_ gnd vdd FILL
XSFILL53800x38050 gnd vdd FILL
XFILL_5__13582_ gnd vdd FILL
XFILL_3__14761_ gnd vdd FILL
XFILL_5__10794_ gnd vdd FILL
XFILL_0__10813_ gnd vdd FILL
XFILL_0__13601_ gnd vdd FILL
XFILL_3__11973_ gnd vdd FILL
XFILL_2__16190_ gnd vdd FILL
XFILL_1__15940_ gnd vdd FILL
XFILL_1__11063_ gnd vdd FILL
XFILL_0__14581_ gnd vdd FILL
XFILL_5__15321_ gnd vdd FILL
XFILL_0__11793_ gnd vdd FILL
XFILL_2__9015_ gnd vdd FILL
XSFILL13800x54050 gnd vdd FILL
XFILL_5__12533_ gnd vdd FILL
XFILL_3__13712_ gnd vdd FILL
XFILL_3__10924_ gnd vdd FILL
X_13988_ _8343_/A _13647_/B _14145_/D _7575_/A gnd _13988_/Y vdd AOI22X1
XFILL_1__10014_ gnd vdd FILL
XFILL_2__15141_ gnd vdd FILL
XFILL_4__11174_ gnd vdd FILL
XFILL_2__12353_ gnd vdd FILL
XFILL_0__16320_ gnd vdd FILL
XFILL_3__14692_ gnd vdd FILL
XFILL_0__13532_ gnd vdd FILL
XFILL_0__10744_ gnd vdd FILL
XFILL_1__15871_ gnd vdd FILL
X_15727_ _8550_/Q gnd _15728_/B vdd INVX1
XFILL_4__10125_ gnd vdd FILL
XFILL_5__15252_ gnd vdd FILL
XFILL_5__12464_ gnd vdd FILL
X_12939_ _12176_/B _8180_/CLK _8937_/R vdd _12939_/D gnd vdd DFFSR
XFILL_3__13643_ gnd vdd FILL
XFILL_2__11304_ gnd vdd FILL
XFILL_4__15982_ gnd vdd FILL
XFILL_1__14822_ gnd vdd FILL
XFILL_2__15072_ gnd vdd FILL
XFILL_0__13463_ gnd vdd FILL
XFILL_2__12284_ gnd vdd FILL
XFILL_0__16251_ gnd vdd FILL
XFILL_5__14203_ gnd vdd FILL
XFILL_5__7956_ gnd vdd FILL
XFILL_0__10675_ gnd vdd FILL
XFILL_5__11415_ gnd vdd FILL
X_15658_ _15658_/A _15656_/Y _15658_/C gnd _15658_/Y vdd NOR3X1
XFILL_6__10966_ gnd vdd FILL
XFILL_5__15183_ gnd vdd FILL
XFILL_1_BUFX2_insert860 gnd vdd FILL
XFILL_2__14023_ gnd vdd FILL
XFILL_5__12395_ gnd vdd FILL
XFILL_3__16362_ gnd vdd FILL
XFILL_4__10056_ gnd vdd FILL
XFILL_4__14933_ gnd vdd FILL
XFILL_0__12414_ gnd vdd FILL
XFILL_0__15202_ gnd vdd FILL
XFILL_1_BUFX2_insert871 gnd vdd FILL
XFILL_3__13574_ gnd vdd FILL
XFILL_2__11235_ gnd vdd FILL
XFILL_3__6971_ gnd vdd FILL
XFILL_0__16182_ gnd vdd FILL
XFILL_3__10786_ gnd vdd FILL
XFILL_1__14753_ gnd vdd FILL
XFILL_5__6907_ gnd vdd FILL
X_14609_ _7230_/A _13619_/B _14572_/C _10862_/Q gnd _14617_/B vdd AOI22X1
XFILL_1__11965_ gnd vdd FILL
XFILL_0__13394_ gnd vdd FILL
XFILL_1_BUFX2_insert882 gnd vdd FILL
XFILL_5__7887_ gnd vdd FILL
XFILL_1_BUFX2_insert893 gnd vdd FILL
XFILL_3__15313_ gnd vdd FILL
XFILL_5__14134_ gnd vdd FILL
X_7540_ _7504_/A _8297_/CLK _7796_/R vdd _7540_/D gnd vdd DFFSR
XFILL_5__11346_ gnd vdd FILL
XFILL_3__12525_ gnd vdd FILL
XFILL_3__8710_ gnd vdd FILL
XFILL_0__9981_ gnd vdd FILL
X_15589_ _15760_/A _15589_/B _15589_/C gnd _15593_/A vdd OAI21X1
XFILL_2__9917_ gnd vdd FILL
XFILL_4__14864_ gnd vdd FILL
XFILL_3__16293_ gnd vdd FILL
XFILL_0__15133_ gnd vdd FILL
XFILL_1__13704_ gnd vdd FILL
XFILL_2__11166_ gnd vdd FILL
XFILL_1__10916_ gnd vdd FILL
XFILL_0__12345_ gnd vdd FILL
XFILL_5__6838_ gnd vdd FILL
XFILL_5__9626_ gnd vdd FILL
XFILL_1__14684_ gnd vdd FILL
XFILL_6__15424_ gnd vdd FILL
XSFILL59160x16050 gnd vdd FILL
XFILL_1__11896_ gnd vdd FILL
XFILL_5__14065_ gnd vdd FILL
XFILL_4__13815_ gnd vdd FILL
XFILL_3__15244_ gnd vdd FILL
X_7471_ _7471_/A gnd _7473_/A vdd INVX1
XFILL_2__10117_ gnd vdd FILL
XFILL_5__11277_ gnd vdd FILL
XSFILL58920x71050 gnd vdd FILL
XFILL_2__9848_ gnd vdd FILL
XFILL_3__12456_ gnd vdd FILL
XFILL_3__8641_ gnd vdd FILL
XFILL_1__13635_ gnd vdd FILL
XFILL_2__15974_ gnd vdd FILL
XFILL_4__14795_ gnd vdd FILL
XFILL_0__15064_ gnd vdd FILL
XFILL_2__11097_ gnd vdd FILL
XFILL_5__13016_ gnd vdd FILL
XFILL_5__9557_ gnd vdd FILL
XFILL_0__12276_ gnd vdd FILL
X_9210_ _9238_/B _9466_/B gnd _9210_/Y vdd NAND2X1
XFILL_3__11407_ gnd vdd FILL
XFILL_0__8863_ gnd vdd FILL
XFILL_4__10958_ gnd vdd FILL
XFILL_3__15175_ gnd vdd FILL
XFILL_2__10048_ gnd vdd FILL
XFILL_4__13746_ gnd vdd FILL
XFILL_0__14015_ gnd vdd FILL
XFILL_2__14925_ gnd vdd FILL
XFILL_5__8508_ gnd vdd FILL
XFILL_3__12387_ gnd vdd FILL
XFILL_1__16354_ gnd vdd FILL
XFILL_3__8572_ gnd vdd FILL
XFILL_0__11227_ gnd vdd FILL
XFILL_2__9779_ gnd vdd FILL
XFILL_1__10778_ gnd vdd FILL
XFILL_1__13566_ gnd vdd FILL
X_9141_ _9195_/Q gnd _9141_/Y vdd INVX1
XFILL_5__9488_ gnd vdd FILL
XFILL_0__7814_ gnd vdd FILL
XFILL_6__11518_ gnd vdd FILL
XFILL_3__14126_ gnd vdd FILL
XFILL_5__10159_ gnd vdd FILL
XFILL_6__15286_ gnd vdd FILL
XFILL_1__15305_ gnd vdd FILL
XFILL_4__13677_ gnd vdd FILL
XSFILL109400x47050 gnd vdd FILL
XFILL_3__11338_ gnd vdd FILL
XFILL_2__14856_ gnd vdd FILL
XFILL_1__12517_ gnd vdd FILL
XFILL_4__10889_ gnd vdd FILL
XFILL_5__8439_ gnd vdd FILL
XFILL_1__16285_ gnd vdd FILL
XFILL_0__11158_ gnd vdd FILL
XFILL_6__14237_ gnd vdd FILL
XFILL_1__13497_ gnd vdd FILL
XFILL_4__12628_ gnd vdd FILL
X_9072_ _9028_/A _7532_/CLK _8816_/R vdd _9072_/D gnd vdd DFFSR
XSFILL79320x29050 gnd vdd FILL
XFILL_0__7745_ gnd vdd FILL
XFILL_4__15416_ gnd vdd FILL
XFILL_2__13807_ gnd vdd FILL
XFILL_3__14057_ gnd vdd FILL
XFILL_5__14967_ gnd vdd FILL
XSFILL63880x9050 gnd vdd FILL
XFILL_1__15236_ gnd vdd FILL
XFILL_3__7454_ gnd vdd FILL
XFILL_4__16396_ gnd vdd FILL
XFILL_0__10109_ gnd vdd FILL
XFILL_3__11269_ gnd vdd FILL
XFILL_1__12448_ gnd vdd FILL
XFILL_2__14787_ gnd vdd FILL
XFILL_2__11999_ gnd vdd FILL
XFILL_0__15966_ gnd vdd FILL
XFILL_0__11089_ gnd vdd FILL
X_8023_ _8023_/Q _8551_/CLK _9959_/R vdd _8023_/D gnd vdd DFFSR
XSFILL64120x71050 gnd vdd FILL
XFILL_3__13008_ gnd vdd FILL
XFILL_5__13918_ gnd vdd FILL
XFILL_4__15347_ gnd vdd FILL
XFILL_0__7676_ gnd vdd FILL
XFILL_2__13738_ gnd vdd FILL
XFILL_5__14898_ gnd vdd FILL
XFILL_1__12379_ gnd vdd FILL
XFILL_1__15167_ gnd vdd FILL
XFILL_0__14917_ gnd vdd FILL
XSFILL3160x57050 gnd vdd FILL
XFILL_0__9415_ gnd vdd FILL
XFILL_6__7094_ gnd vdd FILL
XFILL_0__15897_ gnd vdd FILL
XFILL_5__13849_ gnd vdd FILL
XFILL_3__9124_ gnd vdd FILL
XFILL_6__14099_ gnd vdd FILL
XFILL_4__15278_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1082 gnd vdd FILL
XFILL_1__14118_ gnd vdd FILL
XFILL_2__13669_ gnd vdd FILL
XFILL_0__14848_ gnd vdd FILL
XFILL_1__15098_ gnd vdd FILL
XFILL_4__14229_ gnd vdd FILL
XFILL_0__9346_ gnd vdd FILL
XFILL_2__15408_ gnd vdd FILL
X_9974_ _9974_/A gnd _9974_/Y vdd INVX1
XSFILL69080x3050 gnd vdd FILL
XFILL_2__16388_ gnd vdd FILL
XFILL_1__14049_ gnd vdd FILL
XFILL_3__14959_ gnd vdd FILL
XFILL_5__15519_ gnd vdd FILL
XFILL_0__14779_ gnd vdd FILL
X_8925_ _8925_/Q _7389_/CLK _8285_/R vdd _8845_/Y gnd vdd DFFSR
XFILL_0__9277_ gnd vdd FILL
XFILL_3__8006_ gnd vdd FILL
XFILL_1__8070_ gnd vdd FILL
XFILL_2__15339_ gnd vdd FILL
XFILL_0__8228_ gnd vdd FILL
X_8856_ _8893_/B _8472_/B gnd _8857_/C vdd NAND2X1
XSFILL23720x37050 gnd vdd FILL
XFILL_0__16449_ gnd vdd FILL
X_7807_ _7807_/A gnd _7807_/Y vdd INVX1
XSFILL33880x81050 gnd vdd FILL
XFILL_4__8750_ gnd vdd FILL
XSFILL18840x5050 gnd vdd FILL
X_8787_ _8821_/Q gnd _8789_/A vdd INVX1
XFILL_6__6878_ gnd vdd FILL
XFILL_1__8972_ gnd vdd FILL
X_7738_ _7736_/Y _7672_/B _7737_/Y gnd _7738_/Y vdd OAI21X1
XFILL_4__7701_ gnd vdd FILL
XFILL_3__8908_ gnd vdd FILL
XFILL_3__9888_ gnd vdd FILL
XSFILL64200x51050 gnd vdd FILL
XFILL_6__9597_ gnd vdd FILL
X_7669_ _7669_/Q _9589_/CLK _7285_/R vdd _7669_/D gnd vdd DFFSR
XFILL_3__8839_ gnd vdd FILL
XFILL_4__7632_ gnd vdd FILL
X_9408_ _9406_/Y _9420_/B _9408_/C gnd _9454_/D vdd OAI21X1
XFILL_1__7854_ gnd vdd FILL
XFILL_4__7563_ gnd vdd FILL
X_11270_ _11078_/Y _11270_/B gnd _11270_/Y vdd NOR2X1
X_9339_ _9339_/A _9339_/B _9338_/Y gnd _9339_/Y vdd OAI21X1
XFILL_4_BUFX2_insert233 gnd vdd FILL
XSFILL28840x70050 gnd vdd FILL
XFILL_4_BUFX2_insert244 gnd vdd FILL
X_10221_ _10171_/A _8947_/CLK _8038_/R vdd _10221_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert255 gnd vdd FILL
XFILL_4__7494_ gnd vdd FILL
XFILL_1__9524_ gnd vdd FILL
XFILL_4_BUFX2_insert266 gnd vdd FILL
XFILL_4_BUFX2_insert277 gnd vdd FILL
XFILL_4__9233_ gnd vdd FILL
XFILL_4_BUFX2_insert288 gnd vdd FILL
X_10152_ _10150_/Y _10191_/B _10152_/C gnd _10152_/Y vdd OAI21X1
XFILL_4_BUFX2_insert299 gnd vdd FILL
XFILL_3_BUFX2_insert900 gnd vdd FILL
XSFILL3480x5050 gnd vdd FILL
XFILL_3_BUFX2_insert911 gnd vdd FILL
XSFILL8760x68050 gnd vdd FILL
XFILL_3_BUFX2_insert922 gnd vdd FILL
XSFILL23800x17050 gnd vdd FILL
XFILL_3_BUFX2_insert933 gnd vdd FILL
XFILL_4__9164_ gnd vdd FILL
XSFILL33960x61050 gnd vdd FILL
XFILL_3_BUFX2_insert944 gnd vdd FILL
XFILL_3_BUFX2_insert955 gnd vdd FILL
X_14960_ _9333_/Q gnd _14960_/Y vdd INVX1
X_10083_ _14098_/C _9077_/CLK _7665_/R vdd _10015_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert966 gnd vdd FILL
XFILL_3_BUFX2_insert977 gnd vdd FILL
XSFILL49240x28050 gnd vdd FILL
XFILL_1__9386_ gnd vdd FILL
XFILL_4__8115_ gnd vdd FILL
XFILL_3_BUFX2_insert988 gnd vdd FILL
XFILL_4__9095_ gnd vdd FILL
X_13911_ _9695_/Q gnd _13911_/Y vdd INVX1
XFILL_3_BUFX2_insert999 gnd vdd FILL
XSFILL89640x33050 gnd vdd FILL
XFILL_1__8337_ gnd vdd FILL
X_14891_ _14889_/Y _14891_/B _14891_/C gnd _14907_/B vdd NAND3X1
X_13842_ _7262_/Q gnd _13842_/Y vdd INVX1
XFILL_1__8268_ gnd vdd FILL
XFILL_3_BUFX2_insert1005 gnd vdd FILL
XFILL_2__7061_ gnd vdd FILL
XSFILL13720x69050 gnd vdd FILL
XFILL_3_BUFX2_insert1016 gnd vdd FILL
XFILL_1_BUFX2_insert101 gnd vdd FILL
XSFILL28520x29050 gnd vdd FILL
XFILL_3_BUFX2_insert1027 gnd vdd FILL
XFILL_3_BUFX2_insert1038 gnd vdd FILL
X_13773_ _8924_/Q gnd _13773_/Y vdd INVX1
XFILL_1__7219_ gnd vdd FILL
X_10985_ _10911_/A _12667_/CLK _12689_/R vdd _10985_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert1049 gnd vdd FILL
XFILL_5__7810_ gnd vdd FILL
XFILL_1__8199_ gnd vdd FILL
X_15512_ _15708_/A _15512_/B _15708_/C gnd _15535_/B vdd NOR3X1
X_12724_ _12722_/Y _12723_/A _12724_/C gnd _12724_/Y vdd OAI21X1
XFILL_4__9997_ gnd vdd FILL
XFILL_3__10640_ gnd vdd FILL
XFILL_5__7741_ gnd vdd FILL
XFILL_5__11200_ gnd vdd FILL
X_15443_ _7185_/A gnd _15444_/A vdd INVX1
X_12655_ vdd memoryOutData[29] gnd _12655_/Y vdd NAND2X1
XFILL_5__12180_ gnd vdd FILL
XFILL_4__11930_ gnd vdd FILL
XFILL_0_BUFX2_insert801 gnd vdd FILL
XFILL_2__11020_ gnd vdd FILL
XFILL_0_BUFX2_insert812 gnd vdd FILL
XFILL_3__10571_ gnd vdd FILL
XFILL_0_BUFX2_insert823 gnd vdd FILL
XFILL_2__7963_ gnd vdd FILL
XFILL_1__11750_ gnd vdd FILL
XFILL_0__10391_ gnd vdd FILL
XFILL_5__7672_ gnd vdd FILL
XFILL_0_BUFX2_insert834 gnd vdd FILL
X_11606_ _11587_/C _11574_/B _11606_/C gnd _11608_/B vdd OAI21X1
XFILL_5__11131_ gnd vdd FILL
XFILL_4__8879_ gnd vdd FILL
X_15374_ _15652_/A _9566_/Q _9694_/Q _15652_/D gnd _15381_/A vdd AOI22X1
XFILL_3__12310_ gnd vdd FILL
XFILL_0_BUFX2_insert845 gnd vdd FILL
XFILL_0_BUFX2_insert856 gnd vdd FILL
X_12586_ vdd memoryOutData[6] gnd _12587_/C vdd NAND2X1
XFILL_1_BUFX2_insert1020 gnd vdd FILL
XFILL_2__6914_ gnd vdd FILL
XFILL_6__10682_ gnd vdd FILL
XFILL_4__11861_ gnd vdd FILL
XFILL_3__13290_ gnd vdd FILL
XFILL_1__10701_ gnd vdd FILL
XFILL_1_BUFX2_insert1031 gnd vdd FILL
XFILL_0__12130_ gnd vdd FILL
XFILL_5__9411_ gnd vdd FILL
XFILL_0_BUFX2_insert867 gnd vdd FILL
XFILL_0_BUFX2_insert878 gnd vdd FILL
XFILL_1__11681_ gnd vdd FILL
XFILL_1_BUFX2_insert1042 gnd vdd FILL
XSFILL99480x36050 gnd vdd FILL
X_14325_ _9772_/A gnd _14325_/Y vdd INVX1
XFILL_4__13600_ gnd vdd FILL
XFILL_4__10812_ gnd vdd FILL
XFILL_1_BUFX2_insert1053 gnd vdd FILL
XFILL_0_BUFX2_insert889 gnd vdd FILL
X_11537_ _11537_/A _11550_/C _11295_/Y gnd _11537_/Y vdd OAI21X1
XFILL_5__11062_ gnd vdd FILL
XFILL_4__14580_ gnd vdd FILL
XFILL_1_BUFX2_insert1064 gnd vdd FILL
XFILL_2__9633_ gnd vdd FILL
XFILL_3__12241_ gnd vdd FILL
XSFILL74120x34050 gnd vdd FILL
XFILL_2__6845_ gnd vdd FILL
XFILL_1__10632_ gnd vdd FILL
XFILL_3_BUFX2_insert16 gnd vdd FILL
XFILL_1__13420_ gnd vdd FILL
XFILL_4__11792_ gnd vdd FILL
XFILL_0__12061_ gnd vdd FILL
XFILL_2__12971_ gnd vdd FILL
XFILL_5__9342_ gnd vdd FILL
XFILL_3_BUFX2_insert27 gnd vdd FILL
XFILL_1_BUFX2_insert1086 gnd vdd FILL
XFILL_5__10013_ gnd vdd FILL
XFILL_3_BUFX2_insert38 gnd vdd FILL
X_14256_ _14615_/B _15718_/D _14256_/C _13846_/A gnd _14256_/Y vdd OAI22X1
XFILL_4__13531_ gnd vdd FILL
XFILL_4__10743_ gnd vdd FILL
XFILL_3_BUFX2_insert49 gnd vdd FILL
XFILL_2__14710_ gnd vdd FILL
X_11468_ _11171_/Y _11484_/B _11366_/B _11467_/Y gnd _11470_/C vdd OAI22X1
XFILL_5__15870_ gnd vdd FILL
XFILL_2__11922_ gnd vdd FILL
XFILL_3__12172_ gnd vdd FILL
XFILL_0__11012_ gnd vdd FILL
XFILL_1__13351_ gnd vdd FILL
XFILL_2__15690_ gnd vdd FILL
XFILL_1__10563_ gnd vdd FILL
X_13207_ _13289_/B gnd _13295_/C vdd INVX4
XFILL_5__9273_ gnd vdd FILL
XFILL_6__11303_ gnd vdd FILL
XFILL_5__14821_ gnd vdd FILL
XFILL_6__15071_ gnd vdd FILL
X_10419_ _10426_/B _9267_/B gnd _10419_/Y vdd NAND2X1
X_14187_ _10213_/Q gnd _14187_/Y vdd INVX1
XFILL_4__13462_ gnd vdd FILL
XSFILL13800x49050 gnd vdd FILL
XFILL_2__8515_ gnd vdd FILL
XFILL_3__11123_ gnd vdd FILL
XFILL_4__16250_ gnd vdd FILL
XFILL_2__14641_ gnd vdd FILL
XFILL_1__12302_ gnd vdd FILL
X_11399_ _11096_/C gnd _11400_/C vdd INVX1
XFILL_6_CLKBUF1_insert111 gnd vdd FILL
XFILL_4__10674_ gnd vdd FILL
XFILL_1__13282_ gnd vdd FILL
XFILL_2__9495_ gnd vdd FILL
XFILL_5__8224_ gnd vdd FILL
XFILL_0__15820_ gnd vdd FILL
XFILL_1__16070_ gnd vdd FILL
XFILL_2__11853_ gnd vdd FILL
XFILL_6__14022_ gnd vdd FILL
XFILL_1__10494_ gnd vdd FILL
XFILL_4__12413_ gnd vdd FILL
XFILL_4__15201_ gnd vdd FILL
X_13138_ _13136_/Y _13134_/A _13138_/C gnd _13194_/D vdd OAI21X1
XFILL_4__16181_ gnd vdd FILL
XFILL_5__14752_ gnd vdd FILL
XFILL112280x60050 gnd vdd FILL
XFILL_4__13393_ gnd vdd FILL
XFILL_1__15021_ gnd vdd FILL
XFILL_3__15931_ gnd vdd FILL
XFILL_5__11964_ gnd vdd FILL
XFILL_1__12233_ gnd vdd FILL
XFILL_3__11054_ gnd vdd FILL
XFILL_2__8446_ gnd vdd FILL
XFILL_2__10804_ gnd vdd FILL
XFILL_2__14572_ gnd vdd FILL
XFILL_0__15751_ gnd vdd FILL
XFILL_2__11784_ gnd vdd FILL
XFILL_0__12963_ gnd vdd FILL
XFILL_6__11165_ gnd vdd FILL
XFILL_5__13703_ gnd vdd FILL
XFILL_4__15132_ gnd vdd FILL
XFILL_6_CLKBUF1_insert188 gnd vdd FILL
XFILL_5__10915_ gnd vdd FILL
XFILL_4__12344_ gnd vdd FILL
XFILL_0__7461_ gnd vdd FILL
X_13069_ _6892_/A _13201_/CLK _13201_/R vdd _13069_/D gnd vdd DFFSR
XFILL_2__16311_ gnd vdd FILL
XFILL_3__10005_ gnd vdd FILL
XFILL_2__13523_ gnd vdd FILL
XFILL_5__14683_ gnd vdd FILL
XFILL_2__8377_ gnd vdd FILL
XFILL_3__7170_ gnd vdd FILL
XFILL_5__11895_ gnd vdd FILL
XFILL_1__12164_ gnd vdd FILL
XFILL_0__14702_ gnd vdd FILL
XFILL_5__7106_ gnd vdd FILL
XFILL_3__15862_ gnd vdd FILL
XFILL_0__11914_ gnd vdd FILL
XFILL_0__15682_ gnd vdd FILL
XFILL_0__12894_ gnd vdd FILL
XFILL_5__8086_ gnd vdd FILL
XFILL_5__13634_ gnd vdd FILL
XFILL_4__15063_ gnd vdd FILL
XFILL_2__16242_ gnd vdd FILL
XFILL_3__14813_ gnd vdd FILL
XFILL_2__7328_ gnd vdd FILL
XSFILL43880x44050 gnd vdd FILL
XFILL_4__12275_ gnd vdd FILL
XFILL_1__11115_ gnd vdd FILL
XFILL_2__13454_ gnd vdd FILL
XFILL_3__15793_ gnd vdd FILL
XFILL_0__14633_ gnd vdd FILL
XFILL_1__12095_ gnd vdd FILL
XFILL_2__10666_ gnd vdd FILL
XFILL_5__7037_ gnd vdd FILL
XFILL_0__11845_ gnd vdd FILL
XFILL_4__14014_ gnd vdd FILL
XFILL_0__9131_ gnd vdd FILL
XFILL_5__16353_ gnd vdd FILL
XFILL_4__11226_ gnd vdd FILL
XFILL_2__12405_ gnd vdd FILL
XFILL_5__10777_ gnd vdd FILL
XSFILL34600x28050 gnd vdd FILL
XFILL_5__13565_ gnd vdd FILL
XFILL_3__14744_ gnd vdd FILL
X_6971_ _7021_/Q gnd _6971_/Y vdd INVX1
XFILL_1__15923_ gnd vdd FILL
XFILL_2__16173_ gnd vdd FILL
XFILL_3__11956_ gnd vdd FILL
XFILL_1__11046_ gnd vdd FILL
XSFILL18680x20050 gnd vdd FILL
XFILL_2__13385_ gnd vdd FILL
XFILL_0__14564_ gnd vdd FILL
XFILL_5__15304_ gnd vdd FILL
XSFILL74200x14050 gnd vdd FILL
XFILL_0__11776_ gnd vdd FILL
XFILL_5__12516_ gnd vdd FILL
X_8710_ _8698_/A _9478_/B gnd _8710_/Y vdd NAND2X1
XSFILL18920x82050 gnd vdd FILL
XFILL_3__10907_ gnd vdd FILL
XFILL_5__16284_ gnd vdd FILL
XFILL_4__11157_ gnd vdd FILL
XFILL_2__15124_ gnd vdd FILL
X_9690_ _9602_/A _9707_/CLK _8819_/R vdd _9690_/D gnd vdd DFFSR
XFILL_0__16303_ gnd vdd FILL
XFILL_2__12336_ gnd vdd FILL
XFILL_3__14675_ gnd vdd FILL
XFILL_5__13496_ gnd vdd FILL
XFILL_3__11887_ gnd vdd FILL
XFILL_1__15854_ gnd vdd FILL
XFILL_6_BUFX2_insert306 gnd vdd FILL
XFILL_0__13515_ gnd vdd FILL
XFILL_0__8013_ gnd vdd FILL
XFILL_0__14495_ gnd vdd FILL
XSFILL59000x75050 gnd vdd FILL
XFILL_5__15235_ gnd vdd FILL
XFILL_4__10108_ gnd vdd FILL
XFILL_3__13626_ gnd vdd FILL
XFILL_5__12447_ gnd vdd FILL
XFILL_5__8988_ gnd vdd FILL
XSFILL108920x35050 gnd vdd FILL
XFILL_3__16414_ gnd vdd FILL
X_8641_ _8687_/Q gnd _8641_/Y vdd INVX1
XFILL_1__14805_ gnd vdd FILL
XFILL_6__11998_ gnd vdd FILL
XFILL_2__15055_ gnd vdd FILL
XFILL_4__15965_ gnd vdd FILL
XFILL_3__9811_ gnd vdd FILL
XFILL_4__11088_ gnd vdd FILL
XSFILL99400x80050 gnd vdd FILL
XFILL_0__16234_ gnd vdd FILL
XFILL_0__13446_ gnd vdd FILL
XFILL_2__12267_ gnd vdd FILL
XFILL_0__10658_ gnd vdd FILL
XFILL_1__15785_ gnd vdd FILL
XFILL_1__12997_ gnd vdd FILL
XFILL_5__7939_ gnd vdd FILL
XSFILL78840x17050 gnd vdd FILL
XFILL_4__10039_ gnd vdd FILL
XFILL_3__16345_ gnd vdd FILL
XFILL_2__14006_ gnd vdd FILL
XFILL_5__12378_ gnd vdd FILL
XFILL_5__15166_ gnd vdd FILL
XFILL_4__14916_ gnd vdd FILL
XFILL_1_BUFX2_insert690 gnd vdd FILL
XFILL_3__9742_ gnd vdd FILL
XSFILL23240x54050 gnd vdd FILL
XFILL_3__13557_ gnd vdd FILL
X_8572_ _8572_/A gnd _8574_/A vdd INVX1
XFILL_2__11218_ gnd vdd FILL
XFILL_4__15896_ gnd vdd FILL
XFILL_1__14736_ gnd vdd FILL
XFILL_3__10769_ gnd vdd FILL
XFILL_3__6954_ gnd vdd FILL
XFILL_0__13377_ gnd vdd FILL
XFILL_0__16165_ gnd vdd FILL
XFILL_1__11948_ gnd vdd FILL
XSFILL38840x33050 gnd vdd FILL
XFILL_2__12198_ gnd vdd FILL
XFILL_5__14117_ gnd vdd FILL
XSFILL64120x66050 gnd vdd FILL
XFILL_3__12508_ gnd vdd FILL
X_7523_ _7523_/Q _7530_/CLK _7523_/R vdd _7455_/Y gnd vdd DFFSR
XFILL_5__11329_ gnd vdd FILL
XFILL_4__14847_ gnd vdd FILL
XFILL_5__15097_ gnd vdd FILL
XFILL_3__16276_ gnd vdd FILL
XFILL_3__9673_ gnd vdd FILL
XFILL_0__12328_ gnd vdd FILL
XFILL_6__8402_ gnd vdd FILL
XFILL_2__11149_ gnd vdd FILL
XFILL_3__13488_ gnd vdd FILL
XFILL_0__15116_ gnd vdd FILL
XFILL_5__9609_ gnd vdd FILL
XFILL_3__6885_ gnd vdd FILL
XFILL_0__16096_ gnd vdd FILL
XFILL_1__14667_ gnd vdd FILL
XFILL_6__12619_ gnd vdd FILL
XFILL_1__11879_ gnd vdd FILL
XFILL_0__8915_ gnd vdd FILL
XFILL_3__15227_ gnd vdd FILL
XFILL_5__14048_ gnd vdd FILL
X_7454_ _7430_/A _8606_/B gnd _7454_/Y vdd NAND2X1
XFILL_0__9895_ gnd vdd FILL
XFILL_3__12439_ gnd vdd FILL
XFILL_1__16406_ gnd vdd FILL
XFILL_3__8624_ gnd vdd FILL
XFILL_1__13618_ gnd vdd FILL
XFILL_2__15957_ gnd vdd FILL
XFILL_0__15047_ gnd vdd FILL
XFILL_4__14778_ gnd vdd FILL
XFILL_0__12259_ gnd vdd FILL
XFILL_1__14598_ gnd vdd FILL
XSFILL43960x24050 gnd vdd FILL
XFILL_0__8846_ gnd vdd FILL
X_7385_ _7295_/A _7129_/CLK _9049_/R vdd _7385_/D gnd vdd DFFSR
XSFILL3560x73050 gnd vdd FILL
XSFILL68760x69050 gnd vdd FILL
XFILL_3__15158_ gnd vdd FILL
XFILL_4__13729_ gnd vdd FILL
XFILL_1__16337_ gnd vdd FILL
XFILL_2__14908_ gnd vdd FILL
XFILL_1__13549_ gnd vdd FILL
XFILL_2__15888_ gnd vdd FILL
X_9124_ _9151_/A _9380_/B gnd _9125_/C vdd NAND2X1
XFILL_3__14109_ gnd vdd FILL
XSFILL8600x10050 gnd vdd FILL
XFILL_1__7570_ gnd vdd FILL
XFILL_3__7506_ gnd vdd FILL
XFILL_0__8777_ gnd vdd FILL
XFILL_2__14839_ gnd vdd FILL
XFILL_5__15999_ gnd vdd FILL
XFILL_3__15089_ gnd vdd FILL
XFILL_3__8486_ gnd vdd FILL
XFILL_1__16268_ gnd vdd FILL
XFILL_0__7728_ gnd vdd FILL
X_9055_ _9055_/Q _9823_/CLK _9823_/R vdd _9055_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert229 gnd vdd FILL
XFILL_3__7437_ gnd vdd FILL
XFILL_1__15219_ gnd vdd FILL
XFILL_4__16379_ gnd vdd FILL
XFILL_1__16199_ gnd vdd FILL
XFILL_0__15949_ gnd vdd FILL
XSFILL103560x80050 gnd vdd FILL
XFILL_1__9240_ gnd vdd FILL
X_8006_ _8006_/A _8006_/B _8005_/Y gnd _8006_/Y vdd OAI21X1
XSFILL33880x76050 gnd vdd FILL
XFILL_3__7368_ gnd vdd FILL
XFILL_2_BUFX2_insert907 gnd vdd FILL
XFILL_2_BUFX2_insert918 gnd vdd FILL
XFILL_1__9171_ gnd vdd FILL
XFILL_3__9107_ gnd vdd FILL
XFILL_2_BUFX2_insert929 gnd vdd FILL
XFILL112440x20050 gnd vdd FILL
XFILL_3__7299_ gnd vdd FILL
XSFILL64200x46050 gnd vdd FILL
XFILL_1__8122_ gnd vdd FILL
XFILL_3__9038_ gnd vdd FILL
X_9957_ _9957_/Q _9817_/CLK _7150_/R vdd _9893_/Y gnd vdd DFFSR
XFILL_4__9920_ gnd vdd FILL
XSFILL39000x22050 gnd vdd FILL
X_8908_ _8906_/Y _8893_/B _8908_/C gnd _8946_/D vdd OAI21X1
XSFILL8600x1050 gnd vdd FILL
X_9888_ _9888_/A gnd _9890_/A vdd INVX1
XSFILL3640x53050 gnd vdd FILL
XFILL_4__9851_ gnd vdd FILL
X_10770_ _10773_/A _7186_/B gnd _10771_/C vdd NAND2X1
X_8839_ _8839_/A _8916_/A _8839_/C gnd _8923_/D vdd OAI21X1
XFILL_4__9782_ gnd vdd FILL
XBUFX2_insert906 _10913_/Y gnd _12789_/A vdd BUFX2
XSFILL94280x41050 gnd vdd FILL
XSFILL115160x7050 gnd vdd FILL
XFILL_4__6994_ gnd vdd FILL
XFILL_0_BUFX2_insert108 gnd vdd FILL
XBUFX2_insert917 _15069_/Y gnd _15070_/C vdd BUFX2
XBUFX2_insert928 _12351_/Y gnd _9981_/B vdd BUFX2
XFILL_4__8733_ gnd vdd FILL
XFILL_6_BUFX2_insert884 gnd vdd FILL
XBUFX2_insert939 _13423_/Y gnd _14752_/C vdd BUFX2
X_12440_ _12440_/A vdd gnd _12440_/Y vdd NAND2X1
XFILL_1__8955_ gnd vdd FILL
XSFILL33960x56050 gnd vdd FILL
X_12371_ _12371_/A _12594_/A gnd _12372_/C vdd NAND2X1
XFILL_1__8886_ gnd vdd FILL
XFILL_4__7615_ gnd vdd FILL
X_14110_ _8163_/Q gnd _14111_/A vdd INVX1
X_11322_ _11321_/Y gnd _11325_/B vdd INVX1
XFILL_4__8595_ gnd vdd FILL
X_15090_ _15000_/A _15061_/C _16035_/B gnd _16225_/C vdd NAND3X1
XFILL_1__7837_ gnd vdd FILL
XFILL_4__7546_ gnd vdd FILL
X_14041_ _7394_/Q gnd _14041_/Y vdd INVX1
X_11253_ _11026_/C _11253_/B _11026_/A gnd _11253_/Y vdd AOI21X1
XSFILL48600x80050 gnd vdd FILL
XFILL_4__7477_ gnd vdd FILL
X_10204_ _10120_/A _7269_/CLK _8165_/R vdd _10204_/D gnd vdd DFFSR
XFILL_1__9507_ gnd vdd FILL
X_11184_ _11184_/A _11191_/B gnd _11185_/C vdd NOR2X1
XFILL_2__9280_ gnd vdd FILL
XFILL_4__9216_ gnd vdd FILL
XSFILL3720x33050 gnd vdd FILL
XFILL_1__7699_ gnd vdd FILL
XFILL_3_BUFX2_insert730 gnd vdd FILL
XSFILL94360x6050 gnd vdd FILL
X_10135_ _13994_/A gnd _10137_/A vdd INVX1
XFILL_3_BUFX2_insert741 gnd vdd FILL
X_15992_ _15204_/A _14574_/Y _14582_/Y _15912_/D gnd _15993_/B vdd OAI22X1
XFILL_3_BUFX2_insert752 gnd vdd FILL
XFILL_2__8231_ gnd vdd FILL
XFILL_4__10390_ gnd vdd FILL
XFILL_4__9147_ gnd vdd FILL
XFILL_3_BUFX2_insert763 gnd vdd FILL
XFILL_3_BUFX2_insert774 gnd vdd FILL
XFILL_5__10700_ gnd vdd FILL
XFILL_3_BUFX2_insert785 gnd vdd FILL
X_14943_ _7157_/Q _14847_/C _14481_/C _7029_/Q gnd _14951_/B vdd AOI22X1
X_10066_ _10064_/Y _10066_/B _10065_/Y gnd _10066_/Y vdd OAI21X1
XSFILL69000x38050 gnd vdd FILL
XFILL_5__11680_ gnd vdd FILL
XFILL_3_BUFX2_insert796 gnd vdd FILL
XFILL_1__9369_ gnd vdd FILL
XFILL_2__10520_ gnd vdd FILL
XSFILL79160x82050 gnd vdd FILL
XFILL_4__9078_ gnd vdd FILL
XFILL_5__10631_ gnd vdd FILL
X_14874_ _8525_/A gnd _14875_/D vdd INVX1
XFILL_4__12060_ gnd vdd FILL
XFILL_2__7113_ gnd vdd FILL
XFILL_3__11810_ gnd vdd FILL
XFILL_3__12790_ gnd vdd FILL
XFILL_2__10451_ gnd vdd FILL
XFILL_2__8093_ gnd vdd FILL
XFILL_0__11630_ gnd vdd FILL
XFILL_5__8911_ gnd vdd FILL
X_13825_ _13825_/A _13825_/B gnd _13825_/Y vdd NOR2X1
XFILL_4__11011_ gnd vdd FILL
XFILL_5__13350_ gnd vdd FILL
XFILL_5__9891_ gnd vdd FILL
XSFILL8440x45050 gnd vdd FILL
XFILL_5__10562_ gnd vdd FILL
XFILL_2__7044_ gnd vdd FILL
XFILL_3__11741_ gnd vdd FILL
XFILL_2__10382_ gnd vdd FILL
XFILL_2__13170_ gnd vdd FILL
XFILL_0__11561_ gnd vdd FILL
XFILL_5__8842_ gnd vdd FILL
XSFILL84280x73050 gnd vdd FILL
XFILL_5__12301_ gnd vdd FILL
XFILL_5__13281_ gnd vdd FILL
X_13756_ _10716_/Q gnd _13758_/B vdd INVX1
XFILL_0__13300_ gnd vdd FILL
X_10968_ _12818_/Q _10968_/B gnd _10969_/D vdd NAND2X1
XFILL_3__14460_ gnd vdd FILL
XFILL_2__12121_ gnd vdd FILL
XFILL_5__10493_ gnd vdd FILL
XFILL_0__10512_ gnd vdd FILL
XFILL_3__11672_ gnd vdd FILL
XFILL_1__12851_ gnd vdd FILL
XFILL_0__14280_ gnd vdd FILL
X_12707_ _12707_/A gnd _12709_/A vdd INVX1
XFILL_5__15020_ gnd vdd FILL
XFILL_5__8773_ gnd vdd FILL
XFILL_5__12232_ gnd vdd FILL
XFILL_0__11492_ gnd vdd FILL
XFILL_3__13411_ gnd vdd FILL
XFILL_3__10623_ gnd vdd FILL
X_13687_ _13865_/C _7771_/Q _15268_/A _14956_/D gnd _13698_/A vdd AOI22X1
XFILL_4__15750_ gnd vdd FILL
XFILL_0__13231_ gnd vdd FILL
X_10899_ _10911_/A gnd _10903_/A vdd INVX1
XFILL_4__12962_ gnd vdd FILL
XFILL_2__12052_ gnd vdd FILL
XFILL_3__14391_ gnd vdd FILL
XFILL_1__11802_ gnd vdd FILL
XFILL_0__10443_ gnd vdd FILL
XFILL_2__8995_ gnd vdd FILL
XFILL_1__15570_ gnd vdd FILL
XFILL_5__7724_ gnd vdd FILL
XSFILL109480x16050 gnd vdd FILL
XFILL_1__12782_ gnd vdd FILL
XFILL_0_BUFX2_insert620 gnd vdd FILL
XSFILL8760x7050 gnd vdd FILL
X_15426_ _15415_/Y _15426_/B _15426_/C gnd _15434_/B vdd NAND3X1
X_12638_ _12636_/Y vdd _12638_/C gnd _12686_/D vdd OAI21X1
XFILL_5__12163_ gnd vdd FILL
XFILL_4__14701_ gnd vdd FILL
XFILL_3__16130_ gnd vdd FILL
XFILL_0_BUFX2_insert631 gnd vdd FILL
XFILL_3__13342_ gnd vdd FILL
XFILL_4__11913_ gnd vdd FILL
XSFILL38760x48050 gnd vdd FILL
XFILL_0_BUFX2_insert642 gnd vdd FILL
XSFILL54120x9050 gnd vdd FILL
XFILL_2__11003_ gnd vdd FILL
XFILL_2__7946_ gnd vdd FILL
XFILL_4__15681_ gnd vdd FILL
XFILL_4__12893_ gnd vdd FILL
XFILL_0_BUFX2_insert653 gnd vdd FILL
XFILL_1__14521_ gnd vdd FILL
XFILL_3__10554_ gnd vdd FILL
XFILL112280x55050 gnd vdd FILL
XFILL_0__13162_ gnd vdd FILL
XFILL_1__11733_ gnd vdd FILL
XFILL_0__10374_ gnd vdd FILL
XFILL_5__11114_ gnd vdd FILL
XFILL_0_BUFX2_insert664 gnd vdd FILL
X_15357_ _10763_/A _15357_/B _15916_/B _10717_/Q gnd _15357_/Y vdd AOI22X1
XFILL_0_BUFX2_insert675 gnd vdd FILL
X_12569_ _12567_/Y vdd _12569_/C gnd _12663_/D vdd OAI21X1
XFILL_4__14632_ gnd vdd FILL
XFILL_5__12094_ gnd vdd FILL
XFILL_0__6961_ gnd vdd FILL
XFILL_0_BUFX2_insert686 gnd vdd FILL
XFILL_2__15811_ gnd vdd FILL
XFILL_3__16061_ gnd vdd FILL
XFILL_4__11844_ gnd vdd FILL
XFILL_3__13273_ gnd vdd FILL
XFILL_0__12113_ gnd vdd FILL
XFILL_0_BUFX2_insert697 gnd vdd FILL
XFILL_1__14452_ gnd vdd FILL
XFILL_2__7877_ gnd vdd FILL
XFILL_0__13093_ gnd vdd FILL
X_14308_ _14307_/Y _13574_/C gnd _14309_/C vdd NOR2X1
XFILL_0__8700_ gnd vdd FILL
XFILL_1__11664_ gnd vdd FILL
XFILL_5__15922_ gnd vdd FILL
XFILL_5__7586_ gnd vdd FILL
XFILL_3__15012_ gnd vdd FILL
XFILL_5__11045_ gnd vdd FILL
XFILL_2__9616_ gnd vdd FILL
XFILL_3__12224_ gnd vdd FILL
X_15288_ _15774_/C _13689_/A _15287_/Y _15801_/C gnd _15289_/A vdd OAI22X1
XFILL_0__9680_ gnd vdd FILL
XFILL_4__14563_ gnd vdd FILL
XSFILL79240x62050 gnd vdd FILL
XFILL_1__13403_ gnd vdd FILL
XSFILL43880x39050 gnd vdd FILL
XFILL_0__6892_ gnd vdd FILL
XFILL_2__15742_ gnd vdd FILL
XFILL_4__11775_ gnd vdd FILL
XSFILL114840x69050 gnd vdd FILL
XFILL_0__12044_ gnd vdd FILL
XFILL_1__10615_ gnd vdd FILL
XFILL_2__12954_ gnd vdd FILL
XFILL_1__14383_ gnd vdd FILL
XFILL_1__11595_ gnd vdd FILL
XFILL_0__8631_ gnd vdd FILL
X_14239_ _9382_/A gnd _14240_/D vdd INVX1
XFILL_4__16302_ gnd vdd FILL
X_7170_ _7258_/Q gnd _7172_/A vdd INVX1
XFILL_5__15853_ gnd vdd FILL
XFILL_4__13514_ gnd vdd FILL
XFILL_2__9547_ gnd vdd FILL
XFILL_4__14494_ gnd vdd FILL
XFILL_2__11905_ gnd vdd FILL
XFILL_1__16122_ gnd vdd FILL
XFILL_3__8340_ gnd vdd FILL
XFILL_3__12155_ gnd vdd FILL
XFILL_1__13334_ gnd vdd FILL
XFILL_2__15673_ gnd vdd FILL
XSFILL18680x15050 gnd vdd FILL
XFILL_5__9256_ gnd vdd FILL
XFILL_2__12885_ gnd vdd FILL
XFILL_1__10546_ gnd vdd FILL
XSFILL114440x71050 gnd vdd FILL
XFILL_5__14804_ gnd vdd FILL
XFILL_4__16233_ gnd vdd FILL
XFILL_3__11106_ gnd vdd FILL
XFILL_2__14624_ gnd vdd FILL
XFILL_4__10657_ gnd vdd FILL
XFILL_4__13445_ gnd vdd FILL
XFILL_5__15784_ gnd vdd FILL
XFILL_5__8207_ gnd vdd FILL
XFILL_3__8271_ gnd vdd FILL
XFILL_5__12996_ gnd vdd FILL
XFILL_3__12086_ gnd vdd FILL
XSFILL84360x53050 gnd vdd FILL
XFILL_0__15803_ gnd vdd FILL
XFILL_2__9478_ gnd vdd FILL
XFILL_1__16053_ gnd vdd FILL
XFILL_2__11836_ gnd vdd FILL
XFILL_1__13265_ gnd vdd FILL
XFILL_5__14735_ gnd vdd FILL
XFILL_0__13995_ gnd vdd FILL
XFILL_3__7222_ gnd vdd FILL
XFILL_3__15914_ gnd vdd FILL
XFILL_4__13376_ gnd vdd FILL
XFILL_5__11947_ gnd vdd FILL
XFILL_0__8493_ gnd vdd FILL
XFILL_3__11037_ gnd vdd FILL
XFILL_1__15004_ gnd vdd FILL
XFILL_4__16164_ gnd vdd FILL
XFILL_2__14555_ gnd vdd FILL
XFILL_1__12216_ gnd vdd FILL
XSFILL99400x75050 gnd vdd FILL
XFILL_5__8138_ gnd vdd FILL
XFILL_2__11767_ gnd vdd FILL
XFILL_0__15734_ gnd vdd FILL
XFILL_4__12327_ gnd vdd FILL
XFILL_0__7444_ gnd vdd FILL
XFILL_4__15115_ gnd vdd FILL
XFILL111720x69050 gnd vdd FILL
XFILL_5__14666_ gnd vdd FILL
XFILL_2__13506_ gnd vdd FILL
XFILL_5__11878_ gnd vdd FILL
XFILL_4__16095_ gnd vdd FILL
XFILL_3__15845_ gnd vdd FILL
XFILL_2__14486_ gnd vdd FILL
XFILL_1__12147_ gnd vdd FILL
XFILL_0__15665_ gnd vdd FILL
XFILL_5__16405_ gnd vdd FILL
XSFILL38840x28050 gnd vdd FILL
XFILL_2__11698_ gnd vdd FILL
XFILL_5__8069_ gnd vdd FILL
XFILL_5__13617_ gnd vdd FILL
XFILL_6__8951_ gnd vdd FILL
XFILL112360x35050 gnd vdd FILL
XFILL_0__12877_ gnd vdd FILL
X_9811_ _9811_/A gnd _9811_/Y vdd INVX1
XFILL_5__10829_ gnd vdd FILL
XFILL_2__16225_ gnd vdd FILL
XFILL_0__7375_ gnd vdd FILL
XFILL_6__15956_ gnd vdd FILL
XFILL_4__15046_ gnd vdd FILL
XSFILL24680x34050 gnd vdd FILL
XFILL_4__12258_ gnd vdd FILL
XFILL_5__14597_ gnd vdd FILL
XFILL_2__13437_ gnd vdd FILL
XFILL_0__14616_ gnd vdd FILL
XFILL_1__12078_ gnd vdd FILL
XFILL_2__10649_ gnd vdd FILL
XFILL_3__12988_ gnd vdd FILL
XFILL_3__15776_ gnd vdd FILL
XFILL_3__7084_ gnd vdd FILL
XFILL_0__9114_ gnd vdd FILL
XFILL_0__11828_ gnd vdd FILL
XFILL_5__16336_ gnd vdd FILL
XFILL_0__15596_ gnd vdd FILL
XFILL_6__14907_ gnd vdd FILL
XFILL_4__11209_ gnd vdd FILL
X_9742_ _9742_/A gnd _9742_/Y vdd INVX1
XSFILL89080x65050 gnd vdd FILL
XSFILL109400x60050 gnd vdd FILL
XFILL_5__13548_ gnd vdd FILL
XFILL_1__15906_ gnd vdd FILL
XFILL_4__12189_ gnd vdd FILL
XFILL_3__14727_ gnd vdd FILL
XFILL_3__11939_ gnd vdd FILL
XFILL_1__11029_ gnd vdd FILL
XFILL_2__16156_ gnd vdd FILL
X_6954_ _6955_/B _7594_/B gnd _6954_/Y vdd NAND2X1
XFILL_2__13368_ gnd vdd FILL
XFILL_0__14547_ gnd vdd FILL
XSFILL79320x42050 gnd vdd FILL
XFILL_0__9045_ gnd vdd FILL
XSFILL43960x19050 gnd vdd FILL
XFILL_0__11759_ gnd vdd FILL
XSFILL114920x49050 gnd vdd FILL
XFILL_2__15107_ gnd vdd FILL
XFILL_5__16267_ gnd vdd FILL
XSFILL3560x68050 gnd vdd FILL
X_9673_ _9673_/A _9675_/A _9673_/C gnd _9713_/D vdd OAI21X1
XFILL_2__12319_ gnd vdd FILL
XFILL_5__13479_ gnd vdd FILL
X_6885_ _6885_/A gnd memoryWriteData[15] vdd BUFX2
XFILL_1__15837_ gnd vdd FILL
XFILL_3__14658_ gnd vdd FILL
XFILL_2__16087_ gnd vdd FILL
XFILL_2__13299_ gnd vdd FILL
XFILL_0__14478_ gnd vdd FILL
XFILL_5__15218_ gnd vdd FILL
X_8624_ _8609_/A _8624_/B gnd _8624_/Y vdd NAND2X1
XFILL_6__14769_ gnd vdd FILL
XFILL_3__13609_ gnd vdd FILL
XFILL_5__16198_ gnd vdd FILL
XSFILL114520x51050 gnd vdd FILL
XFILL_2__15038_ gnd vdd FILL
XFILL_4__15948_ gnd vdd FILL
XFILL_3__14589_ gnd vdd FILL
XFILL_0__16217_ gnd vdd FILL
XSFILL44040x28050 gnd vdd FILL
XFILL_0__13429_ gnd vdd FILL
XFILL_1__15768_ gnd vdd FILL
XFILL_6__9503_ gnd vdd FILL
XFILL_3__7986_ gnd vdd FILL
XFILL_5_BUFX2_insert803 gnd vdd FILL
XFILL_5_BUFX2_insert814 gnd vdd FILL
XFILL_5__15149_ gnd vdd FILL
X_8555_ _8555_/Q _9963_/CLK _9963_/R vdd _8503_/Y gnd vdd DFFSR
XFILL_3__16328_ gnd vdd FILL
XFILL_5_BUFX2_insert825 gnd vdd FILL
XFILL_3__6937_ gnd vdd FILL
XFILL_1__14719_ gnd vdd FILL
XFILL_3__9725_ gnd vdd FILL
XFILL_4__15879_ gnd vdd FILL
XFILL_5_BUFX2_insert836 gnd vdd FILL
XBUFX2_insert1000 _12399_/Y gnd _7853_/B vdd BUFX2
XFILL_0__16148_ gnd vdd FILL
XFILL_1__15699_ gnd vdd FILL
XBUFX2_insert1011 _13569_/Y gnd _14283_/C vdd BUFX2
XFILL_5_BUFX2_insert847 gnd vdd FILL
XFILL_1__8740_ gnd vdd FILL
XBUFX2_insert1022 _13340_/Y gnd _9639_/A vdd BUFX2
X_7506_ _7504_/Y _7472_/A _7505_/Y gnd _7540_/D vdd OAI21X1
XFILL_5_BUFX2_insert858 gnd vdd FILL
XBUFX2_insert1033 _13333_/Y gnd _9232_/B vdd BUFX2
XFILL_5_BUFX2_insert869 gnd vdd FILL
XBUFX2_insert1044 _13297_/Y gnd _7744_/B vdd BUFX2
X_8486_ _8550_/Q gnd _8488_/A vdd INVX1
XFILL_3__9656_ gnd vdd FILL
XFILL_3__16259_ gnd vdd FILL
XFILL_3__6868_ gnd vdd FILL
XBUFX2_insert1055 _13527_/Y gnd _13751_/B vdd BUFX2
XFILL111800x49050 gnd vdd FILL
XFILL_0__16079_ gnd vdd FILL
XBUFX2_insert1066 _13327_/Y gnd _8859_/A vdd BUFX2
X_7437_ _7435_/Y _7503_/B _7437_/C gnd _7517_/D vdd OAI21X1
XFILL_0__9878_ gnd vdd FILL
XBUFX2_insert1088 rst gnd BUFX2_insert556/A vdd BUFX2
XSFILL49480x8050 gnd vdd FILL
XFILL_3__8607_ gnd vdd FILL
XFILL_4__8380_ gnd vdd FILL
XSFILL63720x34050 gnd vdd FILL
XFILL112440x15050 gnd vdd FILL
XFILL_1__7622_ gnd vdd FILL
XFILL_6__9296_ gnd vdd FILL
XFILL_0__8829_ gnd vdd FILL
XFILL_4__7331_ gnd vdd FILL
X_7368_ _7336_/B _7496_/B gnd _7369_/C vdd NAND2X1
XFILL_6__8247_ gnd vdd FILL
X_9107_ _9105_/Y _9170_/B _9106_/Y gnd _9107_/Y vdd OAI21X1
XFILL_1__7553_ gnd vdd FILL
X_7299_ _7308_/A _9347_/B gnd _7299_/Y vdd NAND2X1
XFILL_3__8469_ gnd vdd FILL
X_9038_ _8961_/B _8910_/B gnd _9039_/C vdd NAND2X1
XFILL_4__9001_ gnd vdd FILL
XFILL_1__7484_ gnd vdd FILL
XFILL_4__7193_ gnd vdd FILL
XSFILL94280x36050 gnd vdd FILL
XSFILL114600x31050 gnd vdd FILL
XFILL_1__9223_ gnd vdd FILL
XFILL_2_BUFX2_insert704 gnd vdd FILL
XFILL_2_BUFX2_insert715 gnd vdd FILL
XFILL_2_BUFX2_insert726 gnd vdd FILL
X_11940_ _11940_/A _11969_/A _11940_/C gnd _6855_/A vdd OAI21X1
XFILL_2_BUFX2_insert737 gnd vdd FILL
XFILL_2_BUFX2_insert748 gnd vdd FILL
XFILL_1__9154_ gnd vdd FILL
XFILL_2_BUFX2_insert759 gnd vdd FILL
XFILL_1__8105_ gnd vdd FILL
X_11871_ _12113_/A _11865_/Y _11871_/C gnd _16450_/B vdd NOR3X1
XSFILL114280x3050 gnd vdd FILL
XFILL_1__9085_ gnd vdd FILL
XFILL_4__9903_ gnd vdd FILL
X_13610_ _13610_/A _13610_/B _13602_/Y gnd _13611_/B vdd NAND3X1
X_10822_ _10822_/A _10822_/B _10821_/Y gnd _10864_/D vdd OAI21X1
X_14590_ _13467_/A _14588_/Y _13850_/B _14589_/Y gnd _14594_/B vdd OAI22X1
X_13541_ _13467_/A gnd _13541_/Y vdd INVX8
XSFILL8760x81050 gnd vdd FILL
X_10753_ _10753_/A _10789_/B _10752_/Y gnd _10841_/D vdd OAI21X1
XSFILL23800x30050 gnd vdd FILL
XBUFX2_insert703 _11985_/Y gnd _12024_/C vdd BUFX2
XBUFX2_insert714 _15023_/Y gnd _15025_/B vdd BUFX2
XSFILL89240x25050 gnd vdd FILL
XBUFX2_insert725 _13352_/Y gnd _10160_/A vdd BUFX2
XFILL_4__9765_ gnd vdd FILL
XBUFX2_insert736 _15020_/Y gnd _15789_/B vdd BUFX2
XFILL_4__6977_ gnd vdd FILL
X_16260_ _9332_/Q _15892_/B _15380_/C _9936_/A gnd _16260_/Y vdd AOI22X1
XFILL_2__7800_ gnd vdd FILL
X_13472_ _13469_/Y _14643_/B _14643_/C _13468_/Y gnd _13473_/A vdd OAI22X1
XBUFX2_insert747 _13344_/Y gnd _9813_/B vdd BUFX2
X_10684_ _10678_/A _9788_/B gnd _10685_/C vdd NAND2X1
XFILL_1__9987_ gnd vdd FILL
XFILL_2__8780_ gnd vdd FILL
XBUFX2_insert758 _12213_/Y gnd _12300_/C vdd BUFX2
XBUFX2_insert769 _13301_/Y gnd _7821_/B vdd BUFX2
XFILL_4__8716_ gnd vdd FILL
X_15211_ _15211_/A _15646_/D gnd _15215_/A vdd NOR2X1
X_12423_ _12423_/A _12359_/A _12423_/C gnd _12423_/Y vdd OAI21X1
X_16191_ _8946_/Q _16037_/B _16037_/C gnd _16191_/Y vdd NAND3X1
XFILL_2__7731_ gnd vdd FILL
XFILL_5__7440_ gnd vdd FILL
X_15142_ _15142_/A _15139_/Y gnd _15142_/Y vdd NOR2X1
XFILL_4__8647_ gnd vdd FILL
X_12354_ _12352_/Y _12368_/A _12353_/Y gnd _12354_/Y vdd OAI21X1
XFILL_1_CLKBUF1_insert130 gnd vdd FILL
XSFILL13720x82050 gnd vdd FILL
XFILL_1__8869_ gnd vdd FILL
XFILL_1_CLKBUF1_insert141 gnd vdd FILL
XFILL_3__10270_ gnd vdd FILL
XFILL_1_CLKBUF1_insert152 gnd vdd FILL
XFILL_5__7371_ gnd vdd FILL
XFILL_4__8578_ gnd vdd FILL
XFILL_1_CLKBUF1_insert163 gnd vdd FILL
X_11305_ _11304_/Y gnd _11597_/A vdd INVX2
X_15073_ _15322_/D _13444_/A _15073_/C gnd _15073_/Y vdd OAI21X1
XFILL_2__9401_ gnd vdd FILL
XFILL_1_CLKBUF1_insert174 gnd vdd FILL
XFILL_4__11560_ gnd vdd FILL
X_12285_ _6887_/A _12237_/B _12269_/C _12308_/B gnd _12286_/C vdd AOI22X1
XFILL_1_CLKBUF1_insert185 gnd vdd FILL
XFILL_1__10400_ gnd vdd FILL
XFILL_5__9110_ gnd vdd FILL
XFILL_1_CLKBUF1_insert196 gnd vdd FILL
XFILL_2__7593_ gnd vdd FILL
XFILL_1__11380_ gnd vdd FILL
XSFILL94200x80050 gnd vdd FILL
X_14024_ _14024_/A _14024_/B _15651_/C gnd _12985_/B vdd AOI21X1
XFILL_4__10511_ gnd vdd FILL
XFILL_2_BUFX2_insert6 gnd vdd FILL
XSFILL109400x4050 gnd vdd FILL
X_11236_ _12230_/Y _12126_/Y gnd _11236_/Y vdd NOR2X1
XFILL_5__12850_ gnd vdd FILL
XFILL_4__11491_ gnd vdd FILL
XFILL_5__9041_ gnd vdd FILL
XFILL_4__13230_ gnd vdd FILL
XFILL_5__11801_ gnd vdd FILL
XFILL_4__10442_ gnd vdd FILL
XSFILL104600x63050 gnd vdd FILL
X_11167_ _12195_/Y _12322_/Y gnd _11167_/Y vdd NAND2X1
XFILL_5__12781_ gnd vdd FILL
XFILL_2__9263_ gnd vdd FILL
XFILL_2__11621_ gnd vdd FILL
XFILL_3__13960_ gnd vdd FILL
XFILL_1__10262_ gnd vdd FILL
XFILL_3_BUFX2_insert560 gnd vdd FILL
XFILL_0__13780_ gnd vdd FILL
XFILL_5__14520_ gnd vdd FILL
XFILL_3_BUFX2_insert571 gnd vdd FILL
XFILL_0__10992_ gnd vdd FILL
X_10118_ _10106_/A _9478_/B gnd _10119_/C vdd NAND2X1
XFILL_3_BUFX2_insert582 gnd vdd FILL
XFILL_4__13161_ gnd vdd FILL
XFILL_2__8214_ gnd vdd FILL
XFILL_5__11732_ gnd vdd FILL
X_15975_ _15974_/Y _15972_/Y gnd _15975_/Y vdd NOR2X1
XFILL_3__12911_ gnd vdd FILL
XFILL_1__12001_ gnd vdd FILL
XFILL_2__14340_ gnd vdd FILL
X_11098_ _12183_/Y _12306_/Y gnd _11290_/A vdd NOR2X1
XFILL_4__10373_ gnd vdd FILL
XFILL_3_BUFX2_insert593 gnd vdd FILL
XFILL_3__13891_ gnd vdd FILL
XFILL_2__11552_ gnd vdd FILL
XFILL_0__12731_ gnd vdd FILL
XFILL_1__10193_ gnd vdd FILL
XSFILL19080x60050 gnd vdd FILL
XFILL_4__12112_ gnd vdd FILL
XFILL_5__14451_ gnd vdd FILL
X_10049_ _14660_/A gnd _10051_/A vdd INVX1
X_14926_ _8436_/Q _13647_/B _14926_/C _6992_/A gnd _14927_/B vdd AOI22X1
XFILL_3__12842_ gnd vdd FILL
XFILL_3__15630_ gnd vdd FILL
XFILL_4__13092_ gnd vdd FILL
XFILL_5__11663_ gnd vdd FILL
XFILL_2__10503_ gnd vdd FILL
XFILL_2__8145_ gnd vdd FILL
XFILL_2__14271_ gnd vdd FILL
XFILL_0__12662_ gnd vdd FILL
XFILL_0__15450_ gnd vdd FILL
XFILL_2__11483_ gnd vdd FILL
XFILL_5__13402_ gnd vdd FILL
XFILL_6__15741_ gnd vdd FILL
XFILL_2__16010_ gnd vdd FILL
XFILL_0__7160_ gnd vdd FILL
XFILL_5__10614_ gnd vdd FILL
XFILL_4__12043_ gnd vdd FILL
XFILL_2__13222_ gnd vdd FILL
X_14857_ _14857_/A _14857_/B gnd _14858_/C vdd NOR2X1
XFILL_3__15561_ gnd vdd FILL
XFILL_5__14382_ gnd vdd FILL
XFILL_3__12773_ gnd vdd FILL
XFILL_2__8076_ gnd vdd FILL
XFILL_0__14401_ gnd vdd FILL
XFILL_2__10434_ gnd vdd FILL
XFILL_5__11594_ gnd vdd FILL
XFILL_0__11613_ gnd vdd FILL
XFILL_1__13952_ gnd vdd FILL
XFILL_0__12593_ gnd vdd FILL
XFILL_0__15381_ gnd vdd FILL
XFILL_5__16121_ gnd vdd FILL
XFILL_5__13333_ gnd vdd FILL
X_13808_ _10205_/Q gnd _13808_/Y vdd INVX1
XSFILL13800x62050 gnd vdd FILL
XFILL_5__9874_ gnd vdd FILL
XFILL_3__14512_ gnd vdd FILL
XFILL_5__10545_ gnd vdd FILL
XFILL_0__7091_ gnd vdd FILL
XFILL_3__11724_ gnd vdd FILL
X_14788_ _14788_/A _14788_/B gnd _14789_/B vdd NOR2X1
XFILL_2__13153_ gnd vdd FILL
XSFILL79240x57050 gnd vdd FILL
XFILL_1__12903_ gnd vdd FILL
XFILL_3__15492_ gnd vdd FILL
XFILL_6_BUFX2_insert75 gnd vdd FILL
XFILL_0__14332_ gnd vdd FILL
XFILL_0__11544_ gnd vdd FILL
XFILL_2__10365_ gnd vdd FILL
XFILL_1__13883_ gnd vdd FILL
XFILL_6_BUFX2_insert86 gnd vdd FILL
XFILL_5__8825_ gnd vdd FILL
XFILL_4__15802_ gnd vdd FILL
XFILL_5__16052_ gnd vdd FILL
X_13739_ _13714_/Y _13739_/B _15812_/C gnd _12967_/B vdd AOI21X1
XFILL_6__11835_ gnd vdd FILL
XFILL_5__13264_ gnd vdd FILL
XFILL_2__12104_ gnd vdd FILL
XFILL_3__14443_ gnd vdd FILL
XFILL_3__7840_ gnd vdd FILL
XFILL_1__15622_ gnd vdd FILL
XFILL_3__11655_ gnd vdd FILL
XFILL_1__12834_ gnd vdd FILL
XFILL_4__13994_ gnd vdd FILL
XFILL_2__13084_ gnd vdd FILL
XFILL_0__14263_ gnd vdd FILL
XFILL_5__15003_ gnd vdd FILL
XFILL_2__10296_ gnd vdd FILL
XFILL_0__11475_ gnd vdd FILL
XFILL_6__14554_ gnd vdd FILL
XSFILL114440x66050 gnd vdd FILL
XFILL_5__12215_ gnd vdd FILL
XFILL_5__8756_ gnd vdd FILL
XFILL_4__15733_ gnd vdd FILL
XFILL_0__16002_ gnd vdd FILL
XFILL_2__12035_ gnd vdd FILL
XFILL_3__14374_ gnd vdd FILL
XFILL_0__13214_ gnd vdd FILL
XFILL_1__15553_ gnd vdd FILL
XFILL_0__10426_ gnd vdd FILL
XFILL_3__11586_ gnd vdd FILL
XFILL_2__8978_ gnd vdd FILL
XFILL_1__12765_ gnd vdd FILL
XFILL_0__14194_ gnd vdd FILL
XSFILL84360x48050 gnd vdd FILL
XFILL_5__7707_ gnd vdd FILL
XFILL_0_BUFX2_insert450 gnd vdd FILL
XFILL_0__9801_ gnd vdd FILL
XFILL_6__13505_ gnd vdd FILL
X_15409_ _8542_/Q gnd _15409_/Y vdd INVX1
XFILL_0_BUFX2_insert461 gnd vdd FILL
XSFILL48920x4050 gnd vdd FILL
XFILL_3__13325_ gnd vdd FILL
X_16389_ _16387_/Y gnd _16389_/C gnd _16389_/Y vdd OAI21X1
XFILL_3__9510_ gnd vdd FILL
XFILL_3__16113_ gnd vdd FILL
XFILL_0_BUFX2_insert472 gnd vdd FILL
X_8340_ _8340_/A gnd _8342_/A vdd INVX1
XFILL_5__12146_ gnd vdd FILL
XFILL_4__15664_ gnd vdd FILL
XFILL_0__7993_ gnd vdd FILL
XFILL_1__14504_ gnd vdd FILL
XFILL_6__11697_ gnd vdd FILL
XFILL_3__10537_ gnd vdd FILL
XFILL_0__13145_ gnd vdd FILL
XFILL_0_BUFX2_insert483 gnd vdd FILL
XFILL_4__12876_ gnd vdd FILL
XFILL_1__11716_ gnd vdd FILL
XFILL_2__7929_ gnd vdd FILL
XFILL_0_BUFX2_insert494 gnd vdd FILL
XFILL_1__15484_ gnd vdd FILL
XSFILL59160x24050 gnd vdd FILL
XFILL_1__12696_ gnd vdd FILL
XFILL_0__9732_ gnd vdd FILL
X_8271_ _8271_/A _8249_/A _8271_/C gnd _8307_/D vdd OAI21X1
XFILL_3__16044_ gnd vdd FILL
XFILL_4__14615_ gnd vdd FILL
XFILL_0__6944_ gnd vdd FILL
XFILL_5__12077_ gnd vdd FILL
XFILL_3__13256_ gnd vdd FILL
XFILL_4__11827_ gnd vdd FILL
XFILL_1__14435_ gnd vdd FILL
XFILL_4__15595_ gnd vdd FILL
XFILL_2__13986_ gnd vdd FILL
XFILL_1__11647_ gnd vdd FILL
XFILL_5__15905_ gnd vdd FILL
XFILL_0__10288_ gnd vdd FILL
XFILL_5__7569_ gnd vdd FILL
XFILL_5__11028_ gnd vdd FILL
XFILL_6__16155_ gnd vdd FILL
X_7222_ _7181_/B _7222_/B gnd _7222_/Y vdd NAND2X1
XFILL_0__9663_ gnd vdd FILL
XFILL_6__13367_ gnd vdd FILL
XFILL_3__12207_ gnd vdd FILL
XFILL_4__14546_ gnd vdd FILL
XFILL_0__6875_ gnd vdd FILL
XFILL_6__10579_ gnd vdd FILL
XFILL_2__15725_ gnd vdd FILL
XFILL_3__9372_ gnd vdd FILL
XFILL_0__12027_ gnd vdd FILL
XFILL_4__11758_ gnd vdd FILL
XFILL_1__14366_ gnd vdd FILL
XFILL_3__10399_ gnd vdd FILL
XFILL_6__15106_ gnd vdd FILL
XFILL_0__8614_ gnd vdd FILL
XFILL_1__11578_ gnd vdd FILL
XFILL_5__15836_ gnd vdd FILL
X_7153_ _7153_/Q _7786_/CLK _7153_/R vdd _7153_/D gnd vdd DFFSR
XFILL_3__8323_ gnd vdd FILL
XFILL_3__12138_ gnd vdd FILL
XSFILL109400x55050 gnd vdd FILL
XFILL_1__16105_ gnd vdd FILL
XFILL_4__10709_ gnd vdd FILL
XFILL_0__9594_ gnd vdd FILL
XFILL_1__13317_ gnd vdd FILL
XFILL_4__14477_ gnd vdd FILL
XFILL_2__15656_ gnd vdd FILL
XFILL_4__11689_ gnd vdd FILL
XFILL_1__10529_ gnd vdd FILL
XFILL_2__12868_ gnd vdd FILL
XCLKBUF1_insert140 CLKBUF1_insert216/A gnd _7534_/CLK vdd CLKBUF1
XFILL_5__9239_ gnd vdd FILL
XFILL_1__14297_ gnd vdd FILL
XFILL_4__16216_ gnd vdd FILL
XSFILL79320x37050 gnd vdd FILL
XFILL_6__12249_ gnd vdd FILL
XCLKBUF1_insert151 CLKBUF1_insert150/A gnd _8433_/CLK vdd CLKBUF1
XSFILL49080x76050 gnd vdd FILL
XFILL_2__14607_ gnd vdd FILL
XFILL_4__13428_ gnd vdd FILL
X_7084_ _7084_/A gnd _7084_/Y vdd INVX1
XFILL_5__15767_ gnd vdd FILL
XFILL_3__8254_ gnd vdd FILL
XFILL_1__16036_ gnd vdd FILL
XCLKBUF1_insert162 CLKBUF1_insert216/A gnd _8165_/CLK vdd CLKBUF1
XFILL_3__12069_ gnd vdd FILL
XFILL_5__12979_ gnd vdd FILL
XFILL_2__11819_ gnd vdd FILL
XFILL_1__13248_ gnd vdd FILL
XCLKBUF1_insert173 CLKBUF1_insert218/A gnd _9707_/CLK vdd CLKBUF1
XFILL_2__15587_ gnd vdd FILL
XCLKBUF1_insert184 CLKBUF1_insert187/A gnd _13201_/CLK vdd CLKBUF1
XCLKBUF1_insert195 CLKBUF1_insert218/A gnd _7915_/CLK vdd CLKBUF1
XFILL_0__13978_ gnd vdd FILL
XFILL_5__14718_ gnd vdd FILL
XFILL_3__7205_ gnd vdd FILL
XFILL_0__8476_ gnd vdd FILL
XFILL_4__16147_ gnd vdd FILL
XFILL_4__13359_ gnd vdd FILL
XFILL_5__15698_ gnd vdd FILL
XFILL_2__14538_ gnd vdd FILL
XFILL_0__15717_ gnd vdd FILL
XFILL_3__8185_ gnd vdd FILL
XFILL_0__7427_ gnd vdd FILL
XFILL_5__14649_ gnd vdd FILL
XFILL_3__15828_ gnd vdd FILL
XFILL_4__16078_ gnd vdd FILL
XFILL_2__14469_ gnd vdd FILL
XFILL_0__15648_ gnd vdd FILL
XFILL_2__16208_ gnd vdd FILL
XFILL_0__7358_ gnd vdd FILL
XFILL_4__15029_ gnd vdd FILL
XFILL_3__7067_ gnd vdd FILL
XFILL_3__15759_ gnd vdd FILL
X_7986_ _8042_/Q gnd _7988_/A vdd INVX1
XFILL_5__16319_ gnd vdd FILL
XFILL_0__15579_ gnd vdd FILL
X_9725_ _9813_/B _7037_/B gnd _9725_/Y vdd NAND2X1
X_6937_ _6935_/Y _6937_/B _6937_/C gnd _7009_/D vdd OAI21X1
XFILL_2__16139_ gnd vdd FILL
XFILL_0__7289_ gnd vdd FILL
XFILL_4__6900_ gnd vdd FILL
XFILL_4__7880_ gnd vdd FILL
XFILL_0__9028_ gnd vdd FILL
XFILL_1__9910_ gnd vdd FILL
X_9656_ _9708_/Q gnd _9658_/A vdd INVX1
XSFILL23720x45050 gnd vdd FILL
X_6868_ _6868_/A gnd memoryAddress[30] vdd BUFX2
X_8607_ _8607_/A _8607_/B _8606_/Y gnd _8675_/D vdd OAI21X1
XFILL112040x12050 gnd vdd FILL
XFILL_5_BUFX2_insert600 gnd vdd FILL
X_9587_ _9587_/Q _8051_/CLK _8051_/R vdd _9587_/D gnd vdd DFFSR
XFILL_4__9550_ gnd vdd FILL
XFILL_5_BUFX2_insert611 gnd vdd FILL
XFILL_5_BUFX2_insert622 gnd vdd FILL
XFILL_5_BUFX2_insert633 gnd vdd FILL
XFILL_3__7969_ gnd vdd FILL
XFILL_1__9772_ gnd vdd FILL
X_8538_ _8450_/A _8541_/CLK _8285_/R vdd _8452_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert644 gnd vdd FILL
XFILL_4__8501_ gnd vdd FILL
XFILL_5_BUFX2_insert655 gnd vdd FILL
XFILL_1__6984_ gnd vdd FILL
XFILL_4__9481_ gnd vdd FILL
XFILL_5_BUFX2_insert666 gnd vdd FILL
XFILL_5_BUFX2_insert677 gnd vdd FILL
XFILL_5_BUFX2_insert688 gnd vdd FILL
XFILL_1__8723_ gnd vdd FILL
XSFILL114600x26050 gnd vdd FILL
XFILL_5_BUFX2_insert699 gnd vdd FILL
X_8469_ _8469_/A _7061_/B gnd _8470_/C vdd NAND2X1
XFILL_3__9639_ gnd vdd FILL
XFILL_6__9348_ gnd vdd FILL
XFILL_1__8654_ gnd vdd FILL
XFILL_4__8363_ gnd vdd FILL
XFILL_1__7605_ gnd vdd FILL
X_12070_ _12070_/A _12070_/B _12069_/Y gnd _13140_/B vdd NAND3X1
XFILL_2_CLKBUF1_insert203 gnd vdd FILL
XFILL_1__8585_ gnd vdd FILL
XFILL_2_CLKBUF1_insert214 gnd vdd FILL
XFILL_4__7314_ gnd vdd FILL
X_11021_ _11383_/A _11018_/Y _11019_/Y _11020_/Y gnd _11021_/Y vdd OAI22X1
XSFILL104520x78050 gnd vdd FILL
XFILL_4__7245_ gnd vdd FILL
XSFILL23800x25050 gnd vdd FILL
XFILL_1__7467_ gnd vdd FILL
XFILL_2_BUFX2_insert501 gnd vdd FILL
XFILL_4__7176_ gnd vdd FILL
XSFILL33160x50050 gnd vdd FILL
XFILL_2_BUFX2_insert512 gnd vdd FILL
XFILL_2_BUFX2_insert523 gnd vdd FILL
XFILL_1__9206_ gnd vdd FILL
X_15760_ _15760_/A _15760_/B _15760_/C gnd _15762_/A vdd OAI21X1
X_12972_ _6877_/A gnd _12972_/Y vdd INVX1
XFILL_2_BUFX2_insert534 gnd vdd FILL
XFILL_2_BUFX2_insert545 gnd vdd FILL
XFILL_2_BUFX2_insert556 gnd vdd FILL
XFILL_2_BUFX2_insert567 gnd vdd FILL
X_11923_ _12151_/A gnd _11925_/A vdd INVX1
X_14711_ _14711_/A _14711_/B gnd _14711_/Y vdd NOR2X1
XFILL_2_BUFX2_insert578 gnd vdd FILL
X_15691_ _15691_/A _15691_/B _14265_/C gnd _12869_/B vdd AOI21X1
XFILL_1__9137_ gnd vdd FILL
XFILL_2_BUFX2_insert589 gnd vdd FILL
XFILL_5__6940_ gnd vdd FILL
X_14642_ _8638_/A gnd _14642_/Y vdd INVX1
XSFILL74280x5050 gnd vdd FILL
X_11854_ _12467_/B _11853_/Y gnd _11855_/B vdd NOR2X1
XFILL_6_BUFX2_insert1042 gnd vdd FILL
XSFILL13720x77050 gnd vdd FILL
XFILL_6_BUFX2_insert1053 gnd vdd FILL
X_10805_ _10859_/Q gnd _10805_/Y vdd INVX1
XFILL_5__6871_ gnd vdd FILL
X_14573_ _9709_/Q gnd _14573_/Y vdd INVX1
XFILL_1__8019_ gnd vdd FILL
X_11785_ _11785_/A gnd _11787_/A vdd INVX1
XFILL_2__8901_ gnd vdd FILL
XFILL_2__10150_ gnd vdd FILL
XFILL_2__9881_ gnd vdd FILL
XBUFX2_insert500 BUFX2_insert556/A gnd _8688_/R vdd BUFX2
XBUFX2_insert511 BUFX2_insert559/A gnd _7150_/R vdd BUFX2
XFILL_5__8610_ gnd vdd FILL
XFILL_5__9590_ gnd vdd FILL
XFILL_1__10880_ gnd vdd FILL
X_16312_ _16311_/Y _16312_/B gnd _16312_/Y vdd NOR2X1
XFILL_6__11620_ gnd vdd FILL
X_13524_ _7673_/A gnd _13524_/Y vdd INVX1
XBUFX2_insert522 BUFX2_insert607/A gnd _7644_/R vdd BUFX2
X_10736_ _10736_/Q _7268_/CLK _8688_/R vdd _10694_/Y gnd vdd DFFSR
XFILL112040x5050 gnd vdd FILL
XFILL_5__10261_ gnd vdd FILL
XFILL_2__8832_ gnd vdd FILL
XSFILL113880x74050 gnd vdd FILL
XBUFX2_insert533 BUFX2_insert600/A gnd _7140_/R vdd BUFX2
XFILL_3__11440_ gnd vdd FILL
XBUFX2_insert544 BUFX2_insert607/A gnd _8674_/R vdd BUFX2
XFILL_4__10991_ gnd vdd FILL
XBUFX2_insert555 BUFX2_insert496/A gnd _9944_/R vdd BUFX2
XFILL_0__11260_ gnd vdd FILL
X_16243_ _16243_/A _16243_/B _16231_/Y gnd _16244_/B vdd NOR3X1
XBUFX2_insert566 BUFX2_insert570/A gnd _9050_/R vdd BUFX2
XFILL_5__12000_ gnd vdd FILL
XFILL_4__9748_ gnd vdd FILL
X_13455_ _13443_/A _13404_/B _13407_/Y gnd _13455_/Y vdd NAND3X1
XFILL_4__12730_ gnd vdd FILL
XBUFX2_insert577 BUFX2_insert607/A gnd _9046_/R vdd BUFX2
X_10667_ _10665_/Y _10615_/B _10667_/C gnd _10667_/Y vdd OAI21X1
XFILL_5__10192_ gnd vdd FILL
XFILL_2__8763_ gnd vdd FILL
XBUFX2_insert588 BUFX2_insert600/A gnd _7152_/R vdd BUFX2
XFILL_3__11371_ gnd vdd FILL
XBUFX2_insert599 BUFX2_insert520/A gnd _7274_/R vdd BUFX2
X_12406_ _12406_/A gnd _12406_/Y vdd INVX1
XFILL_5__8472_ gnd vdd FILL
XFILL_6__10502_ gnd vdd FILL
XFILL_0__11191_ gnd vdd FILL
XFILL_4__9679_ gnd vdd FILL
X_16174_ _16174_/A _15920_/B _15328_/B _14825_/Y gnd _16175_/C vdd OAI22X1
XFILL_3__13110_ gnd vdd FILL
X_13386_ _13372_/A gnd _13423_/A vdd INVX4
XFILL_2__7714_ gnd vdd FILL
XFILL_3__10322_ gnd vdd FILL
XFILL_6__11482_ gnd vdd FILL
XFILL_4__12661_ gnd vdd FILL
X_10598_ _10534_/A _8038_/CLK _7789_/R vdd _10536_/Y gnd vdd DFFSR
XFILL_2__13840_ gnd vdd FILL
XSFILL59080x39050 gnd vdd FILL
XFILL_3__14090_ gnd vdd FILL
XFILL_1__11501_ gnd vdd FILL
XFILL_5__7423_ gnd vdd FILL
XFILL_2__8694_ gnd vdd FILL
XFILL_0__10142_ gnd vdd FILL
XFILL_1__12481_ gnd vdd FILL
X_15125_ _15119_/Y _15125_/B gnd _15126_/A vdd NAND2X1
XFILL_4__14400_ gnd vdd FILL
X_12337_ _6900_/A _12289_/B _12289_/C _12297_/D gnd _12338_/C vdd AOI22X1
XSFILL74120x42050 gnd vdd FILL
XFILL_4_BUFX2_insert1090 gnd vdd FILL
XFILL_4__11612_ gnd vdd FILL
XFILL_5__13951_ gnd vdd FILL
XFILL_3__13041_ gnd vdd FILL
XFILL_4__12592_ gnd vdd FILL
XFILL_3__10253_ gnd vdd FILL
XFILL_4__15380_ gnd vdd FILL
XFILL_1__14220_ gnd vdd FILL
XFILL_2__13771_ gnd vdd FILL
XFILL_1__11432_ gnd vdd FILL
XFILL_2__10983_ gnd vdd FILL
XFILL_5__7354_ gnd vdd FILL
XFILL_0__14950_ gnd vdd FILL
X_15056_ _15056_/A _15378_/B _15376_/B _13468_/Y gnd _15057_/A vdd OAI22X1
XFILL_5__12902_ gnd vdd FILL
XFILL_2__15510_ gnd vdd FILL
X_12268_ _12248_/A _11879_/B _12248_/C gnd _12270_/B vdd NAND3X1
XFILL_4__14331_ gnd vdd FILL
XFILL_4__11543_ gnd vdd FILL
XFILL_5__13882_ gnd vdd FILL
XFILL_2__12722_ gnd vdd FILL
XFILL_1__14151_ gnd vdd FILL
XFILL_2__7576_ gnd vdd FILL
XFILL_3__10184_ gnd vdd FILL
XFILL_0__13901_ gnd vdd FILL
X_14007_ _14007_/A _14479_/B _13587_/A _15498_/B gnd _14011_/A vdd OAI22X1
XFILL_1__11363_ gnd vdd FILL
XFILL_0__14881_ gnd vdd FILL
XFILL_5__15621_ gnd vdd FILL
X_11219_ _11220_/A _11220_/B _11762_/B gnd _11219_/Y vdd AOI21X1
XFILL_5__12833_ gnd vdd FILL
XSFILL13800x57050 gnd vdd FILL
XFILL_6__10295_ gnd vdd FILL
XFILL_4__14262_ gnd vdd FILL
XFILL_1__13102_ gnd vdd FILL
X_12199_ _11971_/A gnd _12201_/A vdd INVX1
XFILL_4__11474_ gnd vdd FILL
XFILL_2__15441_ gnd vdd FILL
XFILL_2__12653_ gnd vdd FILL
XFILL_1__10314_ gnd vdd FILL
XFILL_5__9024_ gnd vdd FILL
XFILL_0__13832_ gnd vdd FILL
XFILL_3__14992_ gnd vdd FILL
XFILL_1__11294_ gnd vdd FILL
XFILL_1__14082_ gnd vdd FILL
XFILL_4__16001_ gnd vdd FILL
XFILL_0__8330_ gnd vdd FILL
XFILL_6__12034_ gnd vdd FILL
XFILL_4__13213_ gnd vdd FILL
XFILL_5__15552_ gnd vdd FILL
XFILL_4__10425_ gnd vdd FILL
XFILL_5__12764_ gnd vdd FILL
XFILL_4__14193_ gnd vdd FILL
XFILL_2__11604_ gnd vdd FILL
XFILL_2__9246_ gnd vdd FILL
XFILL_2__15372_ gnd vdd FILL
XFILL_1__10245_ gnd vdd FILL
XFILL_3__13943_ gnd vdd FILL
XFILL_1__13033_ gnd vdd FILL
XFILL_2__12584_ gnd vdd FILL
XFILL_3_BUFX2_insert390 gnd vdd FILL
XFILL_0__13763_ gnd vdd FILL
XFILL_5__14503_ gnd vdd FILL
XFILL_0__10975_ gnd vdd FILL
XFILL_4__13144_ gnd vdd FILL
XFILL_0__8261_ gnd vdd FILL
XFILL_5__11715_ gnd vdd FILL
X_15958_ _15957_/Y _15958_/B _15369_/A _14541_/Y gnd _15959_/A vdd OAI22X1
XFILL_2__14323_ gnd vdd FILL
XFILL_5__15483_ gnd vdd FILL
XFILL_5__12695_ gnd vdd FILL
XFILL_2__11535_ gnd vdd FILL
XFILL_0__15502_ gnd vdd FILL
XFILL_0__12714_ gnd vdd FILL
XFILL_1__10176_ gnd vdd FILL
XFILL_3__13874_ gnd vdd FILL
XFILL_0__7212_ gnd vdd FILL
XFILL_0__13694_ gnd vdd FILL
X_14909_ _7376_/A _14738_/A _14909_/C _7156_/Q gnd _14909_/Y vdd AOI22X1
XFILL_5__14434_ gnd vdd FILL
XFILL_0__8192_ gnd vdd FILL
XFILL_2__8128_ gnd vdd FILL
XFILL_3__15613_ gnd vdd FILL
XSFILL43880x52050 gnd vdd FILL
X_7840_ _7840_/A gnd _7842_/A vdd INVX1
XFILL_5__11646_ gnd vdd FILL
XFILL_2__14254_ gnd vdd FILL
XFILL_3__12825_ gnd vdd FILL
XFILL_4__10287_ gnd vdd FILL
X_15889_ _15882_/Y _15888_/Y gnd _15889_/Y vdd NAND2X1
XFILL_0__15433_ gnd vdd FILL
XFILL_2__11466_ gnd vdd FILL
XFILL_0__12645_ gnd vdd FILL
XFILL_1__14984_ gnd vdd FILL
XFILL_5__9926_ gnd vdd FILL
XFILL_3__9990_ gnd vdd FILL
XSFILL59160x19050 gnd vdd FILL
XFILL_4__12026_ gnd vdd FILL
XFILL_5__14365_ gnd vdd FILL
XFILL_3__12756_ gnd vdd FILL
XFILL_3__15544_ gnd vdd FILL
XFILL_2__10417_ gnd vdd FILL
XFILL_2__8059_ gnd vdd FILL
XFILL_5__11577_ gnd vdd FILL
X_7771_ _7771_/Q _8663_/CLK _7131_/R vdd _7771_/D gnd vdd DFFSR
XFILL_2__14185_ gnd vdd FILL
XFILL_1__13935_ gnd vdd FILL
XFILL_0__15364_ gnd vdd FILL
XFILL_5__16104_ gnd vdd FILL
XFILL_2__11397_ gnd vdd FILL
XSFILL74200x22050 gnd vdd FILL
XFILL_5__13316_ gnd vdd FILL
XFILL_0__12576_ gnd vdd FILL
XFILL_5__9857_ gnd vdd FILL
XFILL_6__8650_ gnd vdd FILL
X_9510_ _9574_/Q gnd _9512_/A vdd INVX1
XFILL_0__7074_ gnd vdd FILL
XFILL_5__10528_ gnd vdd FILL
XFILL_6__12867_ gnd vdd FILL
XFILL_3__11707_ gnd vdd FILL
XFILL_2__13136_ gnd vdd FILL
XFILL_5__14296_ gnd vdd FILL
XFILL_3__8872_ gnd vdd FILL
XFILL_0__14315_ gnd vdd FILL
XFILL_3__15475_ gnd vdd FILL
XFILL_1__13866_ gnd vdd FILL
XFILL_0__11527_ gnd vdd FILL
XFILL_6__7601_ gnd vdd FILL
XSFILL59000x83050 gnd vdd FILL
XFILL_5__16035_ gnd vdd FILL
XFILL_0__15295_ gnd vdd FILL
XFILL_5__9788_ gnd vdd FILL
XFILL_5__13247_ gnd vdd FILL
X_9441_ _9367_/A _9188_/CLK _9441_/R vdd _9441_/D gnd vdd DFFSR
XFILL_3__11638_ gnd vdd FILL
XFILL_1__15605_ gnd vdd FILL
XFILL_3__14426_ gnd vdd FILL
XFILL_3__7823_ gnd vdd FILL
XFILL_4_CLKBUF1_insert180 gnd vdd FILL
XFILL_4__13977_ gnd vdd FILL
XFILL_4_CLKBUF1_insert191 gnd vdd FILL
XFILL_0__14246_ gnd vdd FILL
XFILL_2__10279_ gnd vdd FILL
XFILL_0__11458_ gnd vdd FILL
XFILL_5__8739_ gnd vdd FILL
XFILL_1__13797_ gnd vdd FILL
XFILL_4__15716_ gnd vdd FILL
XSFILL3560x50 gnd vdd FILL
XFILL_2__12018_ gnd vdd FILL
X_9372_ _9370_/Y _9372_/B _9371_/Y gnd _9372_/Y vdd OAI21X1
XFILL_3__14357_ gnd vdd FILL
XFILL_3__7754_ gnd vdd FILL
XFILL_1__15536_ gnd vdd FILL
XFILL_0__10409_ gnd vdd FILL
XFILL_3__11569_ gnd vdd FILL
XFILL_1__12748_ gnd vdd FILL
XFILL_0_BUFX2_insert280 gnd vdd FILL
XSFILL109000x52050 gnd vdd FILL
XSFILL38840x41050 gnd vdd FILL
XFILL_0__14177_ gnd vdd FILL
XFILL_0__11389_ gnd vdd FILL
XFILL_0_BUFX2_insert291 gnd vdd FILL
XSFILL64120x74050 gnd vdd FILL
X_8323_ _8333_/B _9859_/B gnd _8324_/C vdd NAND2X1
XFILL_5__12129_ gnd vdd FILL
XFILL_0__7976_ gnd vdd FILL
XFILL_3__13308_ gnd vdd FILL
XFILL_4__15647_ gnd vdd FILL
XFILL_4_BUFX2_insert607 gnd vdd FILL
XFILL_4__12859_ gnd vdd FILL
XFILL_3__14288_ gnd vdd FILL
XFILL_0__13128_ gnd vdd FILL
XFILL_1__15467_ gnd vdd FILL
XFILL_3__7685_ gnd vdd FILL
XFILL_4_BUFX2_insert618 gnd vdd FILL
XFILL_4_BUFX2_insert629 gnd vdd FILL
XFILL_0__6927_ gnd vdd FILL
X_8254_ _8254_/A gnd _8254_/Y vdd INVX1
XFILL_3__13239_ gnd vdd FILL
XFILL_3__16027_ gnd vdd FILL
XFILL_1__14418_ gnd vdd FILL
XFILL_4__15578_ gnd vdd FILL
XFILL_3__9424_ gnd vdd FILL
XFILL_2__13969_ gnd vdd FILL
XFILL_1__15398_ gnd vdd FILL
X_7205_ _7203_/Y _7184_/B _7205_/C gnd _7269_/D vdd OAI21X1
XFILL_0__9646_ gnd vdd FILL
XSFILL3560x81050 gnd vdd FILL
XFILL_0__6858_ gnd vdd FILL
XFILL_4__14529_ gnd vdd FILL
XFILL_2_BUFX2_insert40 gnd vdd FILL
XSFILL68760x77050 gnd vdd FILL
XFILL_3__9355_ gnd vdd FILL
XFILL_2__15708_ gnd vdd FILL
X_8185_ _8185_/A gnd _8185_/Y vdd INVX1
XFILL_2_BUFX2_insert51 gnd vdd FILL
XFILL_1__14349_ gnd vdd FILL
XFILL_2_BUFX2_insert62 gnd vdd FILL
XFILL_2_BUFX2_insert73 gnd vdd FILL
XFILL_5__15819_ gnd vdd FILL
X_7136_ _7060_/A _9578_/CLK _9460_/R vdd _7136_/D gnd vdd DFFSR
XFILL_1__8370_ gnd vdd FILL
XFILL_2_BUFX2_insert84 gnd vdd FILL
XSFILL44040x41050 gnd vdd FILL
XFILL_2_BUFX2_insert95 gnd vdd FILL
XFILL_2__15639_ gnd vdd FILL
XFILL_3__9286_ gnd vdd FILL
XFILL_1__7321_ gnd vdd FILL
XFILL_0__8528_ gnd vdd FILL
X_7067_ _7067_/A _8091_/B gnd _7067_/Y vdd NAND2X1
XSFILL33960x50 gnd vdd FILL
XFILL_1__16019_ gnd vdd FILL
XFILL_4__7030_ gnd vdd FILL
XFILL_3__8237_ gnd vdd FILL
XFILL_0__8459_ gnd vdd FILL
XFILL_1__7252_ gnd vdd FILL
XSFILL18840x8050 gnd vdd FILL
XFILL111800x62050 gnd vdd FILL
XFILL_1__7183_ gnd vdd FILL
XFILL_3__7119_ gnd vdd FILL
XSFILL38920x21050 gnd vdd FILL
XFILL_1_BUFX2_insert508 gnd vdd FILL
XFILL_3__8099_ gnd vdd FILL
XSFILL64200x54050 gnd vdd FILL
XFILL_1_BUFX2_insert519 gnd vdd FILL
XFILL_4__8981_ gnd vdd FILL
X_7969_ _7970_/B _8225_/B gnd _7970_/C vdd NAND2X1
XFILL_4__7932_ gnd vdd FILL
XSFILL39000x30050 gnd vdd FILL
XSFILL27960x45050 gnd vdd FILL
X_9708_ _9708_/Q _7916_/CLK _9964_/R vdd _9708_/D gnd vdd DFFSR
XFILL_4__7863_ gnd vdd FILL
XSFILL3640x61050 gnd vdd FILL
X_11570_ _11570_/A gnd _11570_/Y vdd INVX1
X_9639_ _9639_/A _7847_/B gnd _9640_/C vdd NAND2X1
XFILL_6__8779_ gnd vdd FILL
XFILL_4__9602_ gnd vdd FILL
XSFILL28840x73050 gnd vdd FILL
X_10521_ _10521_/A _10500_/B _10520_/Y gnd _10521_/Y vdd OAI21X1
XFILL_5_BUFX2_insert430 gnd vdd FILL
XFILL_5_BUFX2_insert441 gnd vdd FILL
XFILL_4__9533_ gnd vdd FILL
XFILL_5_BUFX2_insert452 gnd vdd FILL
X_13240_ _13289_/B _13235_/C gnd _13240_/Y vdd NAND2X1
XFILL_5_BUFX2_insert463 gnd vdd FILL
X_10452_ _10395_/A _7380_/B gnd _10452_/Y vdd NAND2X1
XSFILL3480x8050 gnd vdd FILL
XFILL_5_BUFX2_insert474 gnd vdd FILL
XFILL_1__6967_ gnd vdd FILL
XFILL_1__9755_ gnd vdd FILL
XSFILL79400x1050 gnd vdd FILL
XFILL_5_BUFX2_insert485 gnd vdd FILL
XFILL_5_BUFX2_insert496 gnd vdd FILL
XFILL_4__9464_ gnd vdd FILL
XSFILL33960x64050 gnd vdd FILL
X_13171_ _13169_/Y _13173_/A _13171_/C gnd _13205_/D vdd OAI21X1
X_10383_ _10443_/A _7439_/B gnd _10384_/C vdd NAND2X1
XFILL_1__8706_ gnd vdd FILL
XSFILL48760x24050 gnd vdd FILL
XFILL_1__6898_ gnd vdd FILL
XFILL_4__9395_ gnd vdd FILL
X_12122_ _12122_/A _12829_/A gnd _12122_/Y vdd NAND2X1
XFILL_1__8637_ gnd vdd FILL
XFILL_2__7430_ gnd vdd FILL
XFILL_4__8346_ gnd vdd FILL
X_12053_ _12053_/A _12025_/B _12025_/C gnd gnd _12053_/Y vdd AOI22X1
XFILL_1__8568_ gnd vdd FILL
XFILL_2__7361_ gnd vdd FILL
XFILL_4__8277_ gnd vdd FILL
XFILL_5__7070_ gnd vdd FILL
X_11004_ _12230_/Y _12126_/Y gnd _11015_/D vdd OR2X2
XFILL_2__9100_ gnd vdd FILL
XFILL_4__7228_ gnd vdd FILL
XSFILL3720x41050 gnd vdd FILL
XFILL_2__7292_ gnd vdd FILL
XFILL_1__8499_ gnd vdd FILL
X_15812_ _15812_/A _15812_/B _15812_/C gnd _15812_/Y vdd AOI21X1
XFILL_2__9031_ gnd vdd FILL
XFILL_3__10940_ gnd vdd FILL
XFILL_2_BUFX2_insert320 gnd vdd FILL
XSFILL28920x53050 gnd vdd FILL
XFILL_1__10030_ gnd vdd FILL
XFILL_4__11190_ gnd vdd FILL
XFILL_2_BUFX2_insert331 gnd vdd FILL
XFILL_0__10760_ gnd vdd FILL
XFILL_4__7159_ gnd vdd FILL
XFILL_2_BUFX2_insert342 gnd vdd FILL
XFILL_2_BUFX2_insert353 gnd vdd FILL
XFILL_5__11500_ gnd vdd FILL
XFILL_4__10141_ gnd vdd FILL
X_12955_ vdd _12955_/B gnd _12956_/C vdd NAND2X1
X_15743_ _8423_/Q _15978_/B _15978_/C _8551_/Q gnd _15745_/C vdd AOI22X1
XFILL_5__12480_ gnd vdd FILL
XFILL_2_BUFX2_insert364 gnd vdd FILL
XFILL_2__11320_ gnd vdd FILL
XFILL_2_BUFX2_insert375 gnd vdd FILL
XFILL_3__10871_ gnd vdd FILL
XFILL_2_BUFX2_insert386 gnd vdd FILL
XFILL_2_BUFX2_insert397 gnd vdd FILL
X_11906_ _11934_/B _12361_/A gnd _11907_/C vdd NAND2X1
XFILL_0__10691_ gnd vdd FILL
XFILL_3__12610_ gnd vdd FILL
XFILL_5__7972_ gnd vdd FILL
XFILL_5__11431_ gnd vdd FILL
X_15674_ _15674_/A _15394_/B _15394_/C _15673_/Y gnd _15675_/A vdd OAI22X1
X_12886_ _12886_/A gnd _12888_/A vdd INVX1
XFILL_3__13590_ gnd vdd FILL
XFILL_2__11251_ gnd vdd FILL
XFILL_0__12430_ gnd vdd FILL
XFILL_5__6923_ gnd vdd FILL
XFILL_1__11981_ gnd vdd FILL
X_14625_ _14625_/A _14624_/Y gnd _14625_/Y vdd NOR2X1
XFILL_5__14150_ gnd vdd FILL
XFILL_4__13900_ gnd vdd FILL
X_11837_ _12117_/Y _11373_/Y gnd _11837_/Y vdd NOR2X1
XSFILL74120x37050 gnd vdd FILL
XFILL_5__11362_ gnd vdd FILL
XFILL_2__9933_ gnd vdd FILL
XFILL_4__14880_ gnd vdd FILL
XFILL_1__13720_ gnd vdd FILL
XFILL_1__10932_ gnd vdd FILL
XFILL_0__12361_ gnd vdd FILL
XFILL_2__11182_ gnd vdd FILL
XFILL_5__13101_ gnd vdd FILL
XFILL_5__9642_ gnd vdd FILL
XSFILL84280x81050 gnd vdd FILL
X_14556_ _14555_/Y _14552_/Y gnd _14559_/C vdd NOR2X1
XFILL_5__6854_ gnd vdd FILL
XFILL_5__10313_ gnd vdd FILL
XFILL_4__13831_ gnd vdd FILL
XFILL_5__11293_ gnd vdd FILL
XFILL_5__14081_ gnd vdd FILL
XFILL_3__15260_ gnd vdd FILL
X_11768_ _11445_/Y _11768_/B _11767_/Y gnd _11769_/A vdd AOI21X1
XFILL_3__12472_ gnd vdd FILL
XBUFX2_insert330 _12405_/Y gnd _9907_/B vdd BUFX2
XFILL_2__10133_ gnd vdd FILL
XFILL_0__14100_ gnd vdd FILL
XFILL_0__11312_ gnd vdd FILL
XFILL_1__13651_ gnd vdd FILL
XFILL_2__9864_ gnd vdd FILL
XFILL_2__15990_ gnd vdd FILL
XBUFX2_insert341 _12811_/Q gnd _13443_/A vdd BUFX2
XFILL_0__12292_ gnd vdd FILL
XFILL_0__15080_ gnd vdd FILL
XFILL_3__14211_ gnd vdd FILL
XFILL_5__10244_ gnd vdd FILL
XFILL_5__13032_ gnd vdd FILL
X_10719_ _15439_/A _7647_/CLK _9823_/R vdd _10643_/Y gnd vdd DFFSR
XBUFX2_insert352 _13306_/Y gnd _7955_/B vdd BUFX2
X_13507_ _13507_/A _13461_/C _14051_/C _13505_/Y gnd _13511_/A vdd OAI22X1
X_14487_ _9451_/Q gnd _15895_/A vdd INVX1
XFILL_6__12583_ gnd vdd FILL
XBUFX2_insert363 _11352_/Y gnd _11660_/A vdd BUFX2
XFILL_3__11423_ gnd vdd FILL
XFILL_1__12602_ gnd vdd FILL
XFILL_3__15191_ gnd vdd FILL
XFILL_4__13762_ gnd vdd FILL
X_11699_ _11699_/A _11698_/Y gnd _11700_/A vdd NOR2X1
XBUFX2_insert374 _13338_/Y gnd _9514_/A vdd BUFX2
XFILL_4__10974_ gnd vdd FILL
XBUFX2_insert385 _13331_/Y gnd _9151_/A vdd BUFX2
XFILL_1__16370_ gnd vdd FILL
XFILL_0__14031_ gnd vdd FILL
XFILL_2__14941_ gnd vdd FILL
XFILL_0__11243_ gnd vdd FILL
XFILL_2__10064_ gnd vdd FILL
XFILL_5_CLKBUF1_insert220 gnd vdd FILL
XFILL_5__8524_ gnd vdd FILL
XFILL_1__13582_ gnd vdd FILL
XFILL_2__9795_ gnd vdd FILL
X_16226_ _16225_/Y _16226_/B gnd _16231_/A vdd NOR2X1
XBUFX2_insert396 _13293_/Y gnd _7568_/B vdd BUFX2
XFILL_4__15501_ gnd vdd FILL
XFILL_0__7830_ gnd vdd FILL
X_13438_ _13868_/B gnd _13438_/Y vdd INVX8
XFILL_1__10794_ gnd vdd FILL
XFILL_4__12713_ gnd vdd FILL
XFILL_5__10175_ gnd vdd FILL
XFILL_3__14142_ gnd vdd FILL
XSFILL38760x56050 gnd vdd FILL
XFILL_1__15321_ gnd vdd FILL
XFILL_3__11354_ gnd vdd FILL
XFILL_2__14872_ gnd vdd FILL
XFILL112280x63050 gnd vdd FILL
XFILL_1__12533_ gnd vdd FILL
XFILL_2__8746_ gnd vdd FILL
XFILL_4__13693_ gnd vdd FILL
XFILL_0__11174_ gnd vdd FILL
XFILL_5__8455_ gnd vdd FILL
X_16157_ _7921_/Q gnd _16157_/Y vdd INVX1
X_13369_ _13443_/A _13398_/A _13465_/C gnd _14456_/C vdd NAND3X1
XFILL_3__10305_ gnd vdd FILL
XFILL_4__15432_ gnd vdd FILL
XFILL_0__7761_ gnd vdd FILL
XFILL_2__13823_ gnd vdd FILL
XFILL_4__12644_ gnd vdd FILL
XFILL_5__14983_ gnd vdd FILL
XFILL_3__14073_ gnd vdd FILL
XFILL_0__10125_ gnd vdd FILL
XFILL_1__15252_ gnd vdd FILL
XFILL_3__7470_ gnd vdd FILL
XFILL_3__11285_ gnd vdd FILL
XFILL_1__12464_ gnd vdd FILL
XFILL_0__9500_ gnd vdd FILL
XFILL_0__15982_ gnd vdd FILL
XFILL_5__8386_ gnd vdd FILL
X_15108_ _15563_/A _15107_/Y _15563_/C _13517_/D gnd _15108_/Y vdd OAI22X1
XFILL_3__13024_ gnd vdd FILL
X_16088_ _15652_/A _9584_/Q _9712_/Q _15652_/D gnd _16088_/Y vdd AOI22X1
XFILL_5__13934_ gnd vdd FILL
XFILL_0__7692_ gnd vdd FILL
XFILL_1__14203_ gnd vdd FILL
XFILL_4__15363_ gnd vdd FILL
XFILL_2__7628_ gnd vdd FILL
XFILL_3__10236_ gnd vdd FILL
XFILL_4__12575_ gnd vdd FILL
XSFILL114040x58050 gnd vdd FILL
XFILL_2__13754_ gnd vdd FILL
XSFILL43880x47050 gnd vdd FILL
XFILL_1__11415_ gnd vdd FILL
XFILL_2__10966_ gnd vdd FILL
XFILL_1__15183_ gnd vdd FILL
XFILL_5__7337_ gnd vdd FILL
XFILL_0__10056_ gnd vdd FILL
XFILL_0__14933_ gnd vdd FILL
X_15039_ _15220_/B _12812_/Q _16037_/B gnd _15715_/C vdd NAND3X1
XFILL_1__12395_ gnd vdd FILL
XFILL_4__14314_ gnd vdd FILL
XFILL_2__12705_ gnd vdd FILL
XFILL_5__13865_ gnd vdd FILL
XFILL_3__9140_ gnd vdd FILL
XFILL_4__11526_ gnd vdd FILL
XSFILL28840x3050 gnd vdd FILL
XFILL_3__10167_ gnd vdd FILL
XFILL_1__14134_ gnd vdd FILL
XFILL_4__15294_ gnd vdd FILL
XFILL_2__7559_ gnd vdd FILL
XSFILL18680x23050 gnd vdd FILL
XFILL_2__13685_ gnd vdd FILL
XSFILL99560x19050 gnd vdd FILL
XFILL_1__11346_ gnd vdd FILL
XFILL_0__14864_ gnd vdd FILL
XFILL_2__10897_ gnd vdd FILL
XFILL_5__15604_ gnd vdd FILL
XSFILL74200x17050 gnd vdd FILL
XFILL_0__9362_ gnd vdd FILL
XFILL_4__14245_ gnd vdd FILL
XFILL_2__15424_ gnd vdd FILL
XFILL_2__12636_ gnd vdd FILL
XFILL_5__13796_ gnd vdd FILL
XSFILL84360x61050 gnd vdd FILL
X_9990_ _9979_/B _8582_/B gnd _9990_/Y vdd NAND2X1
XFILL_4__11457_ gnd vdd FILL
XFILL_0__13815_ gnd vdd FILL
XFILL_1__14065_ gnd vdd FILL
XFILL_5__9007_ gnd vdd FILL
XFILL_3__14975_ gnd vdd FILL
XFILL_1__11277_ gnd vdd FILL
XFILL_0__8313_ gnd vdd FILL
XSFILL59000x78050 gnd vdd FILL
XFILL_0__14795_ gnd vdd FILL
XFILL_5__15535_ gnd vdd FILL
XFILL_5__7199_ gnd vdd FILL
XFILL_5__12747_ gnd vdd FILL
XFILL_4__10408_ gnd vdd FILL
XFILL_0__9293_ gnd vdd FILL
XFILL_2__9229_ gnd vdd FILL
X_8941_ _8891_/A _9453_/CLK _9453_/R vdd _8893_/Y gnd vdd DFFSR
XFILL_1__13016_ gnd vdd FILL
XFILL_4__14176_ gnd vdd FILL
XFILL_2__15355_ gnd vdd FILL
XFILL_4__11388_ gnd vdd FILL
XFILL_3__13926_ gnd vdd FILL
XSFILL99400x83050 gnd vdd FILL
XFILL_2__12567_ gnd vdd FILL
XFILL_0__13746_ gnd vdd FILL
XFILL_0__10958_ gnd vdd FILL
XFILL_0__8244_ gnd vdd FILL
XFILL_4__13127_ gnd vdd FILL
XFILL_5__15466_ gnd vdd FILL
XFILL_2__14306_ gnd vdd FILL
X_8872_ _8872_/A _8896_/B _8871_/Y gnd _8934_/D vdd OAI21X1
XFILL_2__11518_ gnd vdd FILL
XFILL_3__13857_ gnd vdd FILL
XFILL_2__15286_ gnd vdd FILL
XFILL_2__12498_ gnd vdd FILL
XSFILL38840x36050 gnd vdd FILL
XFILL_1__10159_ gnd vdd FILL
XSFILL38040x17050 gnd vdd FILL
XFILL_0__13677_ gnd vdd FILL
XFILL_6__9751_ gnd vdd FILL
XFILL_5__14417_ gnd vdd FILL
X_7823_ _7872_/B _9487_/B gnd _7824_/C vdd NAND2X1
XFILL112360x43050 gnd vdd FILL
XFILL_0__10889_ gnd vdd FILL
XFILL_5__11629_ gnd vdd FILL
XFILL_5__15397_ gnd vdd FILL
XSFILL64120x69050 gnd vdd FILL
XFILL_2__14237_ gnd vdd FILL
XFILL_2__11449_ gnd vdd FILL
XFILL_0__15416_ gnd vdd FILL
XFILL_5__9909_ gnd vdd FILL
XFILL_0__12628_ gnd vdd FILL
XFILL_3__13788_ gnd vdd FILL
XFILL_1__14967_ gnd vdd FILL
XFILL_6__8702_ gnd vdd FILL
XFILL_0__16396_ gnd vdd FILL
XFILL_4__12009_ gnd vdd FILL
XFILL_5__14348_ gnd vdd FILL
X_7754_ _7794_/Q gnd _7754_/Y vdd INVX1
XFILL_3__15527_ gnd vdd FILL
XFILL_6__6894_ gnd vdd FILL
XFILL_6__13899_ gnd vdd FILL
XFILL_3__12739_ gnd vdd FILL
XFILL_2__14168_ gnd vdd FILL
XFILL_1__13918_ gnd vdd FILL
XFILL_0__15347_ gnd vdd FILL
XFILL_1__14898_ gnd vdd FILL
XFILL_0__7057_ gnd vdd FILL
XSFILL3560x76050 gnd vdd FILL
XFILL_2__13119_ gnd vdd FILL
XFILL_5__14279_ gnd vdd FILL
X_7685_ _7771_/Q gnd _7685_/Y vdd INVX1
XFILL_3__15458_ gnd vdd FILL
XFILL_1__13849_ gnd vdd FILL
XFILL_3__8855_ gnd vdd FILL
XFILL_2__14099_ gnd vdd FILL
XFILL_5__16018_ gnd vdd FILL
XFILL_0__15278_ gnd vdd FILL
X_9424_ _9424_/A gnd _9424_/Y vdd INVX1
XFILL_1__7870_ gnd vdd FILL
XFILL_3__14409_ gnd vdd FILL
XSFILL8600x13050 gnd vdd FILL
XFILL_3__7806_ gnd vdd FILL
XFILL_0__14229_ gnd vdd FILL
XFILL_3__15389_ gnd vdd FILL
XSFILL44040x36050 gnd vdd FILL
XFILL_3__8786_ gnd vdd FILL
X_9355_ _9437_/Q gnd _9355_/Y vdd INVX1
XFILL_6__8495_ gnd vdd FILL
XFILL_1__15519_ gnd vdd FILL
XFILL_4_BUFX2_insert404 gnd vdd FILL
XFILL_3__7737_ gnd vdd FILL
X_8306_ _8266_/A _8306_/CLK _7533_/R vdd _8268_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert415 gnd vdd FILL
XFILL_1__9540_ gnd vdd FILL
XFILL_6__7446_ gnd vdd FILL
XFILL_0__7959_ gnd vdd FILL
XFILL_4_BUFX2_insert426 gnd vdd FILL
XSFILL33880x79050 gnd vdd FILL
XFILL_4_BUFX2_insert437 gnd vdd FILL
X_9286_ _9286_/A _9240_/A _9286_/C gnd _9328_/D vdd OAI21X1
XFILL_4_BUFX2_insert448 gnd vdd FILL
XFILL_4_BUFX2_insert459 gnd vdd FILL
XFILL_1__9471_ gnd vdd FILL
XFILL_4__8200_ gnd vdd FILL
X_8237_ _8237_/A _7853_/B gnd _8238_/C vdd NAND2X1
XFILL_3__9407_ gnd vdd FILL
XSFILL38920x16050 gnd vdd FILL
XFILL_6__9116_ gnd vdd FILL
XFILL112440x23050 gnd vdd FILL
XFILL_3__7599_ gnd vdd FILL
XFILL_0__9629_ gnd vdd FILL
X_8168_ _8168_/Q _8680_/CLK _8034_/R vdd _8168_/D gnd vdd DFFSR
XFILL_4__8131_ gnd vdd FILL
XFILL_3__9338_ gnd vdd FILL
XSFILL39000x25050 gnd vdd FILL
X_7119_ _7117_/Y _7100_/A _7119_/C gnd _7155_/D vdd OAI21X1
XFILL_1__8353_ gnd vdd FILL
XFILL_3__9269_ gnd vdd FILL
X_8099_ _8165_/Q gnd _8101_/A vdd INVX1
XFILL_4__8062_ gnd vdd FILL
XSFILL8600x4050 gnd vdd FILL
XFILL_1__7304_ gnd vdd FILL
XSFILL3640x56050 gnd vdd FILL
XFILL_3_CLKBUF1_insert117 gnd vdd FILL
XFILL_3_CLKBUF1_insert128 gnd vdd FILL
XFILL_5_CLKBUF1_insert1077 gnd vdd FILL
XSFILL28840x68050 gnd vdd FILL
XFILL_3_CLKBUF1_insert139 gnd vdd FILL
XSFILL94280x44050 gnd vdd FILL
XFILL_1__7235_ gnd vdd FILL
X_12740_ _11885_/B gnd _12740_/Y vdd INVX1
XSFILL54280x60050 gnd vdd FILL
XFILL_1_BUFX2_insert305 gnd vdd FILL
XFILL_1_BUFX2_insert316 gnd vdd FILL
XFILL_1__7166_ gnd vdd FILL
XFILL_1_BUFX2_insert327 gnd vdd FILL
XFILL_1_BUFX2_insert338 gnd vdd FILL
XFILL_4__8964_ gnd vdd FILL
XFILL_1_BUFX2_insert349 gnd vdd FILL
X_12671_ _12591_/A _12685_/CLK _12685_/R vdd _12671_/D gnd vdd DFFSR
XSFILL33960x59050 gnd vdd FILL
XFILL_1__7097_ gnd vdd FILL
X_14410_ _14410_/A _14410_/B _13978_/B _14408_/Y gnd _14411_/B vdd OAI22X1
X_11622_ _11621_/Y _11622_/B gnd _11627_/C vdd NOR2X1
XFILL_4__8895_ gnd vdd FILL
X_15390_ _9742_/A _15390_/B gnd _15398_/A vdd NAND2X1
XFILL_2__6930_ gnd vdd FILL
XFILL_4__7846_ gnd vdd FILL
X_14341_ _9516_/A gnd _14341_/Y vdd INVX1
X_11553_ _11552_/A _11553_/B _11553_/C gnd _11856_/B vdd OAI21X1
XFILL_2__6861_ gnd vdd FILL
X_10504_ _15298_/D gnd _10504_/Y vdd INVX1
X_14272_ _14268_/Y _14271_/Y gnd _14275_/C vdd NOR2X1
XFILL_1__9807_ gnd vdd FILL
XFILL_2__8600_ gnd vdd FILL
XFILL_5_BUFX2_insert260 gnd vdd FILL
X_11484_ _11167_/Y _11484_/B _11423_/B _11166_/Y gnd _11485_/A vdd OAI22X1
XFILL_5_BUFX2_insert271 gnd vdd FILL
XFILL_1__7999_ gnd vdd FILL
X_16011_ _16293_/A _7150_/Q _8126_/A _16011_/D gnd _16012_/B vdd AOI22X1
XFILL_5_BUFX2_insert282 gnd vdd FILL
XFILL_4__9516_ gnd vdd FILL
XSFILL3720x36050 gnd vdd FILL
X_13223_ _13289_/B _13231_/B gnd _13225_/D vdd NAND2X1
X_10435_ _10435_/A _10450_/B _10434_/Y gnd _10435_/Y vdd OAI21X1
XSFILL94360x9050 gnd vdd FILL
XFILL_5_BUFX2_insert293 gnd vdd FILL
XFILL_2__8531_ gnd vdd FILL
XFILL_1__9738_ gnd vdd FILL
XFILL_4__10690_ gnd vdd FILL
XSFILL28920x48050 gnd vdd FILL
XFILL_5__8240_ gnd vdd FILL
X_13154_ _13200_/Q gnd _13154_/Y vdd INVX1
X_10366_ _10364_/Y _10363_/B _10366_/C gnd _10366_/Y vdd OAI21X1
XFILL_2__8462_ gnd vdd FILL
XFILL_5__11980_ gnd vdd FILL
XFILL_2__10820_ gnd vdd FILL
XFILL_4_BUFX2_insert960 gnd vdd FILL
XFILL_3__11070_ gnd vdd FILL
XFILL_4_BUFX2_insert971 gnd vdd FILL
XFILL_1__9669_ gnd vdd FILL
X_12105_ _12105_/A _12105_/B _12001_/C gnd gnd _12105_/Y vdd AOI22X1
XSFILL28520x50050 gnd vdd FILL
XFILL_4_BUFX2_insert982 gnd vdd FILL
XFILL_4_BUFX2_insert993 gnd vdd FILL
XFILL_4__9378_ gnd vdd FILL
XFILL_5__10931_ gnd vdd FILL
XFILL_3__10021_ gnd vdd FILL
X_13085_ _13085_/A gnd _13087_/A vdd INVX1
XFILL_4__12360_ gnd vdd FILL
X_10297_ _10280_/B _9785_/B gnd _10297_/Y vdd NAND2X1
XFILL_1__11200_ gnd vdd FILL
XFILL_2__10751_ gnd vdd FILL
XFILL_5__7122_ gnd vdd FILL
XFILL_2__8393_ gnd vdd FILL
XFILL_4__8329_ gnd vdd FILL
XFILL_1__12180_ gnd vdd FILL
XFILL_0__11930_ gnd vdd FILL
X_12036_ _12028_/A _12801_/Q _12024_/C gnd _12036_/Y vdd NAND3X1
XFILL_5__13650_ gnd vdd FILL
XFILL_4__11311_ gnd vdd FILL
XFILL_4__12291_ gnd vdd FILL
XFILL_2__7344_ gnd vdd FILL
XFILL_2__13470_ gnd vdd FILL
XFILL_1__11131_ gnd vdd FILL
XFILL_5__7053_ gnd vdd FILL
XFILL_2__10682_ gnd vdd FILL
XFILL_5__12601_ gnd vdd FILL
XFILL_0__11861_ gnd vdd FILL
XSFILL84280x76050 gnd vdd FILL
XFILL_4__14030_ gnd vdd FILL
XFILL_4__11242_ gnd vdd FILL
XFILL_2__12421_ gnd vdd FILL
XFILL_5__13581_ gnd vdd FILL
XFILL_0__13600_ gnd vdd FILL
XFILL_3__11972_ gnd vdd FILL
XFILL_5__10793_ gnd vdd FILL
XFILL_1__11062_ gnd vdd FILL
XFILL_3__14760_ gnd vdd FILL
XFILL_0__10812_ gnd vdd FILL
XFILL_0__14580_ gnd vdd FILL
XFILL_5__15320_ gnd vdd FILL
XFILL_6__14871_ gnd vdd FILL
XFILL_2__9014_ gnd vdd FILL
XFILL_5__12532_ gnd vdd FILL
XSFILL89320x13050 gnd vdd FILL
XFILL_0__11792_ gnd vdd FILL
XFILL_3__10923_ gnd vdd FILL
XSFILL59080x52050 gnd vdd FILL
XFILL_2__15140_ gnd vdd FILL
XFILL_3__13711_ gnd vdd FILL
XFILL_4__11173_ gnd vdd FILL
XFILL_2__12352_ gnd vdd FILL
X_13987_ _13987_/A _13987_/B _13986_/Y gnd _13998_/B vdd NAND3X1
XFILL_1__10013_ gnd vdd FILL
XFILL_3__14691_ gnd vdd FILL
XFILL_0__13531_ gnd vdd FILL
XSFILL109480x19050 gnd vdd FILL
XFILL_1__15870_ gnd vdd FILL
XFILL_0__10743_ gnd vdd FILL
XFILL_4__10124_ gnd vdd FILL
XFILL_6__13822_ gnd vdd FILL
X_15726_ _15726_/A _14248_/Y _14258_/Y _15197_/C gnd _15729_/B vdd OAI22X1
XFILL_5__15251_ gnd vdd FILL
XFILL_5__12463_ gnd vdd FILL
X_12938_ _12938_/Q _13184_/CLK _8176_/R vdd _12938_/D gnd vdd DFFSR
XFILL_2__11303_ gnd vdd FILL
XFILL_4__15981_ gnd vdd FILL
XFILL_3__13642_ gnd vdd FILL
XFILL_1__14821_ gnd vdd FILL
XFILL_2__15071_ gnd vdd FILL
XFILL112280x58050 gnd vdd FILL
XFILL_0__16250_ gnd vdd FILL
XFILL_2__12283_ gnd vdd FILL
XFILL_5__14202_ gnd vdd FILL
XFILL_0__13462_ gnd vdd FILL
XFILL_0__10674_ gnd vdd FILL
XFILL_5__7955_ gnd vdd FILL
XFILL_5__11414_ gnd vdd FILL
XFILL_5__15182_ gnd vdd FILL
X_15657_ _14177_/Y _15376_/B gnd _15658_/C vdd NOR2X1
XFILL_2__14022_ gnd vdd FILL
XFILL_1_BUFX2_insert850 gnd vdd FILL
XFILL_4__14932_ gnd vdd FILL
XFILL_4__10055_ gnd vdd FILL
XFILL_0__15201_ gnd vdd FILL
X_12869_ vdd _12869_/B gnd _12870_/C vdd NAND2X1
XFILL_5__12394_ gnd vdd FILL
XFILL_3__16361_ gnd vdd FILL
XFILL_3__13573_ gnd vdd FILL
XFILL_2__11234_ gnd vdd FILL
XFILL_0__12413_ gnd vdd FILL
XFILL_3__10785_ gnd vdd FILL
XFILL_3__6970_ gnd vdd FILL
XFILL_1__14752_ gnd vdd FILL
XFILL_1_BUFX2_insert861 gnd vdd FILL
XFILL_0__16181_ gnd vdd FILL
XFILL_1__11964_ gnd vdd FILL
XFILL_1_BUFX2_insert872 gnd vdd FILL
XFILL_5__6906_ gnd vdd FILL
XSFILL13800x70050 gnd vdd FILL
X_14608_ _9918_/A _14867_/C _14213_/A _9838_/Q gnd _14608_/Y vdd AOI22X1
XFILL_5__14133_ gnd vdd FILL
XFILL_0__13393_ gnd vdd FILL
XFILL_1_BUFX2_insert883 gnd vdd FILL
XFILL_5__7886_ gnd vdd FILL
XFILL_1_BUFX2_insert894 gnd vdd FILL
XFILL_3__15312_ gnd vdd FILL
XFILL_6__13684_ gnd vdd FILL
XFILL_5__11345_ gnd vdd FILL
XFILL_2__9916_ gnd vdd FILL
XFILL_4__14863_ gnd vdd FILL
XFILL_3__12524_ gnd vdd FILL
XFILL_1__13703_ gnd vdd FILL
XFILL_0__9980_ gnd vdd FILL
X_15588_ _7325_/A _15114_/B _15114_/C gnd _15589_/C vdd NAND3X1
XFILL_1__10915_ gnd vdd FILL
XSFILL79240x65050 gnd vdd FILL
XFILL_3__16292_ gnd vdd FILL
XFILL_2__11165_ gnd vdd FILL
XFILL_0__15132_ gnd vdd FILL
XFILL_0__12344_ gnd vdd FILL
XFILL_5__9625_ gnd vdd FILL
XFILL_1__14683_ gnd vdd FILL
XFILL_5__6837_ gnd vdd FILL
XFILL_1__11895_ gnd vdd FILL
XFILL_4__13814_ gnd vdd FILL
X_14539_ _8376_/A _13647_/B _14481_/C _7020_/Q gnd _14547_/B vdd AOI22X1
XFILL_5__14064_ gnd vdd FILL
XFILL_2__10116_ gnd vdd FILL
XFILL_3__15243_ gnd vdd FILL
XFILL_3__12455_ gnd vdd FILL
X_7470_ _7470_/A _7470_/B _7469_/Y gnd _7528_/D vdd OAI21X1
XFILL_5__11276_ gnd vdd FILL
XFILL_3__8640_ gnd vdd FILL
XFILL_1__13634_ gnd vdd FILL
XFILL_2__9847_ gnd vdd FILL
XFILL_4__14794_ gnd vdd FILL
XFILL_2__15973_ gnd vdd FILL
XFILL_0__15063_ gnd vdd FILL
XFILL_0__12275_ gnd vdd FILL
XFILL_2__11096_ gnd vdd FILL
XSFILL114680x50 gnd vdd FILL
XSFILL18680x18050 gnd vdd FILL
XFILL_5__13015_ gnd vdd FILL
XFILL_5__9556_ gnd vdd FILL
XSFILL8520x28050 gnd vdd FILL
XFILL_3__11406_ gnd vdd FILL
XFILL_0__8862_ gnd vdd FILL
XFILL_4__13745_ gnd vdd FILL
XFILL_4__10957_ gnd vdd FILL
XFILL_3__15174_ gnd vdd FILL
XFILL_2__10047_ gnd vdd FILL
XFILL_3__12386_ gnd vdd FILL
XFILL_0__14014_ gnd vdd FILL
XFILL_1__16353_ gnd vdd FILL
XFILL_3__8571_ gnd vdd FILL
XFILL_2__14924_ gnd vdd FILL
XFILL_5__8507_ gnd vdd FILL
XSFILL84360x56050 gnd vdd FILL
XFILL_1__13565_ gnd vdd FILL
XFILL_0__11226_ gnd vdd FILL
XFILL_2__9778_ gnd vdd FILL
X_16209_ _16208_/Y _16209_/B gnd _16210_/C vdd NOR2X1
XFILL_1__10777_ gnd vdd FILL
XFILL_0__7813_ gnd vdd FILL
XFILL_5__9487_ gnd vdd FILL
X_9140_ _9140_/A _9112_/A _9139_/Y gnd _9140_/Y vdd OAI21X1
XFILL_1__15304_ gnd vdd FILL
XFILL_3__14125_ gnd vdd FILL
XFILL_5__10158_ gnd vdd FILL
XFILL_3__11337_ gnd vdd FILL
XFILL_2__8729_ gnd vdd FILL
XFILL_4__13676_ gnd vdd FILL
XFILL_1__12516_ gnd vdd FILL
XFILL_2__14855_ gnd vdd FILL
XFILL_1__16284_ gnd vdd FILL
XFILL_4__10888_ gnd vdd FILL
XSFILL59160x32050 gnd vdd FILL
XFILL_0__11157_ gnd vdd FILL
XSFILL99400x78050 gnd vdd FILL
XFILL_5__8438_ gnd vdd FILL
XFILL_1__13496_ gnd vdd FILL
XFILL_0__7744_ gnd vdd FILL
XFILL_4__15415_ gnd vdd FILL
XFILL_4__12627_ gnd vdd FILL
XFILL_3__14056_ gnd vdd FILL
XFILL_5__14966_ gnd vdd FILL
X_9071_ _9025_/A _9823_/CLK _9056_/R vdd _9027_/Y gnd vdd DFFSR
XFILL_4__16395_ gnd vdd FILL
XFILL_2__13806_ gnd vdd FILL
XFILL_1__15235_ gnd vdd FILL
XFILL_3__7453_ gnd vdd FILL
XFILL_0__10108_ gnd vdd FILL
XFILL_3__11268_ gnd vdd FILL
XFILL_1__12447_ gnd vdd FILL
XFILL_2__11998_ gnd vdd FILL
XFILL_0__15965_ gnd vdd FILL
XFILL_2__14786_ gnd vdd FILL
XFILL_0__11088_ gnd vdd FILL
XFILL_6__7162_ gnd vdd FILL
X_8022_ _8022_/Q _8022_/CLK _9046_/R vdd _7928_/Y gnd vdd DFFSR
XFILL111880x31050 gnd vdd FILL
XFILL_3__13007_ gnd vdd FILL
XFILL_5__8369_ gnd vdd FILL
XFILL_5__13917_ gnd vdd FILL
XFILL_4__15346_ gnd vdd FILL
XFILL112360x38050 gnd vdd FILL
XFILL_0__7675_ gnd vdd FILL
XFILL_6__11379_ gnd vdd FILL
XFILL_5__14897_ gnd vdd FILL
XFILL_2__10949_ gnd vdd FILL
XFILL_0__10039_ gnd vdd FILL
XFILL_1__15166_ gnd vdd FILL
XFILL_2__13737_ gnd vdd FILL
XFILL_0__14916_ gnd vdd FILL
XFILL_3__11199_ gnd vdd FILL
XFILL_0__9414_ gnd vdd FILL
XFILL_1__12378_ gnd vdd FILL
XFILL_0__15896_ gnd vdd FILL
XFILL_5__13848_ gnd vdd FILL
XFILL_3__9123_ gnd vdd FILL
XFILL_4__11509_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1083 gnd vdd FILL
XFILL_1__14117_ gnd vdd FILL
XFILL_4__15277_ gnd vdd FILL
XFILL_2__13668_ gnd vdd FILL
XFILL_4__12489_ gnd vdd FILL
XSFILL114600x6050 gnd vdd FILL
XFILL_1__11329_ gnd vdd FILL
XFILL_0__14847_ gnd vdd FILL
XFILL_1__15097_ gnd vdd FILL
XFILL_0__9345_ gnd vdd FILL
XSFILL79320x45050 gnd vdd FILL
XFILL_4__14228_ gnd vdd FILL
XFILL_2__12619_ gnd vdd FILL
XFILL_2__15407_ gnd vdd FILL
XFILL_5__13779_ gnd vdd FILL
X_9973_ _9973_/Q _9205_/CLK _7285_/R vdd _9973_/D gnd vdd DFFSR
XFILL_1__14048_ gnd vdd FILL
XFILL_3__14958_ gnd vdd FILL
XFILL_2__13599_ gnd vdd FILL
XFILL_2__16387_ gnd vdd FILL
XFILL_5__15518_ gnd vdd FILL
XFILL_0__14778_ gnd vdd FILL
X_8924_ _8924_/Q _8926_/CLK _8025_/R vdd _8924_/D gnd vdd DFFSR
XFILL_0__9276_ gnd vdd FILL
XFILL_3__8005_ gnd vdd FILL
XFILL_4__14159_ gnd vdd FILL
XFILL_3__13909_ gnd vdd FILL
XSFILL114520x54050 gnd vdd FILL
XFILL_2__15338_ gnd vdd FILL
XFILL_0__13729_ gnd vdd FILL
XFILL_3__14889_ gnd vdd FILL
XFILL_0__8227_ gnd vdd FILL
XFILL_5__15449_ gnd vdd FILL
X_8855_ _8855_/A gnd _8855_/Y vdd INVX1
XFILL_2__15269_ gnd vdd FILL
XFILL_1__15999_ gnd vdd FILL
X_7806_ _7804_/Y _7814_/A _7806_/C gnd _7806_/Y vdd OAI21X1
XSFILL59240x12050 gnd vdd FILL
X_8786_ _8786_/A _8753_/B _8786_/C gnd _8820_/D vdd OAI21X1
XFILL_0__7109_ gnd vdd FILL
XFILL_0__16379_ gnd vdd FILL
XFILL_0__8089_ gnd vdd FILL
X_7737_ _7684_/B _9785_/B gnd _7737_/Y vdd NAND2X1
XFILL_1__8971_ gnd vdd FILL
XFILL_3__8907_ gnd vdd FILL
XFILL_4__7700_ gnd vdd FILL
XFILL111960x11050 gnd vdd FILL
XFILL_3__9887_ gnd vdd FILL
XFILL112440x18050 gnd vdd FILL
XSFILL23720x53050 gnd vdd FILL
X_7668_ _7632_/A _8297_/CLK _7796_/R vdd _7668_/D gnd vdd DFFSR
XFILL_4__7631_ gnd vdd FILL
XFILL_3__8838_ gnd vdd FILL
X_9407_ _9420_/B _7359_/B gnd _9408_/C vdd NAND2X1
XFILL112040x20050 gnd vdd FILL
XFILL_1__7853_ gnd vdd FILL
XFILL_4__7562_ gnd vdd FILL
X_7599_ _7599_/A gnd _7601_/A vdd INVX1
XFILL_3__8769_ gnd vdd FILL
X_9338_ _9339_/B _9466_/B gnd _9338_/Y vdd NAND2X1
XFILL_4__9301_ gnd vdd FILL
XFILL_4_BUFX2_insert234 gnd vdd FILL
X_10220_ _10220_/Q _8560_/CLK _9313_/R vdd _10170_/Y gnd vdd DFFSR
XFILL_4__7493_ gnd vdd FILL
XFILL_4_BUFX2_insert245 gnd vdd FILL
XSFILL94280x39050 gnd vdd FILL
XFILL_4_BUFX2_insert256 gnd vdd FILL
XFILL_1__9523_ gnd vdd FILL
X_9269_ _9269_/A gnd _9271_/A vdd INVX1
XFILL_4_BUFX2_insert267 gnd vdd FILL
XFILL_4__9232_ gnd vdd FILL
XFILL_4_BUFX2_insert278 gnd vdd FILL
X_10151_ _10191_/B _7847_/B gnd _10152_/C vdd NAND2X1
XFILL_4_BUFX2_insert289 gnd vdd FILL
XFILL_3_BUFX2_insert901 gnd vdd FILL
XFILL_3_BUFX2_insert912 gnd vdd FILL
XSFILL69080x15050 gnd vdd FILL
XFILL_4__9163_ gnd vdd FILL
XFILL_3_BUFX2_insert923 gnd vdd FILL
XFILL_3_BUFX2_insert934 gnd vdd FILL
XFILL_3_BUFX2_insert945 gnd vdd FILL
XFILL_3_BUFX2_insert956 gnd vdd FILL
X_10082_ _10082_/Q _6998_/CLK _7644_/R vdd _10082_/D gnd vdd DFFSR
XFILL_1__8405_ gnd vdd FILL
XFILL_1__9385_ gnd vdd FILL
XFILL_3_BUFX2_insert967 gnd vdd FILL
XFILL_4__8114_ gnd vdd FILL
XFILL_3_BUFX2_insert978 gnd vdd FILL
XFILL_4__9094_ gnd vdd FILL
XFILL_3_BUFX2_insert989 gnd vdd FILL
X_13910_ _7391_/Q _14738_/A _14909_/C _7135_/Q gnd _13918_/B vdd AOI22X1
XFILL_1__8336_ gnd vdd FILL
XSFILL64120x7050 gnd vdd FILL
X_14890_ _7248_/A _14458_/C _14413_/A _8272_/A gnd _14891_/B vdd AOI22X1
X_13841_ _7390_/Q gnd _13843_/D vdd INVX1
XFILL_1__8267_ gnd vdd FILL
XFILL_2__7060_ gnd vdd FILL
XFILL_3_BUFX2_insert1006 gnd vdd FILL
XFILL_3_BUFX2_insert1017 gnd vdd FILL
X_13772_ _13772_/A _13772_/B _13772_/C gnd _13788_/B vdd NAND3X1
XFILL_3_BUFX2_insert1028 gnd vdd FILL
XFILL_1__7218_ gnd vdd FILL
X_10984_ _10984_/Q _12667_/CLK _12689_/R vdd _10984_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert1039 gnd vdd FILL
XFILL_1_BUFX2_insert102 gnd vdd FILL
XFILL_1__8198_ gnd vdd FILL
XSFILL59800x6050 gnd vdd FILL
X_15511_ _15510_/Y _15504_/Y gnd _15536_/A vdd NOR2X1
XFILL_4__9996_ gnd vdd FILL
X_12723_ _12723_/A memoryOutData[9] gnd _12724_/C vdd NAND2X1
XFILL_5__7740_ gnd vdd FILL
XSFILL94360x19050 gnd vdd FILL
X_12654_ _12654_/A gnd _12656_/A vdd INVX1
XFILL_6__10750_ gnd vdd FILL
X_15442_ _7135_/Q gnd _15442_/Y vdd INVX1
XFILL_0_BUFX2_insert802 gnd vdd FILL
XFILL_3__10570_ gnd vdd FILL
XFILL_2__7962_ gnd vdd FILL
XFILL_0_BUFX2_insert813 gnd vdd FILL
X_11605_ _11120_/Y _11573_/C gnd _11606_/C vdd NAND2X1
XFILL_0__10390_ gnd vdd FILL
XFILL_0_BUFX2_insert824 gnd vdd FILL
XFILL_0_BUFX2_insert835 gnd vdd FILL
XFILL_5__7671_ gnd vdd FILL
XFILL_4__8878_ gnd vdd FILL
XFILL_5__11130_ gnd vdd FILL
X_12585_ _12362_/B gnd _12587_/A vdd INVX1
X_15373_ _15373_/A _15373_/B _13274_/A gnd _12845_/B vdd AOI21X1
XFILL_0_BUFX2_insert846 gnd vdd FILL
XFILL_2__6913_ gnd vdd FILL
XFILL_1__10700_ gnd vdd FILL
XFILL_1_BUFX2_insert1010 gnd vdd FILL
XFILL_4__11860_ gnd vdd FILL
XFILL_2__7893_ gnd vdd FILL
XFILL_5__9410_ gnd vdd FILL
XFILL_1_BUFX2_insert1021 gnd vdd FILL
XFILL_0_BUFX2_insert857 gnd vdd FILL
XFILL_1_BUFX2_insert1032 gnd vdd FILL
XFILL_0_BUFX2_insert868 gnd vdd FILL
XFILL_4__7829_ gnd vdd FILL
XFILL_1__11680_ gnd vdd FILL
XFILL_1_BUFX2_insert1043 gnd vdd FILL
XFILL_0_BUFX2_insert879 gnd vdd FILL
X_14324_ _8424_/Q _14037_/B _13884_/C _10796_/A gnd _14324_/Y vdd AOI22X1
X_11536_ _11289_/C _11449_/Y _11536_/C gnd _11537_/A vdd AOI21X1
XSFILL109400x7050 gnd vdd FILL
XFILL_4__10811_ gnd vdd FILL
XFILL_3__12240_ gnd vdd FILL
XFILL_5__11061_ gnd vdd FILL
XFILL_1_BUFX2_insert1054 gnd vdd FILL
XFILL_2__9632_ gnd vdd FILL
XFILL_2__6844_ gnd vdd FILL
XFILL_0__12060_ gnd vdd FILL
XFILL_2__12970_ gnd vdd FILL
XFILL_1__10631_ gnd vdd FILL
XFILL_4__11791_ gnd vdd FILL
XFILL_1_BUFX2_insert1065 gnd vdd FILL
XFILL_3_BUFX2_insert17 gnd vdd FILL
XFILL_5__9341_ gnd vdd FILL
XFILL_1_BUFX2_insert1087 gnd vdd FILL
X_14255_ _8806_/Q gnd _15718_/D vdd INVX1
XFILL_3_BUFX2_insert28 gnd vdd FILL
XFILL_6__12351_ gnd vdd FILL
XFILL_5__10012_ gnd vdd FILL
XFILL_4__13530_ gnd vdd FILL
XFILL_3_BUFX2_insert39 gnd vdd FILL
X_11467_ _11173_/Y gnd _11467_/Y vdd INVX1
XFILL_4__10742_ gnd vdd FILL
XFILL_2__11921_ gnd vdd FILL
XFILL_3__12171_ gnd vdd FILL
XFILL_0__11011_ gnd vdd FILL
XFILL_1__13350_ gnd vdd FILL
X_13206_ _13172_/A _13180_/CLK _13180_/R vdd _13206_/D gnd vdd DFFSR
XFILL_1__10562_ gnd vdd FILL
XFILL_5__14820_ gnd vdd FILL
XFILL_5__9272_ gnd vdd FILL
X_10418_ _10418_/A gnd _10420_/A vdd INVX1
X_14186_ _8421_/Q _13848_/B _13883_/B _9379_/A gnd _14194_/C vdd AOI22X1
XFILL_3__11122_ gnd vdd FILL
XFILL_4__13461_ gnd vdd FILL
XSFILL59080x47050 gnd vdd FILL
XFILL_1__12301_ gnd vdd FILL
XFILL_2__8514_ gnd vdd FILL
X_11398_ _12270_/Y _11278_/B _11687_/A gnd _11400_/B vdd OAI21X1
XFILL_2__14640_ gnd vdd FILL
XFILL_4__10673_ gnd vdd FILL
XFILL_2__9494_ gnd vdd FILL
XFILL_2__11852_ gnd vdd FILL
XFILL_1__13281_ gnd vdd FILL
XFILL_5__8223_ gnd vdd FILL
XFILL_4__15200_ gnd vdd FILL
X_13137_ _13134_/A _13137_/B gnd _13138_/C vdd NAND2X1
XFILL_1__10493_ gnd vdd FILL
X_10349_ _10349_/Q _8429_/CLK _9203_/R vdd _10349_/D gnd vdd DFFSR
XFILL_4__12412_ gnd vdd FILL
XSFILL74120x50050 gnd vdd FILL
XFILL_5__14751_ gnd vdd FILL
XFILL_4__16180_ gnd vdd FILL
XFILL_3__15930_ gnd vdd FILL
XFILL_1__15020_ gnd vdd FILL
XFILL_5__11963_ gnd vdd FILL
XFILL_3__11053_ gnd vdd FILL
XFILL_4_BUFX2_insert790 gnd vdd FILL
XFILL_2__10803_ gnd vdd FILL
XFILL_2__14571_ gnd vdd FILL
XFILL_4__13392_ gnd vdd FILL
XFILL_1__12232_ gnd vdd FILL
XFILL_2__8445_ gnd vdd FILL
XFILL_2__11783_ gnd vdd FILL
XFILL_0__15750_ gnd vdd FILL
XFILL_0__12962_ gnd vdd FILL
XFILL_5__13702_ gnd vdd FILL
XFILL_5__10914_ gnd vdd FILL
X_13068_ _6891_/A _12669_/CLK _12795_/R vdd _13068_/D gnd vdd DFFSR
XFILL_0__7460_ gnd vdd FILL
XFILL_6_CLKBUF1_insert178 gnd vdd FILL
XFILL_3__10004_ gnd vdd FILL
XFILL_4__15131_ gnd vdd FILL
XFILL_4__12343_ gnd vdd FILL
XFILL_2__16310_ gnd vdd FILL
XFILL_5__14682_ gnd vdd FILL
XFILL_2__13522_ gnd vdd FILL
XFILL_2__8376_ gnd vdd FILL
XFILL_5__11894_ gnd vdd FILL
XFILL_0__14701_ gnd vdd FILL
XFILL_3__15861_ gnd vdd FILL
XFILL_0__11913_ gnd vdd FILL
XFILL_1__12163_ gnd vdd FILL
XFILL_5__7105_ gnd vdd FILL
XFILL_0__15681_ gnd vdd FILL
X_12019_ _12047_/A _11912_/B _12011_/C gnd _12019_/Y vdd NAND3X1
XFILL_5__8085_ gnd vdd FILL
XFILL_5__13633_ gnd vdd FILL
XFILL_0__12893_ gnd vdd FILL
XFILL_3__14812_ gnd vdd FILL
XFILL_4__15062_ gnd vdd FILL
XFILL_2__7327_ gnd vdd FILL
XFILL_2__16241_ gnd vdd FILL
XFILL_2__13453_ gnd vdd FILL
XFILL_4__12274_ gnd vdd FILL
XFILL_1__11114_ gnd vdd FILL
XFILL_0__14632_ gnd vdd FILL
XFILL_3__15792_ gnd vdd FILL
XFILL_2__10665_ gnd vdd FILL
XFILL_5__7036_ gnd vdd FILL
XFILL_1__12094_ gnd vdd FILL
XFILL_0__9130_ gnd vdd FILL
XFILL_0__11844_ gnd vdd FILL
XFILL_6__10046_ gnd vdd FILL
XFILL_4__14013_ gnd vdd FILL
XFILL_5__16352_ gnd vdd FILL
XFILL_2__12404_ gnd vdd FILL
XFILL_5__13564_ gnd vdd FILL
XFILL_4__11225_ gnd vdd FILL
XFILL_2__16172_ gnd vdd FILL
XFILL_5__10776_ gnd vdd FILL
X_6970_ _6968_/Y _6937_/B _6969_/Y gnd _6970_/Y vdd OAI21X1
XFILL_3__14743_ gnd vdd FILL
XFILL_1__15922_ gnd vdd FILL
XFILL_3__11955_ gnd vdd FILL
XFILL_2__13384_ gnd vdd FILL
XFILL_1__11045_ gnd vdd FILL
XFILL_0__14563_ gnd vdd FILL
XFILL_5__15303_ gnd vdd FILL
XFILL_5__12515_ gnd vdd FILL
XFILL_0__11775_ gnd vdd FILL
XFILL_4__11156_ gnd vdd FILL
XFILL_2__15123_ gnd vdd FILL
XFILL_5__16283_ gnd vdd FILL
XFILL_3__10906_ gnd vdd FILL
XFILL_0__16302_ gnd vdd FILL
XFILL_2__12335_ gnd vdd FILL
XFILL_5__13495_ gnd vdd FILL
XFILL_3__14674_ gnd vdd FILL
XFILL_2__7189_ gnd vdd FILL
XFILL_0__13514_ gnd vdd FILL
XFILL_3__11886_ gnd vdd FILL
XFILL_0__8012_ gnd vdd FILL
XFILL_1__15853_ gnd vdd FILL
XFILL_0__14494_ gnd vdd FILL
X_15709_ _7910_/Q gnd _15711_/A vdd INVX1
XFILL_5__15234_ gnd vdd FILL
XFILL_4__10107_ gnd vdd FILL
X_8640_ _8638_/Y _8577_/B _8640_/C gnd _8686_/D vdd OAI21X1
XFILL_5__8987_ gnd vdd FILL
XFILL_5__12446_ gnd vdd FILL
XFILL_3__16413_ gnd vdd FILL
XSFILL48920x7050 gnd vdd FILL
XFILL_3__13625_ gnd vdd FILL
XSFILL43880x60050 gnd vdd FILL
XFILL_2__15054_ gnd vdd FILL
XFILL_4__15964_ gnd vdd FILL
XFILL_4__11087_ gnd vdd FILL
XFILL_3__9810_ gnd vdd FILL
XFILL_1__14804_ gnd vdd FILL
XFILL_0__16233_ gnd vdd FILL
XFILL_2__12266_ gnd vdd FILL
XFILL_3__10837_ gnd vdd FILL
XFILL_0__13445_ gnd vdd FILL
XFILL_1__15784_ gnd vdd FILL
XFILL_1__12996_ gnd vdd FILL
XFILL_5__7938_ gnd vdd FILL
XFILL_0__10657_ gnd vdd FILL
XSFILL59160x27050 gnd vdd FILL
XFILL_4__10038_ gnd vdd FILL
XFILL_2__14005_ gnd vdd FILL
XFILL_5__15165_ gnd vdd FILL
XFILL_4__14915_ gnd vdd FILL
XFILL_3__16344_ gnd vdd FILL
XFILL_5__12377_ gnd vdd FILL
XFILL_1_BUFX2_insert680 gnd vdd FILL
X_8571_ _8571_/A _8619_/B _8570_/Y gnd _8663_/D vdd OAI21X1
XFILL_2__11217_ gnd vdd FILL
XFILL_3__10768_ gnd vdd FILL
XFILL_3__9741_ gnd vdd FILL
XFILL_4__15895_ gnd vdd FILL
XFILL_1__14735_ gnd vdd FILL
XFILL_3__13556_ gnd vdd FILL
XFILL_1_BUFX2_insert691 gnd vdd FILL
XFILL_1__11947_ gnd vdd FILL
XSFILL74200x30050 gnd vdd FILL
XFILL_2__12197_ gnd vdd FILL
XFILL_0__16164_ gnd vdd FILL
XFILL_3__6953_ gnd vdd FILL
XFILL_0__13376_ gnd vdd FILL
XFILL_5__14116_ gnd vdd FILL
XFILL_5__7869_ gnd vdd FILL
X_7522_ _7522_/Q _7382_/CLK _8418_/R vdd _7452_/Y gnd vdd DFFSR
XFILL_5__11328_ gnd vdd FILL
XFILL_4__14846_ gnd vdd FILL
XFILL_3__12507_ gnd vdd FILL
XFILL_6__10879_ gnd vdd FILL
XFILL_5__15096_ gnd vdd FILL
XFILL_2__11148_ gnd vdd FILL
XFILL_0__15115_ gnd vdd FILL
XFILL_3__16275_ gnd vdd FILL
XFILL_5__9608_ gnd vdd FILL
XFILL_3__10699_ gnd vdd FILL
XFILL_3__6884_ gnd vdd FILL
XFILL_3__13487_ gnd vdd FILL
XFILL_3__9672_ gnd vdd FILL
XFILL_0__12327_ gnd vdd FILL
XFILL_1__14666_ gnd vdd FILL
XFILL_1__11878_ gnd vdd FILL
XFILL_0__16095_ gnd vdd FILL
XFILL_5__14047_ gnd vdd FILL
XFILL_0__8914_ gnd vdd FILL
XFILL_3__15226_ gnd vdd FILL
X_7453_ _7523_/Q gnd _7455_/A vdd INVX1
XFILL_5__11259_ gnd vdd FILL
XFILL_1__13617_ gnd vdd FILL
XFILL_0__9894_ gnd vdd FILL
XFILL_1__16405_ gnd vdd FILL
XFILL_3__12438_ gnd vdd FILL
XFILL_3__8623_ gnd vdd FILL
XFILL_4__14777_ gnd vdd FILL
XFILL_1__10829_ gnd vdd FILL
XFILL_4__11989_ gnd vdd FILL
XFILL_2__15956_ gnd vdd FILL
XFILL_0__15046_ gnd vdd FILL
XFILL_2__11079_ gnd vdd FILL
XFILL_1__14597_ gnd vdd FILL
XFILL_0__12258_ gnd vdd FILL
XFILL_5__9539_ gnd vdd FILL
XFILL_6__15337_ gnd vdd FILL
XFILL_0__8845_ gnd vdd FILL
XFILL_4__13728_ gnd vdd FILL
XFILL_3__12369_ gnd vdd FILL
XFILL_1__16336_ gnd vdd FILL
XFILL_3__15157_ gnd vdd FILL
X_7384_ _7292_/A _7143_/CLK _7015_/R vdd _7384_/D gnd vdd DFFSR
XFILL_2__14907_ gnd vdd FILL
XFILL_1__13548_ gnd vdd FILL
XFILL_0__11209_ gnd vdd FILL
XFILL_2__15887_ gnd vdd FILL
X_9123_ _9123_/A gnd _9125_/A vdd INVX1
XFILL_0__12189_ gnd vdd FILL
XSFILL64120x82050 gnd vdd FILL
XFILL_3__14108_ gnd vdd FILL
XFILL_0__8776_ gnd vdd FILL
XFILL_4__13659_ gnd vdd FILL
XFILL_3__7505_ gnd vdd FILL
XFILL_5__15998_ gnd vdd FILL
XFILL_2__14838_ gnd vdd FILL
XFILL_3__15088_ gnd vdd FILL
XFILL_1__16267_ gnd vdd FILL
XFILL_3__8485_ gnd vdd FILL
XSFILL113720x2050 gnd vdd FILL
XSFILL74120x2050 gnd vdd FILL
XFILL_1__13479_ gnd vdd FILL
X_9054_ _8974_/A _8537_/CLK _9054_/R vdd _9054_/D gnd vdd DFFSR
XFILL_6__15199_ gnd vdd FILL
XFILL_0__7727_ gnd vdd FILL
XFILL_1__15218_ gnd vdd FILL
XFILL_3__14039_ gnd vdd FILL
XFILL_5__14949_ gnd vdd FILL
XFILL_4__16378_ gnd vdd FILL
XFILL_3__7436_ gnd vdd FILL
XFILL_1__16198_ gnd vdd FILL
XFILL_0__15948_ gnd vdd FILL
XFILL_2__14769_ gnd vdd FILL
XSFILL43960x40050 gnd vdd FILL
X_8005_ _8006_/B _8005_/B gnd _8005_/Y vdd NAND2X1
XFILL_4__15329_ gnd vdd FILL
XFILL_3__7367_ gnd vdd FILL
XFILL_1__15149_ gnd vdd FILL
XFILL_0__15879_ gnd vdd FILL
XFILL_2_BUFX2_insert908 gnd vdd FILL
XFILL_1__9170_ gnd vdd FILL
XFILL_0__7589_ gnd vdd FILL
XFILL_3__9106_ gnd vdd FILL
XFILL_2_BUFX2_insert919 gnd vdd FILL
XFILL_3__7298_ gnd vdd FILL
XFILL_1__8121_ gnd vdd FILL
X_9956_ _9888_/A _7642_/CLK _7258_/R vdd _9890_/Y gnd vdd DFFSR
XFILL_3__9037_ gnd vdd FILL
XSFILL88680x36050 gnd vdd FILL
X_8907_ _8893_/B _8011_/B gnd _8908_/C vdd NAND2X1
XFILL_0__9259_ gnd vdd FILL
X_9887_ _9887_/A _9941_/B _9886_/Y gnd _9955_/D vdd OAI21X1
XFILL_4__9850_ gnd vdd FILL
XSFILL49160x59050 gnd vdd FILL
XSFILL23320x50050 gnd vdd FILL
X_8838_ _8916_/A _6918_/B gnd _8839_/C vdd NAND2X1
XFILL_6__7978_ gnd vdd FILL
XFILL_4__9781_ gnd vdd FILL
XFILL_6__6929_ gnd vdd FILL
XFILL_4__6993_ gnd vdd FILL
XBUFX2_insert907 _10913_/Y gnd _12723_/A vdd BUFX2
XBUFX2_insert918 _15069_/Y gnd _15169_/D vdd BUFX2
XFILL_6_BUFX2_insert863 gnd vdd FILL
XFILL_0_BUFX2_insert109 gnd vdd FILL
X_8769_ _8815_/Q gnd _8771_/A vdd INVX1
XFILL_6_BUFX2_insert874 gnd vdd FILL
XFILL_4__8732_ gnd vdd FILL
XFILL_3__9939_ gnd vdd FILL
XBUFX2_insert929 _12351_/Y gnd _8701_/B vdd BUFX2
XFILL_6__9648_ gnd vdd FILL
XFILL_1__8954_ gnd vdd FILL
X_12370_ _12023_/B gnd _12370_/Y vdd INVX1
XFILL_1__8885_ gnd vdd FILL
XFILL_4__7614_ gnd vdd FILL
XSFILL28840x81050 gnd vdd FILL
X_11321_ _11174_/C _11320_/Y gnd _11321_/Y vdd NOR2X1
XSFILL104280x19050 gnd vdd FILL
XFILL_4__8594_ gnd vdd FILL
XFILL_1__7836_ gnd vdd FILL
X_14040_ _14039_/Y _14200_/C gnd _14040_/Y vdd NOR2X1
XFILL_4__7545_ gnd vdd FILL
X_11252_ _11026_/B gnd _11253_/B vdd INVX1
XSFILL8760x79050 gnd vdd FILL
XSFILL23800x28050 gnd vdd FILL
X_10203_ _13699_/A _8792_/CLK _9048_/R vdd _10203_/D gnd vdd DFFSR
XSFILL33960x72050 gnd vdd FILL
XFILL_4__7476_ gnd vdd FILL
XFILL_1__9506_ gnd vdd FILL
X_11183_ _11181_/Y _11182_/Y _11492_/B gnd _11184_/A vdd OAI21X1
XFILL_4__9215_ gnd vdd FILL
XFILL_1__7698_ gnd vdd FILL
XFILL_3_BUFX2_insert720 gnd vdd FILL
XFILL_3_BUFX2_insert731 gnd vdd FILL
X_10134_ _10134_/A _10193_/A _10133_/Y gnd _10134_/Y vdd OAI21X1
XFILL_2__8230_ gnd vdd FILL
X_15991_ _15989_/Y _15342_/B _15991_/C gnd _15991_/Y vdd OAI21X1
XFILL_3_BUFX2_insert742 gnd vdd FILL
XFILL_3_BUFX2_insert753 gnd vdd FILL
XFILL_3_BUFX2_insert764 gnd vdd FILL
XFILL_4__9146_ gnd vdd FILL
XFILL_3_BUFX2_insert775 gnd vdd FILL
X_14942_ _14942_/A _14389_/B _14942_/C gnd _14951_/A vdd AOI21X1
X_10065_ _10066_/B _8529_/B gnd _10065_/Y vdd NAND2X1
XFILL_3_BUFX2_insert786 gnd vdd FILL
XSFILL74280x8050 gnd vdd FILL
XFILL_1__9368_ gnd vdd FILL
XFILL_3_BUFX2_insert797 gnd vdd FILL
XFILL_2__7112_ gnd vdd FILL
XFILL_5__10630_ gnd vdd FILL
XFILL_1__8319_ gnd vdd FILL
X_14873_ _10355_/Q gnd _14873_/Y vdd INVX1
XFILL_2__8092_ gnd vdd FILL
XFILL_1__9299_ gnd vdd FILL
XFILL_2__10450_ gnd vdd FILL
XFILL_5__8910_ gnd vdd FILL
XFILL_4__11010_ gnd vdd FILL
X_13824_ _13822_/Y _13824_/B _14575_/C _13823_/Y gnd _13825_/B vdd OAI22X1
XFILL_5__9890_ gnd vdd FILL
XFILL_2__7043_ gnd vdd FILL
XFILL_5__10561_ gnd vdd FILL
XFILL_3__11740_ gnd vdd FILL
XFILL_2__10381_ gnd vdd FILL
XFILL_5__8841_ gnd vdd FILL
XFILL_5__12300_ gnd vdd FILL
XFILL_0__11560_ gnd vdd FILL
XFILL_5__13280_ gnd vdd FILL
X_10967_ _12773_/A gnd _10968_/B vdd INVX1
X_13755_ _15331_/D _13868_/B _14643_/C _13755_/D gnd _13759_/A vdd OAI22X1
XFILL_2__12120_ gnd vdd FILL
XFILL_3__11671_ gnd vdd FILL
XFILL_5__10492_ gnd vdd FILL
XFILL_0__10511_ gnd vdd FILL
XFILL_1__12850_ gnd vdd FILL
X_12706_ _12704_/Y _12721_/B _12706_/C gnd _12794_/D vdd OAI21X1
XFILL_5__8772_ gnd vdd FILL
XFILL_5__12231_ gnd vdd FILL
XFILL_0__11491_ gnd vdd FILL
XFILL_4__9979_ gnd vdd FILL
XFILL_3__13410_ gnd vdd FILL
XFILL_3__10622_ gnd vdd FILL
X_10898_ _10987_/Q _10897_/Y gnd _10898_/Y vdd NAND2X1
XFILL_4__12961_ gnd vdd FILL
X_13686_ _13686_/A _13685_/Y _14597_/C gnd _12964_/B vdd AOI21X1
XFILL_2__12051_ gnd vdd FILL
XFILL_1__11801_ gnd vdd FILL
XFILL_0__13230_ gnd vdd FILL
XFILL_3__14390_ gnd vdd FILL
XFILL_1__12781_ gnd vdd FILL
XFILL_0__10442_ gnd vdd FILL
XFILL_2__8994_ gnd vdd FILL
XFILL_0_BUFX2_insert610 gnd vdd FILL
XSFILL48840x12050 gnd vdd FILL
XFILL_6__13521_ gnd vdd FILL
XFILL_5__7723_ gnd vdd FILL
XFILL_4__14700_ gnd vdd FILL
XFILL_0_BUFX2_insert621 gnd vdd FILL
X_15425_ _15423_/Y _15425_/B gnd _15426_/B vdd NOR2X1
X_12637_ vdd memoryOutData[23] gnd _12638_/C vdd NAND2X1
XFILL_4__11912_ gnd vdd FILL
XFILL_5__12162_ gnd vdd FILL
XSFILL49320x19050 gnd vdd FILL
XFILL_2__11002_ gnd vdd FILL
XFILL_0_BUFX2_insert632 gnd vdd FILL
XFILL_3__13341_ gnd vdd FILL
XFILL_4__15680_ gnd vdd FILL
XFILL_1__14520_ gnd vdd FILL
XFILL_3__10553_ gnd vdd FILL
XSFILL74120x45050 gnd vdd FILL
XFILL_2__7945_ gnd vdd FILL
XFILL_4__12892_ gnd vdd FILL
XFILL_0_BUFX2_insert643 gnd vdd FILL
XFILL_1__11732_ gnd vdd FILL
XFILL_0_BUFX2_insert654 gnd vdd FILL
XFILL_0__13161_ gnd vdd FILL
XFILL_0__10373_ gnd vdd FILL
XFILL_0_BUFX2_insert665 gnd vdd FILL
XFILL_5__11113_ gnd vdd FILL
XFILL_4__14631_ gnd vdd FILL
X_12568_ memoryOutData[0] vdd gnd _12569_/C vdd NAND2X1
X_15356_ _10379_/A _15175_/B _15356_/C _10589_/Q gnd _15361_/A vdd AOI22X1
XFILL_0__6960_ gnd vdd FILL
XFILL_3__13272_ gnd vdd FILL
XFILL_5__12093_ gnd vdd FILL
XFILL_2__15810_ gnd vdd FILL
XFILL_3__16060_ gnd vdd FILL
XFILL_0_BUFX2_insert676 gnd vdd FILL
XFILL_4__11843_ gnd vdd FILL
XFILL_1__14451_ gnd vdd FILL
XFILL_0_BUFX2_insert687 gnd vdd FILL
XFILL_0__12112_ gnd vdd FILL
XFILL_6__12403_ gnd vdd FILL
XFILL_2__7876_ gnd vdd FILL
XFILL_1__11663_ gnd vdd FILL
XFILL_0_BUFX2_insert698 gnd vdd FILL
XFILL_6__16171_ gnd vdd FILL
XFILL_0__13092_ gnd vdd FILL
X_14307_ _10215_/Q gnd _14307_/Y vdd INVX1
X_11519_ _11623_/A _11623_/B _11519_/C gnd _11520_/B vdd OAI21X1
XFILL_5__15921_ gnd vdd FILL
XFILL_5__7585_ gnd vdd FILL
XFILL_3__15011_ gnd vdd FILL
XFILL_3__12223_ gnd vdd FILL
XFILL_5__11044_ gnd vdd FILL
XFILL_2__9615_ gnd vdd FILL
XFILL_4__14562_ gnd vdd FILL
XFILL_0__6891_ gnd vdd FILL
XFILL_1__13402_ gnd vdd FILL
X_12499_ _12403_/A gnd _12499_/Y vdd INVX1
X_15287_ _9947_/Q gnd _15287_/Y vdd INVX1
XFILL_1__10614_ gnd vdd FILL
XFILL_4__11774_ gnd vdd FILL
XSFILL109480x32050 gnd vdd FILL
XFILL_2__15741_ gnd vdd FILL
XFILL_0__12043_ gnd vdd FILL
XFILL_2__12953_ gnd vdd FILL
XFILL_1__14382_ gnd vdd FILL
XFILL_6__15122_ gnd vdd FILL
XFILL_0__8630_ gnd vdd FILL
XFILL_4__16301_ gnd vdd FILL
XFILL_1__11594_ gnd vdd FILL
X_14238_ _9702_/Q gnd _14238_/Y vdd INVX1
XFILL_4__13513_ gnd vdd FILL
XSFILL110200x82050 gnd vdd FILL
XFILL_1__16121_ gnd vdd FILL
XFILL_5__15852_ gnd vdd FILL
XFILL_3__12154_ gnd vdd FILL
XFILL_2__9546_ gnd vdd FILL
XFILL_1__13333_ gnd vdd FILL
XFILL112280x71050 gnd vdd FILL
XFILL_4__14493_ gnd vdd FILL
XFILL_2__11904_ gnd vdd FILL
XFILL_2__15672_ gnd vdd FILL
XFILL_1__10545_ gnd vdd FILL
XSFILL54040x12050 gnd vdd FILL
XFILL_2__12884_ gnd vdd FILL
XFILL_5__9255_ gnd vdd FILL
XFILL_4__16232_ gnd vdd FILL
XFILL_5__14803_ gnd vdd FILL
X_14169_ _14169_/A _14168_/Y gnd _14170_/A vdd NAND2X1
XFILL_3__11105_ gnd vdd FILL
XFILL_4__13444_ gnd vdd FILL
XFILL_5__15783_ gnd vdd FILL
XFILL_3__8270_ gnd vdd FILL
XFILL_2__14623_ gnd vdd FILL
XFILL_3__12085_ gnd vdd FILL
XFILL_4__10656_ gnd vdd FILL
XFILL_5__12995_ gnd vdd FILL
XFILL_0__15802_ gnd vdd FILL
XFILL_1__16052_ gnd vdd FILL
XFILL_2__11835_ gnd vdd FILL
XFILL_5__8206_ gnd vdd FILL
XFILL_1__13264_ gnd vdd FILL
XFILL_2__9477_ gnd vdd FILL
XFILL_6__11216_ gnd vdd FILL
XFILL_0__13994_ gnd vdd FILL
XFILL_5__14734_ gnd vdd FILL
XFILL_3__7221_ gnd vdd FILL
XFILL_3__15913_ gnd vdd FILL
XFILL_5__11946_ gnd vdd FILL
XFILL_1__15003_ gnd vdd FILL
XFILL_0__8492_ gnd vdd FILL
XFILL_3__11036_ gnd vdd FILL
XFILL_4__16163_ gnd vdd FILL
XFILL_4__13375_ gnd vdd FILL
XSFILL43880x55050 gnd vdd FILL
XFILL_1__12215_ gnd vdd FILL
XFILL_2__14554_ gnd vdd FILL
XFILL_0__15733_ gnd vdd FILL
XFILL_2__11766_ gnd vdd FILL
XFILL_5__8137_ gnd vdd FILL
XFILL_0__7443_ gnd vdd FILL
XFILL_4__15114_ gnd vdd FILL
XFILL_5__14665_ gnd vdd FILL
XFILL_4__12326_ gnd vdd FILL
XFILL_5__11877_ gnd vdd FILL
XFILL_4__16094_ gnd vdd FILL
XFILL_3__15844_ gnd vdd FILL
XFILL_2__13505_ gnd vdd FILL
XFILL_2__8359_ gnd vdd FILL
XFILL_2__14485_ gnd vdd FILL
XSFILL58920x77050 gnd vdd FILL
XFILL_1__12146_ gnd vdd FILL
XFILL_0__15664_ gnd vdd FILL
XFILL_2__11697_ gnd vdd FILL
XFILL_5__13616_ gnd vdd FILL
XFILL_5__8068_ gnd vdd FILL
XFILL_0__12876_ gnd vdd FILL
XFILL_5__16404_ gnd vdd FILL
X_9810_ _9808_/Y _9785_/A _9809_/Y gnd _9810_/Y vdd OAI21X1
XFILL_0__7374_ gnd vdd FILL
XFILL_5__10828_ gnd vdd FILL
XFILL_4__15045_ gnd vdd FILL
XFILL_6__11078_ gnd vdd FILL
XFILL_5__14596_ gnd vdd FILL
XFILL_2__16224_ gnd vdd FILL
XFILL_4__12257_ gnd vdd FILL
XFILL_2__13436_ gnd vdd FILL
XFILL_0__14615_ gnd vdd FILL
XFILL_2__10648_ gnd vdd FILL
XFILL_3__15775_ gnd vdd FILL
XFILL_3__7083_ gnd vdd FILL
XFILL_1__12077_ gnd vdd FILL
XFILL_0__9113_ gnd vdd FILL
XFILL_3__12987_ gnd vdd FILL
XFILL_0__11827_ gnd vdd FILL
XFILL_5__16335_ gnd vdd FILL
XFILL_0__15595_ gnd vdd FILL
X_9741_ _9741_/A _9741_/B _9740_/Y gnd _9821_/D vdd OAI21X1
XFILL_5__13547_ gnd vdd FILL
XFILL_4__11208_ gnd vdd FILL
XFILL_3__14726_ gnd vdd FILL
XFILL_5__10759_ gnd vdd FILL
X_6953_ _7015_/Q gnd _6955_/A vdd INVX1
XFILL_1__15905_ gnd vdd FILL
XFILL_4__12188_ gnd vdd FILL
XFILL_2__13367_ gnd vdd FILL
XFILL_3__11938_ gnd vdd FILL
XFILL_1__11028_ gnd vdd FILL
XFILL_2__16155_ gnd vdd FILL
XFILL_0__14546_ gnd vdd FILL
XFILL_2__10579_ gnd vdd FILL
XFILL_0__9044_ gnd vdd FILL
XFILL_0__11758_ gnd vdd FILL
XSFILL105080x4050 gnd vdd FILL
XFILL_5__16266_ gnd vdd FILL
X_9672_ _9675_/A _7496_/B gnd _9673_/C vdd NAND2X1
XFILL_4__11139_ gnd vdd FILL
XFILL_2__15106_ gnd vdd FILL
XFILL_5__13478_ gnd vdd FILL
XFILL_2__12318_ gnd vdd FILL
X_6884_ _6884_/A gnd memoryWriteData[14] vdd BUFX2
XFILL_3__14657_ gnd vdd FILL
XFILL_2__16086_ gnd vdd FILL
XFILL_2__13298_ gnd vdd FILL
XFILL_3__11869_ gnd vdd FILL
XFILL_1__15836_ gnd vdd FILL
XFILL_0__10709_ gnd vdd FILL
XSFILL89480x79050 gnd vdd FILL
XFILL_0__14477_ gnd vdd FILL
XFILL_5__15217_ gnd vdd FILL
XSFILL38840x44050 gnd vdd FILL
XFILL_5__12429_ gnd vdd FILL
XFILL112360x51050 gnd vdd FILL
X_8623_ _8681_/Q gnd _8623_/Y vdd INVX1
XFILL_0__11689_ gnd vdd FILL
XSFILL64120x77050 gnd vdd FILL
XFILL_3__13608_ gnd vdd FILL
XFILL_5__16197_ gnd vdd FILL
XFILL_2__15037_ gnd vdd FILL
XFILL_4__15947_ gnd vdd FILL
XFILL_0__16216_ gnd vdd FILL
XFILL_2__12249_ gnd vdd FILL
XFILL_3__14588_ gnd vdd FILL
XFILL_0__13428_ gnd vdd FILL
XFILL_3__7985_ gnd vdd FILL
XFILL_1__15767_ gnd vdd FILL
XFILL_1__12979_ gnd vdd FILL
XFILL_5__15148_ gnd vdd FILL
XFILL_6__7694_ gnd vdd FILL
XFILL_3__16327_ gnd vdd FILL
X_8554_ _8498_/A _9578_/CLK _7793_/R vdd _8554_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert804 gnd vdd FILL
XFILL_5_BUFX2_insert815 gnd vdd FILL
XFILL_3__9724_ gnd vdd FILL
XFILL_3__13539_ gnd vdd FILL
XFILL_4__15878_ gnd vdd FILL
XFILL_3__6936_ gnd vdd FILL
XFILL_1__14718_ gnd vdd FILL
XFILL_5_BUFX2_insert826 gnd vdd FILL
XFILL_0__16147_ gnd vdd FILL
XFILL_0__13359_ gnd vdd FILL
XFILL_1__15698_ gnd vdd FILL
XBUFX2_insert1001 _12399_/Y gnd _9517_/B vdd BUFX2
XFILL_5_BUFX2_insert837 gnd vdd FILL
XBUFX2_insert1012 _13569_/Y gnd _14867_/C vdd BUFX2
XSFILL43960x35050 gnd vdd FILL
X_7505_ _7472_/A _8273_/B gnd _7505_/Y vdd NAND2X1
XFILL_4__14829_ gnd vdd FILL
XFILL_5_BUFX2_insert848 gnd vdd FILL
XFILL_5__15079_ gnd vdd FILL
X_8485_ _8485_/A _8484_/A _8485_/C gnd _8549_/D vdd OAI21X1
XFILL_5_BUFX2_insert859 gnd vdd FILL
XSFILL69080x9050 gnd vdd FILL
XBUFX2_insert1023 _13340_/Y gnd _9628_/B vdd BUFX2
XFILL_3__16258_ gnd vdd FILL
XFILL_3__9655_ gnd vdd FILL
XBUFX2_insert1034 _13333_/Y gnd _9240_/A vdd BUFX2
XFILL_1__14649_ gnd vdd FILL
XFILL_3__6867_ gnd vdd FILL
XFILL_0__16078_ gnd vdd FILL
XBUFX2_insert1045 _13297_/Y gnd _7729_/B vdd BUFX2
XBUFX2_insert1056 _13527_/Y gnd _14712_/B vdd BUFX2
XFILL_6__9364_ gnd vdd FILL
X_7436_ _7503_/B _7948_/B gnd _7437_/C vdd NAND2X1
XFILL_3__15209_ gnd vdd FILL
XSFILL18760x11050 gnd vdd FILL
XFILL_0__9877_ gnd vdd FILL
XFILL_3__8606_ gnd vdd FILL
XBUFX2_insert1067 _13327_/Y gnd _8854_/B vdd BUFX2
XSFILL8600x21050 gnd vdd FILL
XFILL_3__16189_ gnd vdd FILL
XFILL_0__15029_ gnd vdd FILL
XSFILL44040x44050 gnd vdd FILL
XFILL_2__15939_ gnd vdd FILL
XBUFX2_insert1089 rst gnd BUFX2_insert496/A vdd BUFX2
XFILL_6__8315_ gnd vdd FILL
XFILL_1__7621_ gnd vdd FILL
XFILL_0__8828_ gnd vdd FILL
X_7367_ _7367_/A gnd _7367_/Y vdd INVX1
XFILL_4__7330_ gnd vdd FILL
XFILL_1__16319_ gnd vdd FILL
X_9106_ _9170_/B _7186_/B gnd _9106_/Y vdd NAND2X1
XSFILL84280x3050 gnd vdd FILL
XFILL_1__7552_ gnd vdd FILL
XFILL_0__8759_ gnd vdd FILL
X_7298_ _7298_/A gnd _7300_/A vdd INVX1
XFILL_3__8468_ gnd vdd FILL
XFILL111800x65050 gnd vdd FILL
X_9037_ _9075_/Q gnd _9037_/Y vdd INVX1
XFILL_4__9000_ gnd vdd FILL
XFILL_1__7483_ gnd vdd FILL
XFILL_3__7419_ gnd vdd FILL
XFILL_4__7192_ gnd vdd FILL
XFILL112440x31050 gnd vdd FILL
XFILL_3__8399_ gnd vdd FILL
XSFILL64200x57050 gnd vdd FILL
XSFILL79000x17050 gnd vdd FILL
XFILL_1__9222_ gnd vdd FILL
XFILL_2_BUFX2_insert705 gnd vdd FILL
XFILL_2_BUFX2_insert716 gnd vdd FILL
XFILL_2_BUFX2_insert727 gnd vdd FILL
XSFILL39000x33050 gnd vdd FILL
XFILL_1__9153_ gnd vdd FILL
XFILL_6__7059_ gnd vdd FILL
XFILL_2_BUFX2_insert738 gnd vdd FILL
XFILL_2_BUFX2_insert749 gnd vdd FILL
XFILL_1__8104_ gnd vdd FILL
XSFILL3640x64050 gnd vdd FILL
X_11870_ _11356_/A _11868_/Y _11869_/Y gnd _11871_/C vdd NAND3X1
XFILL_1__9084_ gnd vdd FILL
X_9939_ _9973_/Q gnd _9941_/A vdd INVX1
XFILL_4__9902_ gnd vdd FILL
XSFILL28840x76050 gnd vdd FILL
X_10821_ _10822_/B _9797_/B gnd _10821_/Y vdd NAND2X1
XSFILL94280x52050 gnd vdd FILL
X_10752_ _10789_/B _9344_/B gnd _10752_/Y vdd NAND2X1
X_13540_ _13539_/Y _13540_/B gnd _13540_/Y vdd NOR2X1
XSFILL44040x6050 gnd vdd FILL
XBUFX2_insert704 _11985_/Y gnd _12072_/C vdd BUFX2
XBUFX2_insert715 _15023_/Y gnd _15407_/B vdd BUFX2
XSFILL79400x4050 gnd vdd FILL
XFILL_4__9764_ gnd vdd FILL
XBUFX2_insert726 _13352_/Y gnd _10191_/B vdd BUFX2
XFILL_4__6976_ gnd vdd FILL
X_13471_ _13443_/A _13418_/A _13465_/C gnd _13471_/Y vdd NAND3X1
X_10683_ _10683_/A gnd _10685_/A vdd INVX1
XBUFX2_insert737 _12402_/Y gnd _8496_/B vdd BUFX2
XBUFX2_insert748 _13344_/Y gnd _9798_/B vdd BUFX2
XFILL_4__8715_ gnd vdd FILL
XFILL_1__9986_ gnd vdd FILL
XBUFX2_insert759 _12213_/Y gnd _12312_/C vdd BUFX2
X_12422_ _12422_/A _12645_/A gnd _12423_/C vdd NAND2X1
X_15210_ _15652_/A _9562_/Q _9602_/A _15652_/D gnd _15219_/A vdd AOI22X1
X_16190_ _16190_/A _16190_/B gnd _16202_/C vdd NAND2X1
XFILL_2__7730_ gnd vdd FILL
XFILL_4__8646_ gnd vdd FILL
X_12353_ _12368_/A _12576_/A gnd _12353_/Y vdd NAND2X1
X_15141_ _15140_/Y _15581_/C _15756_/D _15141_/D gnd _15142_/A vdd OAI22X1
XFILL_1_CLKBUF1_insert120 gnd vdd FILL
XFILL_1_CLKBUF1_insert131 gnd vdd FILL
XFILL_1_CLKBUF1_insert142 gnd vdd FILL
XFILL_1__8868_ gnd vdd FILL
X_11304_ _11133_/Y _11634_/A _11300_/A gnd _11304_/Y vdd OAI21X1
XFILL_4__8577_ gnd vdd FILL
XFILL_5__7370_ gnd vdd FILL
XFILL_1_CLKBUF1_insert153 gnd vdd FILL
X_15072_ _15000_/A _15044_/C _15024_/C gnd _15072_/Y vdd NAND3X1
XFILL_1_CLKBUF1_insert164 gnd vdd FILL
XFILL_2__9400_ gnd vdd FILL
X_12284_ _12224_/A _12308_/B _12224_/C gnd _12286_/B vdd NAND3X1
XFILL_1__7819_ gnd vdd FILL
XFILL_1_CLKBUF1_insert175 gnd vdd FILL
XFILL_2__7592_ gnd vdd FILL
XFILL_1_CLKBUF1_insert186 gnd vdd FILL
XSFILL38680x79050 gnd vdd FILL
X_14023_ _14023_/A _14023_/B gnd _14024_/A vdd NOR2X1
XFILL_1_CLKBUF1_insert197 gnd vdd FILL
X_11235_ _12230_/Y _12126_/Y gnd _11235_/Y vdd AND2X2
XFILL_4__10510_ gnd vdd FILL
XFILL_2_BUFX2_insert7 gnd vdd FILL
XFILL_4__11490_ gnd vdd FILL
XFILL_5__9040_ gnd vdd FILL
XSFILL94360x32050 gnd vdd FILL
XFILL_4__7459_ gnd vdd FILL
XFILL_6__12050_ gnd vdd FILL
XFILL_5__11800_ gnd vdd FILL
X_11166_ _12195_/Y _12322_/Y gnd _11166_/Y vdd NOR2X1
XFILL_5__12780_ gnd vdd FILL
XFILL_4__10441_ gnd vdd FILL
XFILL_2__11620_ gnd vdd FILL
XFILL_2__9262_ gnd vdd FILL
XFILL_1__10261_ gnd vdd FILL
XFILL_3_BUFX2_insert550 gnd vdd FILL
XFILL_6__11001_ gnd vdd FILL
X_10117_ _13699_/A gnd _10117_/Y vdd INVX1
XFILL_0__10991_ gnd vdd FILL
XFILL_3_BUFX2_insert561 gnd vdd FILL
XFILL_5__11731_ gnd vdd FILL
XFILL_3_BUFX2_insert572 gnd vdd FILL
X_15974_ _16235_/A _14553_/Y _15974_/C _16225_/C gnd _15974_/Y vdd OAI22X1
XFILL_3__12910_ gnd vdd FILL
XFILL_1__12000_ gnd vdd FILL
XFILL_4__10372_ gnd vdd FILL
XFILL_4__13160_ gnd vdd FILL
X_11097_ _11389_/A _11086_/Y _11097_/C gnd _11142_/A vdd AOI21X1
XFILL_2__8213_ gnd vdd FILL
XFILL_3_BUFX2_insert583 gnd vdd FILL
XFILL_2__11551_ gnd vdd FILL
XFILL_0__12730_ gnd vdd FILL
XFILL_3_BUFX2_insert594 gnd vdd FILL
XFILL_3__13890_ gnd vdd FILL
XFILL_4__9129_ gnd vdd FILL
XFILL_1__10192_ gnd vdd FILL
X_10048_ _10048_/A _9975_/B _10047_/Y gnd _10094_/D vdd OAI21X1
XFILL_4__12111_ gnd vdd FILL
X_14925_ _8656_/A _13864_/B _14403_/C _8564_/Q gnd _14925_/Y vdd AOI22X1
XFILL_5__14450_ gnd vdd FILL
XFILL_5__11662_ gnd vdd FILL
XFILL_2__10502_ gnd vdd FILL
XFILL_2__8144_ gnd vdd FILL
XFILL_3__12841_ gnd vdd FILL
XFILL_4__13091_ gnd vdd FILL
XFILL_2__14270_ gnd vdd FILL
XFILL_2__11482_ gnd vdd FILL
XFILL_0__12661_ gnd vdd FILL
XFILL_5__13401_ gnd vdd FILL
XFILL_2__13221_ gnd vdd FILL
X_14856_ _13601_/B _14855_/Y _14174_/C _14854_/Y gnd _14857_/A vdd OAI22X1
XFILL_4__12042_ gnd vdd FILL
XFILL_5__14381_ gnd vdd FILL
XFILL_2__8075_ gnd vdd FILL
XFILL_3__15560_ gnd vdd FILL
XFILL_0__14400_ gnd vdd FILL
XFILL_2__10433_ gnd vdd FILL
XFILL_5__11593_ gnd vdd FILL
XFILL_3__12772_ gnd vdd FILL
XFILL_0__11612_ gnd vdd FILL
XFILL_1__13951_ gnd vdd FILL
XFILL_0__15380_ gnd vdd FILL
XFILL_5__16120_ gnd vdd FILL
XFILL_0__12592_ gnd vdd FILL
XFILL_5__13332_ gnd vdd FILL
X_13807_ _9821_/Q _14470_/B _14878_/C _10589_/Q gnd _13815_/B vdd AOI22X1
XFILL_5__9873_ gnd vdd FILL
XSFILL89320x21050 gnd vdd FILL
XSFILL59080x60050 gnd vdd FILL
XFILL_3__14511_ gnd vdd FILL
XFILL_5__10544_ gnd vdd FILL
XFILL_0__7090_ gnd vdd FILL
XFILL_2__13152_ gnd vdd FILL
XFILL_1__12902_ gnd vdd FILL
X_14787_ _14787_/A _14815_/C gnd _14788_/B vdd NOR2X1
XFILL_3__11723_ gnd vdd FILL
X_11999_ _11999_/A _12352_/A _11999_/C gnd _12002_/A vdd NAND3X1
XFILL_6_BUFX2_insert65 gnd vdd FILL
XFILL_0__14331_ gnd vdd FILL
XSFILL109480x27050 gnd vdd FILL
XFILL_2__10364_ gnd vdd FILL
XFILL_3__15491_ gnd vdd FILL
XFILL_1__13882_ gnd vdd FILL
XFILL_5__8824_ gnd vdd FILL
XFILL_0__11543_ gnd vdd FILL
XFILL_4__15801_ gnd vdd FILL
XFILL_5__16051_ gnd vdd FILL
XFILL_5__13263_ gnd vdd FILL
XFILL_2__12103_ gnd vdd FILL
X_13738_ _13737_/Y _13727_/Y gnd _13739_/B vdd NOR2X1
XFILL_3__14442_ gnd vdd FILL
XFILL112280x66050 gnd vdd FILL
XFILL_1__12833_ gnd vdd FILL
XFILL_1__15621_ gnd vdd FILL
XFILL_4__13993_ gnd vdd FILL
XFILL_2__13083_ gnd vdd FILL
XFILL_3__11654_ gnd vdd FILL
XFILL_2__10295_ gnd vdd FILL
XFILL_0__14262_ gnd vdd FILL
XFILL_5__15002_ gnd vdd FILL
XFILL_5__12214_ gnd vdd FILL
XFILL_5__8755_ gnd vdd FILL
XFILL_0__11474_ gnd vdd FILL
XFILL_4__15732_ gnd vdd FILL
XFILL_0__16001_ gnd vdd FILL
X_13669_ _13668_/Y _14045_/A _14200_/C _13669_/D gnd _13669_/Y vdd OAI22X1
XFILL_2__12034_ gnd vdd FILL
XSFILL94440x12050 gnd vdd FILL
XFILL_0__13213_ gnd vdd FILL
XFILL_1__15552_ gnd vdd FILL
XFILL_3__14373_ gnd vdd FILL
XFILL_3__11585_ gnd vdd FILL
XFILL_1__12764_ gnd vdd FILL
XFILL_5__7706_ gnd vdd FILL
XFILL_0__10425_ gnd vdd FILL
XFILL_2__8977_ gnd vdd FILL
XFILL_0_BUFX2_insert440 gnd vdd FILL
X_15408_ _8670_/Q gnd _15410_/C vdd INVX1
XFILL_0__14193_ gnd vdd FILL
XFILL_0__9800_ gnd vdd FILL
XFILL_0_BUFX2_insert451 gnd vdd FILL
XFILL_3__16112_ gnd vdd FILL
XFILL_5__12145_ gnd vdd FILL
XFILL_3__13324_ gnd vdd FILL
XFILL_4__15663_ gnd vdd FILL
X_16388_ gnd gnd gnd _16389_/C vdd NAND2X1
XFILL_1__14503_ gnd vdd FILL
XFILL_0_BUFX2_insert462 gnd vdd FILL
XFILL_3__10536_ gnd vdd FILL
XSFILL79240x73050 gnd vdd FILL
XFILL_0__7992_ gnd vdd FILL
XFILL_0_BUFX2_insert473 gnd vdd FILL
XFILL_4__12875_ gnd vdd FILL
XFILL_1__11715_ gnd vdd FILL
XFILL_2__7928_ gnd vdd FILL
XFILL_0__13144_ gnd vdd FILL
XFILL_0_BUFX2_insert484 gnd vdd FILL
XFILL_1__15483_ gnd vdd FILL
XFILL_1__12695_ gnd vdd FILL
XFILL_5__7637_ gnd vdd FILL
XFILL_0_BUFX2_insert495 gnd vdd FILL
XFILL_4__14614_ gnd vdd FILL
X_15339_ _9437_/Q _15380_/B gnd _15348_/A vdd NAND2X1
XFILL_0__9731_ gnd vdd FILL
X_8270_ _8249_/A _7502_/B gnd _8271_/C vdd NAND2X1
XFILL_3__16043_ gnd vdd FILL
XFILL_5__12076_ gnd vdd FILL
XFILL_0__6943_ gnd vdd FILL
XFILL_4__11826_ gnd vdd FILL
XFILL_3__13255_ gnd vdd FILL
XSFILL28840x6050 gnd vdd FILL
XFILL_4__15594_ gnd vdd FILL
XFILL_1__14434_ gnd vdd FILL
XFILL_1__11646_ gnd vdd FILL
XFILL_2__7859_ gnd vdd FILL
XSFILL114440x82050 gnd vdd FILL
XFILL_2__13985_ gnd vdd FILL
XFILL_0__10287_ gnd vdd FILL
X_7221_ _7275_/Q gnd _7223_/A vdd INVX1
XFILL_5__7568_ gnd vdd FILL
XFILL_5__15904_ gnd vdd FILL
XFILL_5__11027_ gnd vdd FILL
XFILL_0__9662_ gnd vdd FILL
XFILL_4__14545_ gnd vdd FILL
XFILL_0__6874_ gnd vdd FILL
XFILL_3__12206_ gnd vdd FILL
XSFILL18120x69050 gnd vdd FILL
XFILL_2__15724_ gnd vdd FILL
XFILL_4__11757_ gnd vdd FILL
XSFILL84360x64050 gnd vdd FILL
XFILL_0__12026_ gnd vdd FILL
XFILL_3__9371_ gnd vdd FILL
XFILL_1__14365_ gnd vdd FILL
XFILL_3__10398_ gnd vdd FILL
XFILL_1__11577_ gnd vdd FILL
XFILL_0__8613_ gnd vdd FILL
XFILL_6__9080_ gnd vdd FILL
XFILL_5__7499_ gnd vdd FILL
X_7152_ _7108_/A _8289_/CLK _7152_/R vdd _7152_/D gnd vdd DFFSR
XFILL_5__15835_ gnd vdd FILL
XFILL_4__10708_ gnd vdd FILL
XFILL_1__13316_ gnd vdd FILL
XFILL_4__14476_ gnd vdd FILL
XFILL_3__8322_ gnd vdd FILL
XFILL_3__12137_ gnd vdd FILL
XFILL_1__16104_ gnd vdd FILL
XFILL_2__9529_ gnd vdd FILL
XFILL_0__9593_ gnd vdd FILL
XFILL_2__15655_ gnd vdd FILL
XFILL_1__10528_ gnd vdd FILL
XFILL_4__11688_ gnd vdd FILL
XFILL_2__12867_ gnd vdd FILL
XSFILL59160x40050 gnd vdd FILL
XFILL_5__9238_ gnd vdd FILL
XFILL_1__14296_ gnd vdd FILL
XFILL_4__16215_ gnd vdd FILL
XCLKBUF1_insert130 CLKBUF1_insert193/A gnd _7143_/CLK vdd CLKBUF1
XCLKBUF1_insert141 CLKBUF1_insert216/A gnd _7662_/CLK vdd CLKBUF1
XFILL_4__13427_ gnd vdd FILL
XFILL_4__10639_ gnd vdd FILL
XFILL_2__14606_ gnd vdd FILL
XFILL_1__16035_ gnd vdd FILL
XFILL_3__12068_ gnd vdd FILL
XCLKBUF1_insert152 CLKBUF1_insert150/A gnd _7786_/CLK vdd CLKBUF1
XFILL_5__15766_ gnd vdd FILL
XFILL_5__12978_ gnd vdd FILL
X_7083_ _7081_/Y _7067_/A _7083_/C gnd _7143_/D vdd OAI21X1
XFILL_1__13247_ gnd vdd FILL
XFILL_3__8253_ gnd vdd FILL
XCLKBUF1_insert163 CLKBUF1_insert169/A gnd _7664_/CLK vdd CLKBUF1
XFILL_2__11818_ gnd vdd FILL
XFILL_2__15586_ gnd vdd FILL
XFILL_0__13977_ gnd vdd FILL
XSFILL38840x39050 gnd vdd FILL
XCLKBUF1_insert174 CLKBUF1_insert169/A gnd _8180_/CLK vdd CLKBUF1
XFILL_5__9169_ gnd vdd FILL
XCLKBUF1_insert185 CLKBUF1_insert187/A gnd _12538_/CLK vdd CLKBUF1
XFILL_0__8475_ gnd vdd FILL
XFILL_5__11929_ gnd vdd FILL
XFILL112360x46050 gnd vdd FILL
XFILL_5__14717_ gnd vdd FILL
XFILL_3__11019_ gnd vdd FILL
XFILL_4__16146_ gnd vdd FILL
XCLKBUF1_insert196 CLKBUF1_insert192/A gnd _9817_/CLK vdd CLKBUF1
XFILL_3__7204_ gnd vdd FILL
XFILL_4__13358_ gnd vdd FILL
XFILL_5__15697_ gnd vdd FILL
XFILL_3__8184_ gnd vdd FILL
XFILL_2__14537_ gnd vdd FILL
XFILL_0__15716_ gnd vdd FILL
XFILL_2__11749_ gnd vdd FILL
XFILL_0__7426_ gnd vdd FILL
XFILL_4__12309_ gnd vdd FILL
XSFILL109400x71050 gnd vdd FILL
XFILL_3__15827_ gnd vdd FILL
XFILL_4__16077_ gnd vdd FILL
XFILL_5__14648_ gnd vdd FILL
XFILL_4__13289_ gnd vdd FILL
XFILL_1__12129_ gnd vdd FILL
XFILL_2__14468_ gnd vdd FILL
XFILL_0__15647_ gnd vdd FILL
XFILL_0__12859_ gnd vdd FILL
XFILL_0__7357_ gnd vdd FILL
XSFILL79320x53050 gnd vdd FILL
XFILL_4__15028_ gnd vdd FILL
XFILL_5__14579_ gnd vdd FILL
XFILL_2__16207_ gnd vdd FILL
XSFILL3560x79050 gnd vdd FILL
XFILL_2__13419_ gnd vdd FILL
XFILL_3__7066_ gnd vdd FILL
X_7985_ _7983_/Y _8006_/B _7985_/C gnd _8041_/D vdd OAI21X1
XFILL_3__15758_ gnd vdd FILL
XFILL_2__14399_ gnd vdd FILL
XFILL_0__15578_ gnd vdd FILL
XFILL_5__16318_ gnd vdd FILL
X_9724_ _9816_/Q gnd _9726_/A vdd INVX1
XFILL_0__7288_ gnd vdd FILL
XFILL_3__14709_ gnd vdd FILL
X_6936_ _6937_/B _6936_/B gnd _6937_/C vdd NAND2X1
XFILL_6__15869_ gnd vdd FILL
XSFILL114520x62050 gnd vdd FILL
XSFILL43560x32050 gnd vdd FILL
XSFILL8600x16050 gnd vdd FILL
XFILL_2__16138_ gnd vdd FILL
XFILL_3__15689_ gnd vdd FILL
XFILL_0__14529_ gnd vdd FILL
XSFILL44040x39050 gnd vdd FILL
XFILL_0__9027_ gnd vdd FILL
XSFILL104680x6050 gnd vdd FILL
X_9655_ _9655_/A _9613_/B _9655_/C gnd _9655_/Y vdd OAI21X1
XFILL_5__16249_ gnd vdd FILL
X_6867_ _6867_/A gnd memoryAddress[29] vdd BUFX2
XFILL_1__15819_ gnd vdd FILL
XFILL_2__16069_ gnd vdd FILL
X_8606_ _8607_/B _8606_/B gnd _8606_/Y vdd NAND2X1
X_9586_ _9586_/Q _8942_/CLK _9561_/R vdd _9586_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert601 gnd vdd FILL
XFILL_3__7968_ gnd vdd FILL
XFILL_5_BUFX2_insert612 gnd vdd FILL
XFILL_5_BUFX2_insert623 gnd vdd FILL
XFILL_5_BUFX2_insert634 gnd vdd FILL
X_8537_ _8447_/A _8537_/CLK _8542_/R vdd _8537_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert645 gnd vdd FILL
XFILL_1__9771_ gnd vdd FILL
XFILL_4__8500_ gnd vdd FILL
XFILL_5_BUFX2_insert656 gnd vdd FILL
XFILL_3__6919_ gnd vdd FILL
XFILL_1__6983_ gnd vdd FILL
XSFILL38920x19050 gnd vdd FILL
XFILL_4__9480_ gnd vdd FILL
XFILL112440x26050 gnd vdd FILL
XFILL_5_BUFX2_insert667 gnd vdd FILL
XFILL_1__8722_ gnd vdd FILL
XFILL_0__9929_ gnd vdd FILL
XFILL_5_BUFX2_insert678 gnd vdd FILL
XFILL_5_BUFX2_insert689 gnd vdd FILL
X_8468_ _8544_/Q gnd _8470_/A vdd INVX1
XFILL_3__9638_ gnd vdd FILL
XSFILL23720x61050 gnd vdd FILL
XSFILL39000x28050 gnd vdd FILL
X_7419_ _7417_/Y _7470_/B _7419_/C gnd _7511_/D vdd OAI21X1
XFILL_1__8653_ gnd vdd FILL
X_8399_ _8397_/Y _8360_/B _8399_/C gnd _8399_/Y vdd OAI21X1
XSFILL8600x7050 gnd vdd FILL
XFILL_4__8362_ gnd vdd FILL
XFILL_1__7604_ gnd vdd FILL
XFILL_2_CLKBUF1_insert204 gnd vdd FILL
XFILL_1__8584_ gnd vdd FILL
XFILL_4__7313_ gnd vdd FILL
XFILL_2_CLKBUF1_insert215 gnd vdd FILL
X_11020_ _12242_/Y _12135_/Y gnd _11020_/Y vdd NOR2X1
XSFILL114600x42050 gnd vdd FILL
XFILL_4__7244_ gnd vdd FILL
XFILL_1__7466_ gnd vdd FILL
XFILL_2_BUFX2_insert502 gnd vdd FILL
XFILL_4__7175_ gnd vdd FILL
XFILL_2_BUFX2_insert513 gnd vdd FILL
X_12971_ _12969_/Y vdd _12971_/C gnd _13053_/D vdd OAI21X1
XFILL_2_BUFX2_insert524 gnd vdd FILL
XFILL_2_BUFX2_insert535 gnd vdd FILL
XFILL_2_BUFX2_insert546 gnd vdd FILL
X_14710_ _7536_/Q gnd _14711_/A vdd INVX1
X_11922_ _11920_/Y _11921_/A _11922_/C gnd _6849_/A vdd OAI21X1
XFILL_2_BUFX2_insert557 gnd vdd FILL
X_15690_ _15690_/A _15690_/B gnd _15691_/A vdd NOR2X1
XFILL_2_BUFX2_insert568 gnd vdd FILL
XFILL_1__9136_ gnd vdd FILL
XFILL_2_BUFX2_insert579 gnd vdd FILL
X_14641_ _9022_/A gnd _14641_/Y vdd INVX1
XSFILL23800x41050 gnd vdd FILL
X_11853_ _11754_/A _11800_/A _11853_/C gnd _11853_/Y vdd NAND3X1
XFILL_6_BUFX2_insert1032 gnd vdd FILL
XFILL_5__6870_ gnd vdd FILL
X_10804_ _10804_/A _10822_/B _10803_/Y gnd _10858_/D vdd OAI21X1
X_14572_ _7277_/Q _14458_/C _14572_/C _10861_/Q gnd _14580_/B vdd AOI22X1
XFILL_2__8900_ gnd vdd FILL
XFILL_1__8018_ gnd vdd FILL
X_11784_ _11784_/A _11783_/Y _11784_/C gnd _12458_/B vdd NAND3X1
XFILL_2__9880_ gnd vdd FILL
XSFILL3720x39050 gnd vdd FILL
XBUFX2_insert501 BUFX2_insert559/A gnd _9069_/R vdd BUFX2
X_16311_ _16311_/A _14973_/Y _15025_/B _16310_/Y gnd _16311_/Y vdd OAI22X1
X_13523_ _13523_/A gnd _13525_/D vdd INVX1
XBUFX2_insert512 BUFX2_insert524/A gnd _7515_/R vdd BUFX2
XBUFX2_insert523 BUFX2_insert518/A gnd _9306_/R vdd BUFX2
XFILL_5__10260_ gnd vdd FILL
XSFILL38840x1050 gnd vdd FILL
X_10735_ _14689_/B _7647_/CLK _7775_/R vdd _10691_/Y gnd vdd DFFSR
XFILL_2__8831_ gnd vdd FILL
XBUFX2_insert534 BUFX2_insert570/A gnd _13199_/R vdd BUFX2
XFILL_4__10990_ gnd vdd FILL
XBUFX2_insert545 BUFX2_insert600/A gnd _13180_/R vdd BUFX2
XFILL_6_BUFX2_insert490 gnd vdd FILL
XSFILL94360x27050 gnd vdd FILL
XFILL_4__9747_ gnd vdd FILL
X_16242_ _16242_/A _16242_/B gnd _16243_/A vdd NAND2X1
XBUFX2_insert556 BUFX2_insert556/A gnd _8166_/R vdd BUFX2
XFILL_4__6959_ gnd vdd FILL
XBUFX2_insert567 BUFX2_insert607/A gnd _9692_/R vdd BUFX2
X_13454_ _13372_/A _13407_/Y _13465_/C gnd _13454_/Y vdd NAND3X1
X_10666_ _10615_/B _8874_/B gnd _10667_/C vdd NAND2X1
XFILL_5__10191_ gnd vdd FILL
XBUFX2_insert578 BUFX2_insert570/A gnd _7133_/R vdd BUFX2
XFILL_3__11370_ gnd vdd FILL
XFILL_2__8762_ gnd vdd FILL
XBUFX2_insert589 BUFX2_insert496/A gnd _8664_/R vdd BUFX2
XSFILL78680x81050 gnd vdd FILL
XFILL_0__11190_ gnd vdd FILL
XFILL_4__9678_ gnd vdd FILL
XFILL_5__8471_ gnd vdd FILL
X_12405_ _12403_/Y _12419_/A _12405_/C gnd _12405_/Y vdd OAI21X1
X_16173_ _7282_/Q gnd _16174_/A vdd INVX1
X_13385_ _8790_/Q gnd _14993_/A vdd INVX1
XFILL_3__10321_ gnd vdd FILL
XFILL_4__12660_ gnd vdd FILL
X_10597_ _10531_/A _8046_/CLK _9692_/R vdd _10597_/D gnd vdd DFFSR
XFILL_2__7713_ gnd vdd FILL
XFILL_1__11500_ gnd vdd FILL
XSFILL103720x46050 gnd vdd FILL
XFILL_0__10141_ gnd vdd FILL
XFILL_4__8629_ gnd vdd FILL
XFILL_1__12480_ gnd vdd FILL
XFILL_5__7422_ gnd vdd FILL
X_15124_ _15124_/A _15124_/B gnd _15125_/B vdd NOR2X1
XFILL_3__13040_ gnd vdd FILL
X_12336_ _12216_/B _12297_/D _12300_/C gnd _12338_/B vdd NAND3X1
XFILL_4__11611_ gnd vdd FILL
XFILL_5__13950_ gnd vdd FILL
XFILL_3__10252_ gnd vdd FILL
XFILL_4_BUFX2_insert1091 gnd vdd FILL
XSFILL104360x12050 gnd vdd FILL
XFILL_4__12591_ gnd vdd FILL
XFILL_1__11431_ gnd vdd FILL
XFILL_2__10982_ gnd vdd FILL
XFILL_2__13770_ gnd vdd FILL
XFILL_6__13151_ gnd vdd FILL
XFILL_5__7353_ gnd vdd FILL
X_15055_ _15064_/A _16037_/B _15061_/C gnd _15055_/Y vdd NAND3X1
XFILL_5__12901_ gnd vdd FILL
XFILL_4__14330_ gnd vdd FILL
X_12267_ _12255_/A gnd _12255_/C gnd _12267_/Y vdd NAND3X1
XFILL_5__13881_ gnd vdd FILL
XFILL_4__11542_ gnd vdd FILL
XFILL_2__12721_ gnd vdd FILL
XFILL_1__14150_ gnd vdd FILL
XFILL_3__10183_ gnd vdd FILL
XFILL_0__13900_ gnd vdd FILL
XFILL_2__7575_ gnd vdd FILL
XFILL_1__11362_ gnd vdd FILL
XFILL_0__14880_ gnd vdd FILL
XSFILL74520x56050 gnd vdd FILL
X_14006_ _7703_/A gnd _15498_/B vdd INVX1
X_11218_ _11215_/Y _11218_/B gnd _11762_/B vdd NAND2X1
XFILL_5__15620_ gnd vdd FILL
XFILL_5__12832_ gnd vdd FILL
XFILL_4__14261_ gnd vdd FILL
XFILL_1__13101_ gnd vdd FILL
XSFILL59080x55050 gnd vdd FILL
X_12198_ _12198_/A _12201_/B _12198_/C gnd _12198_/Y vdd OAI21X1
XFILL_2__12652_ gnd vdd FILL
XFILL_1__10313_ gnd vdd FILL
XFILL_2__15440_ gnd vdd FILL
XFILL_4__11473_ gnd vdd FILL
XFILL_0__13831_ gnd vdd FILL
XFILL_5__9023_ gnd vdd FILL
XFILL_3__14991_ gnd vdd FILL
XFILL_1__14081_ gnd vdd FILL
XFILL_4__16000_ gnd vdd FILL
XSFILL99480x60050 gnd vdd FILL
XFILL_1__11293_ gnd vdd FILL
XFILL_4__13212_ gnd vdd FILL
X_11149_ _11149_/A _11133_/Y _11149_/C gnd _11150_/C vdd OAI21X1
XFILL_5__12763_ gnd vdd FILL
XFILL_5__15551_ gnd vdd FILL
XFILL_4__10424_ gnd vdd FILL
XFILL_4__14192_ gnd vdd FILL
XFILL_1__13032_ gnd vdd FILL
XFILL_2__11603_ gnd vdd FILL
XFILL_2__9245_ gnd vdd FILL
XFILL_3__13942_ gnd vdd FILL
XFILL_2__15371_ gnd vdd FILL
XFILL_2__12583_ gnd vdd FILL
XFILL_1__10244_ gnd vdd FILL
XFILL_0__13762_ gnd vdd FILL
XFILL_3_BUFX2_insert380 gnd vdd FILL
XFILL_0__10974_ gnd vdd FILL
XFILL_3_BUFX2_insert391 gnd vdd FILL
XFILL_5__14502_ gnd vdd FILL
XFILL_0__8260_ gnd vdd FILL
XFILL_5__11714_ gnd vdd FILL
XFILL_4__13143_ gnd vdd FILL
X_15957_ _7916_/Q gnd _15957_/Y vdd INVX1
XFILL_5__15482_ gnd vdd FILL
XFILL_0__15501_ gnd vdd FILL
XFILL_2__14322_ gnd vdd FILL
XFILL_2__11534_ gnd vdd FILL
XFILL_3__13873_ gnd vdd FILL
XFILL_0__12713_ gnd vdd FILL
XFILL_1__10175_ gnd vdd FILL
XFILL_0__7211_ gnd vdd FILL
XFILL_0__13693_ gnd vdd FILL
X_14908_ _7632_/A _14145_/D _14739_/C _16246_/A gnd _14908_/Y vdd AOI22X1
XFILL_5__14433_ gnd vdd FILL
XFILL_0__8191_ gnd vdd FILL
XSFILL13800x73050 gnd vdd FILL
XFILL_3__15612_ gnd vdd FILL
XFILL_5__11645_ gnd vdd FILL
XFILL_2__8127_ gnd vdd FILL
XFILL_3__12824_ gnd vdd FILL
X_15888_ _15884_/Y _15887_/Y gnd _15888_/Y vdd NOR2X1
XFILL_2__14253_ gnd vdd FILL
XFILL_4__10286_ gnd vdd FILL
XFILL_0__15432_ gnd vdd FILL
XFILL_2__11465_ gnd vdd FILL
XFILL_0__12644_ gnd vdd FILL
XFILL_5__9925_ gnd vdd FILL
XFILL_1__14983_ gnd vdd FILL
X_14839_ _10189_/A gnd _14839_/Y vdd INVX1
XFILL_4__12025_ gnd vdd FILL
XFILL_5__14364_ gnd vdd FILL
X_7770_ _7682_/A _9818_/CLK _9441_/R vdd _7770_/D gnd vdd DFFSR
XFILL_3__15543_ gnd vdd FILL
XFILL_2__10416_ gnd vdd FILL
XFILL_5__11576_ gnd vdd FILL
XFILL_3__12755_ gnd vdd FILL
XFILL_2__14184_ gnd vdd FILL
XFILL_2__8058_ gnd vdd FILL
XFILL_0__15363_ gnd vdd FILL
XFILL_2__11396_ gnd vdd FILL
XFILL_1__13934_ gnd vdd FILL
XFILL_5__13315_ gnd vdd FILL
XFILL_5__9856_ gnd vdd FILL
XFILL_0__12575_ gnd vdd FILL
XFILL_5__16103_ gnd vdd FILL
XFILL_6__15654_ gnd vdd FILL
XFILL_0__7073_ gnd vdd FILL
XFILL_5__10527_ gnd vdd FILL
XFILL_2__13135_ gnd vdd FILL
XFILL_3__11706_ gnd vdd FILL
XFILL_5__14295_ gnd vdd FILL
XFILL_0__14314_ gnd vdd FILL
XFILL_3__15474_ gnd vdd FILL
XFILL_3__8871_ gnd vdd FILL
XSFILL84360x59050 gnd vdd FILL
XFILL_0__11526_ gnd vdd FILL
XFILL_1__13865_ gnd vdd FILL
XFILL_6__14605_ gnd vdd FILL
XFILL_5__16034_ gnd vdd FILL
XFILL_0__15294_ gnd vdd FILL
XFILL_5__9787_ gnd vdd FILL
XFILL_5__13246_ gnd vdd FILL
X_9440_ _9440_/Q _7535_/CLK _7648_/R vdd _9366_/Y gnd vdd DFFSR
XFILL_3__14425_ gnd vdd FILL
XFILL_3__7822_ gnd vdd FILL
XFILL_4__13976_ gnd vdd FILL
XFILL_4_CLKBUF1_insert170 gnd vdd FILL
XFILL_3__11637_ gnd vdd FILL
XFILL_1__15604_ gnd vdd FILL
XFILL_4_CLKBUF1_insert181 gnd vdd FILL
XFILL_0__14245_ gnd vdd FILL
XFILL_2__10278_ gnd vdd FILL
XFILL_1__13796_ gnd vdd FILL
XFILL_5__8738_ gnd vdd FILL
XFILL_0__11457_ gnd vdd FILL
XFILL_4_CLKBUF1_insert192 gnd vdd FILL
XFILL_4__15715_ gnd vdd FILL
XFILL_2__12017_ gnd vdd FILL
X_9371_ _9372_/B _9371_/B gnd _9371_/Y vdd NAND2X1
XFILL_6__11748_ gnd vdd FILL
XFILL_3__14356_ gnd vdd FILL
XFILL_5__10389_ gnd vdd FILL
XFILL_1__12747_ gnd vdd FILL
XFILL_0__10408_ gnd vdd FILL
XFILL_1__15535_ gnd vdd FILL
XFILL_3__11568_ gnd vdd FILL
XFILL_3__7753_ gnd vdd FILL
XFILL_0_BUFX2_insert270 gnd vdd FILL
XFILL_0__14176_ gnd vdd FILL
X_8322_ _8410_/Q gnd _8322_/Y vdd INVX1
XFILL_0_BUFX2_insert281 gnd vdd FILL
XFILL_5__12128_ gnd vdd FILL
XFILL_0__11388_ gnd vdd FILL
XFILL_3__13307_ gnd vdd FILL
XFILL_0_BUFX2_insert292 gnd vdd FILL
XFILL_6__14467_ gnd vdd FILL
XFILL_4__15646_ gnd vdd FILL
XFILL_0__7975_ gnd vdd FILL
XFILL_3__10519_ gnd vdd FILL
XFILL_4__12858_ gnd vdd FILL
XFILL_4_BUFX2_insert608 gnd vdd FILL
XFILL_0__13127_ gnd vdd FILL
XFILL_3__14287_ gnd vdd FILL
XFILL_6__16206_ gnd vdd FILL
XFILL_3__7684_ gnd vdd FILL
XFILL_3__11499_ gnd vdd FILL
XFILL_1__15466_ gnd vdd FILL
XFILL_6__13418_ gnd vdd FILL
XFILL_4_BUFX2_insert619 gnd vdd FILL
XFILL_0__6926_ gnd vdd FILL
X_8253_ _8251_/Y _8249_/A _8253_/C gnd _8253_/Y vdd OAI21X1
XFILL_3__16026_ gnd vdd FILL
XFILL_5__12059_ gnd vdd FILL
XFILL_4__11809_ gnd vdd FILL
XFILL_3__13238_ gnd vdd FILL
XFILL_3__9423_ gnd vdd FILL
XFILL_4__15577_ gnd vdd FILL
XFILL_4__12789_ gnd vdd FILL
XFILL_1__11629_ gnd vdd FILL
XFILL_1__14417_ gnd vdd FILL
XFILL_1__15397_ gnd vdd FILL
XSFILL114600x9050 gnd vdd FILL
XFILL_2__13968_ gnd vdd FILL
X_7204_ _7184_/B _8868_/B gnd _7205_/C vdd NAND2X1
XSFILL79320x48050 gnd vdd FILL
XFILL_4__14528_ gnd vdd FILL
XFILL_0__9645_ gnd vdd FILL
XFILL_2__15707_ gnd vdd FILL
X_8184_ _8182_/Y _8232_/B _8184_/C gnd _8278_/D vdd OAI21X1
XFILL_0__6857_ gnd vdd FILL
XFILL_3__9354_ gnd vdd FILL
XFILL_2_BUFX2_insert30 gnd vdd FILL
XFILL_3__13169_ gnd vdd FILL
XFILL_0__12009_ gnd vdd FILL
XFILL_1__14348_ gnd vdd FILL
XFILL_2_BUFX2_insert41 gnd vdd FILL
XFILL_2_BUFX2_insert52 gnd vdd FILL
XFILL_2__13899_ gnd vdd FILL
XFILL_5__15818_ gnd vdd FILL
XFILL_2_BUFX2_insert63 gnd vdd FILL
XFILL_6__16068_ gnd vdd FILL
X_7135_ _7135_/Q _7156_/CLK _7775_/R vdd _7059_/Y gnd vdd DFFSR
XFILL_2_BUFX2_insert74 gnd vdd FILL
XFILL_4__14459_ gnd vdd FILL
XSFILL114520x57050 gnd vdd FILL
XFILL_2__15638_ gnd vdd FILL
XFILL_6__8014_ gnd vdd FILL
XFILL_2_BUFX2_insert85 gnd vdd FILL
XFILL_3__9285_ gnd vdd FILL
XFILL_1__14279_ gnd vdd FILL
XFILL_2_BUFX2_insert96 gnd vdd FILL
XFILL_1__7320_ gnd vdd FILL
XFILL_0__8527_ gnd vdd FILL
X_7066_ _7138_/Q gnd _7066_/Y vdd INVX1
XFILL_5__15749_ gnd vdd FILL
XFILL_1__16018_ gnd vdd FILL
XFILL_3__8236_ gnd vdd FILL
XFILL_2__15569_ gnd vdd FILL
XFILL_4__16129_ gnd vdd FILL
XFILL_1__7251_ gnd vdd FILL
XFILL_0__8458_ gnd vdd FILL
XSFILL59240x15050 gnd vdd FILL
XFILL_1__7182_ gnd vdd FILL
XFILL_0__8389_ gnd vdd FILL
XFILL_3__7118_ gnd vdd FILL
XFILL111960x14050 gnd vdd FILL
XFILL_3__8098_ gnd vdd FILL
XFILL_4__8980_ gnd vdd FILL
XFILL_1_BUFX2_insert509 gnd vdd FILL
XFILL_6__9896_ gnd vdd FILL
X_7968_ _8036_/Q gnd _7970_/A vdd INVX1
XSFILL23720x56050 gnd vdd FILL
XFILL_3__7049_ gnd vdd FILL
XFILL_4__7931_ gnd vdd FILL
XFILL_6__8847_ gnd vdd FILL
X_9707_ _9653_/A _9707_/CLK _8819_/R vdd _9655_/Y gnd vdd DFFSR
X_6919_ _6919_/A _6955_/B _6918_/Y gnd _6919_/Y vdd OAI21X1
X_7899_ _7813_/A _8792_/CLK _7896_/R vdd _7815_/Y gnd vdd DFFSR
XFILL_4__7862_ gnd vdd FILL
XFILL_4__9601_ gnd vdd FILL
X_9638_ _9702_/Q gnd _9640_/A vdd INVX1
XSFILL100120x5050 gnd vdd FILL
XSFILL64200x70050 gnd vdd FILL
X_10520_ _10500_/B _8600_/B gnd _10520_/Y vdd NAND2X1
XSFILL114600x37050 gnd vdd FILL
XFILL_5_BUFX2_insert420 gnd vdd FILL
X_9569_ _9569_/Q _9707_/CLK _8801_/R vdd _9497_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert431 gnd vdd FILL
XFILL_4__9532_ gnd vdd FILL
XFILL_5_BUFX2_insert442 gnd vdd FILL
XFILL_5_BUFX2_insert453 gnd vdd FILL
X_10451_ _14942_/A gnd _10451_/Y vdd INVX1
XFILL_5_BUFX2_insert464 gnd vdd FILL
XFILL_1__9754_ gnd vdd FILL
XFILL_5_BUFX2_insert475 gnd vdd FILL
XSFILL69080x18050 gnd vdd FILL
XFILL_1__6966_ gnd vdd FILL
XFILL_4__9463_ gnd vdd FILL
XFILL_5_BUFX2_insert486 gnd vdd FILL
X_13170_ _13173_/A _12110_/Y gnd _13171_/C vdd NAND2X1
XFILL_5_BUFX2_insert497 gnd vdd FILL
XFILL_1__8705_ gnd vdd FILL
X_10382_ _10462_/Q gnd _10382_/Y vdd INVX1
XSFILL109480x2050 gnd vdd FILL
XSFILL84120x21050 gnd vdd FILL
XFILL_1__9685_ gnd vdd FILL
X_12121_ _13085_/A gnd _12123_/A vdd INVX1
XSFILL104280x27050 gnd vdd FILL
XFILL_1__6897_ gnd vdd FILL
XFILL_4__9394_ gnd vdd FILL
XFILL_1__8636_ gnd vdd FILL
XFILL_4__8345_ gnd vdd FILL
X_12052_ _12028_/A _11882_/B _12024_/C gnd _12054_/B vdd NAND3X1
XFILL_2__7360_ gnd vdd FILL
XSFILL23800x36050 gnd vdd FILL
XFILL_1__8567_ gnd vdd FILL
X_11003_ _12230_/Y _12126_/Y gnd _11003_/Y vdd NAND2X1
XSFILL63400x22050 gnd vdd FILL
XSFILL33960x80050 gnd vdd FILL
XFILL_4__8276_ gnd vdd FILL
XFILL_2__7291_ gnd vdd FILL
XSFILL74040x73050 gnd vdd FILL
XFILL_4__7227_ gnd vdd FILL
XFILL_1__8498_ gnd vdd FILL
X_15811_ _15811_/A _15788_/Y _15811_/C gnd _15812_/B vdd NOR3X1
XFILL_2__9030_ gnd vdd FILL
XFILL_2_BUFX2_insert310 gnd vdd FILL
XFILL_2_BUFX2_insert321 gnd vdd FILL
XFILL_1__7449_ gnd vdd FILL
XFILL_4__7158_ gnd vdd FILL
XFILL_2_BUFX2_insert332 gnd vdd FILL
XFILL_2_BUFX2_insert343 gnd vdd FILL
X_15742_ _7271_/Q _15177_/B _15742_/C gnd _15742_/Y vdd AOI21X1
XFILL_4__10140_ gnd vdd FILL
XFILL_2_BUFX2_insert354 gnd vdd FILL
X_12954_ _6871_/A gnd _12954_/Y vdd INVX1
XFILL_2_BUFX2_insert365 gnd vdd FILL
XFILL_3__10870_ gnd vdd FILL
XFILL_2_BUFX2_insert376 gnd vdd FILL
XFILL_5__7971_ gnd vdd FILL
X_11905_ _13097_/A gnd _11907_/A vdd INVX1
XFILL_2_BUFX2_insert387 gnd vdd FILL
XFILL_4__7089_ gnd vdd FILL
XFILL_5__11430_ gnd vdd FILL
XFILL_0__10690_ gnd vdd FILL
XFILL_6__10981_ gnd vdd FILL
X_15673_ _10659_/A gnd _15673_/Y vdd INVX1
XFILL_2_BUFX2_insert398 gnd vdd FILL
XFILL_1__9119_ gnd vdd FILL
XFILL_2__11250_ gnd vdd FILL
X_12885_ _12883_/Y vdd _12885_/C gnd _12939_/D vdd OAI21X1
XFILL_5__6922_ gnd vdd FILL
XFILL_1__11980_ gnd vdd FILL
X_14624_ _14623_/Y _13882_/B _13633_/C _14622_/Y gnd _14624_/Y vdd OAI22X1
XFILL_5__11361_ gnd vdd FILL
X_11836_ _11835_/A _11427_/A _11836_/C gnd _11836_/Y vdd OAI21X1
XFILL_2__9932_ gnd vdd FILL
XFILL_1__10931_ gnd vdd FILL
XFILL_2__11181_ gnd vdd FILL
XFILL_5__13100_ gnd vdd FILL
XFILL_0__12360_ gnd vdd FILL
XFILL_5__9641_ gnd vdd FILL
XFILL_5__6853_ gnd vdd FILL
XFILL_5__10312_ gnd vdd FILL
X_14555_ _14553_/Y _14555_/B _14555_/C _14554_/Y gnd _14555_/Y vdd OAI22X1
XFILL_4__13830_ gnd vdd FILL
XFILL_5__14080_ gnd vdd FILL
XFILL_5__11292_ gnd vdd FILL
XFILL_2__10132_ gnd vdd FILL
X_11767_ _11253_/Y gnd _11767_/Y vdd INVX1
XFILL_1__13650_ gnd vdd FILL
XBUFX2_insert320 _15000_/Y gnd _15394_/C vdd BUFX2
XFILL_3__12471_ gnd vdd FILL
XFILL_2__9863_ gnd vdd FILL
XFILL_0__11311_ gnd vdd FILL
XBUFX2_insert331 _12405_/Y gnd _9779_/B vdd BUFX2
XFILL_5__13031_ gnd vdd FILL
XFILL_0__12291_ gnd vdd FILL
XBUFX2_insert342 _12396_/Y gnd _7594_/B vdd BUFX2
X_13506_ _8023_/Q gnd _13507_/A vdd INVX1
XBUFX2_insert353 _13306_/Y gnd _7937_/B vdd BUFX2
X_10718_ _10638_/A _7790_/CLK _9561_/R vdd _10718_/D gnd vdd DFFSR
XFILL_3__14210_ gnd vdd FILL
XFILL_5__10243_ gnd vdd FILL
XFILL_1__12601_ gnd vdd FILL
X_14486_ _14484_/Y _14567_/A _14849_/B _14485_/Y gnd _14486_/Y vdd OAI22X1
XFILL_4__13761_ gnd vdd FILL
XFILL_3__11422_ gnd vdd FILL
XFILL_4__10973_ gnd vdd FILL
XFILL_2__10063_ gnd vdd FILL
XFILL_3__15190_ gnd vdd FILL
XFILL_0__14030_ gnd vdd FILL
XBUFX2_insert364 _13487_/Y gnd _14847_/C vdd BUFX2
XFILL_2__14940_ gnd vdd FILL
X_11698_ _11698_/A _11695_/Y _11697_/Y gnd _11698_/Y vdd NAND3X1
XFILL_5__8523_ gnd vdd FILL
XBUFX2_insert375 _13338_/Y gnd _9529_/A vdd BUFX2
XFILL_1__13581_ gnd vdd FILL
XFILL_2__9794_ gnd vdd FILL
XFILL_0__11242_ gnd vdd FILL
X_16225_ _16224_/Y _15972_/B _16225_/C _14873_/Y gnd _16225_/Y vdd OAI22X1
XSFILL99480x55050 gnd vdd FILL
XFILL_4__15500_ gnd vdd FILL
XBUFX2_insert386 _13331_/Y gnd _9164_/B vdd BUFX2
XFILL_5_CLKBUF1_insert210 gnd vdd FILL
XFILL_1__10793_ gnd vdd FILL
XFILL_6__11533_ gnd vdd FILL
XBUFX2_insert397 _13293_/Y gnd _7592_/B vdd BUFX2
XFILL_4__12712_ gnd vdd FILL
X_13437_ _13423_/A _13404_/B _13407_/Y gnd _13868_/B vdd NAND3X1
XSFILL49320x27050 gnd vdd FILL
XFILL_5_CLKBUF1_insert221 gnd vdd FILL
XFILL_5__10174_ gnd vdd FILL
XSFILL74120x53050 gnd vdd FILL
XFILL_3__14141_ gnd vdd FILL
X_10649_ _10649_/A _10658_/B _10649_/C gnd _10721_/D vdd OAI21X1
XFILL_1__15320_ gnd vdd FILL
XFILL_1__12532_ gnd vdd FILL
XFILL_2__8745_ gnd vdd FILL
XFILL_4__13692_ gnd vdd FILL
XFILL_3__11353_ gnd vdd FILL
XFILL_2__14871_ gnd vdd FILL
XFILL_5__8454_ gnd vdd FILL
XFILL_0__11173_ gnd vdd FILL
XFILL_6__14252_ gnd vdd FILL
XFILL_4__15431_ gnd vdd FILL
X_16156_ _16156_/A _16156_/B gnd _16162_/B vdd NOR2X1
XFILL_3__10304_ gnd vdd FILL
XFILL_4__12643_ gnd vdd FILL
X_13368_ _11881_/A _12809_/Q gnd _13398_/A vdd AND2X2
XFILL_0__7760_ gnd vdd FILL
XFILL_2__13822_ gnd vdd FILL
XFILL_1__15251_ gnd vdd FILL
XFILL_5__14982_ gnd vdd FILL
XFILL_3__14072_ gnd vdd FILL
XFILL_3__11284_ gnd vdd FILL
XFILL_0__10124_ gnd vdd FILL
XFILL_1__12463_ gnd vdd FILL
XFILL_0__15981_ gnd vdd FILL
X_15107_ _7127_/Q gnd _15107_/Y vdd INVX1
X_12319_ _12327_/A gnd _12319_/C gnd _12322_/A vdd NAND3X1
XFILL_5__8385_ gnd vdd FILL
XSFILL99160x8050 gnd vdd FILL
XSFILL53960x11050 gnd vdd FILL
XFILL_0__7691_ gnd vdd FILL
XFILL_1__14202_ gnd vdd FILL
XFILL_4__15362_ gnd vdd FILL
XFILL_3__13023_ gnd vdd FILL
XFILL_6__11395_ gnd vdd FILL
XFILL_3__10235_ gnd vdd FILL
XFILL_5__13933_ gnd vdd FILL
X_16087_ _16086_/Y _16087_/B _14402_/C gnd _12899_/B vdd AOI21X1
X_13299_ _13299_/A gnd _13300_/B vdd INVX2
XFILL_4__12574_ gnd vdd FILL
XFILL_2__7627_ gnd vdd FILL
XSFILL109480x40050 gnd vdd FILL
XFILL_1__11414_ gnd vdd FILL
XFILL_1__15182_ gnd vdd FILL
XFILL_2__13753_ gnd vdd FILL
XFILL_2__10965_ gnd vdd FILL
XFILL_5__7336_ gnd vdd FILL
XFILL_1__12394_ gnd vdd FILL
XFILL_0__14932_ gnd vdd FILL
XFILL_0__10055_ gnd vdd FILL
X_15038_ _15244_/C _16037_/B _15061_/C gnd _15038_/Y vdd NAND3X1
XFILL_4__14313_ gnd vdd FILL
XFILL_4__11525_ gnd vdd FILL
XFILL_2__12704_ gnd vdd FILL
XFILL_3__10166_ gnd vdd FILL
XFILL_5__13864_ gnd vdd FILL
XFILL_1__14133_ gnd vdd FILL
XFILL_4__15293_ gnd vdd FILL
XFILL_2__7558_ gnd vdd FILL
XFILL_1__11345_ gnd vdd FILL
XFILL_0__14863_ gnd vdd FILL
XSFILL113960x65050 gnd vdd FILL
XFILL_2__13684_ gnd vdd FILL
XFILL_2__10896_ gnd vdd FILL
XFILL_5__15603_ gnd vdd FILL
XFILL_4__14244_ gnd vdd FILL
XFILL_0__9361_ gnd vdd FILL
XFILL_5__13795_ gnd vdd FILL
XFILL_4__11456_ gnd vdd FILL
XFILL_2__15423_ gnd vdd FILL
XFILL_2__12635_ gnd vdd FILL
XFILL_0__13814_ gnd vdd FILL
XFILL_1__14064_ gnd vdd FILL
XFILL_5__9006_ gnd vdd FILL
XFILL_3__14974_ gnd vdd FILL
XFILL_1__11276_ gnd vdd FILL
XFILL_2__7489_ gnd vdd FILL
XFILL_0__14794_ gnd vdd FILL
XFILL_0__8312_ gnd vdd FILL
XFILL_4__10407_ gnd vdd FILL
XFILL_5__12746_ gnd vdd FILL
XFILL_5__15534_ gnd vdd FILL
XFILL_0__9292_ gnd vdd FILL
XFILL_5__7198_ gnd vdd FILL
XFILL_4__14175_ gnd vdd FILL
XFILL_2__9228_ gnd vdd FILL
XFILL_1__13015_ gnd vdd FILL
XSFILL43880x63050 gnd vdd FILL
X_8940_ _8888_/A _9958_/CLK _8929_/R vdd _8940_/D gnd vdd DFFSR
XFILL_3__8021_ gnd vdd FILL
XFILL_3__13925_ gnd vdd FILL
XFILL_2__15354_ gnd vdd FILL
XFILL_4__11387_ gnd vdd FILL
XFILL_0__13745_ gnd vdd FILL
XFILL_0__10957_ gnd vdd FILL
XFILL_0__8243_ gnd vdd FILL
XFILL_4__13126_ gnd vdd FILL
X_8871_ _8896_/B _7847_/B gnd _8871_/Y vdd NAND2X1
XFILL_2__14305_ gnd vdd FILL
XFILL_5__15465_ gnd vdd FILL
XFILL_3__13856_ gnd vdd FILL
XFILL_2__11517_ gnd vdd FILL
XFILL_2__9159_ gnd vdd FILL
XFILL_2__12497_ gnd vdd FILL
XFILL_1__10158_ gnd vdd FILL
XFILL_2__15285_ gnd vdd FILL
XFILL_0__13676_ gnd vdd FILL
XSFILL74200x33050 gnd vdd FILL
X_7822_ _7902_/Q gnd _7822_/Y vdd INVX1
XFILL_0__10888_ gnd vdd FILL
XFILL_5__11628_ gnd vdd FILL
XFILL_5__14416_ gnd vdd FILL
XFILL_5__15396_ gnd vdd FILL
XFILL_2__14236_ gnd vdd FILL
XFILL_4__10269_ gnd vdd FILL
XFILL_2__11448_ gnd vdd FILL
XFILL_0__15415_ gnd vdd FILL
XFILL_0__12627_ gnd vdd FILL
XFILL_3__13787_ gnd vdd FILL
XFILL_0__16395_ gnd vdd FILL
XFILL_0__7125_ gnd vdd FILL
XFILL_1__14966_ gnd vdd FILL
XFILL_5__9908_ gnd vdd FILL
XFILL_3__10999_ gnd vdd FILL
XFILL_4__12008_ gnd vdd FILL
XFILL_5__14347_ gnd vdd FILL
XFILL_6__12918_ gnd vdd FILL
XFILL_3__15526_ gnd vdd FILL
XFILL_5__11559_ gnd vdd FILL
X_7753_ _7753_/A _7753_/B _7753_/C gnd _7753_/Y vdd OAI21X1
XFILL_3__12738_ gnd vdd FILL
XFILL_0__15346_ gnd vdd FILL
XFILL_2__14167_ gnd vdd FILL
XFILL112440x3050 gnd vdd FILL
XFILL_1__13917_ gnd vdd FILL
XFILL_2__11379_ gnd vdd FILL
XFILL_0__7056_ gnd vdd FILL
XSFILL78840x36050 gnd vdd FILL
XFILL_1__14897_ gnd vdd FILL
XFILL_5__14278_ gnd vdd FILL
X_7684_ _7682_/Y _7684_/B _7684_/C gnd _7770_/D vdd OAI21X1
XFILL_2__13118_ gnd vdd FILL
XFILL_3__15457_ gnd vdd FILL
XFILL_3__8854_ gnd vdd FILL
XFILL_0__11509_ gnd vdd FILL
XFILL_2__14098_ gnd vdd FILL
XFILL_1__13848_ gnd vdd FILL
XFILL_0__15277_ gnd vdd FILL
XFILL_5__13229_ gnd vdd FILL
XFILL_5__16017_ gnd vdd FILL
X_9423_ _9421_/Y _9356_/A _9422_/Y gnd _9459_/D vdd OAI21X1
XFILL_0__12489_ gnd vdd FILL
XFILL_3__14408_ gnd vdd FILL
XFILL_3__7805_ gnd vdd FILL
XFILL_4__13959_ gnd vdd FILL
XFILL_3__15388_ gnd vdd FILL
XFILL_0__14228_ gnd vdd FILL
XSFILL74120x5050 gnd vdd FILL
XFILL_3__8785_ gnd vdd FILL
XFILL_1__13779_ gnd vdd FILL
X_9354_ _9354_/A _9420_/B _9354_/C gnd _9436_/D vdd OAI21X1
XFILL_3__14339_ gnd vdd FILL
XFILL_1__15518_ gnd vdd FILL
XFILL_3__7736_ gnd vdd FILL
XFILL_0__14159_ gnd vdd FILL
XFILL_4_BUFX2_insert405 gnd vdd FILL
XSFILL43960x43050 gnd vdd FILL
X_8305_ _8305_/Q _9205_/CLK _8433_/R vdd _8305_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert416 gnd vdd FILL
XFILL_4__15629_ gnd vdd FILL
X_9285_ _9240_/A _8005_/B gnd _9286_/C vdd NAND2X1
XFILL_4_BUFX2_insert427 gnd vdd FILL
XFILL_0__7958_ gnd vdd FILL
XFILL_4_BUFX2_insert438 gnd vdd FILL
XFILL_1__15449_ gnd vdd FILL
XFILL_4_BUFX2_insert449 gnd vdd FILL
XFILL_3__16009_ gnd vdd FILL
X_8236_ _8236_/A gnd _8238_/A vdd INVX1
XFILL_0__6909_ gnd vdd FILL
XFILL_3__9406_ gnd vdd FILL
XFILL_1__9470_ gnd vdd FILL
XSFILL44040x52050 gnd vdd FILL
XFILL_0__7889_ gnd vdd FILL
XFILL_3__7598_ gnd vdd FILL
XFILL_0__9628_ gnd vdd FILL
X_8167_ _8167_/Q _8679_/CLK _9959_/R vdd _8167_/D gnd vdd DFFSR
XFILL112440x50 gnd vdd FILL
XFILL_4__8130_ gnd vdd FILL
XFILL_3__9337_ gnd vdd FILL
X_7118_ _7100_/A _8910_/B gnd _7119_/C vdd NAND2X1
XFILL_1__8352_ gnd vdd FILL
XSFILL23880x10050 gnd vdd FILL
XFILL112040x18050 gnd vdd FILL
X_8098_ _8098_/A _8098_/B _8097_/Y gnd _8098_/Y vdd OAI21X1
XFILL_3__9268_ gnd vdd FILL
XFILL_4__8061_ gnd vdd FILL
XFILL111800x73050 gnd vdd FILL
XFILL_1__7303_ gnd vdd FILL
X_7049_ _7068_/B _9993_/B gnd _7050_/C vdd NAND2X1
XSFILL90040x55050 gnd vdd FILL
XFILL_3__8219_ gnd vdd FILL
XFILL_3_CLKBUF1_insert118 gnd vdd FILL
XSFILL64200x65050 gnd vdd FILL
XFILL_3_CLKBUF1_insert129 gnd vdd FILL
XFILL_5_CLKBUF1_insert1078 gnd vdd FILL
XFILL_1__7234_ gnd vdd FILL
XSFILL39000x41050 gnd vdd FILL
XFILL_1_BUFX2_insert306 gnd vdd FILL
XFILL_1__7165_ gnd vdd FILL
XFILL_1_BUFX2_insert317 gnd vdd FILL
XFILL_1_BUFX2_insert328 gnd vdd FILL
XFILL_4__8963_ gnd vdd FILL
XFILL_1_BUFX2_insert339 gnd vdd FILL
X_12670_ _12588_/A _12692_/CLK _12692_/R vdd _12670_/D gnd vdd DFFSR
XFILL_1__7096_ gnd vdd FILL
XFILL_4__8894_ gnd vdd FILL
XSFILL94280x60050 gnd vdd FILL
X_11621_ _11300_/A _11484_/B _11621_/C _11133_/Y gnd _11621_/Y vdd OAI22X1
XFILL_4__7845_ gnd vdd FILL
X_14340_ _14340_/A _14340_/B gnd _14340_/Y vdd NOR2X1
X_11552_ _11552_/A _11553_/B gnd _11856_/A vdd AND2X2
XFILL_2__6860_ gnd vdd FILL
X_10503_ _10503_/A _10539_/B _10503_/C gnd _10587_/D vdd OAI21X1
XFILL_1__9806_ gnd vdd FILL
X_11483_ _11174_/C _11226_/B _11483_/C gnd _11483_/Y vdd OAI21X1
X_14271_ _14270_/Y _14068_/C _14030_/C _14271_/D gnd _14271_/Y vdd OAI22X1
XFILL_5_BUFX2_insert250 gnd vdd FILL
XFILL_5_BUFX2_insert261 gnd vdd FILL
XFILL_4__9515_ gnd vdd FILL
XFILL_1__7998_ gnd vdd FILL
X_16010_ _15652_/A _9534_/A _9710_/Q _15652_/D gnd _16010_/Y vdd AOI22X1
XSFILL23400x33050 gnd vdd FILL
XFILL_5_BUFX2_insert272 gnd vdd FILL
X_13222_ _13209_/Y _13222_/B gnd _13244_/A vdd NOR2X1
XFILL_5_BUFX2_insert283 gnd vdd FILL
X_10434_ _10450_/B _6978_/B gnd _10434_/Y vdd NAND2X1
XSFILL89640x47050 gnd vdd FILL
XFILL_5_BUFX2_insert294 gnd vdd FILL
XFILL_1__9737_ gnd vdd FILL
XFILL_2__8530_ gnd vdd FILL
XFILL_1__6949_ gnd vdd FILL
X_13153_ _13151_/Y _13153_/B _13152_/Y gnd _13199_/D vdd OAI21X1
X_10365_ _10363_/B _8701_/B gnd _10366_/C vdd NAND2X1
XFILL_4_BUFX2_insert950 gnd vdd FILL
XFILL_2__8461_ gnd vdd FILL
XFILL_1__9668_ gnd vdd FILL
XFILL_4_BUFX2_insert961 gnd vdd FILL
XFILL_4_BUFX2_insert972 gnd vdd FILL
X_12104_ _12084_/A _11974_/A _12084_/C gnd _12106_/B vdd NAND3X1
XFILL_4__9377_ gnd vdd FILL
XFILL_5__10930_ gnd vdd FILL
XFILL_4_BUFX2_insert983 gnd vdd FILL
XFILL_3__10020_ gnd vdd FILL
X_13084_ _13082_/Y _13155_/A _13084_/C gnd _13176_/D vdd OAI21X1
XFILL_6__11180_ gnd vdd FILL
XFILL_4_BUFX2_insert994 gnd vdd FILL
X_10296_ _10348_/Q gnd _10298_/A vdd INVX1
XFILL_1__8619_ gnd vdd FILL
XSFILL3720x52050 gnd vdd FILL
XFILL_2__10750_ gnd vdd FILL
XFILL_1__9599_ gnd vdd FILL
XFILL_4__8328_ gnd vdd FILL
XFILL_5__7121_ gnd vdd FILL
XFILL_2__8392_ gnd vdd FILL
X_12035_ _12031_/A _12035_/B _12031_/C gnd _12038_/A vdd NAND3X1
XFILL_4__11310_ gnd vdd FILL
XSFILL28920x64050 gnd vdd FILL
XSFILL28120x45050 gnd vdd FILL
XFILL_2__7343_ gnd vdd FILL
XFILL_4__12290_ gnd vdd FILL
XFILL_1__11130_ gnd vdd FILL
XFILL_2__10681_ gnd vdd FILL
XFILL_5__12600_ gnd vdd FILL
XFILL_5__7052_ gnd vdd FILL
XFILL_0__11860_ gnd vdd FILL
XFILL_4__8259_ gnd vdd FILL
XFILL_6__10062_ gnd vdd FILL
XFILL_5__13580_ gnd vdd FILL
XFILL_4__11241_ gnd vdd FILL
XFILL_5__10792_ gnd vdd FILL
XFILL_2__12420_ gnd vdd FILL
XFILL_0__10811_ gnd vdd FILL
XFILL_3__11971_ gnd vdd FILL
XFILL_1__11061_ gnd vdd FILL
XSFILL29000x73050 gnd vdd FILL
XFILL_5__12531_ gnd vdd FILL
XFILL_0__11791_ gnd vdd FILL
XFILL_2__9013_ gnd vdd FILL
XFILL_3__13710_ gnd vdd FILL
XFILL_3__10922_ gnd vdd FILL
XFILL_2__12351_ gnd vdd FILL
X_13986_ _13986_/A _13982_/Y gnd _13986_/Y vdd NOR2X1
XFILL_1__10012_ gnd vdd FILL
XFILL_4__11172_ gnd vdd FILL
XFILL_3__14690_ gnd vdd FILL
XFILL_0__13530_ gnd vdd FILL
XFILL_0__10742_ gnd vdd FILL
X_15725_ _15724_/Y _15725_/B gnd _15725_/Y vdd NOR2X1
XFILL_5__15250_ gnd vdd FILL
XFILL_4__10123_ gnd vdd FILL
XFILL_5__12462_ gnd vdd FILL
X_12937_ _12170_/B _8176_/CLK _8176_/R vdd _12937_/D gnd vdd DFFSR
XFILL_2__11302_ gnd vdd FILL
XFILL_3__13641_ gnd vdd FILL
XSFILL74120x48050 gnd vdd FILL
XFILL_4__15980_ gnd vdd FILL
XFILL_1__14820_ gnd vdd FILL
XFILL_2__15070_ gnd vdd FILL
XFILL_2__12282_ gnd vdd FILL
XFILL_5__14201_ gnd vdd FILL
XFILL_0__13461_ gnd vdd FILL
XFILL_0__10673_ gnd vdd FILL
XFILL_5__7954_ gnd vdd FILL
XFILL_5__11413_ gnd vdd FILL
XFILL_5__15181_ gnd vdd FILL
X_15656_ _15656_/A _15656_/B _15656_/C gnd _15656_/Y vdd NOR3X1
XFILL_0__15200_ gnd vdd FILL
XFILL_5__12393_ gnd vdd FILL
X_12868_ _12934_/Q gnd _12868_/Y vdd INVX1
XFILL_2__14021_ gnd vdd FILL
XFILL_4__10054_ gnd vdd FILL
XFILL_4__14931_ gnd vdd FILL
XFILL_3__16360_ gnd vdd FILL
XFILL_1_BUFX2_insert840 gnd vdd FILL
XFILL_2__11233_ gnd vdd FILL
XFILL_0__12412_ gnd vdd FILL
XFILL_1_BUFX2_insert851 gnd vdd FILL
XFILL_3__13572_ gnd vdd FILL
XFILL_1_BUFX2_insert862 gnd vdd FILL
XFILL_0__16180_ gnd vdd FILL
XFILL_3__10784_ gnd vdd FILL
XFILL_1__11963_ gnd vdd FILL
XFILL_1__14751_ gnd vdd FILL
XFILL_5__6905_ gnd vdd FILL
X_14607_ _14607_/A _14607_/B _14604_/Y gnd _14618_/A vdd NAND3X1
XFILL_0__13392_ gnd vdd FILL
XFILL_5__14132_ gnd vdd FILL
XFILL_5__7885_ gnd vdd FILL
XFILL_3__15311_ gnd vdd FILL
XFILL_1_BUFX2_insert873 gnd vdd FILL
XFILL_5__11344_ gnd vdd FILL
X_11819_ _11818_/Y _11819_/B gnd _11820_/C vdd AND2X2
XFILL_2__9915_ gnd vdd FILL
XFILL_4__14862_ gnd vdd FILL
XFILL_3__12523_ gnd vdd FILL
XFILL_1_BUFX2_insert884 gnd vdd FILL
X_15587_ _16141_/A _14101_/A _16141_/C gnd _15609_/B vdd NOR3X1
X_12799_ _12719_/A _12685_/CLK _12799_/R vdd _12799_/D gnd vdd DFFSR
XFILL_1__10914_ gnd vdd FILL
XFILL_1_BUFX2_insert895 gnd vdd FILL
XFILL_3__16291_ gnd vdd FILL
XFILL_2__11164_ gnd vdd FILL
XFILL_1__13702_ gnd vdd FILL
XFILL_0__15131_ gnd vdd FILL
XFILL_0__12343_ gnd vdd FILL
XFILL_5__9624_ gnd vdd FILL
XFILL_5__6836_ gnd vdd FILL
XFILL_1__11894_ gnd vdd FILL
XFILL_1__14682_ gnd vdd FILL
XFILL_6__12634_ gnd vdd FILL
XFILL_4__13813_ gnd vdd FILL
X_14538_ _7404_/Q _13818_/A _14847_/C _7148_/Q gnd _14547_/A vdd AOI22X1
XFILL_5__14063_ gnd vdd FILL
XFILL_2__10115_ gnd vdd FILL
XFILL_3__15242_ gnd vdd FILL
XFILL_5__11275_ gnd vdd FILL
XFILL112280x74050 gnd vdd FILL
XFILL_4__14793_ gnd vdd FILL
XFILL_2__9846_ gnd vdd FILL
XFILL_3__12454_ gnd vdd FILL
XFILL_2__15972_ gnd vdd FILL
XFILL_1__13633_ gnd vdd FILL
XFILL_0__15062_ gnd vdd FILL
XFILL_2__11095_ gnd vdd FILL
XSFILL54040x15050 gnd vdd FILL
XFILL_5__13014_ gnd vdd FILL
XFILL_5__9555_ gnd vdd FILL
XFILL_0__12274_ gnd vdd FILL
XSFILL79640x79050 gnd vdd FILL
XSFILL28200x25050 gnd vdd FILL
X_14469_ _14468_/Y _14865_/C gnd _14469_/Y vdd NOR2X1
XSFILL53800x70050 gnd vdd FILL
XFILL_4__13744_ gnd vdd FILL
XFILL_0__8861_ gnd vdd FILL
XFILL_3__11405_ gnd vdd FILL
XSFILL94440x20050 gnd vdd FILL
XFILL_4__10956_ gnd vdd FILL
XFILL_2__10046_ gnd vdd FILL
XFILL_3__15173_ gnd vdd FILL
XFILL_0__14013_ gnd vdd FILL
XFILL_2__14923_ gnd vdd FILL
XFILL_5__8506_ gnd vdd FILL
XFILL_3__12385_ gnd vdd FILL
XFILL_2__9777_ gnd vdd FILL
XFILL_1__16352_ gnd vdd FILL
XFILL_3__8570_ gnd vdd FILL
XFILL_1__13564_ gnd vdd FILL
XFILL_0__11225_ gnd vdd FILL
XFILL_2__6989_ gnd vdd FILL
X_16208_ _16207_/Y _16208_/B _15204_/A _14840_/Y gnd _16208_/Y vdd OAI22X1
XFILL_1__10776_ gnd vdd FILL
XFILL_5__9486_ gnd vdd FILL
XFILL_0__7812_ gnd vdd FILL
XFILL_3__14124_ gnd vdd FILL
XFILL_5__10157_ gnd vdd FILL
XFILL_4__13675_ gnd vdd FILL
XFILL_2__8728_ gnd vdd FILL
XSFILL43880x58050 gnd vdd FILL
XFILL_1__15303_ gnd vdd FILL
XFILL_1__12515_ gnd vdd FILL
XFILL_3__11336_ gnd vdd FILL
XFILL_2__14854_ gnd vdd FILL
XFILL_4__10887_ gnd vdd FILL
XFILL_0__11156_ gnd vdd FILL
XFILL_1__13495_ gnd vdd FILL
XFILL_1__16283_ gnd vdd FILL
XFILL_4__15414_ gnd vdd FILL
X_16139_ _16132_/Y _16139_/B _16139_/C gnd _16139_/Y vdd NAND3X1
XFILL_0__7743_ gnd vdd FILL
XFILL_4__12626_ gnd vdd FILL
X_9070_ _9022_/A _8165_/CLK _8165_/R vdd _9024_/Y gnd vdd DFFSR
XFILL_2__13805_ gnd vdd FILL
XFILL_3__14055_ gnd vdd FILL
XFILL_5__14965_ gnd vdd FILL
XFILL_4__16394_ gnd vdd FILL
XFILL_1__15234_ gnd vdd FILL
XFILL_1__12446_ gnd vdd FILL
XFILL_3__7452_ gnd vdd FILL
XSFILL18680x34050 gnd vdd FILL
XFILL_0__10107_ gnd vdd FILL
XFILL_3__11267_ gnd vdd FILL
XFILL_2__8659_ gnd vdd FILL
XSFILL8520x44050 gnd vdd FILL
XFILL_2__14785_ gnd vdd FILL
XFILL_2__11997_ gnd vdd FILL
XFILL_0__15964_ gnd vdd FILL
X_8021_ _8021_/A _7997_/B _8021_/C gnd _8053_/D vdd OAI21X1
XFILL_5__8368_ gnd vdd FILL
XSFILL74200x28050 gnd vdd FILL
XFILL_0__11087_ gnd vdd FILL
XFILL_4__15345_ gnd vdd FILL
XFILL_3__13006_ gnd vdd FILL
XFILL_5__13916_ gnd vdd FILL
XSFILL59560x46050 gnd vdd FILL
XFILL_0__7674_ gnd vdd FILL
XFILL_1__15165_ gnd vdd FILL
XFILL_2__13736_ gnd vdd FILL
XFILL_5__14896_ gnd vdd FILL
XFILL_3__11198_ gnd vdd FILL
XFILL_2__10948_ gnd vdd FILL
XFILL_0__10038_ gnd vdd FILL
XFILL_1__12377_ gnd vdd FILL
XFILL_5__7319_ gnd vdd FILL
XFILL_0__14915_ gnd vdd FILL
XFILL_0__9413_ gnd vdd FILL
XFILL_0__15895_ gnd vdd FILL
XFILL_4__11508_ gnd vdd FILL
XFILL_5__13847_ gnd vdd FILL
XFILL_3__9122_ gnd vdd FILL
XFILL_4__15276_ gnd vdd FILL
XFILL_3__10149_ gnd vdd FILL
XFILL_4__12488_ gnd vdd FILL
XFILL_1__11328_ gnd vdd FILL
XFILL_1__14116_ gnd vdd FILL
XFILL_2__13667_ gnd vdd FILL
XFILL_1__15096_ gnd vdd FILL
XFILL_0__14846_ gnd vdd FILL
XFILL_2__10879_ gnd vdd FILL
XFILL_0__9344_ gnd vdd FILL
XFILL_4__14227_ gnd vdd FILL
XSFILL109560x15050 gnd vdd FILL
XFILL_2__15406_ gnd vdd FILL
XFILL_4__11439_ gnd vdd FILL
XFILL_2__12618_ gnd vdd FILL
XFILL_5__13778_ gnd vdd FILL
XFILL_1__14047_ gnd vdd FILL
XFILL_3__14957_ gnd vdd FILL
X_9972_ _9936_/A _9194_/CLK _7914_/R vdd _9972_/D gnd vdd DFFSR
XFILL_2__16386_ gnd vdd FILL
XFILL_1__11259_ gnd vdd FILL
XFILL_2__13598_ gnd vdd FILL
XSFILL38840x47050 gnd vdd FILL
XFILL_0__14777_ gnd vdd FILL
XFILL_0__11989_ gnd vdd FILL
XFILL112360x54050 gnd vdd FILL
XFILL_5__15517_ gnd vdd FILL
XFILL_5__12729_ gnd vdd FILL
XFILL_0__9275_ gnd vdd FILL
XFILL_4__14158_ gnd vdd FILL
XFILL_3__8004_ gnd vdd FILL
X_8923_ _8837_/A _8792_/CLK _7896_/R vdd _8923_/D gnd vdd DFFSR
XFILL_3__13908_ gnd vdd FILL
XFILL_2__15337_ gnd vdd FILL
XFILL_3__14888_ gnd vdd FILL
XFILL_6__9802_ gnd vdd FILL
XFILL_0__13728_ gnd vdd FILL
XFILL_0__8226_ gnd vdd FILL
XFILL_4__13109_ gnd vdd FILL
XFILL_6__7994_ gnd vdd FILL
XFILL_5__15448_ gnd vdd FILL
XFILL_3__13839_ gnd vdd FILL
XFILL_6__14999_ gnd vdd FILL
X_8854_ _8854_/A _8854_/B _8853_/Y gnd _8854_/Y vdd OAI21X1
XFILL_4__14089_ gnd vdd FILL
XFILL_2__15268_ gnd vdd FILL
XFILL_0__13659_ gnd vdd FILL
XFILL_1__15998_ gnd vdd FILL
XSFILL79320x61050 gnd vdd FILL
XFILL_6__6945_ gnd vdd FILL
XSFILL43960x38050 gnd vdd FILL
X_7805_ _7814_/A _8701_/B gnd _7806_/C vdd NAND2X1
XFILL_5__15379_ gnd vdd FILL
XFILL_2__14219_ gnd vdd FILL
X_8785_ _8753_/B _7889_/B gnd _8786_/C vdd NAND2X1
XFILL_2__15199_ gnd vdd FILL
XFILL_1__14949_ gnd vdd FILL
XFILL_0__16378_ gnd vdd FILL
XFILL_0__7108_ gnd vdd FILL
XFILL_0__8088_ gnd vdd FILL
XFILL_3__15509_ gnd vdd FILL
X_7736_ _7736_/A gnd _7736_/Y vdd INVX1
XSFILL18760x14050 gnd vdd FILL
XSFILL114520x70050 gnd vdd FILL
XFILL_1__8970_ gnd vdd FILL
XFILL_3__8906_ gnd vdd FILL
XSFILL8600x24050 gnd vdd FILL
XFILL_0__15329_ gnd vdd FILL
XFILL_3__9886_ gnd vdd FILL
XFILL_0__7039_ gnd vdd FILL
XSFILL84440x52050 gnd vdd FILL
X_7667_ _7629_/A _7661_/CLK _7789_/R vdd _7667_/D gnd vdd DFFSR
XFILL_4__7630_ gnd vdd FILL
XFILL_3__8837_ gnd vdd FILL
XSFILL84280x6050 gnd vdd FILL
X_9406_ _9454_/Q gnd _9406_/Y vdd INVX1
XFILL_1__7852_ gnd vdd FILL
X_7598_ _7596_/Y _7598_/B _7598_/C gnd _7598_/Y vdd OAI21X1
XFILL_3__8768_ gnd vdd FILL
XFILL_4__7561_ gnd vdd FILL
XSFILL73480x76050 gnd vdd FILL
XFILL_4__9300_ gnd vdd FILL
X_9337_ _9431_/Q gnd _9339_/A vdd INVX1
XFILL_3__7719_ gnd vdd FILL
XFILL112440x34050 gnd vdd FILL
XFILL_4__7492_ gnd vdd FILL
XFILL_4_BUFX2_insert235 gnd vdd FILL
XFILL_3__8699_ gnd vdd FILL
XFILL_4_BUFX2_insert246 gnd vdd FILL
XFILL_1__9522_ gnd vdd FILL
XSFILL79800x39050 gnd vdd FILL
X_9268_ _9268_/A _9240_/A _9267_/Y gnd _9268_/Y vdd OAI21X1
XFILL_4__9231_ gnd vdd FILL
XFILL_4_BUFX2_insert257 gnd vdd FILL
XFILL_4_BUFX2_insert268 gnd vdd FILL
X_10150_ _10214_/Q gnd _10150_/Y vdd INVX1
XFILL_4_BUFX2_insert279 gnd vdd FILL
X_8219_ _8232_/B _9371_/B gnd _8220_/C vdd NAND2X1
XFILL_3_BUFX2_insert902 gnd vdd FILL
X_9199_ _9199_/Q _7274_/CLK _7274_/R vdd _9155_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert913 gnd vdd FILL
XFILL_4__9162_ gnd vdd FILL
XFILL_3_BUFX2_insert924 gnd vdd FILL
XFILL_3_BUFX2_insert935 gnd vdd FILL
X_10081_ _14016_/A _9953_/CLK _7276_/R vdd _10009_/Y gnd vdd DFFSR
XFILL_1__8404_ gnd vdd FILL
XFILL_3_BUFX2_insert946 gnd vdd FILL
XFILL_1__9384_ gnd vdd FILL
XFILL_4__8113_ gnd vdd FILL
XFILL_3_BUFX2_insert957 gnd vdd FILL
XFILL_3_BUFX2_insert968 gnd vdd FILL
XSFILL28840x79050 gnd vdd FILL
XFILL_3_BUFX2_insert979 gnd vdd FILL
XFILL_4__9093_ gnd vdd FILL
XSFILL94280x55050 gnd vdd FILL
XSFILL114600x50050 gnd vdd FILL
XFILL_1__8335_ gnd vdd FILL
XSFILL84520x32050 gnd vdd FILL
X_13840_ _13840_/A _13840_/B _13274_/A gnd _12973_/B vdd AOI21X1
XSFILL69080x31050 gnd vdd FILL
XFILL_1__8266_ gnd vdd FILL
XSFILL44040x9050 gnd vdd FILL
XSFILL103640x74050 gnd vdd FILL
XFILL_3_BUFX2_insert1007 gnd vdd FILL
XFILL_3_BUFX2_insert1018 gnd vdd FILL
X_13771_ _14180_/C _15298_/D _8540_/Q _13771_/D gnd _13772_/B vdd AOI22X1
XFILL_1__7217_ gnd vdd FILL
X_10983_ _10983_/A vdd _10982_/Y gnd _10983_/Y vdd OAI21X1
XFILL_3_BUFX2_insert1029 gnd vdd FILL
XFILL_1_BUFX2_insert103 gnd vdd FILL
XFILL_1__8197_ gnd vdd FILL
X_15510_ _15508_/Y _15509_/Y _15510_/C gnd _15510_/Y vdd NAND3X1
XFILL_4__9995_ gnd vdd FILL
X_12722_ _12800_/Q gnd _12722_/Y vdd INVX1
XSFILL34040x79050 gnd vdd FILL
X_15441_ _13909_/A _15680_/B _15680_/C gnd _15441_/Y vdd NAND3X1
X_12653_ _12651_/Y vdd _12652_/Y gnd _12691_/D vdd OAI21X1
XFILL_1__7079_ gnd vdd FILL
XFILL_2__7961_ gnd vdd FILL
XFILL_0_BUFX2_insert803 gnd vdd FILL
XFILL_0_BUFX2_insert814 gnd vdd FILL
XFILL_5__7670_ gnd vdd FILL
XFILL_4__8877_ gnd vdd FILL
X_11604_ _11582_/C _11604_/B _11604_/C gnd _11612_/A vdd AOI21X1
XFILL_0_BUFX2_insert825 gnd vdd FILL
X_15372_ _15372_/A _15371_/Y gnd _15373_/A vdd NOR2X1
XFILL_2__6912_ gnd vdd FILL
X_12584_ _12582_/Y vdd _12584_/C gnd _12584_/Y vdd OAI21X1
XFILL_0_BUFX2_insert836 gnd vdd FILL
XFILL_1_BUFX2_insert1000 gnd vdd FILL
XSFILL3720x47050 gnd vdd FILL
XFILL_1_BUFX2_insert1011 gnd vdd FILL
XFILL_0_BUFX2_insert847 gnd vdd FILL
XFILL_4__7828_ gnd vdd FILL
XFILL_0_BUFX2_insert858 gnd vdd FILL
XFILL_2__7892_ gnd vdd FILL
XFILL_1_BUFX2_insert1022 gnd vdd FILL
XFILL_0_BUFX2_insert869 gnd vdd FILL
X_14323_ _8236_/A _14323_/B _14065_/C _15806_/A gnd _14323_/Y vdd AOI22X1
XFILL_1_BUFX2_insert1033 gnd vdd FILL
XFILL_4__10810_ gnd vdd FILL
XFILL_5__11060_ gnd vdd FILL
X_11535_ _11099_/Y _11527_/C _11534_/Y gnd _11535_/Y vdd NAND3X1
XFILL_1_BUFX2_insert1044 gnd vdd FILL
XFILL_2__9631_ gnd vdd FILL
XSFILL28920x59050 gnd vdd FILL
XFILL_1_BUFX2_insert1055 gnd vdd FILL
XFILL_2__6843_ gnd vdd FILL
XFILL_1__10630_ gnd vdd FILL
XFILL_4__11790_ gnd vdd FILL
XSFILL94360x35050 gnd vdd FILL
XFILL_1_BUFX2_insert1066 gnd vdd FILL
XFILL_5__9340_ gnd vdd FILL
XFILL_4__7759_ gnd vdd FILL
XFILL_3_BUFX2_insert18 gnd vdd FILL
XFILL_5__10011_ gnd vdd FILL
XFILL_3_BUFX2_insert29 gnd vdd FILL
X_14254_ _10214_/Q gnd _14256_/C vdd INVX1
XFILL_1_BUFX2_insert1088 gnd vdd FILL
X_11466_ _11415_/C _11466_/B _11465_/Y gnd _11466_/Y vdd NAND3X1
XFILL_2__11920_ gnd vdd FILL
XFILL_3__12170_ gnd vdd FILL
XFILL_0__11010_ gnd vdd FILL
XFILL_1__10561_ gnd vdd FILL
XFILL_5__9271_ gnd vdd FILL
X_13205_ _12108_/B _13180_/CLK _13180_/R vdd _13205_/D gnd vdd DFFSR
XSFILL69160x11050 gnd vdd FILL
X_10417_ _10415_/Y _10426_/B _10417_/C gnd _10473_/D vdd OAI21X1
X_14185_ _7653_/Q _14185_/B _14184_/Y gnd _14194_/A vdd AOI21X1
XFILL_4__13460_ gnd vdd FILL
XFILL_1__12300_ gnd vdd FILL
XFILL_3__11121_ gnd vdd FILL
XFILL_2__8513_ gnd vdd FILL
X_11397_ _11278_/Y _11279_/Y _11089_/Y gnd _11687_/A vdd OAI21X1
XFILL_4__10672_ gnd vdd FILL
XFILL_1__13280_ gnd vdd FILL
XFILL_4__9429_ gnd vdd FILL
XFILL_2__9493_ gnd vdd FILL
XFILL_5__8222_ gnd vdd FILL
XFILL_2__11851_ gnd vdd FILL
XFILL_1__10492_ gnd vdd FILL
XFILL_4__12411_ gnd vdd FILL
X_13136_ _13194_/Q gnd _13136_/Y vdd INVX1
XFILL_5__11962_ gnd vdd FILL
XFILL_4_BUFX2_insert780 gnd vdd FILL
X_10348_ _10348_/Q _7020_/CLK _8053_/R vdd _10298_/Y gnd vdd DFFSR
XFILL_5__14750_ gnd vdd FILL
XFILL_3__11052_ gnd vdd FILL
XSFILL104360x20050 gnd vdd FILL
XFILL_4__13391_ gnd vdd FILL
XFILL_1__12231_ gnd vdd FILL
XFILL_2__8444_ gnd vdd FILL
XFILL_4_BUFX2_insert791 gnd vdd FILL
XFILL_2__10802_ gnd vdd FILL
XFILL_2__14570_ gnd vdd FILL
XFILL_6_CLKBUF1_insert157 gnd vdd FILL
XFILL_0__12961_ gnd vdd FILL
XFILL_2__11782_ gnd vdd FILL
XFILL_6_CLKBUF1_insert168 gnd vdd FILL
XFILL_4__15130_ gnd vdd FILL
XFILL_5__13701_ gnd vdd FILL
XFILL_5__10913_ gnd vdd FILL
X_10279_ _10280_/B _7079_/B gnd _10279_/Y vdd NAND2X1
XFILL_4__12342_ gnd vdd FILL
XFILL_3__10003_ gnd vdd FILL
X_13067_ _6890_/A _8169_/CLK _8937_/R vdd _13013_/Y gnd vdd DFFSR
XFILL_5__11893_ gnd vdd FILL
XFILL_5__14681_ gnd vdd FILL
XFILL_2__13521_ gnd vdd FILL
XFILL_3__15860_ gnd vdd FILL
XSFILL8840x80050 gnd vdd FILL
XFILL_2__8375_ gnd vdd FILL
XFILL_5__7104_ gnd vdd FILL
XFILL_0__11912_ gnd vdd FILL
XFILL_1__12162_ gnd vdd FILL
XFILL_0__14700_ gnd vdd FILL
XFILL_0__15680_ gnd vdd FILL
XFILL_6__10114_ gnd vdd FILL
XFILL_0__12892_ gnd vdd FILL
X_12018_ _12018_/A _12018_/B _12017_/Y gnd _13101_/B vdd NAND3X1
XFILL_5__8084_ gnd vdd FILL
XFILL_5__13632_ gnd vdd FILL
XFILL_6__15971_ gnd vdd FILL
XSFILL59080x63050 gnd vdd FILL
XFILL_3__14811_ gnd vdd FILL
XFILL_4__15061_ gnd vdd FILL
XFILL_2__16240_ gnd vdd FILL
XFILL_4__12273_ gnd vdd FILL
XFILL_2__7326_ gnd vdd FILL
XFILL_1__11113_ gnd vdd FILL
XFILL_0__14631_ gnd vdd FILL
XFILL_2__10664_ gnd vdd FILL
XFILL_2__13452_ gnd vdd FILL
XFILL_3__15791_ gnd vdd FILL
XFILL_1__12093_ gnd vdd FILL
XFILL_5__7035_ gnd vdd FILL
XFILL_0__11843_ gnd vdd FILL
XFILL_4__14012_ gnd vdd FILL
XFILL_6__14922_ gnd vdd FILL
XSFILL3800x27050 gnd vdd FILL
XFILL_5__16351_ gnd vdd FILL
XFILL_5__13563_ gnd vdd FILL
XFILL_4__11224_ gnd vdd FILL
XFILL_2__12403_ gnd vdd FILL
XFILL_5__10775_ gnd vdd FILL
XFILL_3__14742_ gnd vdd FILL
XFILL_1__15921_ gnd vdd FILL
XFILL_2__16171_ gnd vdd FILL
XFILL_3__11954_ gnd vdd FILL
XFILL_1__11044_ gnd vdd FILL
XFILL112280x69050 gnd vdd FILL
XFILL_0__14562_ gnd vdd FILL
XFILL_2__13383_ gnd vdd FILL
XFILL_5__15302_ gnd vdd FILL
XFILL_0__11774_ gnd vdd FILL
XFILL_5__12514_ gnd vdd FILL
XFILL_3__10905_ gnd vdd FILL
XFILL_5__13494_ gnd vdd FILL
XFILL_4__11155_ gnd vdd FILL
X_13969_ _14946_/A _13969_/B _14506_/C _15464_/C gnd _13970_/A vdd OAI22X1
XSFILL94440x15050 gnd vdd FILL
XFILL_2__15122_ gnd vdd FILL
XFILL_5__16282_ gnd vdd FILL
XFILL_0__16301_ gnd vdd FILL
XFILL_2__12334_ gnd vdd FILL
XFILL_3__14673_ gnd vdd FILL
XFILL_0__13513_ gnd vdd FILL
XFILL_3__11885_ gnd vdd FILL
XFILL_1__15852_ gnd vdd FILL
XFILL_2__7188_ gnd vdd FILL
XFILL_0__14493_ gnd vdd FILL
X_15708_ _15708_/A _15708_/B _15708_/C gnd _15708_/Y vdd NOR3X1
XFILL_0__8011_ gnd vdd FILL
XSFILL13800x81050 gnd vdd FILL
XFILL_5__15233_ gnd vdd FILL
XFILL_5__12445_ gnd vdd FILL
XFILL_5__8986_ gnd vdd FILL
XFILL_4__10106_ gnd vdd FILL
XFILL_3__16412_ gnd vdd FILL
XFILL_3__13624_ gnd vdd FILL
XFILL_6__14784_ gnd vdd FILL
XSFILL79240x76050 gnd vdd FILL
XFILL_0__16232_ gnd vdd FILL
XFILL_1__14803_ gnd vdd FILL
XFILL_2__15053_ gnd vdd FILL
XFILL_4__15963_ gnd vdd FILL
XFILL_4__11086_ gnd vdd FILL
XFILL_3__10836_ gnd vdd FILL
XFILL_0__13444_ gnd vdd FILL
XFILL_2__12265_ gnd vdd FILL
XFILL_5__7937_ gnd vdd FILL
XFILL_0__10656_ gnd vdd FILL
XFILL_1__15783_ gnd vdd FILL
X_15639_ _15915_/C _15639_/B _15912_/D _14125_/A gnd _15640_/B vdd OAI22X1
XFILL_1__12995_ gnd vdd FILL
XFILL_6__13735_ gnd vdd FILL
XFILL_4__10037_ gnd vdd FILL
XFILL_3__16343_ gnd vdd FILL
XFILL_1_BUFX2_insert670 gnd vdd FILL
XFILL_5__12376_ gnd vdd FILL
XFILL_2__14004_ gnd vdd FILL
XFILL_5__15164_ gnd vdd FILL
X_8570_ _8619_/B _9978_/B gnd _8570_/Y vdd NAND2X1
XFILL_4__14914_ gnd vdd FILL
XFILL_3__9740_ gnd vdd FILL
XFILL_1_BUFX2_insert681 gnd vdd FILL
XFILL_3__13555_ gnd vdd FILL
XSFILL28840x9050 gnd vdd FILL
XFILL_2__11216_ gnd vdd FILL
XFILL_3__6952_ gnd vdd FILL
XFILL_3__10767_ gnd vdd FILL
XFILL_4__15894_ gnd vdd FILL
XFILL_1__14734_ gnd vdd FILL
XFILL_2__12196_ gnd vdd FILL
XSFILL18680x29050 gnd vdd FILL
XFILL_0__16163_ gnd vdd FILL
XFILL_1_BUFX2_insert692 gnd vdd FILL
XFILL_0__13375_ gnd vdd FILL
XFILL_1__11946_ gnd vdd FILL
XSFILL8520x39050 gnd vdd FILL
XFILL_5__7868_ gnd vdd FILL
X_7521_ _7447_/A _8560_/CLK _8676_/R vdd _7521_/D gnd vdd DFFSR
XFILL_5__14115_ gnd vdd FILL
XFILL_5__11327_ gnd vdd FILL
XFILL_3__12506_ gnd vdd FILL
XFILL_5__15095_ gnd vdd FILL
XFILL_4__14845_ gnd vdd FILL
XFILL_2__11147_ gnd vdd FILL
XFILL_0__15114_ gnd vdd FILL
XFILL_3__16274_ gnd vdd FILL
XSFILL84360x67050 gnd vdd FILL
XFILL_3__13486_ gnd vdd FILL
XFILL_3__9671_ gnd vdd FILL
XFILL_0__12326_ gnd vdd FILL
XFILL_3__10698_ gnd vdd FILL
XFILL_0__16094_ gnd vdd FILL
XFILL_5__9607_ gnd vdd FILL
XFILL_3__6883_ gnd vdd FILL
XFILL_1__14665_ gnd vdd FILL
XFILL_1__11877_ gnd vdd FILL
XFILL_5__14046_ gnd vdd FILL
XFILL_0__8913_ gnd vdd FILL
XFILL_6__16385_ gnd vdd FILL
XFILL_5__7799_ gnd vdd FILL
XFILL_3__15225_ gnd vdd FILL
X_7452_ _7450_/Y _7416_/B _7452_/C gnd _7452_/Y vdd OAI21X1
XFILL_5__11258_ gnd vdd FILL
XFILL_6__13597_ gnd vdd FILL
XFILL_3__12437_ gnd vdd FILL
XFILL_0__9893_ gnd vdd FILL
XFILL_3__8622_ gnd vdd FILL
XFILL_1__16404_ gnd vdd FILL
XSFILL94760x7050 gnd vdd FILL
XFILL_1__13616_ gnd vdd FILL
XFILL_0__15045_ gnd vdd FILL
XFILL_4__11988_ gnd vdd FILL
XFILL_2__15955_ gnd vdd FILL
XFILL_2__11078_ gnd vdd FILL
XFILL_4__14776_ gnd vdd FILL
XFILL_1__10828_ gnd vdd FILL
XFILL_0__12257_ gnd vdd FILL
XFILL_5__9538_ gnd vdd FILL
XFILL_1__14596_ gnd vdd FILL
XFILL_0__8844_ gnd vdd FILL
XFILL_4__10939_ gnd vdd FILL
XFILL_2__10029_ gnd vdd FILL
XFILL_3__15156_ gnd vdd FILL
XFILL_5__11189_ gnd vdd FILL
XFILL_4__13727_ gnd vdd FILL
XFILL_2__14906_ gnd vdd FILL
X_7383_ _7383_/Q _9447_/CLK _9447_/R vdd _7383_/D gnd vdd DFFSR
XFILL_3__12368_ gnd vdd FILL
XFILL_1__16335_ gnd vdd FILL
XFILL_0__11208_ gnd vdd FILL
XFILL_1__10759_ gnd vdd FILL
XFILL_1__13547_ gnd vdd FILL
XFILL_2__15886_ gnd vdd FILL
XFILL_0__12188_ gnd vdd FILL
X_9122_ _9120_/Y _9164_/B _9121_/Y gnd _9188_/D vdd OAI21X1
XFILL111880x42050 gnd vdd FILL
XFILL_6__8262_ gnd vdd FILL
XFILL_5__9469_ gnd vdd FILL
XFILL_3__14107_ gnd vdd FILL
XFILL_4__13658_ gnd vdd FILL
XFILL112360x49050 gnd vdd FILL
XFILL_6__12479_ gnd vdd FILL
XFILL_3__11319_ gnd vdd FILL
XFILL_3__7504_ gnd vdd FILL
XFILL_0__8775_ gnd vdd FILL
XFILL_2__14837_ gnd vdd FILL
XFILL_5__15997_ gnd vdd FILL
XFILL_3__15087_ gnd vdd FILL
XFILL_3__8484_ gnd vdd FILL
XFILL_6__7213_ gnd vdd FILL
XFILL_3__12299_ gnd vdd FILL
XFILL_0__11139_ gnd vdd FILL
XFILL_1__16266_ gnd vdd FILL
XFILL_1__13478_ gnd vdd FILL
X_9053_ _8971_/A _8171_/CLK _8171_/R vdd _8973_/Y gnd vdd DFFSR
XFILL_4__12609_ gnd vdd FILL
XFILL_0__7726_ gnd vdd FILL
XSFILL109400x74050 gnd vdd FILL
XFILL_3__14038_ gnd vdd FILL
XFILL_5__14948_ gnd vdd FILL
XFILL_3__7435_ gnd vdd FILL
XFILL_4__13589_ gnd vdd FILL
XFILL_1__15217_ gnd vdd FILL
XFILL_4__16377_ gnd vdd FILL
XFILL_1__12429_ gnd vdd FILL
XFILL_2__14768_ gnd vdd FILL
XSFILL8680x2050 gnd vdd FILL
XFILL_1__16197_ gnd vdd FILL
XFILL_0__15947_ gnd vdd FILL
X_8004_ _8048_/Q gnd _8006_/A vdd INVX1
XSFILL79320x56050 gnd vdd FILL
XSFILL54040x4050 gnd vdd FILL
XFILL_4__15328_ gnd vdd FILL
XSFILL89400x2050 gnd vdd FILL
XFILL_5__14879_ gnd vdd FILL
XFILL_2__13719_ gnd vdd FILL
XFILL_3__7366_ gnd vdd FILL
XFILL_1__15148_ gnd vdd FILL
XFILL_2__14699_ gnd vdd FILL
XFILL_0__15878_ gnd vdd FILL
XFILL_4__15259_ gnd vdd FILL
XFILL_3__9105_ gnd vdd FILL
XFILL_2_BUFX2_insert909 gnd vdd FILL
XFILL_0__7588_ gnd vdd FILL
XSFILL8600x19050 gnd vdd FILL
XFILL_3__7297_ gnd vdd FILL
XFILL_3__15989_ gnd vdd FILL
XFILL_0__14829_ gnd vdd FILL
XFILL_1__15079_ gnd vdd FILL
XFILL_1__8120_ gnd vdd FILL
XSFILL33800x12050 gnd vdd FILL
XFILL_3__9036_ gnd vdd FILL
X_9955_ _9955_/Q _9077_/CLK _7665_/R vdd _9955_/D gnd vdd DFFSR
XFILL_2__16369_ gnd vdd FILL
X_8906_ _8946_/Q gnd _8906_/Y vdd INVX1
XFILL_0__9258_ gnd vdd FILL
X_9886_ _9941_/B _9374_/B gnd _9886_/Y vdd NAND2X1
XFILL_0__8209_ gnd vdd FILL
X_8837_ _8837_/A gnd _8839_/A vdd INVX1
XFILL111960x22050 gnd vdd FILL
XFILL112440x29050 gnd vdd FILL
XFILL_4__9780_ gnd vdd FILL
XFILL_4__6992_ gnd vdd FILL
XBUFX2_insert908 _10913_/Y gnd _10944_/C vdd BUFX2
XFILL_6_BUFX2_insert853 gnd vdd FILL
X_8768_ _8766_/Y _8740_/A _8768_/C gnd _8768_/Y vdd OAI21X1
XSFILL23720x64050 gnd vdd FILL
XFILL_4__8731_ gnd vdd FILL
XBUFX2_insert919 _15069_/Y gnd _16314_/D vdd BUFX2
XFILL_3__9938_ gnd vdd FILL
XFILL112040x31050 gnd vdd FILL
X_7719_ _7744_/B _7847_/B gnd _7719_/Y vdd NAND2X1
XFILL_1__8953_ gnd vdd FILL
XFILL_3__9869_ gnd vdd FILL
X_8699_ _8699_/A _8698_/A _8699_/C gnd _8699_/Y vdd OAI21X1
XFILL_4__7613_ gnd vdd FILL
XFILL_1__8884_ gnd vdd FILL
X_11320_ _11461_/A gnd _11320_/Y vdd INVX2
XFILL_4__8593_ gnd vdd FILL
XSFILL114600x45050 gnd vdd FILL
XFILL_1__7835_ gnd vdd FILL
XFILL_4__7544_ gnd vdd FILL
X_11251_ _11247_/Y _11251_/B gnd _11251_/Y vdd NOR2X1
X_10202_ _10114_/A _9306_/CLK _9306_/R vdd _10202_/D gnd vdd DFFSR
XFILL_4__7475_ gnd vdd FILL
XFILL_1__9505_ gnd vdd FILL
XSFILL29080x42050 gnd vdd FILL
X_11182_ _12189_/Y _12314_/Y gnd _11182_/Y vdd NOR2X1
XFILL_4__9214_ gnd vdd FILL
XFILL_1__7697_ gnd vdd FILL
XFILL_3_BUFX2_insert710 gnd vdd FILL
X_10133_ _10193_/A _7445_/B gnd _10133_/Y vdd NAND2X1
XFILL_3_BUFX2_insert721 gnd vdd FILL
X_15990_ _9453_/Q _15202_/B _15995_/C gnd _15991_/C vdd NAND3X1
XFILL_3_BUFX2_insert732 gnd vdd FILL
XFILL_3_BUFX2_insert743 gnd vdd FILL
XFILL_4__9145_ gnd vdd FILL
XFILL_3_BUFX2_insert754 gnd vdd FILL
XFILL_3_BUFX2_insert765 gnd vdd FILL
X_14941_ _14941_/A _14830_/B gnd _14942_/C vdd NOR2X1
X_10064_ _10100_/Q gnd _10064_/Y vdd INVX1
XFILL_3_BUFX2_insert776 gnd vdd FILL
XFILL_1__9367_ gnd vdd FILL
XFILL_3_BUFX2_insert787 gnd vdd FILL
XFILL_3_BUFX2_insert798 gnd vdd FILL
XSFILL89240x39050 gnd vdd FILL
XFILL112120x11050 gnd vdd FILL
X_14872_ _13587_/A _14871_/Y _14872_/C _14870_/Y gnd _14876_/B vdd OAI22X1
XFILL_2__7111_ gnd vdd FILL
XFILL_1__8318_ gnd vdd FILL
XFILL_2__8091_ gnd vdd FILL
XFILL_1__9298_ gnd vdd FILL
X_13823_ _9565_/Q gnd _13823_/Y vdd INVX1
XFILL_5__10560_ gnd vdd FILL
XSFILL38840x4050 gnd vdd FILL
XFILL_1__8249_ gnd vdd FILL
XFILL_2__7042_ gnd vdd FILL
XFILL_2__10380_ gnd vdd FILL
XFILL_5__8840_ gnd vdd FILL
X_13754_ _8200_/A gnd _15331_/D vdd INVX1
XFILL_6__11850_ gnd vdd FILL
X_10966_ _10957_/Y _10948_/Y gnd _10970_/B vdd NOR2X1
XFILL_5__10491_ gnd vdd FILL
XFILL_0__10510_ gnd vdd FILL
XFILL_3__11670_ gnd vdd FILL
X_12705_ _12721_/B memoryOutData[3] gnd _12706_/C vdd NAND2X1
XFILL_5__12230_ gnd vdd FILL
XFILL_6__10801_ gnd vdd FILL
XFILL_5__8771_ gnd vdd FILL
XFILL_0__11490_ gnd vdd FILL
XFILL_4__9978_ gnd vdd FILL
XFILL_4__12960_ gnd vdd FILL
X_13685_ _13674_/Y _13684_/Y gnd _13685_/Y vdd NOR2X1
XFILL_2__12050_ gnd vdd FILL
XFILL_3__10621_ gnd vdd FILL
X_10897_ _10906_/A gnd _10897_/Y vdd INVX2
XFILL_1__11800_ gnd vdd FILL
XFILL_1__12780_ gnd vdd FILL
XFILL_2__8993_ gnd vdd FILL
XFILL_0__10441_ gnd vdd FILL
XFILL_5__7722_ gnd vdd FILL
XFILL_0_BUFX2_insert600 gnd vdd FILL
X_15424_ _16261_/A _13912_/Y _13911_/Y _16261_/D gnd _15425_/B vdd OAI22X1
X_12636_ _12413_/B gnd _12636_/Y vdd INVX1
XFILL_4__11911_ gnd vdd FILL
XFILL_5__12161_ gnd vdd FILL
XFILL_0_BUFX2_insert611 gnd vdd FILL
XFILL_2__11001_ gnd vdd FILL
XFILL_3__13340_ gnd vdd FILL
XFILL_0_BUFX2_insert622 gnd vdd FILL
XFILL_2__7944_ gnd vdd FILL
XFILL_0_BUFX2_insert633 gnd vdd FILL
XFILL_3__10552_ gnd vdd FILL
XFILL_4__12891_ gnd vdd FILL
XSFILL104360x15050 gnd vdd FILL
XFILL_0_BUFX2_insert644 gnd vdd FILL
XFILL_0__13160_ gnd vdd FILL
XFILL_1__11731_ gnd vdd FILL
XFILL_0__10372_ gnd vdd FILL
XFILL_5__11112_ gnd vdd FILL
X_15355_ _15355_/A _15355_/B gnd _15373_/B vdd NOR2X1
XFILL_0_BUFX2_insert655 gnd vdd FILL
X_12567_ _12663_/Q gnd _12567_/Y vdd INVX1
XFILL_4__14630_ gnd vdd FILL
XFILL_5__12092_ gnd vdd FILL
XFILL_0_BUFX2_insert666 gnd vdd FILL
XFILL_4__11842_ gnd vdd FILL
XFILL_3__13271_ gnd vdd FILL
XFILL_0_BUFX2_insert677 gnd vdd FILL
XFILL_0__12111_ gnd vdd FILL
XFILL_0_BUFX2_insert688 gnd vdd FILL
XFILL_1__11662_ gnd vdd FILL
XFILL_2__7875_ gnd vdd FILL
XFILL_1__14450_ gnd vdd FILL
XSFILL8840x75050 gnd vdd FILL
XFILL_0__13091_ gnd vdd FILL
X_14306_ _13865_/C _7721_/A _7081_/A _14344_/C gnd _14306_/Y vdd AOI22X1
XFILL_5__15920_ gnd vdd FILL
XFILL_5__7584_ gnd vdd FILL
XFILL_3__15010_ gnd vdd FILL
XFILL_5__11043_ gnd vdd FILL
X_11518_ _11118_/Y gnd _11518_/Y vdd INVX1
XFILL_0_BUFX2_insert699 gnd vdd FILL
XFILL_2__9614_ gnd vdd FILL
XFILL_4__14561_ gnd vdd FILL
XSFILL59080x58050 gnd vdd FILL
XFILL_6__13382_ gnd vdd FILL
X_15286_ _15802_/A _13708_/D _15286_/C _15802_/D gnd _15286_/Y vdd OAI22X1
XSFILL89320x19050 gnd vdd FILL
XFILL_3__12222_ gnd vdd FILL
XFILL_1__13401_ gnd vdd FILL
X_12498_ _12496_/Y vdd _12498_/C gnd _12554_/D vdd OAI21X1
XFILL_2__15740_ gnd vdd FILL
XFILL_4__11773_ gnd vdd FILL
XFILL_0__6890_ gnd vdd FILL
XFILL_2__12952_ gnd vdd FILL
XFILL_0__12042_ gnd vdd FILL
XFILL_1__14381_ gnd vdd FILL
XSFILL99480x63050 gnd vdd FILL
XFILL_1__11593_ gnd vdd FILL
X_14237_ _14237_/A _14237_/B _13876_/C _14237_/D gnd _14237_/Y vdd OAI22X1
XFILL_4__16300_ gnd vdd FILL
XFILL_4__13512_ gnd vdd FILL
XSFILL74120x61050 gnd vdd FILL
XFILL_5__15851_ gnd vdd FILL
X_11449_ _11447_/Y _11256_/Y _11448_/Y gnd _11449_/Y vdd OAI21X1
XFILL_4__14492_ gnd vdd FILL
XFILL_1__16120_ gnd vdd FILL
XFILL_2__11903_ gnd vdd FILL
XFILL_3__12153_ gnd vdd FILL
XFILL_2__9545_ gnd vdd FILL
XFILL_1__13332_ gnd vdd FILL
XFILL_2__15671_ gnd vdd FILL
XFILL_1__10544_ gnd vdd FILL
XFILL_5__9254_ gnd vdd FILL
XFILL_2__12883_ gnd vdd FILL
XFILL_5__14802_ gnd vdd FILL
XFILL_4__16231_ gnd vdd FILL
XFILL_4__13443_ gnd vdd FILL
X_14168_ _14168_/A _14164_/Y gnd _14168_/Y vdd NOR2X1
XFILL_6__12264_ gnd vdd FILL
XFILL_3__11104_ gnd vdd FILL
XFILL_2__14622_ gnd vdd FILL
XFILL_5__15782_ gnd vdd FILL
XFILL_4__10655_ gnd vdd FILL
XFILL_2__9476_ gnd vdd FILL
XFILL_1__13263_ gnd vdd FILL
XFILL_5__8205_ gnd vdd FILL
XFILL_3__12084_ gnd vdd FILL
XFILL_5__12994_ gnd vdd FILL
XFILL_0__15801_ gnd vdd FILL
XFILL_1__16051_ gnd vdd FILL
XFILL_2__11834_ gnd vdd FILL
XFILL_0__13993_ gnd vdd FILL
X_13119_ _13155_/A _13119_/B gnd _13120_/C vdd NAND2X1
XSFILL13800x76050 gnd vdd FILL
XFILL_5__14733_ gnd vdd FILL
XFILL_4__16162_ gnd vdd FILL
XFILL_3__15912_ gnd vdd FILL
XFILL_1__15002_ gnd vdd FILL
XFILL_4__13374_ gnd vdd FILL
XFILL_5__11945_ gnd vdd FILL
XFILL_1__12214_ gnd vdd FILL
XFILL_0__8491_ gnd vdd FILL
X_14099_ _14099_/A gnd _14101_/A vdd INVX1
XFILL_3__7220_ gnd vdd FILL
XFILL_3__11035_ gnd vdd FILL
XFILL_2__14553_ gnd vdd FILL
XSFILL64520x5050 gnd vdd FILL
XFILL_0__15732_ gnd vdd FILL
XFILL_5__8136_ gnd vdd FILL
XSFILL94840x31050 gnd vdd FILL
XFILL_2__11765_ gnd vdd FILL
XSFILL13800x1050 gnd vdd FILL
XFILL_4__15113_ gnd vdd FILL
XSFILL38760x80050 gnd vdd FILL
XFILL_0__7442_ gnd vdd FILL
XFILL_4__12325_ gnd vdd FILL
XFILL_4__16093_ gnd vdd FILL
XFILL_5__14664_ gnd vdd FILL
XFILL_2__13504_ gnd vdd FILL
XFILL_2__8358_ gnd vdd FILL
XFILL_5__11876_ gnd vdd FILL
XFILL_3__15843_ gnd vdd FILL
XFILL_1__12145_ gnd vdd FILL
XFILL_2__14484_ gnd vdd FILL
XFILL_0__15663_ gnd vdd FILL
XFILL_5__8067_ gnd vdd FILL
XFILL_0__12875_ gnd vdd FILL
XFILL_2__11696_ gnd vdd FILL
XFILL_5__16403_ gnd vdd FILL
XFILL_5__13615_ gnd vdd FILL
XFILL_4__15044_ gnd vdd FILL
XFILL_2__16223_ gnd vdd FILL
XFILL_2__7309_ gnd vdd FILL
XFILL_0__7373_ gnd vdd FILL
XFILL_5__10827_ gnd vdd FILL
XFILL_4__12256_ gnd vdd FILL
XFILL_5__14595_ gnd vdd FILL
XFILL_2__13435_ gnd vdd FILL
XFILL_3__15774_ gnd vdd FILL
XFILL_0__14614_ gnd vdd FILL
XFILL_1__12076_ gnd vdd FILL
XFILL_2__10647_ gnd vdd FILL
XFILL_3__12986_ gnd vdd FILL
XFILL_3__7082_ gnd vdd FILL
XFILL_0__11826_ gnd vdd FILL
XFILL_0__9112_ gnd vdd FILL
XFILL_5__16334_ gnd vdd FILL
XFILL_0__15594_ gnd vdd FILL
XFILL_4__11207_ gnd vdd FILL
X_6952_ _6950_/Y _6951_/A _6952_/C gnd _7014_/D vdd OAI21X1
XSFILL43880x71050 gnd vdd FILL
X_9740_ _9741_/B _7564_/B gnd _9740_/Y vdd NAND2X1
XFILL_3__14725_ gnd vdd FILL
XFILL_5__13546_ gnd vdd FILL
XFILL_5__10758_ gnd vdd FILL
XFILL_1__15904_ gnd vdd FILL
XFILL_4__12187_ gnd vdd FILL
XFILL_3__11937_ gnd vdd FILL
XSFILL74600x39050 gnd vdd FILL
XFILL_1__11027_ gnd vdd FILL
XFILL_2__16154_ gnd vdd FILL
XSFILL98920x77050 gnd vdd FILL
XFILL_2__13366_ gnd vdd FILL
XFILL_0__14545_ gnd vdd FILL
XFILL_2__10578_ gnd vdd FILL
XFILL_0__11757_ gnd vdd FILL
XFILL_0__9043_ gnd vdd FILL
XFILL_4__11138_ gnd vdd FILL
XFILL_2__15105_ gnd vdd FILL
XFILL_5__16265_ gnd vdd FILL
X_9671_ _9671_/A gnd _9673_/A vdd INVX1
X_6883_ _6883_/A gnd memoryWriteData[13] vdd BUFX2
XFILL_3__14656_ gnd vdd FILL
XFILL_5__10689_ gnd vdd FILL
XFILL_5__13477_ gnd vdd FILL
XFILL_2__12317_ gnd vdd FILL
XFILL_1__15835_ gnd vdd FILL
XFILL_3__11868_ gnd vdd FILL
XFILL_0__10708_ gnd vdd FILL
XFILL_2__16085_ gnd vdd FILL
XFILL_2__13297_ gnd vdd FILL
XFILL_0__14476_ gnd vdd FILL
XFILL_5__15216_ gnd vdd FILL
XFILL_0__11688_ gnd vdd FILL
XFILL_3__13607_ gnd vdd FILL
XFILL_5__12428_ gnd vdd FILL
XFILL_5__8969_ gnd vdd FILL
X_8622_ _8620_/Y _8567_/B _8622_/C gnd _8680_/D vdd OAI21X1
XFILL_5__16196_ gnd vdd FILL
XFILL_2__15036_ gnd vdd FILL
XFILL_4__15946_ gnd vdd FILL
XFILL_3__10819_ gnd vdd FILL
XFILL_4__11069_ gnd vdd FILL
XFILL_0__16215_ gnd vdd FILL
XFILL_3__14587_ gnd vdd FILL
XFILL_0__13427_ gnd vdd FILL
XFILL_2__12248_ gnd vdd FILL
XFILL_0__10639_ gnd vdd FILL
XFILL_3__7984_ gnd vdd FILL
XFILL_1__15766_ gnd vdd FILL
XFILL_3__11799_ gnd vdd FILL
XFILL_1__12978_ gnd vdd FILL
XSFILL108920x62050 gnd vdd FILL
XFILL_5__12359_ gnd vdd FILL
XFILL_3__16326_ gnd vdd FILL
XFILL_5__15147_ gnd vdd FILL
XFILL_5_BUFX2_insert805 gnd vdd FILL
X_8553_ _8495_/A _7786_/CLK _7153_/R vdd _8553_/D gnd vdd DFFSR
XFILL_3__13538_ gnd vdd FILL
XFILL_3__9723_ gnd vdd FILL
XSFILL109400x69050 gnd vdd FILL
XFILL_3__6935_ gnd vdd FILL
XFILL_1__14717_ gnd vdd FILL
XFILL_4__15877_ gnd vdd FILL
XFILL_5_BUFX2_insert816 gnd vdd FILL
XFILL_0__13358_ gnd vdd FILL
XFILL_2__12179_ gnd vdd FILL
XFILL_1__11929_ gnd vdd FILL
XFILL_0__16146_ gnd vdd FILL
XFILL_5_BUFX2_insert827 gnd vdd FILL
XFILL_1__15697_ gnd vdd FILL
XFILL_5_BUFX2_insert838 gnd vdd FILL
XBUFX2_insert1002 _12399_/Y gnd _9005_/B vdd BUFX2
X_7504_ _7504_/A gnd _7504_/Y vdd INVX1
X_8484_ _8484_/A _7972_/B gnd _8485_/C vdd NAND2X1
XFILL_4__14828_ gnd vdd FILL
XBUFX2_insert1013 _13569_/Y gnd _13751_/C vdd BUFX2
XFILL_5__15078_ gnd vdd FILL
XFILL_3__16257_ gnd vdd FILL
XFILL_5_BUFX2_insert849 gnd vdd FILL
XFILL_3__9654_ gnd vdd FILL
XFILL_3__13469_ gnd vdd FILL
XBUFX2_insert1024 _13340_/Y gnd _9675_/A vdd BUFX2
XFILL_0__12309_ gnd vdd FILL
XBUFX2_insert1035 _12390_/Y gnd _8228_/B vdd BUFX2
XSFILL38840x60050 gnd vdd FILL
XFILL_3__6866_ gnd vdd FILL
XFILL_0__16077_ gnd vdd FILL
XFILL_1__14648_ gnd vdd FILL
XFILL_0__13289_ gnd vdd FILL
X_7435_ _7435_/A gnd _7435_/Y vdd INVX1
XFILL_3__15208_ gnd vdd FILL
XFILL_5__14029_ gnd vdd FILL
XBUFX2_insert1046 _13297_/Y gnd _7723_/B vdd BUFX2
XBUFX2_insert1057 _15051_/Y gnd _16037_/C vdd BUFX2
XFILL_0__9876_ gnd vdd FILL
XFILL_3__8605_ gnd vdd FILL
XFILL_3__16188_ gnd vdd FILL
XBUFX2_insert1068 _13327_/Y gnd _8893_/B vdd BUFX2
XFILL_0__15028_ gnd vdd FILL
XFILL_2__15938_ gnd vdd FILL
XFILL_4__14759_ gnd vdd FILL
XFILL_1__14579_ gnd vdd FILL
XFILL_1__7620_ gnd vdd FILL
XFILL_0__8827_ gnd vdd FILL
X_7366_ _7366_/A _7366_/B _7365_/Y gnd _7366_/Y vdd OAI21X1
XFILL_3__15139_ gnd vdd FILL
XFILL_1__16318_ gnd vdd FILL
XFILL_2__15869_ gnd vdd FILL
XSFILL43960x51050 gnd vdd FILL
X_9105_ _9105_/A gnd _9105_/Y vdd INVX1
XFILL_1__7551_ gnd vdd FILL
XFILL_0__8758_ gnd vdd FILL
X_7297_ _7297_/A _7297_/B _7297_/C gnd _7385_/D vdd OAI21X1
XFILL_3__8467_ gnd vdd FILL
XFILL_1__16249_ gnd vdd FILL
X_9036_ _9036_/A _8969_/A _9036_/C gnd _9036_/Y vdd OAI21X1
XFILL_0__7709_ gnd vdd FILL
XSFILL44040x60050 gnd vdd FILL
XFILL_1__7482_ gnd vdd FILL
XSFILL99560x3050 gnd vdd FILL
XFILL_3__7418_ gnd vdd FILL
XFILL_3__8398_ gnd vdd FILL
XFILL_4__7191_ gnd vdd FILL
XFILL_1__9221_ gnd vdd FILL
XFILL_3__7349_ gnd vdd FILL
XFILL_2_BUFX2_insert706 gnd vdd FILL
XFILL_2_BUFX2_insert717 gnd vdd FILL
XFILL_1__9152_ gnd vdd FILL
XFILL_2_BUFX2_insert728 gnd vdd FILL
XFILL_2_BUFX2_insert739 gnd vdd FILL
XFILL_1__8103_ gnd vdd FILL
XFILL_3__9019_ gnd vdd FILL
XFILL_1__9083_ gnd vdd FILL
X_9938_ _9936_/Y _9937_/A _9938_/C gnd _9972_/D vdd OAI21X1
XFILL_4__9901_ gnd vdd FILL
X_10820_ _16107_/A gnd _10822_/A vdd INVX1
XSFILL79000x33050 gnd vdd FILL
X_9869_ _9869_/A _9917_/B _9868_/Y gnd _9869_/Y vdd OAI21X1
X_10751_ _10751_/A gnd _10753_/A vdd INVX1
XFILL_4__9763_ gnd vdd FILL
XBUFX2_insert705 _11985_/Y gnd _12096_/C vdd BUFX2
XSFILL3640x80050 gnd vdd FILL
XFILL_4__6975_ gnd vdd FILL
XBUFX2_insert716 _13418_/Y gnd _14174_/C vdd BUFX2
XBUFX2_insert727 _13352_/Y gnd _10127_/A vdd BUFX2
X_13470_ _13423_/A _13398_/A _13423_/B gnd _13470_/Y vdd NAND3X1
XSFILL109480x5050 gnd vdd FILL
X_10682_ _10680_/Y _10681_/A _10682_/C gnd _10732_/D vdd OAI21X1
XBUFX2_insert738 _12402_/Y gnd _8624_/B vdd BUFX2
XSFILL84120x24050 gnd vdd FILL
XFILL_1__9985_ gnd vdd FILL
XFILL_4__8714_ gnd vdd FILL
XBUFX2_insert749 _13344_/Y gnd _9764_/A vdd BUFX2
XFILL_6_BUFX2_insert694 gnd vdd FILL
X_12421_ _12091_/B gnd _12423_/A vdd INVX1
XFILL_4__8645_ gnd vdd FILL
X_15140_ _7804_/A gnd _15140_/Y vdd INVX1
X_12352_ _12352_/A gnd _12352_/Y vdd INVX1
XSFILL23800x39050 gnd vdd FILL
XFILL_1_CLKBUF1_insert121 gnd vdd FILL
XFILL_1__8867_ gnd vdd FILL
XFILL_1_CLKBUF1_insert132 gnd vdd FILL
XSFILL33960x83050 gnd vdd FILL
XFILL_4__8576_ gnd vdd FILL
XFILL_1_CLKBUF1_insert143 gnd vdd FILL
X_11303_ _11536_/C _11303_/B gnd _11433_/C vdd NOR2X1
X_15071_ _9334_/A _15202_/B _15071_/C gnd _15073_/C vdd NAND3X1
XFILL_1_CLKBUF1_insert154 gnd vdd FILL
XFILL_1__7818_ gnd vdd FILL
XFILL_1_CLKBUF1_insert165 gnd vdd FILL
X_12283_ _12227_/A gnd _12307_/C gnd _12283_/Y vdd NAND3X1
XFILL_2__7591_ gnd vdd FILL
XFILL_1_CLKBUF1_insert176 gnd vdd FILL
XFILL_1_CLKBUF1_insert187 gnd vdd FILL
X_14022_ _14022_/A _14022_/B _14022_/C gnd _14023_/B vdd NAND3X1
XFILL_1_CLKBUF1_insert198 gnd vdd FILL
X_11234_ _11376_/B _11376_/A gnd _11234_/Y vdd NOR2X1
XFILL_2_BUFX2_insert8 gnd vdd FILL
XFILL_1__7749_ gnd vdd FILL
XFILL_4__7458_ gnd vdd FILL
XFILL_4__10440_ gnd vdd FILL
X_11165_ _11569_/C _11404_/A _11408_/A gnd _11185_/B vdd OAI21X1
XFILL_2__9261_ gnd vdd FILL
XFILL_1__10260_ gnd vdd FILL
XFILL_3_BUFX2_insert540 gnd vdd FILL
X_10116_ _10114_/Y _10166_/A _10116_/C gnd _10202_/D vdd OAI21X1
XFILL_0__10990_ gnd vdd FILL
XFILL_3_BUFX2_insert551 gnd vdd FILL
X_15973_ _10349_/Q gnd _15974_/C vdd INVX1
XFILL_3_BUFX2_insert562 gnd vdd FILL
XFILL_1__9419_ gnd vdd FILL
X_11096_ _11663_/C _11096_/B _11096_/C gnd _11097_/C vdd OAI21X1
XFILL_2__8212_ gnd vdd FILL
XFILL_5__11730_ gnd vdd FILL
XSFILL3720x60050 gnd vdd FILL
XFILL_3_BUFX2_insert573 gnd vdd FILL
XFILL_4__10371_ gnd vdd FILL
XFILL_4__9128_ gnd vdd FILL
XFILL_2__11550_ gnd vdd FILL
XFILL_1__10191_ gnd vdd FILL
XFILL_3_BUFX2_insert584 gnd vdd FILL
XSFILL29160x17050 gnd vdd FILL
XFILL_3_BUFX2_insert595 gnd vdd FILL
X_10047_ _9975_/B _8511_/B gnd _10047_/Y vdd NAND2X1
XFILL_4__12110_ gnd vdd FILL
X_14924_ _14920_/Y _14924_/B gnd _14924_/Y vdd NOR2X1
XFILL_5__11661_ gnd vdd FILL
XFILL_2__8143_ gnd vdd FILL
XSFILL28920x72050 gnd vdd FILL
XFILL_4__13090_ gnd vdd FILL
XFILL_2__10501_ gnd vdd FILL
XFILL_3__12840_ gnd vdd FILL
XFILL_0__12660_ gnd vdd FILL
XFILL_2__11481_ gnd vdd FILL
XFILL_5__13400_ gnd vdd FILL
XFILL_5__9941_ gnd vdd FILL
X_14855_ _9293_/A gnd _14855_/Y vdd INVX1
XFILL_4__12041_ gnd vdd FILL
XFILL_2__13220_ gnd vdd FILL
XFILL_5__14380_ gnd vdd FILL
XFILL_5__11592_ gnd vdd FILL
XFILL_3__12771_ gnd vdd FILL
XFILL_2__10432_ gnd vdd FILL
XFILL_2__8074_ gnd vdd FILL
XFILL_0__11611_ gnd vdd FILL
XFILL_1__13950_ gnd vdd FILL
XSFILL29000x81050 gnd vdd FILL
XFILL_0__12591_ gnd vdd FILL
X_13806_ _10379_/A _14389_/B _13883_/B _9437_/Q gnd _13815_/A vdd AOI22X1
XFILL_5__13331_ gnd vdd FILL
XFILL_5__9872_ gnd vdd FILL
XFILL_3__14510_ gnd vdd FILL
XFILL_5__10543_ gnd vdd FILL
XFILL_6__12882_ gnd vdd FILL
X_14786_ _9543_/A gnd _14787_/A vdd INVX1
XFILL_3__11722_ gnd vdd FILL
XSFILL85000x7050 gnd vdd FILL
XFILL_2__13151_ gnd vdd FILL
X_11998_ _11998_/A _11998_/B _11998_/C gnd _13086_/B vdd NAND3X1
XFILL_1__12901_ gnd vdd FILL
XFILL_0__14330_ gnd vdd FILL
XFILL_2__10363_ gnd vdd FILL
XFILL_3__15490_ gnd vdd FILL
XFILL_6_BUFX2_insert55 gnd vdd FILL
XFILL_0__11542_ gnd vdd FILL
XFILL_1__13881_ gnd vdd FILL
XFILL_5__8823_ gnd vdd FILL
XFILL_5__13262_ gnd vdd FILL
XSFILL99480x58050 gnd vdd FILL
XFILL_4__15800_ gnd vdd FILL
XFILL_5__16050_ gnd vdd FILL
X_13737_ _13737_/A _13736_/Y _13737_/C gnd _13737_/Y vdd NAND3X1
X_10949_ _10940_/Y _10941_/Y _10948_/Y gnd _10950_/C vdd OAI21X1
XFILL_2__12102_ gnd vdd FILL
XFILL_3__14441_ gnd vdd FILL
XFILL_1__15620_ gnd vdd FILL
XFILL_3__11653_ gnd vdd FILL
XFILL_2__10294_ gnd vdd FILL
XFILL_0__14261_ gnd vdd FILL
XFILL_1__12832_ gnd vdd FILL
XFILL_4__13992_ gnd vdd FILL
XFILL_2__13082_ gnd vdd FILL
XFILL_5__15001_ gnd vdd FILL
XFILL_5__12213_ gnd vdd FILL
XFILL_5__8754_ gnd vdd FILL
XFILL_0__11473_ gnd vdd FILL
XFILL_4__15731_ gnd vdd FILL
X_13668_ _7258_/Q gnd _13668_/Y vdd INVX1
XFILL_0__13212_ gnd vdd FILL
XFILL_0__16000_ gnd vdd FILL
XSFILL49720x51050 gnd vdd FILL
XFILL_2__12033_ gnd vdd FILL
XFILL_3__14372_ gnd vdd FILL
XFILL_2__8976_ gnd vdd FILL
XFILL_5__7705_ gnd vdd FILL
XFILL_1__15551_ gnd vdd FILL
XFILL_0__10424_ gnd vdd FILL
XFILL_3__11584_ gnd vdd FILL
XFILL_1__12763_ gnd vdd FILL
X_15407_ _15407_/A _15407_/B _15407_/C _13867_/Y gnd _15411_/A vdd OAI22X1
XFILL_0__14192_ gnd vdd FILL
XFILL_0_BUFX2_insert430 gnd vdd FILL
X_12619_ vdd memoryOutData[17] gnd _12620_/C vdd NAND2X1
XFILL_3__16111_ gnd vdd FILL
XSFILL38920x50 gnd vdd FILL
XSFILL53960x14050 gnd vdd FILL
XFILL_0_BUFX2_insert441 gnd vdd FILL
XFILL_5__12144_ gnd vdd FILL
XFILL_3__13323_ gnd vdd FILL
X_16387_ _16439_/Q gnd _16387_/Y vdd INVX1
XFILL_0_BUFX2_insert452 gnd vdd FILL
XFILL_0__7991_ gnd vdd FILL
XFILL_3__10535_ gnd vdd FILL
X_13599_ _9215_/A gnd _13599_/Y vdd INVX1
XFILL_4__15662_ gnd vdd FILL
XFILL_1__14502_ gnd vdd FILL
XFILL_0_BUFX2_insert463 gnd vdd FILL
XFILL_4__12874_ gnd vdd FILL
XFILL_2__7927_ gnd vdd FILL
XFILL_0__13143_ gnd vdd FILL
XSFILL109480x43050 gnd vdd FILL
XFILL_1__11714_ gnd vdd FILL
XFILL_6__16222_ gnd vdd FILL
XFILL_5__7636_ gnd vdd FILL
XFILL_1__15482_ gnd vdd FILL
XFILL_0_BUFX2_insert474 gnd vdd FILL
X_15338_ _15338_/A _15338_/B _15338_/C gnd _12842_/B vdd AOI21X1
XFILL_0__9730_ gnd vdd FILL
XFILL_6__13434_ gnd vdd FILL
XFILL_0_BUFX2_insert485 gnd vdd FILL
XFILL_0_BUFX2_insert496 gnd vdd FILL
XFILL_3__16042_ gnd vdd FILL
XFILL_4__14613_ gnd vdd FILL
XFILL_5__12075_ gnd vdd FILL
XFILL_0__6942_ gnd vdd FILL
XFILL_4__11825_ gnd vdd FILL
XFILL_6__10646_ gnd vdd FILL
XFILL_3__13254_ gnd vdd FILL
XFILL_4__15593_ gnd vdd FILL
XSFILL54040x23050 gnd vdd FILL
XFILL_2__7858_ gnd vdd FILL
XFILL_1__14433_ gnd vdd FILL
XFILL_2__13984_ gnd vdd FILL
XFILL_1__11645_ gnd vdd FILL
XFILL_5__7567_ gnd vdd FILL
XFILL_5__15903_ gnd vdd FILL
XFILL_0__10286_ gnd vdd FILL
X_7220_ _7220_/A _7250_/B _7220_/C gnd _7274_/D vdd OAI21X1
XFILL_5__11026_ gnd vdd FILL
XFILL_0__9661_ gnd vdd FILL
XFILL_3__12205_ gnd vdd FILL
X_15269_ _15268_/Y _16151_/B _16225_/C _13701_/B gnd _15269_/Y vdd OAI22X1
XFILL_0__6873_ gnd vdd FILL
XFILL_2__15723_ gnd vdd FILL
XFILL_4__14544_ gnd vdd FILL
XFILL_4__11756_ gnd vdd FILL
XFILL_0__12025_ gnd vdd FILL
XFILL_3__9370_ gnd vdd FILL
XFILL_1__14364_ gnd vdd FILL
XFILL_3__10397_ gnd vdd FILL
XFILL_1__11576_ gnd vdd FILL
XFILL_0__8612_ gnd vdd FILL
XFILL_6__12316_ gnd vdd FILL
XFILL_5__7498_ gnd vdd FILL
XFILL_5__15834_ gnd vdd FILL
XFILL_4__10707_ gnd vdd FILL
X_7151_ _7105_/A _7791_/CLK _9711_/R vdd _7151_/D gnd vdd DFFSR
XFILL_6__16084_ gnd vdd FILL
XFILL_3__8321_ gnd vdd FILL
XFILL_4__14475_ gnd vdd FILL
XFILL_3__12136_ gnd vdd FILL
XFILL_0__9592_ gnd vdd FILL
XFILL_1__16103_ gnd vdd FILL
XFILL_2__9528_ gnd vdd FILL
XFILL_1__13315_ gnd vdd FILL
XSFILL43880x66050 gnd vdd FILL
XFILL_2__15654_ gnd vdd FILL
XFILL_4__11687_ gnd vdd FILL
XFILL_1__10527_ gnd vdd FILL
XFILL_2__12866_ gnd vdd FILL
XFILL_5__9237_ gnd vdd FILL
XCLKBUF1_insert120 CLKBUF1_insert206/A gnd _7642_/CLK vdd CLKBUF1
XFILL_6__15035_ gnd vdd FILL
XFILL_1__14295_ gnd vdd FILL
XCLKBUF1_insert131 CLKBUF1_insert192/A gnd _8537_/CLK vdd CLKBUF1
XFILL_4__16214_ gnd vdd FILL
XFILL_4__13426_ gnd vdd FILL
XFILL_4__10638_ gnd vdd FILL
XCLKBUF1_insert142 CLKBUF1_insert192/A gnd _7021_/CLK vdd CLKBUF1
XFILL_2__14605_ gnd vdd FILL
XFILL_5__15765_ gnd vdd FILL
X_7082_ _7067_/A _9898_/B gnd _7083_/C vdd NAND2X1
XFILL_3__8252_ gnd vdd FILL
XFILL_5__12977_ gnd vdd FILL
XFILL_1__16034_ gnd vdd FILL
XFILL_3__12067_ gnd vdd FILL
XSFILL18680x42050 gnd vdd FILL
XFILL_2__11817_ gnd vdd FILL
XFILL_1__13246_ gnd vdd FILL
XCLKBUF1_insert153 CLKBUF1_insert187/A gnd _13180_/CLK vdd CLKBUF1
XFILL_2__15585_ gnd vdd FILL
XCLKBUF1_insert164 CLKBUF1_insert193/A gnd _8663_/CLK vdd CLKBUF1
XFILL_5__9168_ gnd vdd FILL
XSFILL98520x74050 gnd vdd FILL
XFILL_0__13976_ gnd vdd FILL
XFILL_5__14716_ gnd vdd FILL
XCLKBUF1_insert175 CLKBUF1_insert216/A gnd _8022_/CLK vdd CLKBUF1
XFILL_4__13357_ gnd vdd FILL
XFILL_3__7203_ gnd vdd FILL
XCLKBUF1_insert186 CLKBUF1_insert218/A gnd _9453_/CLK vdd CLKBUF1
XFILL_0__8474_ gnd vdd FILL
XFILL_5__11928_ gnd vdd FILL
XFILL_3__11018_ gnd vdd FILL
XFILL_4__16145_ gnd vdd FILL
XSFILL84360x80050 gnd vdd FILL
XFILL_5__15696_ gnd vdd FILL
XFILL_2__14536_ gnd vdd FILL
XFILL_4__10569_ gnd vdd FILL
XFILL_5__8119_ gnd vdd FILL
XFILL_0__15715_ gnd vdd FILL
XFILL_3__8183_ gnd vdd FILL
XFILL_2__11748_ gnd vdd FILL
XCLKBUF1_insert197 CLKBUF1_insert150/A gnd _9578_/CLK vdd CLKBUF1
XFILL_1__10389_ gnd vdd FILL
XFILL_5__9099_ gnd vdd FILL
XFILL_0__7425_ gnd vdd FILL
XFILL_4__12308_ gnd vdd FILL
XFILL_6__11129_ gnd vdd FILL
XSFILL49000x12050 gnd vdd FILL
XFILL_5__14647_ gnd vdd FILL
XFILL_4__16076_ gnd vdd FILL
XFILL_4__13288_ gnd vdd FILL
XFILL_1__12128_ gnd vdd FILL
XFILL_3__15826_ gnd vdd FILL
XFILL_5__11859_ gnd vdd FILL
XFILL_2__14467_ gnd vdd FILL
XFILL112440x6050 gnd vdd FILL
XFILL_0__15646_ gnd vdd FILL
XFILL_2__11679_ gnd vdd FILL
XFILL_0__12858_ gnd vdd FILL
XFILL_2__16206_ gnd vdd FILL
XFILL_0__7356_ gnd vdd FILL
XFILL_4__15027_ gnd vdd FILL
XFILL_4__12239_ gnd vdd FILL
XSFILL109560x23050 gnd vdd FILL
XFILL_5__14578_ gnd vdd FILL
XFILL_2__13418_ gnd vdd FILL
XFILL_1__12059_ gnd vdd FILL
XFILL_3__7065_ gnd vdd FILL
XFILL_3__12969_ gnd vdd FILL
X_7984_ _8006_/B _9008_/B gnd _7985_/C vdd NAND2X1
XFILL_3__15757_ gnd vdd FILL
XSFILL38840x55050 gnd vdd FILL
XFILL_2__14398_ gnd vdd FILL
XFILL_0__11809_ gnd vdd FILL
XFILL_0__12789_ gnd vdd FILL
XFILL_5__16317_ gnd vdd FILL
XFILL_0__15577_ gnd vdd FILL
XFILL112360x62050 gnd vdd FILL
XFILL_5__13529_ gnd vdd FILL
X_9723_ _9721_/Y _9770_/A _9723_/C gnd _9815_/D vdd OAI21X1
XFILL_0__7287_ gnd vdd FILL
XFILL_3__14708_ gnd vdd FILL
X_6935_ _6935_/A gnd _6935_/Y vdd INVX1
XFILL_2__16137_ gnd vdd FILL
XFILL_2__13349_ gnd vdd FILL
XFILL_3__15688_ gnd vdd FILL
XFILL_0__14528_ gnd vdd FILL
XFILL_0__9026_ gnd vdd FILL
XSFILL74120x8050 gnd vdd FILL
XSFILL113720x8050 gnd vdd FILL
XFILL_5__16248_ gnd vdd FILL
X_9654_ _9613_/B _8630_/B gnd _9655_/C vdd NAND2X1
XFILL_3__14639_ gnd vdd FILL
X_6866_ _6866_/A gnd memoryAddress[28] vdd BUFX2
XFILL_1__15818_ gnd vdd FILL
XFILL_2__16068_ gnd vdd FILL
XFILL_0__14459_ gnd vdd FILL
XFILL_6__7745_ gnd vdd FILL
X_8605_ _8675_/Q gnd _8607_/A vdd INVX1
XFILL_4__15929_ gnd vdd FILL
XFILL_5__16179_ gnd vdd FILL
XFILL_2__15019_ gnd vdd FILL
X_9585_ _9543_/A _7537_/CLK _7537_/R vdd _9585_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert602 gnd vdd FILL
XFILL_3__7967_ gnd vdd FILL
XFILL_1__15749_ gnd vdd FILL
XFILL_5_BUFX2_insert613 gnd vdd FILL
XFILL_5_BUFX2_insert624 gnd vdd FILL
XSFILL18760x22050 gnd vdd FILL
XFILL_1__9770_ gnd vdd FILL
XSFILL8600x32050 gnd vdd FILL
XFILL_3__16309_ gnd vdd FILL
X_8536_ _8536_/Q _7143_/CLK _7015_/R vdd _8446_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert635 gnd vdd FILL
XSFILL44040x55050 gnd vdd FILL
XFILL_1__6982_ gnd vdd FILL
XFILL_3__6918_ gnd vdd FILL
XFILL_5_BUFX2_insert646 gnd vdd FILL
XFILL_0__16129_ gnd vdd FILL
XFILL_5_BUFX2_insert657 gnd vdd FILL
XFILL_6__9415_ gnd vdd FILL
XFILL_5_BUFX2_insert668 gnd vdd FILL
XFILL_1__8721_ gnd vdd FILL
XFILL_0__9928_ gnd vdd FILL
XFILL_5_BUFX2_insert679 gnd vdd FILL
XFILL_3__9637_ gnd vdd FILL
X_8467_ _8465_/Y _8469_/A _8467_/C gnd _8543_/D vdd OAI21X1
XFILL_3__6849_ gnd vdd FILL
XFILL_1__8652_ gnd vdd FILL
XFILL_0__9859_ gnd vdd FILL
XSFILL23880x13050 gnd vdd FILL
X_7418_ _7470_/B _9082_/B gnd _7419_/C vdd NAND2X1
X_8398_ _8360_/B _8654_/B gnd _8399_/C vdd NAND2X1
XFILL_4__8361_ gnd vdd FILL
XFILL111800x76050 gnd vdd FILL
XFILL_1__7603_ gnd vdd FILL
X_7349_ _7403_/Q gnd _7351_/A vdd INVX1
XFILL_4__7312_ gnd vdd FILL
XFILL_3__8519_ gnd vdd FILL
XSFILL38920x35050 gnd vdd FILL
XFILL_1__8583_ gnd vdd FILL
XFILL_2_CLKBUF1_insert205 gnd vdd FILL
XFILL112440x42050 gnd vdd FILL
XSFILL53880x50 gnd vdd FILL
XFILL_2_CLKBUF1_insert216 gnd vdd FILL
XSFILL64200x68050 gnd vdd FILL
XFILL_3__9499_ gnd vdd FILL
XFILL_4__7243_ gnd vdd FILL
XSFILL39000x44050 gnd vdd FILL
X_9019_ _9069_/Q gnd _9019_/Y vdd INVX1
XFILL_1__7465_ gnd vdd FILL
XFILL_4__7174_ gnd vdd FILL
XFILL_2_BUFX2_insert503 gnd vdd FILL
XSFILL3640x75050 gnd vdd FILL
X_12970_ vdd _12970_/B gnd _12971_/C vdd NAND2X1
XFILL_2_BUFX2_insert514 gnd vdd FILL
XFILL_2_BUFX2_insert525 gnd vdd FILL
XFILL_2_BUFX2_insert536 gnd vdd FILL
XFILL_2_BUFX2_insert547 gnd vdd FILL
XSFILL94280x63050 gnd vdd FILL
X_11921_ _11921_/A _12031_/B gnd _11922_/C vdd NAND2X1
XFILL_2_BUFX2_insert558 gnd vdd FILL
XFILL_1__9135_ gnd vdd FILL
XFILL_2_BUFX2_insert569 gnd vdd FILL
X_14640_ _13467_/A _14638_/Y _14640_/C _16024_/D gnd _14644_/B vdd OAI22X1
X_11852_ _12005_/A _12449_/B _11852_/C gnd _11853_/C vdd NOR3X1
XFILL_6_BUFX2_insert1022 gnd vdd FILL
X_10803_ _10822_/B _9267_/B gnd _10803_/Y vdd NAND2X1
XSFILL33960x78050 gnd vdd FILL
X_14571_ _13865_/C _7739_/A _7611_/A _13848_/C gnd _14580_/A vdd AOI22X1
XFILL_1__8017_ gnd vdd FILL
X_11783_ _11781_/Y _11782_/Y gnd _11783_/Y vdd OR2X2
X_16310_ _8437_/Q gnd _16310_/Y vdd INVX1
XFILL_6_BUFX2_insert1088 gnd vdd FILL
XBUFX2_insert502 BUFX2_insert520/A gnd _9823_/R vdd BUFX2
X_13522_ _13520_/Y _14030_/A _13467_/A _13522_/D gnd _13526_/B vdd OAI22X1
X_10734_ _14598_/A _8942_/CLK _8942_/R vdd _10688_/Y gnd vdd DFFSR
XFILL_2__8830_ gnd vdd FILL
XBUFX2_insert513 BUFX2_insert496/A gnd _7131_/R vdd BUFX2
XBUFX2_insert524 BUFX2_insert524/A gnd _7911_/R vdd BUFX2
XBUFX2_insert535 BUFX2_insert559/A gnd _9566_/R vdd BUFX2
XFILL_6_BUFX2_insert480 gnd vdd FILL
X_16241_ _16238_/Y _16240_/Y gnd _16242_/B vdd NOR2X1
XBUFX2_insert546 BUFX2_insert556/A gnd _9441_/R vdd BUFX2
XFILL_4__6958_ gnd vdd FILL
XFILL_4__9746_ gnd vdd FILL
X_13453_ _9974_/A gnd _13453_/Y vdd INVX1
XBUFX2_insert557 BUFX2_insert524/A gnd _7413_/R vdd BUFX2
XFILL_5__10190_ gnd vdd FILL
X_10665_ _10727_/Q gnd _10665_/Y vdd INVX1
XBUFX2_insert568 BUFX2_insert518/A gnd _8819_/R vdd BUFX2
XFILL_2__8761_ gnd vdd FILL
XSFILL18760x3050 gnd vdd FILL
XBUFX2_insert579 BUFX2_insert600/A gnd _8176_/R vdd BUFX2
XFILL_4__9677_ gnd vdd FILL
X_12404_ _12371_/A _12683_/Q gnd _12405_/C vdd NAND2X1
XFILL_5__8470_ gnd vdd FILL
X_16172_ _16172_/A _16172_/B _16172_/C gnd _16179_/B vdd NAND3X1
XFILL_4__6889_ gnd vdd FILL
XSFILL58920x8050 gnd vdd FILL
XFILL_2__7712_ gnd vdd FILL
X_13384_ _9302_/Q gnd _15056_/A vdd INVX1
XFILL_3__10320_ gnd vdd FILL
X_10596_ _10596_/Q _9188_/CLK _8801_/R vdd _10530_/Y gnd vdd DFFSR
XFILL_0__10140_ gnd vdd FILL
XFILL_5__7421_ gnd vdd FILL
XFILL_4__8628_ gnd vdd FILL
XFILL_1__9899_ gnd vdd FILL
XSFILL53480x31050 gnd vdd FILL
X_15123_ _16306_/A _15123_/B _15558_/D _13525_/D gnd _15124_/B vdd OAI22X1
X_12335_ _12327_/A gnd _12311_/C gnd _12338_/A vdd NAND3X1
XFILL_4__11610_ gnd vdd FILL
XFILL_4_BUFX2_insert1070 gnd vdd FILL
XFILL_4__12590_ gnd vdd FILL
XFILL_3__10251_ gnd vdd FILL
XSFILL28920x67050 gnd vdd FILL
XFILL_1__11430_ gnd vdd FILL
XSFILL94360x43050 gnd vdd FILL
XFILL_4_BUFX2_insert1092 gnd vdd FILL
XFILL_2__10981_ gnd vdd FILL
XFILL_5__7352_ gnd vdd FILL
X_15054_ _14986_/A _16037_/B _14981_/Y gnd _15054_/Y vdd NAND3X1
XFILL_6__10362_ gnd vdd FILL
XFILL_5__12900_ gnd vdd FILL
X_12266_ _12263_/Y _12266_/B _12266_/C gnd _12266_/Y vdd NAND3X1
XFILL_4__11541_ gnd vdd FILL
XFILL_2__12720_ gnd vdd FILL
XFILL_5__13880_ gnd vdd FILL
XFILL_3__10182_ gnd vdd FILL
XFILL_2__7574_ gnd vdd FILL
XFILL_1__11361_ gnd vdd FILL
XFILL_6__12101_ gnd vdd FILL
X_14005_ _7831_/A gnd _14007_/A vdd INVX1
X_11217_ gnd _11216_/Y gnd _11218_/B vdd NOR2X1
XFILL_4__14260_ gnd vdd FILL
XFILL_5__12831_ gnd vdd FILL
XFILL_1__13100_ gnd vdd FILL
XFILL_1__10312_ gnd vdd FILL
X_12197_ _12201_/B _12946_/Q gnd _12198_/C vdd NAND2X1
XFILL_4__11472_ gnd vdd FILL
XFILL_2__12651_ gnd vdd FILL
XFILL_3__14990_ gnd vdd FILL
XFILL_5__9022_ gnd vdd FILL
XFILL_1__14080_ gnd vdd FILL
XFILL_0__13830_ gnd vdd FILL
XFILL_1__11292_ gnd vdd FILL
XFILL_4__13211_ gnd vdd FILL
XFILL_4__10423_ gnd vdd FILL
XFILL_5__15550_ gnd vdd FILL
X_11148_ _12282_/Y _11617_/A gnd _11149_/C vdd NOR2X1
XFILL_5__12762_ gnd vdd FILL
XFILL_4__14191_ gnd vdd FILL
XFILL_2__9244_ gnd vdd FILL
XFILL_1__13031_ gnd vdd FILL
XFILL_2__11602_ gnd vdd FILL
XFILL_3__13941_ gnd vdd FILL
XFILL_2__15370_ gnd vdd FILL
XFILL_1__10243_ gnd vdd FILL
XFILL_2__12582_ gnd vdd FILL
XFILL_3_BUFX2_insert370 gnd vdd FILL
XFILL_0__10973_ gnd vdd FILL
XFILL_3_BUFX2_insert381 gnd vdd FILL
XFILL_5__14501_ gnd vdd FILL
XFILL_0__13761_ gnd vdd FILL
XSFILL74280x10050 gnd vdd FILL
XFILL_4__13142_ gnd vdd FILL
XFILL_3_BUFX2_insert392 gnd vdd FILL
XFILL_5__11713_ gnd vdd FILL
X_15956_ _15644_/D _14533_/Y _15170_/D _14544_/Y gnd _15956_/Y vdd OAI22X1
XFILL_2__14321_ gnd vdd FILL
X_11079_ _12141_/Y _11078_/Y gnd _11079_/Y vdd NAND2X1
XFILL_5__15481_ gnd vdd FILL
XSFILL48440x20050 gnd vdd FILL
XFILL_3__13872_ gnd vdd FILL
XFILL_0__15500_ gnd vdd FILL
XFILL_2__11533_ gnd vdd FILL
XFILL_1__10174_ gnd vdd FILL
XFILL_0__12712_ gnd vdd FILL
XSFILL84120x3050 gnd vdd FILL
XFILL_0__13692_ gnd vdd FILL
XFILL_0__7210_ gnd vdd FILL
XSFILL59080x71050 gnd vdd FILL
XSFILL89320x32050 gnd vdd FILL
XFILL_5__14432_ gnd vdd FILL
X_14907_ _14907_/A _14907_/B gnd _14929_/B vdd NOR2X1
XFILL_2__8126_ gnd vdd FILL
XFILL_3__15611_ gnd vdd FILL
XFILL_3__12823_ gnd vdd FILL
XFILL_5__11644_ gnd vdd FILL
XFILL_0__8190_ gnd vdd FILL
X_15887_ _16106_/A _15885_/Y _15726_/A _15886_/Y gnd _15887_/Y vdd OAI22X1
XFILL_2__14252_ gnd vdd FILL
XFILL_4__10285_ gnd vdd FILL
XFILL_0__12643_ gnd vdd FILL
XFILL_0__15431_ gnd vdd FILL
XFILL_2__11464_ gnd vdd FILL
XFILL_1__14982_ gnd vdd FILL
XFILL_5__9924_ gnd vdd FILL
XFILL_4__12024_ gnd vdd FILL
X_14838_ _8819_/Q _13853_/B _14838_/C gnd _14838_/Y vdd AOI21X1
XFILL_3__15542_ gnd vdd FILL
XSFILL3800x35050 gnd vdd FILL
XFILL_5__14363_ gnd vdd FILL
XFILL_5__11575_ gnd vdd FILL
XFILL_3__12754_ gnd vdd FILL
XFILL_2__10415_ gnd vdd FILL
XFILL_2__8057_ gnd vdd FILL
XFILL112280x77050 gnd vdd FILL
XSFILL13400x68050 gnd vdd FILL
XFILL_2__14183_ gnd vdd FILL
XFILL_1__13933_ gnd vdd FILL
XSFILL54040x18050 gnd vdd FILL
XFILL_0__12574_ gnd vdd FILL
XFILL_0__15362_ gnd vdd FILL
XFILL_5__16102_ gnd vdd FILL
XFILL_2__11395_ gnd vdd FILL
XFILL_5__13314_ gnd vdd FILL
XFILL_5__9855_ gnd vdd FILL
XFILL_0__7072_ gnd vdd FILL
XFILL_3__11705_ gnd vdd FILL
XFILL_5__10526_ gnd vdd FILL
X_14769_ _10737_/Q gnd _16127_/B vdd INVX1
XFILL_2__13134_ gnd vdd FILL
XFILL_5__14294_ gnd vdd FILL
XFILL_3__15473_ gnd vdd FILL
XFILL_3__8870_ gnd vdd FILL
XFILL_0__14313_ gnd vdd FILL
XFILL_0__11525_ gnd vdd FILL
XFILL_1__13864_ gnd vdd FILL
XFILL_0__15293_ gnd vdd FILL
XFILL_5__16033_ gnd vdd FILL
XFILL_5__13245_ gnd vdd FILL
XFILL_5__9786_ gnd vdd FILL
XFILL_3__14424_ gnd vdd FILL
XFILL_3__7821_ gnd vdd FILL
XFILL_3__11636_ gnd vdd FILL
XFILL_1__15603_ gnd vdd FILL
XFILL_4_CLKBUF1_insert160 gnd vdd FILL
XFILL_2__10277_ gnd vdd FILL
XFILL_0__14244_ gnd vdd FILL
XFILL_4__13975_ gnd vdd FILL
XFILL_4_CLKBUF1_insert171 gnd vdd FILL
XFILL_0__11456_ gnd vdd FILL
XFILL_1__13795_ gnd vdd FILL
XFILL_5__8737_ gnd vdd FILL
XFILL_4_CLKBUF1_insert182 gnd vdd FILL
XFILL_4_CLKBUF1_insert193 gnd vdd FILL
XFILL_4__15714_ gnd vdd FILL
X_16439_ _16439_/Q _9453_/CLK _9453_/R vdd _16389_/Y gnd vdd DFFSR
XFILL_2__12016_ gnd vdd FILL
X_9370_ _9442_/Q gnd _9370_/Y vdd INVX1
XFILL_3__14355_ gnd vdd FILL
XFILL_5__10388_ gnd vdd FILL
XFILL_2__8959_ gnd vdd FILL
XFILL_0__10407_ gnd vdd FILL
XFILL_1__15534_ gnd vdd FILL
XFILL_3__11567_ gnd vdd FILL
XFILL_3__7752_ gnd vdd FILL
XFILL_1__12746_ gnd vdd FILL
XFILL_0__14175_ gnd vdd FILL
XSFILL18680x37050 gnd vdd FILL
XFILL_0_BUFX2_insert260 gnd vdd FILL
XFILL_6__7461_ gnd vdd FILL
XFILL_0_BUFX2_insert271 gnd vdd FILL
XFILL_0__11387_ gnd vdd FILL
XFILL_3__13306_ gnd vdd FILL
X_8321_ _8319_/Y _8321_/B _8320_/Y gnd _8409_/D vdd OAI21X1
XFILL_0_BUFX2_insert282 gnd vdd FILL
XFILL_5__12127_ gnd vdd FILL
XFILL_0__7974_ gnd vdd FILL
XFILL_4__15645_ gnd vdd FILL
XFILL_3__10518_ gnd vdd FILL
XFILL_0__13126_ gnd vdd FILL
XFILL_4__12857_ gnd vdd FILL
XSFILL33720x40050 gnd vdd FILL
XFILL_0_BUFX2_insert293 gnd vdd FILL
XFILL_3__14286_ gnd vdd FILL
XSFILL84360x75050 gnd vdd FILL
XFILL_3__7683_ gnd vdd FILL
XFILL_3__11498_ gnd vdd FILL
XFILL_1__15465_ gnd vdd FILL
XFILL_5__7619_ gnd vdd FILL
XFILL_4_BUFX2_insert609 gnd vdd FILL
X_8252_ _8249_/A _8636_/B gnd _8253_/C vdd NAND2X1
XFILL_3__16025_ gnd vdd FILL
XFILL_0__6925_ gnd vdd FILL
XFILL_5__8599_ gnd vdd FILL
XFILL_5__12058_ gnd vdd FILL
XFILL_3__13237_ gnd vdd FILL
XFILL_3__9422_ gnd vdd FILL
XSFILL74600x52050 gnd vdd FILL
XFILL_4__11808_ gnd vdd FILL
XFILL_3__10449_ gnd vdd FILL
XFILL_4__15576_ gnd vdd FILL
XFILL_1__14416_ gnd vdd FILL
XFILL_4__12788_ gnd vdd FILL
XSFILL59160x51050 gnd vdd FILL
XSFILL89400x12050 gnd vdd FILL
XFILL_1__11628_ gnd vdd FILL
XFILL_2__13967_ gnd vdd FILL
XFILL_6__9131_ gnd vdd FILL
X_7203_ _7269_/Q gnd _7203_/Y vdd INVX1
XFILL_1__15396_ gnd vdd FILL
XFILL_0__10269_ gnd vdd FILL
XFILL_5__11009_ gnd vdd FILL
XFILL_0__9644_ gnd vdd FILL
X_8183_ _8183_/A _8232_/B gnd _8184_/C vdd NAND2X1
XFILL_0__6856_ gnd vdd FILL
XFILL_4__14527_ gnd vdd FILL
XSFILL109560x18050 gnd vdd FILL
XFILL_3__13168_ gnd vdd FILL
XFILL_2__15706_ gnd vdd FILL
XFILL_3__9353_ gnd vdd FILL
XFILL_2_BUFX2_insert20 gnd vdd FILL
XFILL_0__12008_ gnd vdd FILL
XFILL_2__12918_ gnd vdd FILL
XFILL_4__11739_ gnd vdd FILL
XFILL_2_BUFX2_insert31 gnd vdd FILL
XFILL_1__14347_ gnd vdd FILL
XFILL_2_BUFX2_insert42 gnd vdd FILL
XFILL_2__13898_ gnd vdd FILL
XFILL_1__11559_ gnd vdd FILL
X_7134_ _7054_/A _8926_/CLK _7262_/R vdd _7134_/D gnd vdd DFFSR
XFILL_5__15817_ gnd vdd FILL
XFILL_2_BUFX2_insert53 gnd vdd FILL
XFILL112360x57050 gnd vdd FILL
XFILL_3__12119_ gnd vdd FILL
XFILL_4__14458_ gnd vdd FILL
XFILL_2__15637_ gnd vdd FILL
XFILL_2_BUFX2_insert64 gnd vdd FILL
XFILL_2_BUFX2_insert75 gnd vdd FILL
XFILL_2__12849_ gnd vdd FILL
XFILL_3__13099_ gnd vdd FILL
XFILL_3__9284_ gnd vdd FILL
XFILL_2_BUFX2_insert86 gnd vdd FILL
XFILL_1__14278_ gnd vdd FILL
XFILL_0__8526_ gnd vdd FILL
XFILL_2_BUFX2_insert97 gnd vdd FILL
XFILL_4__13409_ gnd vdd FILL
X_7065_ _7065_/A _7064_/A _7065_/C gnd _7137_/D vdd OAI21X1
XFILL_5__15748_ gnd vdd FILL
XFILL_1__16017_ gnd vdd FILL
XFILL_3__8235_ gnd vdd FILL
XFILL_1__13229_ gnd vdd FILL
XFILL_2__15568_ gnd vdd FILL
XFILL_4__14389_ gnd vdd FILL
XFILL_0__13959_ gnd vdd FILL
XFILL_0__8457_ gnd vdd FILL
XFILL_4__16128_ gnd vdd FILL
XFILL_1__7250_ gnd vdd FILL
XFILL_5__15679_ gnd vdd FILL
XFILL_2__14519_ gnd vdd FILL
XFILL_2__15499_ gnd vdd FILL
XSFILL18760x17050 gnd vdd FILL
XFILL_3__7117_ gnd vdd FILL
XFILL_1__7181_ gnd vdd FILL
XFILL_0__8388_ gnd vdd FILL
XFILL_3__15809_ gnd vdd FILL
XFILL_4__16059_ gnd vdd FILL
XSFILL114520x73050 gnd vdd FILL
XSFILL8600x27050 gnd vdd FILL
XFILL_0__15629_ gnd vdd FILL
XFILL_3__8097_ gnd vdd FILL
XFILL_0__7339_ gnd vdd FILL
XFILL_3__7048_ gnd vdd FILL
X_7967_ _7967_/A _7955_/B _7966_/Y gnd _7967_/Y vdd OAI21X1
XFILL_4__7930_ gnd vdd FILL
X_9706_ _9650_/A _9578_/CLK _7153_/R vdd _9652_/Y gnd vdd DFFSR
XSFILL59240x31050 gnd vdd FILL
X_6918_ _6955_/B _6918_/B gnd _6918_/Y vdd NAND2X1
XFILL_4__7861_ gnd vdd FILL
X_7898_ _7810_/A _7915_/CLK _7915_/R vdd _7898_/D gnd vdd DFFSR
XFILL_0__9009_ gnd vdd FILL
X_9637_ _9635_/Y _9615_/A _9637_/C gnd _9637_/Y vdd OAI21X1
XFILL_4__9600_ gnd vdd FILL
X_6849_ _6849_/A gnd memoryAddress[11] vdd BUFX2
XFILL111960x30050 gnd vdd FILL
XFILL_3__8999_ gnd vdd FILL
XFILL112440x37050 gnd vdd FILL
XFILL_5_BUFX2_insert410 gnd vdd FILL
XFILL_4__9531_ gnd vdd FILL
XFILL_5_BUFX2_insert421 gnd vdd FILL
X_9568_ _9492_/A _9568_/CLK _8431_/R vdd _9494_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert432 gnd vdd FILL
XFILL_5_BUFX2_insert443 gnd vdd FILL
XSFILL39000x39050 gnd vdd FILL
X_10450_ _10450_/A _10450_/B _10449_/Y gnd _10484_/D vdd OAI21X1
XFILL_5_BUFX2_insert454 gnd vdd FILL
XFILL_1__9753_ gnd vdd FILL
X_8519_ _8519_/A gnd _8519_/Y vdd INVX1
XFILL_1__6965_ gnd vdd FILL
XFILL_5_BUFX2_insert465 gnd vdd FILL
XFILL_4__9462_ gnd vdd FILL
X_9499_ _9466_/A _9371_/B gnd _9500_/C vdd NAND2X1
XFILL_5_BUFX2_insert476 gnd vdd FILL
XFILL_5_BUFX2_insert487 gnd vdd FILL
XFILL_1__8704_ gnd vdd FILL
XFILL_5_BUFX2_insert498 gnd vdd FILL
X_10381_ _10379_/Y _10423_/B _10381_/C gnd _10461_/D vdd OAI21X1
XFILL_1__9684_ gnd vdd FILL
XFILL_1__6896_ gnd vdd FILL
XFILL_4__9393_ gnd vdd FILL
X_12120_ _12120_/A _12123_/B _12119_/Y gnd _12120_/Y vdd OAI21X1
XFILL_1__8635_ gnd vdd FILL
XSFILL94280x58050 gnd vdd FILL
XFILL_4__8344_ gnd vdd FILL
X_12051_ _12007_/A _11936_/B _12031_/C gnd _12051_/Y vdd NAND3X1
XSFILL69080x34050 gnd vdd FILL
XFILL_1__8566_ gnd vdd FILL
XFILL_4__8275_ gnd vdd FILL
X_11002_ _12226_/Y _11002_/B gnd _11006_/A vdd NOR2X1
XFILL_4__7226_ gnd vdd FILL
XFILL_1__8497_ gnd vdd FILL
XFILL_2__7290_ gnd vdd FILL
XSFILL104280x43050 gnd vdd FILL
X_15810_ _15810_/A _15803_/Y gnd _15811_/C vdd NAND2X1
XFILL_2_BUFX2_insert300 gnd vdd FILL
XFILL_1__7448_ gnd vdd FILL
XFILL_2_BUFX2_insert311 gnd vdd FILL
XFILL_2_BUFX2_insert322 gnd vdd FILL
XFILL_2_BUFX2_insert333 gnd vdd FILL
X_15741_ _14301_/A _15565_/B _15569_/C _14270_/Y gnd _15742_/C vdd OAI22X1
XSFILL23800x52050 gnd vdd FILL
X_12953_ _12951_/Y vdd _12953_/C gnd _13047_/D vdd OAI21X1
XFILL_2_BUFX2_insert344 gnd vdd FILL
XFILL_2_BUFX2_insert355 gnd vdd FILL
XFILL_1__7379_ gnd vdd FILL
XFILL_2_BUFX2_insert366 gnd vdd FILL
XFILL_5__7970_ gnd vdd FILL
X_11904_ _11902_/Y _11900_/A _11903_/Y gnd _6843_/A vdd OAI21X1
XFILL_4__7088_ gnd vdd FILL
XFILL_2_BUFX2_insert377 gnd vdd FILL
XFILL_2_BUFX2_insert388 gnd vdd FILL
X_15672_ _15670_/Y _15392_/B _15392_/C _15672_/D gnd _15672_/Y vdd OAI22X1
XFILL_1__9118_ gnd vdd FILL
X_12884_ vdd _12884_/B gnd _12885_/C vdd NAND2X1
XFILL_2_BUFX2_insert399 gnd vdd FILL
XFILL_5__6921_ gnd vdd FILL
X_14623_ _8046_/Q gnd _14623_/Y vdd INVX1
XFILL_5__11360_ gnd vdd FILL
X_11835_ _11835_/A _11427_/A _11835_/C gnd _11836_/C vdd AOI21X1
XFILL_2__9931_ gnd vdd FILL
XFILL_2__11180_ gnd vdd FILL
XFILL_1__10930_ gnd vdd FILL
XFILL_5__9640_ gnd vdd FILL
XFILL_5__6852_ gnd vdd FILL
XSFILL94360x38050 gnd vdd FILL
XFILL_5__10311_ gnd vdd FILL
X_14554_ _7021_/Q gnd _14554_/Y vdd INVX1
XFILL_5__11291_ gnd vdd FILL
XFILL_2__10131_ gnd vdd FILL
X_11766_ _11019_/Y gnd _11766_/Y vdd INVX1
XFILL_3__12470_ gnd vdd FILL
XFILL_2__9862_ gnd vdd FILL
XFILL_0__11310_ gnd vdd FILL
XBUFX2_insert310 _11222_/Y gnd _11223_/B vdd BUFX2
XBUFX2_insert321 _13345_/Y gnd _9865_/A vdd BUFX2
XFILL_0__12290_ gnd vdd FILL
XSFILL69160x14050 gnd vdd FILL
X_13505_ _9431_/Q gnd _13505_/Y vdd INVX1
X_10717_ _10717_/Q _9963_/CLK _9963_/R vdd _10717_/D gnd vdd DFFSR
XFILL_5__10242_ gnd vdd FILL
XFILL_5__13030_ gnd vdd FILL
XBUFX2_insert332 _12405_/Y gnd _9267_/B vdd BUFX2
X_14485_ _7989_/A gnd _14485_/Y vdd INVX1
XBUFX2_insert343 _12396_/Y gnd _9770_/B vdd BUFX2
XFILL_3__11421_ gnd vdd FILL
XBUFX2_insert354 _13306_/Y gnd _7948_/A vdd BUFX2
XFILL_1__12600_ gnd vdd FILL
XFILL_2__10062_ gnd vdd FILL
XFILL_4__10972_ gnd vdd FILL
XFILL_4__13760_ gnd vdd FILL
X_11697_ _11046_/Y _11676_/B _11696_/Y gnd _11697_/Y vdd OAI21X1
XBUFX2_insert365 _13487_/Y gnd _13592_/D vdd BUFX2
XFILL_5__8522_ gnd vdd FILL
XFILL_2__9793_ gnd vdd FILL
XFILL_0__11241_ gnd vdd FILL
XFILL_4__9729_ gnd vdd FILL
X_16224_ _10867_/Q gnd _16224_/Y vdd INVX1
XFILL_1__10792_ gnd vdd FILL
XFILL_1__13580_ gnd vdd FILL
XBUFX2_insert376 _12211_/Y gnd _12255_/C vdd BUFX2
XFILL_5_CLKBUF1_insert200 gnd vdd FILL
XFILL_5_CLKBUF1_insert211 gnd vdd FILL
XSFILL115080x5050 gnd vdd FILL
X_13436_ _14410_/A gnd _13865_/C vdd INVX8
XFILL_5__10173_ gnd vdd FILL
XFILL_4__12711_ gnd vdd FILL
X_10648_ _10700_/B _9624_/B gnd _10649_/C vdd NAND2X1
XFILL_3__14140_ gnd vdd FILL
XBUFX2_insert387 _13331_/Y gnd _9116_/B vdd BUFX2
XFILL_2__8744_ gnd vdd FILL
XBUFX2_insert398 _13293_/Y gnd _7562_/B vdd BUFX2
XFILL_5_CLKBUF1_insert222 gnd vdd FILL
XFILL_3__11352_ gnd vdd FILL
XFILL_4__13691_ gnd vdd FILL
XSFILL104360x23050 gnd vdd FILL
XFILL_2__14870_ gnd vdd FILL
XFILL_1__12531_ gnd vdd FILL
XSFILL104520x6050 gnd vdd FILL
XFILL_5__8453_ gnd vdd FILL
XFILL_0__11172_ gnd vdd FILL
XSFILL33640x55050 gnd vdd FILL
X_16155_ _15774_/C _14751_/Y _16155_/C _16155_/D gnd _16156_/B vdd OAI22X1
XFILL_3__10303_ gnd vdd FILL
X_13367_ _13371_/B _12807_/Q gnd _13465_/C vdd AND2X2
XFILL_4__15430_ gnd vdd FILL
XFILL_2__13821_ gnd vdd FILL
XFILL_4__12642_ gnd vdd FILL
XFILL_5__14981_ gnd vdd FILL
XFILL_3__14071_ gnd vdd FILL
X_10579_ _16305_/A gnd _10579_/Y vdd INVX1
XFILL_0__10123_ gnd vdd FILL
XFILL_1__15250_ gnd vdd FILL
XFILL_3__11283_ gnd vdd FILL
XFILL_1__12462_ gnd vdd FILL
X_15106_ _15801_/A _15106_/B _15801_/C _13510_/D gnd _15109_/B vdd OAI22X1
XFILL_0__15980_ gnd vdd FILL
XFILL_5__8384_ gnd vdd FILL
X_12318_ _12318_/A _12318_/B _12318_/C gnd _12318_/Y vdd NAND3X1
XFILL_3__13022_ gnd vdd FILL
XSFILL89320x27050 gnd vdd FILL
XFILL_5__13932_ gnd vdd FILL
X_16086_ _16086_/A _16086_/B gnd _16086_/Y vdd NOR2X1
X_13298_ _13215_/B _13326_/A _13259_/C gnd _13299_/A vdd OAI21X1
XFILL_0__7690_ gnd vdd FILL
XFILL_1__14201_ gnd vdd FILL
XFILL_4__12573_ gnd vdd FILL
XSFILL59080x66050 gnd vdd FILL
XFILL_4__15361_ gnd vdd FILL
XFILL_2__7626_ gnd vdd FILL
XFILL_3__10234_ gnd vdd FILL
XFILL_2__13752_ gnd vdd FILL
XFILL_1__11413_ gnd vdd FILL
XFILL_2__10964_ gnd vdd FILL
XFILL_1__15181_ gnd vdd FILL
XFILL_5__7335_ gnd vdd FILL
XFILL_1__12393_ gnd vdd FILL
XFILL_0__10054_ gnd vdd FILL
XFILL_0__14931_ gnd vdd FILL
X_15037_ _15031_/B _15014_/C _15037_/C gnd _15245_/B vdd OAI21X1
X_12249_ _6878_/A _12249_/B _12249_/C _12713_/A gnd _12250_/C vdd AOI22X1
XFILL_4__11524_ gnd vdd FILL
XFILL_4__14312_ gnd vdd FILL
XFILL_2__12703_ gnd vdd FILL
XFILL_5__13863_ gnd vdd FILL
XFILL_4__15292_ gnd vdd FILL
XFILL_3__10165_ gnd vdd FILL
XFILL_1__14132_ gnd vdd FILL
XFILL_2__7557_ gnd vdd FILL
XFILL_2__13683_ gnd vdd FILL
XFILL_1__11344_ gnd vdd FILL
XFILL_0__14862_ gnd vdd FILL
XFILL_2__10895_ gnd vdd FILL
XFILL_5__15602_ gnd vdd FILL
XFILL_0__9360_ gnd vdd FILL
XSFILL109080x35050 gnd vdd FILL
XFILL_4__14243_ gnd vdd FILL
XFILL_4__11455_ gnd vdd FILL
XFILL_2__15422_ gnd vdd FILL
XSFILL94440x18050 gnd vdd FILL
XFILL_2__12634_ gnd vdd FILL
XFILL_5__13794_ gnd vdd FILL
XFILL_5__9005_ gnd vdd FILL
XFILL_0__13813_ gnd vdd FILL
XFILL_2__7488_ gnd vdd FILL
XFILL_1__14063_ gnd vdd FILL
XFILL_3__14973_ gnd vdd FILL
XFILL_1__11275_ gnd vdd FILL
XFILL_0__8311_ gnd vdd FILL
XFILL_4__10406_ gnd vdd FILL
XSFILL13000x65050 gnd vdd FILL
XFILL_0__14793_ gnd vdd FILL
XFILL_5__15533_ gnd vdd FILL
XFILL_5__7197_ gnd vdd FILL
XFILL_5__12745_ gnd vdd FILL
XFILL_2__9227_ gnd vdd FILL
XFILL_4__14174_ gnd vdd FILL
XFILL_0__9291_ gnd vdd FILL
XFILL_3__8020_ gnd vdd FILL
XFILL_1__13014_ gnd vdd FILL
XFILL_2__15353_ gnd vdd FILL
XFILL_4__11386_ gnd vdd FILL
XFILL_3__13924_ gnd vdd FILL
XFILL_0__13744_ gnd vdd FILL
XSFILL94280x4050 gnd vdd FILL
XFILL_0__10956_ gnd vdd FILL
XFILL_4__13125_ gnd vdd FILL
XFILL_0__8242_ gnd vdd FILL
X_15939_ _14522_/A _15357_/B _16166_/A _10348_/Q gnd _15939_/Y vdd AOI22X1
XFILL_2__14304_ gnd vdd FILL
XFILL_5__15464_ gnd vdd FILL
X_8870_ _8870_/A gnd _8872_/A vdd INVX1
XFILL_2__11516_ gnd vdd FILL
XFILL_2__9158_ gnd vdd FILL
XFILL_3__13855_ gnd vdd FILL
XFILL_1__10157_ gnd vdd FILL
XFILL_2__15284_ gnd vdd FILL
XFILL_2__12496_ gnd vdd FILL
XFILL_0__13675_ gnd vdd FILL
XFILL_0__10887_ gnd vdd FILL
XFILL_5__14415_ gnd vdd FILL
X_7821_ _7819_/Y _7821_/B _7821_/C gnd _7821_/Y vdd OAI21X1
XFILL_2__8109_ gnd vdd FILL
XFILL_5__11627_ gnd vdd FILL
XFILL_6__13966_ gnd vdd FILL
XFILL_5__15395_ gnd vdd FILL
XFILL_2__14235_ gnd vdd FILL
XFILL_4__10268_ gnd vdd FILL
XFILL_2__9089_ gnd vdd FILL
XFILL_0__15414_ gnd vdd FILL
XFILL_3__13786_ gnd vdd FILL
XFILL_2__11447_ gnd vdd FILL
XFILL_0__12626_ gnd vdd FILL
XFILL_5__9907_ gnd vdd FILL
XFILL_1__14965_ gnd vdd FILL
XFILL_3__10998_ gnd vdd FILL
XFILL_6__15705_ gnd vdd FILL
XFILL_4__12007_ gnd vdd FILL
XFILL_0__7124_ gnd vdd FILL
XFILL_0__16394_ gnd vdd FILL
XFILL_5__14346_ gnd vdd FILL
XFILL_3__12737_ gnd vdd FILL
XFILL_3__15525_ gnd vdd FILL
XFILL_5__11558_ gnd vdd FILL
X_7752_ _7753_/B _7752_/B gnd _7753_/C vdd NAND2X1
XFILL_2__14166_ gnd vdd FILL
XFILL_1__13916_ gnd vdd FILL
XFILL_0__15345_ gnd vdd FILL
XFILL_2__11378_ gnd vdd FILL
XFILL_1__14896_ gnd vdd FILL
XFILL_0__7055_ gnd vdd FILL
XFILL_5__10509_ gnd vdd FILL
XFILL_2__13117_ gnd vdd FILL
XFILL_5__14277_ gnd vdd FILL
X_7683_ _7759_/B _9859_/B gnd _7684_/C vdd NAND2X1
XFILL_3__8853_ gnd vdd FILL
XFILL_5__11489_ gnd vdd FILL
XFILL_3__15456_ gnd vdd FILL
XFILL_1__13847_ gnd vdd FILL
XFILL_0__11508_ gnd vdd FILL
XFILL_2__14097_ gnd vdd FILL
XFILL_5__16016_ gnd vdd FILL
XFILL_0__12488_ gnd vdd FILL
XFILL_0__15276_ gnd vdd FILL
XFILL_5__13228_ gnd vdd FILL
X_9422_ _9356_/A _8526_/B gnd _9422_/Y vdd NAND2X1
XFILL_6__15567_ gnd vdd FILL
XFILL_5__9769_ gnd vdd FILL
XFILL_6__12779_ gnd vdd FILL
XFILL_3__14407_ gnd vdd FILL
XFILL_3__11619_ gnd vdd FILL
XFILL_3__15387_ gnd vdd FILL
XFILL_3__7804_ gnd vdd FILL
XFILL_4__13958_ gnd vdd FILL
XFILL_0__14227_ gnd vdd FILL
XFILL_3__12599_ gnd vdd FILL
XFILL_0__11439_ gnd vdd FILL
XFILL_3__8784_ gnd vdd FILL
XFILL_1__13778_ gnd vdd FILL
XFILL_6__14518_ gnd vdd FILL
X_9353_ _9420_/B _9353_/B gnd _9354_/C vdd NAND2X1
XFILL_5__13159_ gnd vdd FILL
XFILL_4__12909_ gnd vdd FILL
XFILL_3__14338_ gnd vdd FILL
XFILL_3__7735_ gnd vdd FILL
XFILL_1__15517_ gnd vdd FILL
XFILL_1__12729_ gnd vdd FILL
XFILL_4__13889_ gnd vdd FILL
XFILL_0__14158_ gnd vdd FILL
XSFILL8680x5050 gnd vdd FILL
X_8304_ _8304_/Q _8289_/CLK _7152_/R vdd _8304_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert406 gnd vdd FILL
XFILL_4__15628_ gnd vdd FILL
XFILL_0__7957_ gnd vdd FILL
X_9284_ _9284_/A gnd _9286_/A vdd INVX1
XFILL_4_BUFX2_insert417 gnd vdd FILL
XFILL_3__14269_ gnd vdd FILL
XFILL_4_BUFX2_insert428 gnd vdd FILL
XFILL_0__13109_ gnd vdd FILL
XFILL_1__15448_ gnd vdd FILL
XFILL_4_BUFX2_insert439 gnd vdd FILL
XFILL_2__14999_ gnd vdd FILL
XFILL_0__14089_ gnd vdd FILL
XFILL_0__6908_ gnd vdd FILL
XFILL_3__16008_ gnd vdd FILL
X_8235_ _8233_/Y _8237_/A _8235_/C gnd _8295_/D vdd OAI21X1
XFILL_3__9405_ gnd vdd FILL
XFILL_4__15559_ gnd vdd FILL
XFILL_0__7888_ gnd vdd FILL
XSFILL114520x68050 gnd vdd FILL
XFILL_1__15379_ gnd vdd FILL
XFILL_6__16119_ gnd vdd FILL
XFILL_3__7597_ gnd vdd FILL
XFILL_0__9627_ gnd vdd FILL
XFILL_0__6839_ gnd vdd FILL
XSFILL33800x15050 gnd vdd FILL
X_8166_ _8166_/Q _7282_/CLK _8166_/R vdd _8104_/Y gnd vdd DFFSR
XFILL_3__9336_ gnd vdd FILL
XSFILL115160x34050 gnd vdd FILL
X_7117_ _7155_/Q gnd _7117_/Y vdd INVX1
XFILL_1__8351_ gnd vdd FILL
X_8097_ _8098_/B _7713_/B gnd _8097_/Y vdd NAND2X1
XFILL_3__9267_ gnd vdd FILL
XFILL_4__8060_ gnd vdd FILL
XFILL_0__8509_ gnd vdd FILL
XFILL_1__7302_ gnd vdd FILL
X_7048_ _7048_/A gnd _7048_/Y vdd INVX1
XFILL_3__8218_ gnd vdd FILL
XFILL_0__9489_ gnd vdd FILL
XFILL111960x25050 gnd vdd FILL
XFILL_3_CLKBUF1_insert119 gnd vdd FILL
XFILL_1__7233_ gnd vdd FILL
XFILL_5_CLKBUF1_insert1079 gnd vdd FILL
XFILL_3__8149_ gnd vdd FILL
XFILL112040x34050 gnd vdd FILL
XFILL_1__7164_ gnd vdd FILL
XFILL_1_BUFX2_insert307 gnd vdd FILL
X_8999_ _8961_/B _7847_/B gnd _9000_/C vdd NAND2X1
XFILL_1_BUFX2_insert318 gnd vdd FILL
XFILL_4__8962_ gnd vdd FILL
XFILL_1_BUFX2_insert329 gnd vdd FILL
XFILL_1__7095_ gnd vdd FILL
XSFILL64200x81050 gnd vdd FILL
XFILL_4__8893_ gnd vdd FILL
X_11620_ _11366_/B _11620_/B _11614_/A _11778_/B gnd _11622_/B vdd OAI22X1
XSFILL114600x48050 gnd vdd FILL
XSFILL114520x1050 gnd vdd FILL
XFILL_4__7844_ gnd vdd FILL
X_11551_ _11551_/A _11116_/Y _11311_/Y gnd _11552_/A vdd OAI21X1
XSFILL69080x29050 gnd vdd FILL
X_10502_ _10539_/B _9094_/B gnd _10503_/C vdd NAND2X1
X_14270_ _8745_/A gnd _14270_/Y vdd INVX1
XFILL_1__9805_ gnd vdd FILL
XFILL_5_BUFX2_insert240 gnd vdd FILL
X_11482_ _11166_/Y _11223_/B gnd _11483_/C vdd NAND2X1
XFILL_5_BUFX2_insert251 gnd vdd FILL
XFILL_1__7997_ gnd vdd FILL
XFILL_5_BUFX2_insert262 gnd vdd FILL
XFILL_4__9514_ gnd vdd FILL
XFILL_5_BUFX2_insert273 gnd vdd FILL
X_13221_ _13305_/A _13266_/A gnd _13222_/B vdd NOR2X1
X_10433_ _16070_/A gnd _10435_/A vdd INVX1
XFILL_5_BUFX2_insert284 gnd vdd FILL
XFILL_5_BUFX2_insert295 gnd vdd FILL
XFILL_1__6948_ gnd vdd FILL
XFILL_1__9736_ gnd vdd FILL
X_13152_ _13153_/B _13152_/B gnd _13152_/Y vdd NAND2X1
XSFILL78520x6050 gnd vdd FILL
XSFILL23800x47050 gnd vdd FILL
XFILL_4_BUFX2_insert940 gnd vdd FILL
X_10364_ _10364_/A gnd _10364_/Y vdd INVX1
XFILL_2__8460_ gnd vdd FILL
XFILL_1__9667_ gnd vdd FILL
XFILL_4_BUFX2_insert951 gnd vdd FILL
XFILL_1__6879_ gnd vdd FILL
XFILL_4_BUFX2_insert962 gnd vdd FILL
X_12103_ _11999_/A _12430_/A _11999_/C gnd _12103_/Y vdd NAND3X1
XFILL_4__9376_ gnd vdd FILL
XFILL112120x14050 gnd vdd FILL
XFILL_4_BUFX2_insert973 gnd vdd FILL
X_13083_ _13155_/A _13083_/B gnd _13084_/C vdd NAND2X1
XFILL_1__8618_ gnd vdd FILL
XFILL_4_BUFX2_insert984 gnd vdd FILL
XFILL_4_BUFX2_insert995 gnd vdd FILL
X_10295_ _10295_/A _10294_/A _10295_/C gnd _10347_/D vdd OAI21X1
XFILL_1__9598_ gnd vdd FILL
XFILL_4__8327_ gnd vdd FILL
XFILL_5__7120_ gnd vdd FILL
XFILL_2__8391_ gnd vdd FILL
X_12034_ _12034_/A _12032_/Y _12033_/Y gnd _12034_/Y vdd NAND3X1
XFILL_6__10130_ gnd vdd FILL
XSFILL38840x7050 gnd vdd FILL
XFILL_2__7342_ gnd vdd FILL
XFILL_5__7051_ gnd vdd FILL
XFILL_2__10680_ gnd vdd FILL
XFILL_4__8258_ gnd vdd FILL
XFILL_4__11240_ gnd vdd FILL
XFILL_5__10791_ gnd vdd FILL
XFILL_3__11970_ gnd vdd FILL
XFILL_1__11060_ gnd vdd FILL
XFILL_4__7209_ gnd vdd FILL
XFILL_0__10810_ gnd vdd FILL
XFILL_4__8189_ gnd vdd FILL
XFILL_0__11790_ gnd vdd FILL
XFILL_5__12530_ gnd vdd FILL
XFILL_2__9012_ gnd vdd FILL
XFILL_3__10921_ gnd vdd FILL
X_13985_ _13985_/A _13879_/B _14456_/C _13985_/D gnd _13986_/A vdd OAI22X1
XFILL_1__10011_ gnd vdd FILL
XFILL_4__11171_ gnd vdd FILL
XFILL_2__12350_ gnd vdd FILL
XSFILL84200x12050 gnd vdd FILL
XFILL_4__10122_ gnd vdd FILL
X_15724_ _15724_/A _15972_/B _15899_/A _15724_/D gnd _15724_/Y vdd OAI22X1
X_12936_ _12936_/Q _8176_/CLK _7408_/R vdd _12876_/Y gnd vdd DFFSR
XSFILL28920x80050 gnd vdd FILL
XFILL_3__13640_ gnd vdd FILL
XFILL_5__12461_ gnd vdd FILL
XFILL_2__11301_ gnd vdd FILL
XSFILL104360x18050 gnd vdd FILL
XFILL_0__13460_ gnd vdd FILL
XFILL_2__12281_ gnd vdd FILL
XFILL_5__14200_ gnd vdd FILL
XFILL_0__10672_ gnd vdd FILL
XFILL_6__13751_ gnd vdd FILL
XFILL_5__7953_ gnd vdd FILL
XFILL_5__11412_ gnd vdd FILL
XFILL_5__15180_ gnd vdd FILL
X_15655_ _9379_/A gnd _15656_/A vdd INVX1
XFILL_2__14020_ gnd vdd FILL
X_12867_ _12865_/Y vdd _12867_/C gnd _12933_/D vdd OAI21X1
XFILL_4__14930_ gnd vdd FILL
XFILL_4__10053_ gnd vdd FILL
XFILL_1_BUFX2_insert830 gnd vdd FILL
XFILL_5__12392_ gnd vdd FILL
XFILL_3__13571_ gnd vdd FILL
XFILL_1_BUFX2_insert841 gnd vdd FILL
XFILL_2__11232_ gnd vdd FILL
XFILL_0__12411_ gnd vdd FILL
XFILL_1__14750_ gnd vdd FILL
XFILL_3__10783_ gnd vdd FILL
XFILL_1_BUFX2_insert852 gnd vdd FILL
XFILL_6__12702_ gnd vdd FILL
XFILL_0__13391_ gnd vdd FILL
XFILL_5__6904_ gnd vdd FILL
XFILL_1__11962_ gnd vdd FILL
X_14606_ _7150_/Q _13592_/D _13853_/C _6974_/A gnd _14607_/B vdd AOI22X1
XFILL_5__14131_ gnd vdd FILL
XFILL_1_BUFX2_insert863 gnd vdd FILL
X_11818_ _11005_/Y _11816_/Y _11818_/C gnd _11818_/Y vdd OAI21X1
XFILL_5__7884_ gnd vdd FILL
XFILL_3__15310_ gnd vdd FILL
XFILL_1_BUFX2_insert874 gnd vdd FILL
XFILL_3__12522_ gnd vdd FILL
X_15586_ _15586_/A _15586_/B gnd _15610_/A vdd NOR2X1
XFILL_5__11343_ gnd vdd FILL
XFILL_4__14861_ gnd vdd FILL
X_12798_ _12716_/A _7005_/CLK _12799_/R vdd _12798_/D gnd vdd DFFSR
XFILL_2__9914_ gnd vdd FILL
XFILL_3__16290_ gnd vdd FILL
XFILL_6__10894_ gnd vdd FILL
XFILL_1_BUFX2_insert885 gnd vdd FILL
XFILL_1__13701_ gnd vdd FILL
XFILL_1__10913_ gnd vdd FILL
XFILL_0__12342_ gnd vdd FILL
XFILL_2__11163_ gnd vdd FILL
XFILL_0__15130_ gnd vdd FILL
XFILL_5__9623_ gnd vdd FILL
XFILL_1_BUFX2_insert896 gnd vdd FILL
XFILL_1__14681_ gnd vdd FILL
XSFILL64040x2050 gnd vdd FILL
XSFILL99480x66050 gnd vdd FILL
XFILL_1__11893_ gnd vdd FILL
X_14537_ _14528_/Y _14529_/Y _14537_/C gnd _14537_/Y vdd NAND3X1
XSFILL74120x64050 gnd vdd FILL
XFILL_4__13812_ gnd vdd FILL
XFILL_3__15241_ gnd vdd FILL
XFILL_5__14062_ gnd vdd FILL
XFILL_5__11274_ gnd vdd FILL
X_11749_ _11745_/Y _11748_/Y _11749_/C gnd _11752_/C vdd AOI21X1
XFILL_2__10114_ gnd vdd FILL
XFILL_3__12453_ gnd vdd FILL
XFILL_1__13632_ gnd vdd FILL
XFILL_4__14792_ gnd vdd FILL
XFILL_2__15971_ gnd vdd FILL
XFILL_0__15061_ gnd vdd FILL
XFILL_0__12273_ gnd vdd FILL
XFILL_2__11094_ gnd vdd FILL
XFILL_6__15352_ gnd vdd FILL
XFILL_5__9554_ gnd vdd FILL
XFILL_5__13013_ gnd vdd FILL
X_14468_ _7531_/Q gnd _14468_/Y vdd INVX1
XFILL_0__8860_ gnd vdd FILL
XFILL_3__11404_ gnd vdd FILL
XFILL_4__13743_ gnd vdd FILL
XFILL_3__15172_ gnd vdd FILL
XFILL_4__10955_ gnd vdd FILL
XFILL_2__10045_ gnd vdd FILL
XFILL_0__14012_ gnd vdd FILL
XFILL_3__12384_ gnd vdd FILL
XFILL_1__16351_ gnd vdd FILL
XFILL_0__11224_ gnd vdd FILL
XFILL_2__14922_ gnd vdd FILL
XFILL_2__6988_ gnd vdd FILL
XFILL_5__8505_ gnd vdd FILL
XFILL_2__9776_ gnd vdd FILL
XFILL_6__14303_ gnd vdd FILL
XFILL_1__13563_ gnd vdd FILL
XFILL_0__7811_ gnd vdd FILL
X_16207_ _8819_/Q gnd _16207_/Y vdd INVX1
X_13419_ _13377_/Y _13407_/Y gnd _13419_/Y vdd NAND2X1
XFILL_1__10775_ gnd vdd FILL
XSFILL53960x22050 gnd vdd FILL
XFILL_5__9485_ gnd vdd FILL
XFILL_3__14123_ gnd vdd FILL
XFILL_5__10156_ gnd vdd FILL
XFILL_1__15302_ gnd vdd FILL
XFILL_6__12495_ gnd vdd FILL
X_14399_ _8367_/A _13647_/B _13864_/B _8681_/Q gnd _14399_/Y vdd AOI22X1
XFILL_3__11335_ gnd vdd FILL
XFILL_2__14853_ gnd vdd FILL
XFILL_2__8727_ gnd vdd FILL
XFILL_4__13674_ gnd vdd FILL
XSFILL109480x51050 gnd vdd FILL
XFILL_1__12514_ gnd vdd FILL
XFILL_4__10886_ gnd vdd FILL
XFILL_0__11155_ gnd vdd FILL
XSFILL64520x8050 gnd vdd FILL
XFILL_1__16282_ gnd vdd FILL
XFILL_1__13494_ gnd vdd FILL
X_16138_ _16137_/Y _16138_/B gnd _16139_/C vdd NOR2X1
XFILL_0__7742_ gnd vdd FILL
XFILL_4__15413_ gnd vdd FILL
XSFILL13800x4050 gnd vdd FILL
XFILL_6__11446_ gnd vdd FILL
XFILL_4__12625_ gnd vdd FILL
XFILL_2__13804_ gnd vdd FILL
XFILL_3__14054_ gnd vdd FILL
XFILL_5__14964_ gnd vdd FILL
XFILL_4__16393_ gnd vdd FILL
XFILL_1__15233_ gnd vdd FILL
XFILL_3__7451_ gnd vdd FILL
XFILL_0__10106_ gnd vdd FILL
XFILL_3__11266_ gnd vdd FILL
XFILL_2__8658_ gnd vdd FILL
XFILL_1__12445_ gnd vdd FILL
XFILL_2__14784_ gnd vdd FILL
XFILL_2__11996_ gnd vdd FILL
XFILL_0__15963_ gnd vdd FILL
XFILL_5__8367_ gnd vdd FILL
XFILL_0__11086_ gnd vdd FILL
XFILL_6__14165_ gnd vdd FILL
X_8020_ _7997_/B _7508_/B gnd _8021_/C vdd NAND2X1
XFILL_3__13005_ gnd vdd FILL
X_16069_ _15524_/A _14662_/D _16069_/C _15521_/C gnd _16069_/Y vdd OAI22X1
XFILL_5__13915_ gnd vdd FILL
XFILL_2__7609_ gnd vdd FILL
XFILL_4__15344_ gnd vdd FILL
XFILL_0__7673_ gnd vdd FILL
XFILL_2__13735_ gnd vdd FILL
XFILL_5__14895_ gnd vdd FILL
XFILL_2__10947_ gnd vdd FILL
XFILL_2__8589_ gnd vdd FILL
XFILL_0__10037_ gnd vdd FILL
XFILL_1__15164_ gnd vdd FILL
XFILL_5__7318_ gnd vdd FILL
XFILL_3__11197_ gnd vdd FILL
XFILL_0__14914_ gnd vdd FILL
XFILL_0__9412_ gnd vdd FILL
XFILL_1__12376_ gnd vdd FILL
XSFILL115080x49050 gnd vdd FILL
XFILL_0__15894_ gnd vdd FILL
XFILL_5__13846_ gnd vdd FILL
XFILL_3__9121_ gnd vdd FILL
XFILL_4__11507_ gnd vdd FILL
XSFILL43880x74050 gnd vdd FILL
XFILL_3__10148_ gnd vdd FILL
XFILL_4__12487_ gnd vdd FILL
XFILL_1__14115_ gnd vdd FILL
XFILL_4__15275_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1074 gnd vdd FILL
XFILL_2__13666_ gnd vdd FILL
XFILL_1__11327_ gnd vdd FILL
XFILL_0__14845_ gnd vdd FILL
XFILL_2__10878_ gnd vdd FILL
XFILL_5__7249_ gnd vdd FILL
XFILL_1__15095_ gnd vdd FILL
XFILL_0__9343_ gnd vdd FILL
XFILL_2__15405_ gnd vdd FILL
XFILL_4__14226_ gnd vdd FILL
XFILL_6__10259_ gnd vdd FILL
XFILL_4__11438_ gnd vdd FILL
XFILL_2__12617_ gnd vdd FILL
X_9971_ _9933_/A _9963_/CLK _7789_/R vdd _9971_/D gnd vdd DFFSR
XFILL_5__13777_ gnd vdd FILL
XSFILL18680x50050 gnd vdd FILL
XSFILL48920x11050 gnd vdd FILL
XFILL_2__16385_ gnd vdd FILL
XFILL_1__14046_ gnd vdd FILL
XFILL_5__10989_ gnd vdd FILL
XFILL_3__14956_ gnd vdd FILL
XFILL_2__13597_ gnd vdd FILL
XSFILL74200x44050 gnd vdd FILL
XFILL_1__11258_ gnd vdd FILL
XFILL_5__15516_ gnd vdd FILL
XFILL_0__14776_ gnd vdd FILL
XFILL_5__12728_ gnd vdd FILL
X_8922_ _8834_/A _7389_/CLK _8285_/R vdd _8922_/D gnd vdd DFFSR
XFILL_0__9274_ gnd vdd FILL
XFILL_0__11988_ gnd vdd FILL
XFILL_3__8003_ gnd vdd FILL
XFILL_2__15336_ gnd vdd FILL
XFILL_4__14157_ gnd vdd FILL
XFILL_3__13907_ gnd vdd FILL
XFILL_4__11369_ gnd vdd FILL
XFILL_1__11189_ gnd vdd FILL
XFILL_0__13727_ gnd vdd FILL
XFILL_3__14887_ gnd vdd FILL
XFILL_0__10939_ gnd vdd FILL
XFILL_0__8225_ gnd vdd FILL
XFILL_4__13108_ gnd vdd FILL
XFILL_5__15447_ gnd vdd FILL
XFILL_5__12659_ gnd vdd FILL
XSFILL108920x65050 gnd vdd FILL
X_8853_ _8854_/B _8853_/B gnd _8853_/Y vdd NAND2X1
XFILL_4__14088_ gnd vdd FILL
XFILL_3__13838_ gnd vdd FILL
XFILL_2__15267_ gnd vdd FILL
XFILL_2__12479_ gnd vdd FILL
XFILL_1__15997_ gnd vdd FILL
XFILL_0__13658_ gnd vdd FILL
XFILL_4__13039_ gnd vdd FILL
X_7804_ _7804_/A gnd _7804_/Y vdd INVX1
XFILL_2__14218_ gnd vdd FILL
XFILL_5__15378_ gnd vdd FILL
X_8784_ _8820_/Q gnd _8786_/A vdd INVX1
XFILL_2__15198_ gnd vdd FILL
XSFILL38840x63050 gnd vdd FILL
XFILL_0__12609_ gnd vdd FILL
XFILL_3__13769_ gnd vdd FILL
XFILL_1__14948_ gnd vdd FILL
XFILL_0__16377_ gnd vdd FILL
XFILL_0__7107_ gnd vdd FILL
XFILL_6__9663_ gnd vdd FILL
XFILL_0__13589_ gnd vdd FILL
XFILL112360x70050 gnd vdd FILL
XSFILL54120x11050 gnd vdd FILL
XFILL_5__14329_ gnd vdd FILL
X_7735_ _7735_/A _7759_/B _7734_/Y gnd _7735_/Y vdd OAI21X1
XFILL_0__8087_ gnd vdd FILL
XFILL_3__15508_ gnd vdd FILL
XFILL_2__14149_ gnd vdd FILL
XFILL_3__8905_ gnd vdd FILL
XFILL_0__15328_ gnd vdd FILL
XFILL_6__8614_ gnd vdd FILL
XFILL_1__14879_ gnd vdd FILL
XFILL_3__9885_ gnd vdd FILL
XFILL_0__7038_ gnd vdd FILL
X_7666_ _7626_/A _8562_/CLK _9430_/R vdd _7666_/D gnd vdd DFFSR
XFILL_3__15439_ gnd vdd FILL
XFILL_3__8836_ gnd vdd FILL
XFILL_5_BUFX2_insert90 gnd vdd FILL
XFILL_0__15259_ gnd vdd FILL
XSFILL114120x65050 gnd vdd FILL
X_9405_ _9403_/Y _9356_/A _9405_/C gnd _9405_/Y vdd OAI21X1
XFILL_1__7851_ gnd vdd FILL
XFILL_4__7560_ gnd vdd FILL
X_7597_ _7598_/B _9005_/B gnd _7598_/C vdd NAND2X1
XFILL_3__8767_ gnd vdd FILL
XSFILL58200x57050 gnd vdd FILL
XSFILL18760x30050 gnd vdd FILL
X_9336_ _9336_/A _9420_/B _9335_/Y gnd _9430_/D vdd OAI21X1
XSFILL8600x40050 gnd vdd FILL
XFILL_0__8989_ gnd vdd FILL
XFILL_3__7718_ gnd vdd FILL
XSFILL44040x63050 gnd vdd FILL
XSFILL99560x6050 gnd vdd FILL
XFILL_4_BUFX2_insert225 gnd vdd FILL
XFILL_4__7491_ gnd vdd FILL
XFILL_3__8698_ gnd vdd FILL
XFILL_1__9521_ gnd vdd FILL
XSFILL48840x2050 gnd vdd FILL
XFILL_4_BUFX2_insert236 gnd vdd FILL
XFILL_4__9230_ gnd vdd FILL
XFILL_4_BUFX2_insert247 gnd vdd FILL
X_9267_ _9240_/A _9267_/B gnd _9267_/Y vdd NAND2X1
XFILL_4_BUFX2_insert258 gnd vdd FILL
XFILL_4_BUFX2_insert269 gnd vdd FILL
XFILL_6__7358_ gnd vdd FILL
X_8218_ _8290_/Q gnd _8218_/Y vdd INVX1
XSFILL23880x21050 gnd vdd FILL
XFILL_3_BUFX2_insert903 gnd vdd FILL
X_9198_ _9198_/Q _8046_/CLK _9692_/R vdd _9198_/D gnd vdd DFFSR
XFILL_4__9161_ gnd vdd FILL
XFILL_3_BUFX2_insert914 gnd vdd FILL
XFILL_1__8403_ gnd vdd FILL
XFILL_3_BUFX2_insert925 gnd vdd FILL
XFILL_3_BUFX2_insert936 gnd vdd FILL
X_10080_ _15475_/A _7530_/CLK _7523_/R vdd _10080_/D gnd vdd DFFSR
XFILL_1__9383_ gnd vdd FILL
XFILL_3_BUFX2_insert947 gnd vdd FILL
X_8149_ _8149_/A _8098_/B _8149_/C gnd _8149_/Y vdd OAI21X1
XFILL_4__8112_ gnd vdd FILL
XFILL_4__9092_ gnd vdd FILL
XFILL112440x50050 gnd vdd FILL
XFILL_3_BUFX2_insert958 gnd vdd FILL
XFILL_3_BUFX2_insert969 gnd vdd FILL
XSFILL64200x76050 gnd vdd FILL
XFILL_1__8334_ gnd vdd FILL
XSFILL99000x8050 gnd vdd FILL
XSFILL39000x52050 gnd vdd FILL
XFILL_1__8265_ gnd vdd FILL
XSFILL3640x83050 gnd vdd FILL
XSFILL68840x79050 gnd vdd FILL
X_13770_ _13865_/C _7688_/A _7560_/A _14185_/B gnd _13772_/A vdd AOI22X1
XFILL_1__7216_ gnd vdd FILL
XFILL_3_BUFX2_insert1008 gnd vdd FILL
X_10982_ vdd _10971_/Y gnd _10982_/Y vdd NAND2X1
XFILL_3_BUFX2_insert1019 gnd vdd FILL
XFILL_1__8196_ gnd vdd FILL
XFILL_1_BUFX2_insert104 gnd vdd FILL
XSFILL18840x10050 gnd vdd FILL
X_12721_ _12721_/A _12721_/B _12721_/C gnd _12799_/D vdd OAI21X1
XSFILL94280x71050 gnd vdd FILL
XFILL_4__9994_ gnd vdd FILL
XSFILL68440x81050 gnd vdd FILL
X_15440_ _15440_/A _15440_/B _15437_/Y gnd _15440_/Y vdd NAND3X1
X_12652_ vdd memoryOutData[28] gnd _12652_/Y vdd NAND2X1
XFILL_1__7078_ gnd vdd FILL
XFILL_2__7960_ gnd vdd FILL
X_11603_ _11571_/A _11587_/Y gnd _11604_/C vdd NAND2X1
XFILL_0_BUFX2_insert804 gnd vdd FILL
X_15371_ _15371_/A _15370_/Y _15371_/C gnd _15371_/Y vdd NAND3X1
XFILL_0_BUFX2_insert815 gnd vdd FILL
XFILL_4__8876_ gnd vdd FILL
XFILL_2__6911_ gnd vdd FILL
X_12583_ vdd memoryOutData[5] gnd _12584_/C vdd NAND2X1
XFILL_0_BUFX2_insert826 gnd vdd FILL
XFILL_0_BUFX2_insert837 gnd vdd FILL
XFILL_1_BUFX2_insert1001 gnd vdd FILL
XFILL_2__7891_ gnd vdd FILL
XFILL_1_BUFX2_insert1012 gnd vdd FILL
X_14322_ _14322_/A _14322_/B _14321_/Y gnd _14333_/A vdd NAND3X1
XFILL_4__7827_ gnd vdd FILL
XFILL_0_BUFX2_insert848 gnd vdd FILL
XFILL_0_BUFX2_insert859 gnd vdd FILL
X_11534_ _11534_/A _11312_/Y _11542_/A gnd _11534_/Y vdd OAI21X1
XFILL_1_BUFX2_insert1023 gnd vdd FILL
XFILL_1_BUFX2_insert1034 gnd vdd FILL
XFILL_2__6842_ gnd vdd FILL
XFILL_2__9630_ gnd vdd FILL
XFILL_1_BUFX2_insert1045 gnd vdd FILL
XFILL_5__10010_ gnd vdd FILL
XFILL_1_BUFX2_insert1056 gnd vdd FILL
XFILL_4__7758_ gnd vdd FILL
XSFILL49640x74050 gnd vdd FILL
X_14253_ _14253_/A _14253_/B _14250_/Y gnd _14253_/Y vdd NAND3X1
XFILL_1_BUFX2_insert1067 gnd vdd FILL
XFILL_3_BUFX2_insert19 gnd vdd FILL
X_11465_ _11464_/Y _11194_/Y _11320_/Y gnd _11465_/Y vdd OAI21X1
XFILL_1_BUFX2_insert1089 gnd vdd FILL
XSFILL89240x60050 gnd vdd FILL
XSFILL53880x37050 gnd vdd FILL
XFILL_1__10560_ gnd vdd FILL
XFILL_5__9270_ gnd vdd FILL
X_13204_ _11974_/A _12538_/CLK _12795_/R vdd _13204_/D gnd vdd DFFSR
XFILL_4__7689_ gnd vdd FILL
X_10416_ _10426_/B _7856_/B gnd _10417_/C vdd NAND2X1
XFILL_2__8512_ gnd vdd FILL
X_14184_ _14184_/A _14640_/C gnd _14184_/Y vdd NOR2X1
XFILL_6__12280_ gnd vdd FILL
XFILL_3__11120_ gnd vdd FILL
XSFILL13880x53050 gnd vdd FILL
XFILL_1__9719_ gnd vdd FILL
XFILL_4__10671_ gnd vdd FILL
X_11396_ _11055_/B _11392_/Y _11395_/Y gnd _11401_/B vdd AOI21X1
XFILL_2__9492_ gnd vdd FILL
XFILL_5__8221_ gnd vdd FILL
XFILL_2__11850_ gnd vdd FILL
XFILL_4__9428_ gnd vdd FILL
XFILL_1__10491_ gnd vdd FILL
X_13135_ _13135_/A _13134_/A _13135_/C gnd _13193_/D vdd OAI21X1
XFILL_6__11231_ gnd vdd FILL
XFILL_4__12410_ gnd vdd FILL
X_10347_ _10293_/A _7147_/CLK _7531_/R vdd _10347_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert770 gnd vdd FILL
XFILL_5__11961_ gnd vdd FILL
XFILL_4__13390_ gnd vdd FILL
XFILL_2__10801_ gnd vdd FILL
XFILL_3__11051_ gnd vdd FILL
XFILL_2__8443_ gnd vdd FILL
XFILL_3_CLKBUF1_insert1080 gnd vdd FILL
XSFILL28920x75050 gnd vdd FILL
XFILL_1__12230_ gnd vdd FILL
XFILL_4_BUFX2_insert781 gnd vdd FILL
XSFILL94360x51050 gnd vdd FILL
XFILL_4_BUFX2_insert792 gnd vdd FILL
XFILL_6_CLKBUF1_insert147 gnd vdd FILL
XFILL_2__11781_ gnd vdd FILL
XFILL_4__9359_ gnd vdd FILL
XFILL_0__12960_ gnd vdd FILL
XFILL_5__13700_ gnd vdd FILL
XFILL_5__10912_ gnd vdd FILL
XFILL_4__12341_ gnd vdd FILL
X_13066_ _6889_/A _8169_/CLK _7408_/R vdd _13066_/D gnd vdd DFFSR
XFILL_3__10002_ gnd vdd FILL
X_10278_ _14221_/A gnd _10280_/A vdd INVX1
XFILL_5__14680_ gnd vdd FILL
XFILL_2__13520_ gnd vdd FILL
XFILL_2__8374_ gnd vdd FILL
XFILL_5__7103_ gnd vdd FILL
XFILL_5__11892_ gnd vdd FILL
XFILL_0__11911_ gnd vdd FILL
XFILL_1__12161_ gnd vdd FILL
X_12017_ _12461_/B _12073_/B _12073_/C gnd gnd _12017_/Y vdd AOI22X1
XFILL_5__8083_ gnd vdd FILL
XFILL_5__13631_ gnd vdd FILL
XFILL_0__12891_ gnd vdd FILL
XFILL_3__14810_ gnd vdd FILL
XFILL_4__15060_ gnd vdd FILL
XFILL_4__12272_ gnd vdd FILL
XFILL_6__11093_ gnd vdd FILL
XFILL_2__7325_ gnd vdd FILL
XFILL_2__13451_ gnd vdd FILL
XFILL_1__11112_ gnd vdd FILL
XFILL_0__14630_ gnd vdd FILL
XFILL_2__10663_ gnd vdd FILL
XFILL_1__12092_ gnd vdd FILL
XFILL_3__15790_ gnd vdd FILL
XFILL_5__7034_ gnd vdd FILL
XFILL_0__11842_ gnd vdd FILL
XFILL_4__14011_ gnd vdd FILL
XFILL_5__16350_ gnd vdd FILL
XFILL_4__11223_ gnd vdd FILL
XFILL_2__12402_ gnd vdd FILL
XFILL_5__13562_ gnd vdd FILL
XFILL_1__15920_ gnd vdd FILL
XSFILL74120x59050 gnd vdd FILL
XFILL_2__16170_ gnd vdd FILL
XFILL_3__11953_ gnd vdd FILL
XFILL_3__14741_ gnd vdd FILL
XFILL_1__11043_ gnd vdd FILL
XFILL_5__10774_ gnd vdd FILL
XFILL_2__13382_ gnd vdd FILL
XFILL_0__14561_ gnd vdd FILL
XFILL_5__15301_ gnd vdd FILL
XFILL_5__12513_ gnd vdd FILL
XFILL_0__11773_ gnd vdd FILL
XFILL_3__10904_ gnd vdd FILL
XFILL_4__11154_ gnd vdd FILL
XFILL_2__15121_ gnd vdd FILL
XFILL_5__16281_ gnd vdd FILL
XFILL_0__16300_ gnd vdd FILL
XFILL_2__12333_ gnd vdd FILL
XFILL_5__13493_ gnd vdd FILL
X_13968_ _9696_/Q gnd _15464_/C vdd INVX1
XFILL_3__11884_ gnd vdd FILL
XFILL_1__15851_ gnd vdd FILL
XFILL_2__7187_ gnd vdd FILL
XFILL_3__14672_ gnd vdd FILL
XFILL_0__13512_ gnd vdd FILL
XFILL_0__8010_ gnd vdd FILL
XFILL_0__14492_ gnd vdd FILL
XFILL_5__15232_ gnd vdd FILL
X_15707_ _14262_/A gnd _15708_/B vdd INVX1
XSFILL89320x40050 gnd vdd FILL
XFILL_4__10105_ gnd vdd FILL
XFILL_5__8985_ gnd vdd FILL
X_12919_ _12823_/A _8560_/CLK _8033_/R vdd _12919_/D gnd vdd DFFSR
XFILL_5__12444_ gnd vdd FILL
XFILL_3__16411_ gnd vdd FILL
XSFILL53960x17050 gnd vdd FILL
XFILL_3__13623_ gnd vdd FILL
XFILL_1__14802_ gnd vdd FILL
XFILL_4__15962_ gnd vdd FILL
XFILL_2__15052_ gnd vdd FILL
XFILL_4__11085_ gnd vdd FILL
X_13899_ _14712_/B _9745_/A _9105_/A _14868_/D gnd _13907_/B vdd AOI22X1
XFILL_3__10835_ gnd vdd FILL
XFILL_0__16231_ gnd vdd FILL
XSFILL109480x46050 gnd vdd FILL
XFILL_2__12264_ gnd vdd FILL
XFILL_0__13443_ gnd vdd FILL
XFILL_1__15782_ gnd vdd FILL
XFILL_0__10655_ gnd vdd FILL
XFILL_5__7936_ gnd vdd FILL
XFILL_1__12994_ gnd vdd FILL
XFILL_6__10946_ gnd vdd FILL
X_15638_ _10596_/Q gnd _15639_/B vdd INVX1
XFILL_1_BUFX2_insert660 gnd vdd FILL
XFILL_2__14003_ gnd vdd FILL
XFILL_4__10036_ gnd vdd FILL
XFILL_5__15163_ gnd vdd FILL
XFILL_4__14913_ gnd vdd FILL
XFILL_3__16342_ gnd vdd FILL
XFILL_5__12375_ gnd vdd FILL
XFILL_3__13554_ gnd vdd FILL
XFILL_2__11215_ gnd vdd FILL
XFILL_3__6951_ gnd vdd FILL
XFILL_3__10766_ gnd vdd FILL
XFILL_4__15893_ gnd vdd FILL
XFILL_1_BUFX2_insert671 gnd vdd FILL
XFILL_1__14733_ gnd vdd FILL
XFILL_1__11945_ gnd vdd FILL
XFILL_2__12195_ gnd vdd FILL
XFILL_1_BUFX2_insert682 gnd vdd FILL
XFILL_0__16162_ gnd vdd FILL
XFILL_0__13374_ gnd vdd FILL
XFILL_1_BUFX2_insert693 gnd vdd FILL
XFILL_5__14114_ gnd vdd FILL
XFILL_5__7867_ gnd vdd FILL
XFILL_3__12505_ gnd vdd FILL
XFILL_5__11326_ gnd vdd FILL
X_7520_ _7520_/Q _9716_/CLK _8682_/R vdd _7520_/D gnd vdd DFFSR
XFILL_4__14844_ gnd vdd FILL
X_15569_ _15681_/B _14044_/Y _15569_/C _14067_/Y gnd _15569_/Y vdd OAI22X1
XFILL_5__15094_ gnd vdd FILL
XFILL_2__11146_ gnd vdd FILL
XFILL_3__13485_ gnd vdd FILL
XFILL_0__15113_ gnd vdd FILL
XFILL_3__16273_ gnd vdd FILL
XFILL_3__9670_ gnd vdd FILL
XFILL_3__6882_ gnd vdd FILL
XFILL_5__9606_ gnd vdd FILL
XFILL_1__14664_ gnd vdd FILL
XFILL_3__10697_ gnd vdd FILL
XFILL_0__12325_ gnd vdd FILL
XFILL_1__11876_ gnd vdd FILL
XFILL_0__16093_ gnd vdd FILL
XFILL_5__14045_ gnd vdd FILL
XFILL_0__8912_ gnd vdd FILL
XFILL_0__9892_ gnd vdd FILL
XFILL_5__7798_ gnd vdd FILL
XFILL_3__12436_ gnd vdd FILL
X_7451_ _7416_/B _7451_/B gnd _7452_/C vdd NAND2X1
XFILL_3__15224_ gnd vdd FILL
XFILL_1__16403_ gnd vdd FILL
XFILL_5__11257_ gnd vdd FILL
XFILL_1__13615_ gnd vdd FILL
XSFILL43880x69050 gnd vdd FILL
XFILL_3__8621_ gnd vdd FILL
XFILL_4__14775_ gnd vdd FILL
XFILL_1__10827_ gnd vdd FILL
XFILL_4__11987_ gnd vdd FILL
XFILL_0__15044_ gnd vdd FILL
XFILL_2__15954_ gnd vdd FILL
XFILL_0__12256_ gnd vdd FILL
XFILL_2__11077_ gnd vdd FILL
XFILL_1__14595_ gnd vdd FILL
XFILL_6__8330_ gnd vdd FILL
XFILL_5__9537_ gnd vdd FILL
XFILL_0__8843_ gnd vdd FILL
XSFILL74040x50 gnd vdd FILL
XFILL_3__15155_ gnd vdd FILL
XFILL_5__11188_ gnd vdd FILL
XFILL_4__13726_ gnd vdd FILL
XFILL_4__10938_ gnd vdd FILL
XFILL_3__12367_ gnd vdd FILL
XFILL_1__16334_ gnd vdd FILL
X_7382_ _7286_/A _7382_/CLK _8674_/R vdd _7382_/D gnd vdd DFFSR
XFILL_2__10028_ gnd vdd FILL
XFILL_2__14905_ gnd vdd FILL
XSFILL18680x45050 gnd vdd FILL
XFILL_1__13546_ gnd vdd FILL
XFILL_2__9759_ gnd vdd FILL
XFILL_0__11207_ gnd vdd FILL
XFILL_0__12187_ gnd vdd FILL
XSFILL8520x55050 gnd vdd FILL
XFILL_1__10758_ gnd vdd FILL
XFILL_2__15885_ gnd vdd FILL
X_9121_ _9164_/B _9633_/B gnd _9121_/Y vdd NAND2X1
XFILL_5__9468_ gnd vdd FILL
XFILL_3__7503_ gnd vdd FILL
XFILL_0__8774_ gnd vdd FILL
XFILL_3__11318_ gnd vdd FILL
XFILL_5__10139_ gnd vdd FILL
XFILL_3__14106_ gnd vdd FILL
XFILL_5__15996_ gnd vdd FILL
XFILL_4__13657_ gnd vdd FILL
XFILL_3__15086_ gnd vdd FILL
XSFILL84360x83050 gnd vdd FILL
XFILL_2__14836_ gnd vdd FILL
XFILL_3__8483_ gnd vdd FILL
XFILL_0__11138_ gnd vdd FILL
XFILL_1__16265_ gnd vdd FILL
XFILL_3__12298_ gnd vdd FILL
XFILL_1__13477_ gnd vdd FILL
XSFILL99160x43050 gnd vdd FILL
XFILL_0__7725_ gnd vdd FILL
XFILL_1__10689_ gnd vdd FILL
XSFILL49000x15050 gnd vdd FILL
XFILL_5__9399_ gnd vdd FILL
XFILL_4__12608_ gnd vdd FILL
X_9052_ _8968_/A _7662_/CLK _9454_/R vdd _9052_/D gnd vdd DFFSR
XFILL_3__14037_ gnd vdd FILL
XFILL_5__14947_ gnd vdd FILL
XFILL_3__7434_ gnd vdd FILL
XFILL_1__15216_ gnd vdd FILL
XFILL_4__16376_ gnd vdd FILL
XFILL_3__11249_ gnd vdd FILL
XFILL_4__13588_ gnd vdd FILL
XFILL_1__12428_ gnd vdd FILL
XFILL_2__14767_ gnd vdd FILL
XFILL_1__16196_ gnd vdd FILL
XFILL_0__15946_ gnd vdd FILL
XFILL_2__11979_ gnd vdd FILL
XFILL_0__11069_ gnd vdd FILL
XFILL112440x9050 gnd vdd FILL
X_8003_ _8001_/Y _7955_/B _8002_/Y gnd _8003_/Y vdd OAI21X1
XFILL_4__15327_ gnd vdd FILL
XFILL_5__14878_ gnd vdd FILL
XFILL_2__13718_ gnd vdd FILL
XFILL_3__7365_ gnd vdd FILL
XFILL_1__15147_ gnd vdd FILL
XFILL_1__12359_ gnd vdd FILL
XFILL_2__14698_ gnd vdd FILL
XSFILL38840x58050 gnd vdd FILL
XFILL_6__7074_ gnd vdd FILL
XFILL_0__15877_ gnd vdd FILL
XFILL_3__9104_ gnd vdd FILL
XFILL_5__13829_ gnd vdd FILL
XFILL112360x65050 gnd vdd FILL
XFILL_0__7587_ gnd vdd FILL
XFILL_4__15258_ gnd vdd FILL
XFILL_2__13649_ gnd vdd FILL
XFILL_3__7296_ gnd vdd FILL
XFILL_3__15988_ gnd vdd FILL
XFILL_0__14828_ gnd vdd FILL
XFILL_1__15078_ gnd vdd FILL
XSFILL39480x24050 gnd vdd FILL
XFILL_4__14209_ gnd vdd FILL
XSFILL79080x10050 gnd vdd FILL
XFILL_3__9035_ gnd vdd FILL
X_9954_ _9954_/Q _6998_/CLK _9430_/R vdd _9884_/Y gnd vdd DFFSR
XFILL_4__15189_ gnd vdd FILL
XFILL_1__14029_ gnd vdd FILL
XFILL_3__14939_ gnd vdd FILL
XFILL_2__16368_ gnd vdd FILL
XFILL_0__14759_ gnd vdd FILL
XSFILL79320x72050 gnd vdd FILL
XSFILL43960x49050 gnd vdd FILL
X_8905_ _8903_/Y _8859_/A _8905_/C gnd _8945_/D vdd OAI21X1
XFILL_0__9257_ gnd vdd FILL
XFILL_2__15319_ gnd vdd FILL
X_9885_ _9955_/Q gnd _9887_/A vdd INVX1
XFILL_2__16299_ gnd vdd FILL
XFILL_0__8208_ gnd vdd FILL
X_8836_ _8836_/A _8845_/B _8835_/Y gnd _8922_/D vdd OAI21X1
XSFILL114520x81050 gnd vdd FILL
XSFILL8600x35050 gnd vdd FILL
XSFILL44040x58050 gnd vdd FILL
XFILL_4__6991_ gnd vdd FILL
XFILL_0__8139_ gnd vdd FILL
XSFILL84440x63050 gnd vdd FILL
X_8767_ _8740_/A _8255_/B gnd _8768_/C vdd NAND2X1
XFILL_6_BUFX2_insert843 gnd vdd FILL
XBUFX2_insert909 _10913_/Y gnd _12721_/B vdd BUFX2
XFILL_4__8730_ gnd vdd FILL
XFILL_3__9937_ gnd vdd FILL
X_7718_ _7782_/Q gnd _7718_/Y vdd INVX1
XFILL_6__6858_ gnd vdd FILL
XFILL_1__8952_ gnd vdd FILL
XSFILL23880x16050 gnd vdd FILL
X_8698_ _8698_/A _8314_/B gnd _8699_/C vdd NAND2X1
XFILL_3__9868_ gnd vdd FILL
XFILL_4__8661_ gnd vdd FILL
X_7649_ _7575_/A _8289_/CLK _7649_/R vdd _7577_/Y gnd vdd DFFSR
XFILL_1__8883_ gnd vdd FILL
XFILL_4__7612_ gnd vdd FILL
XSFILL38920x38050 gnd vdd FILL
XFILL_4__8592_ gnd vdd FILL
XFILL112440x45050 gnd vdd FILL
XFILL_3__9799_ gnd vdd FILL
XFILL_1__7834_ gnd vdd FILL
XSFILL23720x80050 gnd vdd FILL
XFILL_4__7543_ gnd vdd FILL
XSFILL38520x40050 gnd vdd FILL
X_11250_ _11787_/C _11249_/Y gnd _11251_/B vdd NAND2X1
XFILL_6__8459_ gnd vdd FILL
XSFILL39000x47050 gnd vdd FILL
X_9319_ _9257_/A _7912_/CLK _7911_/R vdd _9259_/Y gnd vdd DFFSR
XFILL_1__7765_ gnd vdd FILL
X_10201_ _10201_/Q _7021_/CLK _9069_/R vdd _10113_/Y gnd vdd DFFSR
XFILL_4__7474_ gnd vdd FILL
XSFILL3640x78050 gnd vdd FILL
XFILL_1__9504_ gnd vdd FILL
X_11181_ _11179_/Y _11180_/Y gnd _11181_/Y vdd NOR2X1
XSFILL3720x6050 gnd vdd FILL
XFILL_1__7696_ gnd vdd FILL
XFILL_4__9213_ gnd vdd FILL
XFILL_3_BUFX2_insert700 gnd vdd FILL
XFILL_3_BUFX2_insert711 gnd vdd FILL
X_10132_ _13932_/A gnd _10134_/A vdd INVX1
XSFILL94280x66050 gnd vdd FILL
XSFILL114600x61050 gnd vdd FILL
XFILL_3_BUFX2_insert722 gnd vdd FILL
XSFILL68440x76050 gnd vdd FILL
XFILL_4__9144_ gnd vdd FILL
XFILL_3_BUFX2_insert733 gnd vdd FILL
XFILL_3_BUFX2_insert744 gnd vdd FILL
XFILL_3_BUFX2_insert755 gnd vdd FILL
X_10063_ _10061_/Y _9985_/B _10063_/C gnd _10099_/D vdd OAI21X1
XFILL_3_BUFX2_insert766 gnd vdd FILL
X_14940_ _9683_/A gnd _14941_/A vdd INVX1
XFILL_1__9366_ gnd vdd FILL
XFILL_3_BUFX2_insert777 gnd vdd FILL
XFILL_3_BUFX2_insert788 gnd vdd FILL
XFILL_3_BUFX2_insert799 gnd vdd FILL
XFILL_2__7110_ gnd vdd FILL
XFILL_1__8317_ gnd vdd FILL
X_14871_ _7757_/A gnd _14871_/Y vdd INVX1
XFILL_2__8090_ gnd vdd FILL
XFILL_1__9297_ gnd vdd FILL
X_13822_ _9611_/A gnd _13822_/Y vdd INVX1
XFILL_2__7041_ gnd vdd FILL
XFILL_1__8248_ gnd vdd FILL
X_13753_ _8968_/A gnd _13755_/D vdd INVX1
X_10965_ _10898_/Y _10938_/A gnd _10965_/Y vdd OR2X2
XFILL_5__10490_ gnd vdd FILL
XSFILL18760x6050 gnd vdd FILL
X_12704_ _12704_/A gnd _12704_/Y vdd INVX1
XFILL_5__8770_ gnd vdd FILL
XFILL_4__9977_ gnd vdd FILL
X_13684_ _13684_/A _13683_/Y _13684_/C gnd _13684_/Y vdd NAND3X1
XFILL_3__10620_ gnd vdd FILL
XSFILL13880x48050 gnd vdd FILL
X_10896_ _10896_/A _10890_/Y _10877_/Y gnd _10896_/Y vdd OAI21X1
XFILL_0__10440_ gnd vdd FILL
XFILL_2__8992_ gnd vdd FILL
XFILL_5__7721_ gnd vdd FILL
X_12635_ _12635_/A vdd _12635_/C gnd _12685_/D vdd OAI21X1
X_15423_ _15172_/A _15423_/B _16155_/D _15423_/D gnd _15423_/Y vdd OAI22X1
XFILL_0_BUFX2_insert601 gnd vdd FILL
XFILL_4__11910_ gnd vdd FILL
XFILL_5__12160_ gnd vdd FILL
XFILL_0_BUFX2_insert612 gnd vdd FILL
XFILL_2__11000_ gnd vdd FILL
XFILL_3__10551_ gnd vdd FILL
XFILL_0_BUFX2_insert623 gnd vdd FILL
XFILL_4__12890_ gnd vdd FILL
XFILL_2__7943_ gnd vdd FILL
XFILL_1__11730_ gnd vdd FILL
XFILL_0_BUFX2_insert634 gnd vdd FILL
XFILL_0__10371_ gnd vdd FILL
XSFILL94360x46050 gnd vdd FILL
X_15354_ _15354_/A _15354_/B _15353_/Y gnd _15355_/A vdd NAND3X1
XFILL_4__8859_ gnd vdd FILL
XFILL_0_BUFX2_insert645 gnd vdd FILL
XFILL_5__11111_ gnd vdd FILL
XFILL_0_BUFX2_insert656 gnd vdd FILL
XFILL_6__10662_ gnd vdd FILL
XFILL_5__12091_ gnd vdd FILL
X_12566_ _12436_/A _13201_/CLK _13201_/R vdd _12566_/D gnd vdd DFFSR
XFILL_3__13270_ gnd vdd FILL
XFILL_0__12110_ gnd vdd FILL
XFILL_4__11841_ gnd vdd FILL
XFILL_0_BUFX2_insert667 gnd vdd FILL
XFILL_2__7874_ gnd vdd FILL
XFILL_0__13090_ gnd vdd FILL
XFILL_1__11661_ gnd vdd FILL
XFILL_0_BUFX2_insert678 gnd vdd FILL
XFILL_0_BUFX2_insert689 gnd vdd FILL
X_14305_ _14305_/A _14305_/B gnd _14310_/C vdd NOR2X1
X_11517_ _11527_/B gnd _11517_/Y vdd INVX1
XFILL_5__7583_ gnd vdd FILL
XFILL_5__11042_ gnd vdd FILL
X_15285_ _15285_/A _15285_/B gnd _15295_/A vdd NAND2X1
XFILL_3__12221_ gnd vdd FILL
XFILL_2__9613_ gnd vdd FILL
XFILL_4__14560_ gnd vdd FILL
XFILL_1__13400_ gnd vdd FILL
X_12497_ vdd _12065_/A gnd _12498_/C vdd NAND2X1
XFILL_0__12041_ gnd vdd FILL
XFILL_2__12951_ gnd vdd FILL
XFILL_4__11772_ gnd vdd FILL
XFILL_1__14380_ gnd vdd FILL
X_14236_ _9190_/Q gnd _14237_/A vdd INVX1
XFILL_1__11592_ gnd vdd FILL
XFILL_5__15850_ gnd vdd FILL
X_11448_ _11448_/A _11448_/B gnd _11448_/Y vdd AND2X2
XFILL_4__13511_ gnd vdd FILL
XFILL_2__11902_ gnd vdd FILL
XFILL_3__12152_ gnd vdd FILL
XSFILL104360x31050 gnd vdd FILL
XFILL_1__13331_ gnd vdd FILL
XFILL_4__14491_ gnd vdd FILL
XFILL_2__15670_ gnd vdd FILL
XFILL_2__9544_ gnd vdd FILL
XFILL_2__12882_ gnd vdd FILL
XFILL_1__10543_ gnd vdd FILL
XFILL_5__9253_ gnd vdd FILL
XFILL_5__14801_ gnd vdd FILL
XFILL_4__16230_ gnd vdd FILL
XSFILL33640x63050 gnd vdd FILL
X_14167_ _15611_/B _13836_/B _14862_/C _15646_/C gnd _14168_/A vdd OAI22X1
XFILL_3__11103_ gnd vdd FILL
XSFILL74280x13050 gnd vdd FILL
XFILL_2__14621_ gnd vdd FILL
XFILL_4__13442_ gnd vdd FILL
XFILL_5__15781_ gnd vdd FILL
XFILL_4__10654_ gnd vdd FILL
X_11379_ _11377_/Y _11379_/B _11379_/C gnd _11379_/Y vdd OAI21X1
XFILL_2__9475_ gnd vdd FILL
XFILL_3__12083_ gnd vdd FILL
XFILL_5__12993_ gnd vdd FILL
XFILL_0__15800_ gnd vdd FILL
XFILL_1__16050_ gnd vdd FILL
XFILL_2__11833_ gnd vdd FILL
XFILL_1__13262_ gnd vdd FILL
XSFILL8040x72050 gnd vdd FILL
XFILL_5__8204_ gnd vdd FILL
X_13118_ _13188_/Q gnd _13118_/Y vdd INVX1
XFILL_0__13992_ gnd vdd FILL
XFILL_5__14732_ gnd vdd FILL
XFILL_3__15911_ gnd vdd FILL
XFILL_1__15001_ gnd vdd FILL
XFILL_5__11944_ gnd vdd FILL
XSFILL89320x35050 gnd vdd FILL
XFILL_0__8490_ gnd vdd FILL
X_14098_ _14273_/C _8477_/A _14098_/C _14214_/C gnd _14106_/C vdd AOI22X1
XFILL_4__16161_ gnd vdd FILL
XFILL_3__11034_ gnd vdd FILL
XFILL_2__14552_ gnd vdd FILL
XFILL_1__12213_ gnd vdd FILL
XFILL_4__13373_ gnd vdd FILL
XFILL_0__15731_ gnd vdd FILL
XFILL_5__8135_ gnd vdd FILL
XFILL_2__11764_ gnd vdd FILL
XFILL_0__7441_ gnd vdd FILL
XFILL_4__15112_ gnd vdd FILL
X_13049_ _6872_/A _8169_/CLK _8937_/R vdd _12959_/Y gnd vdd DFFSR
XFILL_4__12324_ gnd vdd FILL
XFILL_5__14663_ gnd vdd FILL
XFILL_2__13503_ gnd vdd FILL
XFILL_5__11875_ gnd vdd FILL
XFILL_2__8357_ gnd vdd FILL
XSFILL12920x64050 gnd vdd FILL
XFILL_4__16092_ gnd vdd FILL
XFILL_3__15842_ gnd vdd FILL
XFILL_2__14483_ gnd vdd FILL
XFILL_1__12144_ gnd vdd FILL
XFILL_0__15662_ gnd vdd FILL
XFILL_5__8066_ gnd vdd FILL
XFILL_2__11695_ gnd vdd FILL
XFILL_5__16402_ gnd vdd FILL
XFILL_5__13614_ gnd vdd FILL
XFILL_0__12874_ gnd vdd FILL
XFILL_0__7372_ gnd vdd FILL
XFILL_2__7308_ gnd vdd FILL
XFILL_2__16222_ gnd vdd FILL
XFILL_5__10826_ gnd vdd FILL
XFILL_4__15043_ gnd vdd FILL
XFILL_5__14594_ gnd vdd FILL
XFILL_2__13434_ gnd vdd FILL
XFILL_4__12255_ gnd vdd FILL
XSFILL94440x26050 gnd vdd FILL
XFILL_0__14613_ gnd vdd FILL
XFILL_3__15773_ gnd vdd FILL
XFILL_2__10646_ gnd vdd FILL
XFILL_3__7081_ gnd vdd FILL
XFILL_1__12075_ gnd vdd FILL
XFILL_0__9111_ gnd vdd FILL
XFILL_3__12985_ gnd vdd FILL
XFILL_0__11825_ gnd vdd FILL
XFILL_5__16333_ gnd vdd FILL
XFILL_0__15593_ gnd vdd FILL
XFILL_5__13545_ gnd vdd FILL
XFILL_4__11206_ gnd vdd FILL
X_6951_ _6951_/A _7847_/B gnd _6952_/C vdd NAND2X1
XFILL_4__12186_ gnd vdd FILL
XFILL_3__14724_ gnd vdd FILL
XFILL_5__10757_ gnd vdd FILL
XFILL_2__7239_ gnd vdd FILL
XFILL_2__16153_ gnd vdd FILL
XFILL_6__15884_ gnd vdd FILL
XFILL_2__13365_ gnd vdd FILL
XFILL_1__15903_ gnd vdd FILL
XFILL_3__11936_ gnd vdd FILL
XFILL_1__11026_ gnd vdd FILL
XFILL_0__14544_ gnd vdd FILL
XFILL_2__10577_ gnd vdd FILL
XFILL_0__9042_ gnd vdd FILL
XFILL_0__11756_ gnd vdd FILL
XFILL_6__14835_ gnd vdd FILL
XFILL_4__11137_ gnd vdd FILL
XFILL_2__15104_ gnd vdd FILL
XFILL_5__16264_ gnd vdd FILL
XFILL_5__13476_ gnd vdd FILL
X_9670_ _9668_/Y _9625_/B _9670_/C gnd _9712_/D vdd OAI21X1
XFILL_2__12316_ gnd vdd FILL
XFILL_5__10688_ gnd vdd FILL
X_6882_ _6882_/A gnd memoryWriteData[12] vdd BUFX2
XFILL_1__15834_ gnd vdd FILL
XFILL_3__14655_ gnd vdd FILL
XFILL_2__16084_ gnd vdd FILL
XFILL_2__13296_ gnd vdd FILL
XFILL_6_BUFX2_insert106 gnd vdd FILL
XFILL_3__11867_ gnd vdd FILL
XFILL_0__10707_ gnd vdd FILL
XFILL_0__14475_ gnd vdd FILL
XFILL_5__15215_ gnd vdd FILL
XSFILL104440x11050 gnd vdd FILL
XFILL_5__12427_ gnd vdd FILL
XFILL_5__8968_ gnd vdd FILL
X_8621_ _8567_/B _9517_/B gnd _8622_/C vdd NAND2X1
XFILL_0__11687_ gnd vdd FILL
XFILL_6__7761_ gnd vdd FILL
XFILL_3__13606_ gnd vdd FILL
XFILL_5__16195_ gnd vdd FILL
XFILL_2__15035_ gnd vdd FILL
XFILL_4__15945_ gnd vdd FILL
XFILL_6__11978_ gnd vdd FILL
XFILL_4__11068_ gnd vdd FILL
XSFILL83880x71050 gnd vdd FILL
XFILL_0__16214_ gnd vdd FILL
XFILL_2__12247_ gnd vdd FILL
XFILL_3__10818_ gnd vdd FILL
XSFILL84360x78050 gnd vdd FILL
XFILL_3__14586_ gnd vdd FILL
XFILL_0__13426_ gnd vdd FILL
XFILL_1__15765_ gnd vdd FILL
XFILL_3__11798_ gnd vdd FILL
XFILL_0__10638_ gnd vdd FILL
XFILL_1__12977_ gnd vdd FILL
XFILL_3__7983_ gnd vdd FILL
XFILL_4__10019_ gnd vdd FILL
XFILL_5__15146_ gnd vdd FILL
XFILL_5__12358_ gnd vdd FILL
XFILL_1_BUFX2_insert490 gnd vdd FILL
XFILL_6__14697_ gnd vdd FILL
X_8552_ _8492_/A _7400_/CLK _9704_/R vdd _8494_/Y gnd vdd DFFSR
XFILL_3__16325_ gnd vdd FILL
XFILL_5__8899_ gnd vdd FILL
XFILL_1__14716_ gnd vdd FILL
XFILL_3__10749_ gnd vdd FILL
XFILL_3__13537_ gnd vdd FILL
XFILL_3__9722_ gnd vdd FILL
XFILL_4__15876_ gnd vdd FILL
XFILL_2__12178_ gnd vdd FILL
XFILL_5_BUFX2_insert806 gnd vdd FILL
XFILL_1__11928_ gnd vdd FILL
XFILL_3__6934_ gnd vdd FILL
XSFILL89400x15050 gnd vdd FILL
XFILL_0__16145_ gnd vdd FILL
XFILL_0__13357_ gnd vdd FILL
XFILL_1__15696_ gnd vdd FILL
XFILL_5_BUFX2_insert817 gnd vdd FILL
X_7503_ _7503_/A _7503_/B _7502_/Y gnd _7503_/Y vdd OAI21X1
XFILL_6__13648_ gnd vdd FILL
XFILL_5_BUFX2_insert828 gnd vdd FILL
XFILL_5__11309_ gnd vdd FILL
XFILL_0__10569_ gnd vdd FILL
XBUFX2_insert1003 _12399_/Y gnd _9901_/B vdd BUFX2
XFILL_4__14827_ gnd vdd FILL
XFILL_5__15077_ gnd vdd FILL
XFILL_5_BUFX2_insert839 gnd vdd FILL
X_8483_ _8549_/Q gnd _8485_/A vdd INVX1
XFILL_5__12289_ gnd vdd FILL
XFILL_2__11129_ gnd vdd FILL
XFILL_3__16256_ gnd vdd FILL
XFILL_3__9653_ gnd vdd FILL
XFILL_1__14647_ gnd vdd FILL
XBUFX2_insert1014 _15054_/Y gnd _15376_/B vdd BUFX2
XFILL_3__13468_ gnd vdd FILL
XFILL_3__6865_ gnd vdd FILL
XFILL_0__12308_ gnd vdd FILL
XBUFX2_insert1025 _13340_/Y gnd _9615_/A vdd BUFX2
XFILL_1__11859_ gnd vdd FILL
XFILL_0__16076_ gnd vdd FILL
XFILL_0__13288_ gnd vdd FILL
XBUFX2_insert1036 _12390_/Y gnd _9380_/B vdd BUFX2
XFILL111880x53050 gnd vdd FILL
XFILL_5__14028_ gnd vdd FILL
XFILL_3__15207_ gnd vdd FILL
X_7434_ _7434_/A _7460_/A _7433_/Y gnd _7434_/Y vdd OAI21X1
XBUFX2_insert1047 _13297_/Y gnd _7684_/B vdd BUFX2
XFILL_3__12419_ gnd vdd FILL
XFILL_3__8604_ gnd vdd FILL
XFILL_0__9875_ gnd vdd FILL
XFILL_4__14758_ gnd vdd FILL
XFILL_3__16187_ gnd vdd FILL
XFILL_0__15027_ gnd vdd FILL
XFILL_3__13399_ gnd vdd FILL
XFILL_2__15937_ gnd vdd FILL
XBUFX2_insert1058 _15051_/Y gnd _15764_/C vdd BUFX2
XFILL_1__14578_ gnd vdd FILL
XFILL_0__12239_ gnd vdd FILL
XBUFX2_insert1069 _13327_/Y gnd _8902_/B vdd BUFX2
XFILL_6__16298_ gnd vdd FILL
XFILL_0__8826_ gnd vdd FILL
XFILL_4__13709_ gnd vdd FILL
X_7365_ _7366_/B _9797_/B gnd _7365_/Y vdd NAND2X1
XFILL_1__16317_ gnd vdd FILL
XFILL_3__15138_ gnd vdd FILL
XFILL_4__14689_ gnd vdd FILL
XFILL_1__13529_ gnd vdd FILL
XFILL_2__15868_ gnd vdd FILL
X_9104_ _9104_/A _9163_/A _9104_/C gnd _9182_/D vdd OAI21X1
XSFILL79320x67050 gnd vdd FILL
XFILL_0__8757_ gnd vdd FILL
XFILL_1__7550_ gnd vdd FILL
X_7296_ _7297_/B _7424_/B gnd _7297_/C vdd NAND2X1
XFILL_5__15979_ gnd vdd FILL
XFILL_2__14819_ gnd vdd FILL
XFILL_3__15069_ gnd vdd FILL
XFILL_3__8466_ gnd vdd FILL
XFILL_1__16248_ gnd vdd FILL
XFILL_0__7708_ gnd vdd FILL
XFILL_2__15799_ gnd vdd FILL
X_9035_ _8969_/A _7243_/B gnd _9036_/C vdd NAND2X1
XFILL_4__16359_ gnd vdd FILL
XFILL_1__7481_ gnd vdd FILL
XSFILL114520x76050 gnd vdd FILL
XFILL_3__7417_ gnd vdd FILL
XFILL_3__8397_ gnd vdd FILL
XFILL_0__15929_ gnd vdd FILL
XFILL_1__16179_ gnd vdd FILL
XFILL_4__7190_ gnd vdd FILL
XFILL_1__9220_ gnd vdd FILL
XSFILL33800x23050 gnd vdd FILL
XFILL_3__7348_ gnd vdd FILL
XSFILL99240x18050 gnd vdd FILL
XFILL_2_BUFX2_insert707 gnd vdd FILL
XFILL_1__9151_ gnd vdd FILL
XFILL_2_BUFX2_insert718 gnd vdd FILL
XSFILL28760x1050 gnd vdd FILL
XFILL_2_BUFX2_insert729 gnd vdd FILL
XFILL_1__8102_ gnd vdd FILL
XFILL_1__9082_ gnd vdd FILL
X_9937_ _9937_/A _8401_/B gnd _9938_/C vdd NAND2X1
XFILL_3__9018_ gnd vdd FILL
XFILL_4__9900_ gnd vdd FILL
XFILL111960x33050 gnd vdd FILL
X_9868_ _9868_/A _7564_/B gnd _9868_/Y vdd NAND2X1
XSFILL23720x75050 gnd vdd FILL
X_10750_ _10750_/A _10809_/A _10749_/Y gnd _10750_/Y vdd OAI21X1
X_8819_ _8819_/Q _9707_/CLK _8819_/R vdd _8819_/D gnd vdd DFFSR
XFILL112040x42050 gnd vdd FILL
X_9799_ _9841_/Q gnd _9801_/A vdd INVX1
XFILL_4__9762_ gnd vdd FILL
XBUFX2_insert706 _11985_/Y gnd _12084_/C vdd BUFX2
XSFILL79400x47050 gnd vdd FILL
XFILL_4__6974_ gnd vdd FILL
XBUFX2_insert717 _13418_/Y gnd _14778_/B vdd BUFX2
X_10681_ _10681_/A _9785_/B gnd _10682_/C vdd NAND2X1
XBUFX2_insert728 _12411_/Y gnd _9785_/B vdd BUFX2
XFILL_1__9984_ gnd vdd FILL
XFILL_4__8713_ gnd vdd FILL
XFILL_6_BUFX2_insert684 gnd vdd FILL
XBUFX2_insert739 _12402_/Y gnd _7856_/B vdd BUFX2
X_12420_ _12418_/Y _12419_/A _12420_/C gnd _12420_/Y vdd OAI21X1
XFILL_4__8644_ gnd vdd FILL
X_12351_ _12349_/Y _12419_/A _12351_/C gnd _12351_/Y vdd OAI21X1
XSFILL69080x37050 gnd vdd FILL
XFILL_1_CLKBUF1_insert111 gnd vdd FILL
XFILL_1__8866_ gnd vdd FILL
XFILL_1_CLKBUF1_insert122 gnd vdd FILL
XFILL_1_CLKBUF1_insert133 gnd vdd FILL
X_11302_ _11301_/Y _11298_/Y gnd _11536_/C vdd NAND2X1
XFILL_4__8575_ gnd vdd FILL
X_15070_ _13417_/Y _15328_/B _15070_/C _13457_/Y gnd _15074_/B vdd OAI22X1
XFILL_1_CLKBUF1_insert144 gnd vdd FILL
X_12282_ _12279_/Y _12282_/B _12282_/C gnd _12282_/Y vdd NAND3X1
XFILL_1__7817_ gnd vdd FILL
XFILL_1_CLKBUF1_insert155 gnd vdd FILL
XFILL_2__7590_ gnd vdd FILL
XFILL_1_CLKBUF1_insert166 gnd vdd FILL
X_14021_ _14868_/D _9185_/Q _15509_/A _14877_/D gnd _14022_/B vdd AOI22X1
XFILL_1_CLKBUF1_insert177 gnd vdd FILL
XFILL_1_CLKBUF1_insert188 gnd vdd FILL
X_11233_ _12226_/Y _11013_/B gnd _11376_/B vdd NOR2X1
XFILL_1_CLKBUF1_insert199 gnd vdd FILL
XFILL_1__7748_ gnd vdd FILL
XFILL_2_BUFX2_insert9 gnd vdd FILL
XFILL_4__7457_ gnd vdd FILL
XSFILL73960x83050 gnd vdd FILL
X_11164_ _11143_/A _11159_/Y _11163_/Y gnd _11408_/A vdd AOI21X1
XSFILL94600x7050 gnd vdd FILL
XSFILL23800x55050 gnd vdd FILL
XFILL_2__9260_ gnd vdd FILL
XFILL_1__7679_ gnd vdd FILL
XFILL_3_BUFX2_insert530 gnd vdd FILL
X_10115_ _10166_/A _9859_/B gnd _10116_/C vdd NAND2X1
XFILL_3_BUFX2_insert541 gnd vdd FILL
XFILL112120x22050 gnd vdd FILL
XFILL_2__8211_ gnd vdd FILL
X_15972_ _15972_/A _15972_/B _15972_/C _14566_/Y gnd _15972_/Y vdd OAI22X1
XFILL_1__9418_ gnd vdd FILL
XFILL_4__10370_ gnd vdd FILL
X_11095_ _11092_/Y _11061_/C _11094_/Y gnd _11096_/C vdd AOI21X1
XFILL_3_BUFX2_insert552 gnd vdd FILL
XFILL_3_BUFX2_insert563 gnd vdd FILL
XFILL_1__10190_ gnd vdd FILL
XFILL_4__9127_ gnd vdd FILL
XFILL_3_BUFX2_insert574 gnd vdd FILL
XFILL_3_BUFX2_insert585 gnd vdd FILL
X_10046_ _10094_/Q gnd _10048_/A vdd INVX1
X_14923_ _14721_/A _16263_/A _14545_/B _14923_/D gnd _14924_/B vdd OAI22X1
XFILL_2__8142_ gnd vdd FILL
XFILL_3_BUFX2_insert596 gnd vdd FILL
XFILL_2__10500_ gnd vdd FILL
XFILL_5__11660_ gnd vdd FILL
XFILL_1__9349_ gnd vdd FILL
XSFILL93880x34050 gnd vdd FILL
XFILL_2__11480_ gnd vdd FILL
XFILL_5__9940_ gnd vdd FILL
XFILL_4__12040_ gnd vdd FILL
XSFILL104040x3050 gnd vdd FILL
X_14854_ _16408_/A gnd _14854_/Y vdd INVX1
XFILL_2__8073_ gnd vdd FILL
XFILL_3__12770_ gnd vdd FILL
XFILL_2__10431_ gnd vdd FILL
XSFILL53880x50050 gnd vdd FILL
XFILL_5__11591_ gnd vdd FILL
XFILL_0__11610_ gnd vdd FILL
XFILL_4__8009_ gnd vdd FILL
XFILL_6__11901_ gnd vdd FILL
XFILL_0__12590_ gnd vdd FILL
XFILL_5__13330_ gnd vdd FILL
XFILL_5__9871_ gnd vdd FILL
X_13805_ _13804_/Y _13805_/B gnd _13805_/Y vdd NAND2X1
XSFILL69160x17050 gnd vdd FILL
XFILL_5__10542_ gnd vdd FILL
XFILL_2__13150_ gnd vdd FILL
X_11997_ _11997_/A _12093_/B _12061_/C gnd gnd _11998_/C vdd AOI22X1
XFILL_3__11721_ gnd vdd FILL
XFILL_1__12900_ gnd vdd FILL
X_14785_ _14784_/Y _14949_/C gnd _14788_/A vdd NOR2X1
XFILL_6_BUFX2_insert45 gnd vdd FILL
XFILL_2__10362_ gnd vdd FILL
XFILL_1__13880_ gnd vdd FILL
XFILL_5__8822_ gnd vdd FILL
XFILL_0__11541_ gnd vdd FILL
XSFILL84200x20050 gnd vdd FILL
XFILL_6__14620_ gnd vdd FILL
XFILL_5__13261_ gnd vdd FILL
X_10948_ _10930_/Y _10948_/B gnd _10948_/Y vdd NAND2X1
XFILL_2__12101_ gnd vdd FILL
X_13736_ _15275_/A _14344_/B _14283_/C _9947_/Q gnd _13736_/Y vdd AOI22X1
XSFILL104360x26050 gnd vdd FILL
XFILL_3__11652_ gnd vdd FILL
XFILL_3__14440_ gnd vdd FILL
XFILL_2__13081_ gnd vdd FILL
XFILL_4__13991_ gnd vdd FILL
XFILL_1__12831_ gnd vdd FILL
XFILL_2__10293_ gnd vdd FILL
XFILL_0__14260_ gnd vdd FILL
XFILL_5__15000_ gnd vdd FILL
XSFILL104520x9050 gnd vdd FILL
XFILL_0__11472_ gnd vdd FILL
XFILL_5__12212_ gnd vdd FILL
XFILL_5__8753_ gnd vdd FILL
XFILL_4__15730_ gnd vdd FILL
XFILL_6__11763_ gnd vdd FILL
X_13667_ _7130_/Q gnd _13669_/D vdd INVX1
XFILL_2__12032_ gnd vdd FILL
X_10879_ _12695_/A _12792_/Q gnd _10879_/Y vdd NOR2X1
XFILL_3__14371_ gnd vdd FILL
XFILL_0__13211_ gnd vdd FILL
XFILL_1__15550_ gnd vdd FILL
XFILL_3__11583_ gnd vdd FILL
XFILL_0__10423_ gnd vdd FILL
XFILL_1__12762_ gnd vdd FILL
XFILL_2__8975_ gnd vdd FILL
XFILL_5__7704_ gnd vdd FILL
XFILL_0_BUFX2_insert420 gnd vdd FILL
X_15406_ _8414_/Q gnd _15407_/A vdd INVX1
XFILL_0__14191_ gnd vdd FILL
XFILL_0_BUFX2_insert431 gnd vdd FILL
X_12618_ _12618_/A gnd _12618_/Y vdd INVX1
XFILL_6__14482_ gnd vdd FILL
XFILL_3__16110_ gnd vdd FILL
XFILL_5__12143_ gnd vdd FILL
XFILL_0__7990_ gnd vdd FILL
XFILL_3__10534_ gnd vdd FILL
XFILL_3__13322_ gnd vdd FILL
X_16386_ _16386_/A gnd _16385_/Y gnd _16386_/Y vdd OAI21X1
XSFILL59080x69050 gnd vdd FILL
X_13598_ _13597_/Y _13860_/B _13857_/C _13596_/Y gnd _13602_/B vdd OAI22X1
XFILL_4__15661_ gnd vdd FILL
XFILL_1__14501_ gnd vdd FILL
XFILL_0_BUFX2_insert442 gnd vdd FILL
XFILL_0_BUFX2_insert453 gnd vdd FILL
XFILL_2__7926_ gnd vdd FILL
XFILL_4__12873_ gnd vdd FILL
XFILL_1__11713_ gnd vdd FILL
XFILL_0__13142_ gnd vdd FILL
XFILL_0_BUFX2_insert464 gnd vdd FILL
XFILL_1__15481_ gnd vdd FILL
XFILL_0_BUFX2_insert475 gnd vdd FILL
XFILL_5__7635_ gnd vdd FILL
XFILL_4__14612_ gnd vdd FILL
X_15337_ _15324_/Y _15337_/B gnd _15338_/B vdd NOR2X1
X_12549_ _12385_/A _12537_/CLK _9060_/R vdd _12549_/D gnd vdd DFFSR
XFILL_0__6941_ gnd vdd FILL
XFILL_3__13253_ gnd vdd FILL
XSFILL74120x72050 gnd vdd FILL
XFILL_3__16041_ gnd vdd FILL
XFILL_5__12074_ gnd vdd FILL
XFILL_0_BUFX2_insert486 gnd vdd FILL
XFILL_4__11824_ gnd vdd FILL
XFILL_0_BUFX2_insert497 gnd vdd FILL
XFILL_4__15592_ gnd vdd FILL
XFILL_1__14432_ gnd vdd FILL
XFILL_2__13983_ gnd vdd FILL
XFILL_2__7857_ gnd vdd FILL
XFILL_1__11644_ gnd vdd FILL
XFILL_0__10285_ gnd vdd FILL
XFILL_0__9660_ gnd vdd FILL
XFILL_5__7566_ gnd vdd FILL
XFILL_5__15902_ gnd vdd FILL
XFILL_3__12204_ gnd vdd FILL
XFILL_5__11025_ gnd vdd FILL
XFILL_4__14543_ gnd vdd FILL
X_15268_ _15268_/A gnd _15268_/Y vdd INVX1
XFILL_0__6872_ gnd vdd FILL
XFILL_2__15722_ gnd vdd FILL
XFILL_4__11755_ gnd vdd FILL
XFILL_0__12024_ gnd vdd FILL
XFILL_3__10396_ gnd vdd FILL
XFILL_1__14363_ gnd vdd FILL
XFILL_0__8611_ gnd vdd FILL
XFILL_1__11575_ gnd vdd FILL
X_14219_ _8166_/Q gnd _14219_/Y vdd INVX1
XSFILL53960x30050 gnd vdd FILL
XFILL_6__13295_ gnd vdd FILL
XFILL_3__8320_ gnd vdd FILL
X_7150_ _7150_/Q _7902_/CLK _7150_/R vdd _7104_/Y gnd vdd DFFSR
X_15199_ _6911_/A gnd _15200_/B vdd INVX1
XFILL_3__12135_ gnd vdd FILL
XFILL_0__9591_ gnd vdd FILL
XFILL_5__7497_ gnd vdd FILL
XFILL_1__16102_ gnd vdd FILL
XFILL_5__15833_ gnd vdd FILL
XFILL_4__10706_ gnd vdd FILL
XFILL_1__13314_ gnd vdd FILL
XFILL_2__9527_ gnd vdd FILL
XFILL_4__14474_ gnd vdd FILL
XFILL_2__15653_ gnd vdd FILL
XFILL_2__12865_ gnd vdd FILL
XFILL_4__11686_ gnd vdd FILL
XFILL_1__10526_ gnd vdd FILL
XFILL_1__14294_ gnd vdd FILL
XFILL_5__9236_ gnd vdd FILL
XFILL_4__16213_ gnd vdd FILL
XFILL_4__13425_ gnd vdd FILL
XCLKBUF1_insert121 CLKBUF1_insert220/A gnd _7010_/CLK vdd CLKBUF1
XFILL_5__15764_ gnd vdd FILL
X_7081_ _7081_/A gnd _7081_/Y vdd INVX1
XFILL_4__10637_ gnd vdd FILL
XFILL_3__8251_ gnd vdd FILL
XFILL_5__12976_ gnd vdd FILL
XFILL_2__14604_ gnd vdd FILL
XFILL_1__16033_ gnd vdd FILL
XFILL_3__12066_ gnd vdd FILL
XCLKBUF1_insert132 CLKBUF1_insert220/A gnd _8818_/CLK vdd CLKBUF1
XFILL_2__11816_ gnd vdd FILL
XFILL_1__13245_ gnd vdd FILL
XCLKBUF1_insert143 CLKBUF1_insert187/A gnd _12537_/CLK vdd CLKBUF1
XSFILL83720x8050 gnd vdd FILL
XCLKBUF1_insert154 CLKBUF1_insert169/A gnd _7647_/CLK vdd CLKBUF1
XFILL_2__15584_ gnd vdd FILL
XFILL_5__9167_ gnd vdd FILL
XFILL_5__14715_ gnd vdd FILL
XFILL_0__13975_ gnd vdd FILL
XFILL_0__8473_ gnd vdd FILL
XFILL_3__7202_ gnd vdd FILL
XFILL_5__11927_ gnd vdd FILL
XCLKBUF1_insert165 CLKBUF1_insert182/A gnd _9568_/CLK vdd CLKBUF1
XFILL_6__12177_ gnd vdd FILL
XFILL_3__11017_ gnd vdd FILL
XFILL_4__16144_ gnd vdd FILL
XFILL_4__13356_ gnd vdd FILL
XFILL_5__15695_ gnd vdd FILL
XCLKBUF1_insert176 CLKBUF1_insert220/A gnd _6998_/CLK vdd CLKBUF1
XCLKBUF1_insert187 CLKBUF1_insert187/A gnd _12685_/CLK vdd CLKBUF1
XFILL_0__15714_ gnd vdd FILL
XFILL_3__8182_ gnd vdd FILL
XFILL_2__14535_ gnd vdd FILL
XFILL_2__11747_ gnd vdd FILL
XFILL_4__10568_ gnd vdd FILL
XFILL_5__8118_ gnd vdd FILL
XFILL_2__9389_ gnd vdd FILL
XCLKBUF1_insert198 CLKBUF1_insert169/A gnd _7532_/CLK vdd CLKBUF1
XFILL_0__7424_ gnd vdd FILL
XFILL_1__10388_ gnd vdd FILL
XFILL_5__14646_ gnd vdd FILL
XFILL_5__9098_ gnd vdd FILL
XFILL_4__12307_ gnd vdd FILL
XSFILL43880x82050 gnd vdd FILL
XFILL_3__15825_ gnd vdd FILL
XFILL_4__16075_ gnd vdd FILL
XFILL_5__11858_ gnd vdd FILL
XFILL_4__13287_ gnd vdd FILL
XFILL_2__14466_ gnd vdd FILL
XFILL_4__10499_ gnd vdd FILL
XFILL_1__12127_ gnd vdd FILL
XFILL_0__15645_ gnd vdd FILL
XFILL_2__11678_ gnd vdd FILL
XFILL_0__12857_ gnd vdd FILL
XFILL_0__7355_ gnd vdd FILL
XFILL_4__15026_ gnd vdd FILL
XFILL_5__10809_ gnd vdd FILL
XFILL_5__14577_ gnd vdd FILL
XFILL_2__16205_ gnd vdd FILL
XFILL_2__13417_ gnd vdd FILL
XFILL_4__12238_ gnd vdd FILL
XFILL_3__7064_ gnd vdd FILL
X_7983_ _8041_/Q gnd _7983_/Y vdd INVX1
XFILL_2__10629_ gnd vdd FILL
XFILL_5__11789_ gnd vdd FILL
XFILL_3__15756_ gnd vdd FILL
XFILL_1__12058_ gnd vdd FILL
XFILL_2__14397_ gnd vdd FILL
XFILL_0__11808_ gnd vdd FILL
XFILL_3__12968_ gnd vdd FILL
XFILL_5__16316_ gnd vdd FILL
XFILL_0__15576_ gnd vdd FILL
XFILL_0__12788_ gnd vdd FILL
XFILL111880x48050 gnd vdd FILL
XFILL_6__8862_ gnd vdd FILL
XFILL_5__13528_ gnd vdd FILL
X_9722_ _9770_/A _9082_/B gnd _9723_/C vdd NAND2X1
XFILL_0__7286_ gnd vdd FILL
XFILL_3__14707_ gnd vdd FILL
X_6934_ _6932_/Y _6985_/B _6934_/C gnd _7008_/D vdd OAI21X1
XFILL_2__13348_ gnd vdd FILL
XFILL_3__11919_ gnd vdd FILL
XFILL_4__12169_ gnd vdd FILL
XFILL_2__16136_ gnd vdd FILL
XFILL_1__11009_ gnd vdd FILL
XFILL_3__15687_ gnd vdd FILL
XFILL_0__14527_ gnd vdd FILL
XFILL_6__7813_ gnd vdd FILL
XFILL_0__9025_ gnd vdd FILL
XFILL_0__11739_ gnd vdd FILL
XFILL_3__12899_ gnd vdd FILL
XFILL_5__16247_ gnd vdd FILL
X_9653_ _9653_/A gnd _9655_/A vdd INVX1
XFILL_5__13459_ gnd vdd FILL
XFILL_3__14638_ gnd vdd FILL
X_6865_ _6865_/A gnd memoryAddress[27] vdd BUFX2
XFILL_2__16067_ gnd vdd FILL
XFILL_2__13279_ gnd vdd FILL
XFILL_1__15817_ gnd vdd FILL
XFILL_0__14458_ gnd vdd FILL
XSFILL8680x8050 gnd vdd FILL
X_8604_ _8604_/A _8567_/B _8604_/C gnd _8604_/Y vdd OAI21X1
XFILL_4__15928_ gnd vdd FILL
XFILL_5__16178_ gnd vdd FILL
XFILL_2__15018_ gnd vdd FILL
X_9584_ _9584_/Q _9953_/CLK _7276_/R vdd _9584_/D gnd vdd DFFSR
XFILL_3__14569_ gnd vdd FILL
XFILL_0__13409_ gnd vdd FILL
XSFILL38840x71050 gnd vdd FILL
XFILL_1__15748_ gnd vdd FILL
XFILL_3__7966_ gnd vdd FILL
XSFILL39320x78050 gnd vdd FILL
XFILL_5_BUFX2_insert603 gnd vdd FILL
XFILL_0__14389_ gnd vdd FILL
XFILL_5__15129_ gnd vdd FILL
XFILL_5_BUFX2_insert614 gnd vdd FILL
XFILL_3__16308_ gnd vdd FILL
X_8535_ _8441_/A _9205_/CLK _9447_/R vdd _8535_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert625 gnd vdd FILL
XFILL_1__6981_ gnd vdd FILL
XFILL_4__15859_ gnd vdd FILL
XFILL_5_BUFX2_insert636 gnd vdd FILL
XFILL_0__16128_ gnd vdd FILL
XFILL_3__6917_ gnd vdd FILL
XFILL_1__15679_ gnd vdd FILL
XFILL_5_BUFX2_insert647 gnd vdd FILL
XFILL_1__8720_ gnd vdd FILL
XFILL_5_BUFX2_insert658 gnd vdd FILL
XSFILL83960x46050 gnd vdd FILL
XFILL_0__9927_ gnd vdd FILL
XFILL_3__16239_ gnd vdd FILL
XFILL_5_BUFX2_insert669 gnd vdd FILL
X_8466_ _8469_/A _8466_/B gnd _8467_/C vdd NAND2X1
XSFILL33800x18050 gnd vdd FILL
XFILL_3__9636_ gnd vdd FILL
XFILL_3__6848_ gnd vdd FILL
XSFILL49720x9050 gnd vdd FILL
XFILL_0__16059_ gnd vdd FILL
XSFILL43960x62050 gnd vdd FILL
XFILL_1__8651_ gnd vdd FILL
X_7417_ _7511_/Q gnd _7417_/Y vdd INVX1
XFILL_0__9858_ gnd vdd FILL
XSFILL18600x79050 gnd vdd FILL
XFILL_4__8360_ gnd vdd FILL
X_8397_ _8435_/Q gnd _8397_/Y vdd INVX1
XFILL_1__7602_ gnd vdd FILL
XFILL_1__8582_ gnd vdd FILL
X_7348_ _7346_/Y _7354_/B _7347_/Y gnd _7402_/D vdd OAI21X1
XFILL_0__9789_ gnd vdd FILL
XFILL_4__7311_ gnd vdd FILL
XSFILL44040x71050 gnd vdd FILL
XFILL_3__8518_ gnd vdd FILL
XFILL111960x28050 gnd vdd FILL
XFILL_2_CLKBUF1_insert206 gnd vdd FILL
XFILL_3__9498_ gnd vdd FILL
XFILL_2_CLKBUF1_insert217 gnd vdd FILL
XFILL_4__7242_ gnd vdd FILL
X_7279_ _7279_/Q _7535_/CLK _8682_/R vdd _7279_/D gnd vdd DFFSR
XFILL_3__8449_ gnd vdd FILL
X_9018_ _9016_/Y _9017_/A _9018_/C gnd _9068_/D vdd OAI21X1
XFILL_1__7464_ gnd vdd FILL
XFILL112040x37050 gnd vdd FILL
XFILL_4__7173_ gnd vdd FILL
XSFILL23320x72050 gnd vdd FILL
XSFILL38120x32050 gnd vdd FILL
XFILL_2_BUFX2_insert504 gnd vdd FILL
XFILL_2_BUFX2_insert515 gnd vdd FILL
XFILL_2_BUFX2_insert526 gnd vdd FILL
XFILL_2_BUFX2_insert537 gnd vdd FILL
X_11920_ _13186_/Q gnd _11920_/Y vdd INVX1
XFILL_1__9134_ gnd vdd FILL
XFILL_2_BUFX2_insert548 gnd vdd FILL
XFILL_2_BUFX2_insert559 gnd vdd FILL
XSFILL39000x60050 gnd vdd FILL
X_11851_ _11830_/A _11850_/Y gnd _11852_/C vdd NAND2X1
XFILL_6_BUFX2_insert1001 gnd vdd FILL
XFILL_6_BUFX2_insert1012 gnd vdd FILL
X_10802_ _10802_/A gnd _10804_/A vdd INVX1
X_14570_ _14570_/A _14570_/B gnd _14570_/Y vdd NOR2X1
XFILL_1__8016_ gnd vdd FILL
X_11782_ _11769_/A _11776_/A _11360_/C gnd _11782_/Y vdd OAI21X1
X_10733_ _10683_/A _8038_/CLK _8038_/R vdd _10733_/D gnd vdd DFFSR
X_13521_ _8441_/A gnd _13522_/D vdd INVX1
XBUFX2_insert503 BUFX2_insert559/A gnd _9049_/R vdd BUFX2
XBUFX2_insert514 BUFX2_insert520/A gnd _7796_/R vdd BUFX2
XBUFX2_insert525 BUFX2_insert520/A gnd _7408_/R vdd BUFX2
XFILL_4__9745_ gnd vdd FILL
X_16240_ _15915_/C _16239_/Y _15912_/D _14839_/Y gnd _16240_/Y vdd OAI22X1
X_13452_ _13452_/A gnd _15062_/A vdd INVX1
XBUFX2_insert536 BUFX2_insert600/A gnd _8033_/R vdd BUFX2
XFILL_4__6957_ gnd vdd FILL
XBUFX2_insert547 BUFX2_insert518/A gnd _7533_/R vdd BUFX2
X_10664_ _10664_/A _10700_/B _10664_/C gnd _10726_/D vdd OAI21X1
XBUFX2_insert558 BUFX2_insert518/A gnd _8669_/R vdd BUFX2
XFILL_2__8760_ gnd vdd FILL
XBUFX2_insert569 BUFX2_insert600/A gnd _9060_/R vdd BUFX2
X_12403_ _12403_/A gnd _12403_/Y vdd INVX1
XFILL_4__9676_ gnd vdd FILL
X_16171_ _16171_/A _16171_/B gnd _16172_/C vdd NOR2X1
X_13383_ _10358_/A _14389_/B _14626_/A _7286_/A gnd _13401_/B vdd AOI22X1
XFILL_4__6888_ gnd vdd FILL
XFILL_2__7711_ gnd vdd FILL
X_10595_ _10595_/Q _9077_/CLK _7921_/R vdd _10527_/Y gnd vdd DFFSR
XFILL_5__7420_ gnd vdd FILL
XFILL_4__8627_ gnd vdd FILL
XFILL_1__9898_ gnd vdd FILL
X_12334_ _12331_/Y _12332_/Y _12334_/C gnd _12334_/Y vdd NAND3X1
X_15122_ _15122_/A gnd _15123_/B vdd INVX1
XFILL_4_BUFX2_insert1060 gnd vdd FILL
XFILL_3__10250_ gnd vdd FILL
XFILL_4_BUFX2_insert1071 gnd vdd FILL
XFILL_1__8849_ gnd vdd FILL
XFILL_2__10980_ gnd vdd FILL
XFILL_4_BUFX2_insert1093 gnd vdd FILL
XFILL_5__7351_ gnd vdd FILL
X_15053_ _16036_/A _13403_/Y _15321_/C _13402_/Y gnd _15057_/B vdd OAI22X1
X_12265_ _6882_/A _12249_/B _12249_/C _12801_/Q gnd _12266_/C vdd AOI22X1
XFILL_4__11540_ gnd vdd FILL
XFILL_3__10181_ gnd vdd FILL
XFILL_2__7573_ gnd vdd FILL
X_14004_ _9879_/A _13645_/C _14004_/C gnd _14012_/B vdd AOI21X1
XFILL_4__7509_ gnd vdd FILL
XFILL_1__11360_ gnd vdd FILL
X_11216_ _10896_/Y gnd _11216_/Y vdd INVX1
XFILL_4__8489_ gnd vdd FILL
XFILL_5__12830_ gnd vdd FILL
X_12196_ _13202_/Q gnd _12198_/A vdd INVX1
XFILL_2__12650_ gnd vdd FILL
XFILL_1__10311_ gnd vdd FILL
XFILL_4__11471_ gnd vdd FILL
XFILL_5__9021_ gnd vdd FILL
XFILL_1__11291_ gnd vdd FILL
XFILL_4__13210_ gnd vdd FILL
X_11147_ _12168_/Y gnd _11147_/Y vdd INVX1
XSFILL84200x15050 gnd vdd FILL
XFILL_4__10422_ gnd vdd FILL
XFILL_5__12761_ gnd vdd FILL
XFILL_2__11601_ gnd vdd FILL
XSFILL28920x83050 gnd vdd FILL
XFILL_4__14190_ gnd vdd FILL
XFILL_2__9243_ gnd vdd FILL
XFILL_1__13030_ gnd vdd FILL
XFILL_3__13940_ gnd vdd FILL
XFILL_2__12581_ gnd vdd FILL
XFILL_1__10242_ gnd vdd FILL
XFILL_3_BUFX2_insert360 gnd vdd FILL
XFILL_5__14500_ gnd vdd FILL
XFILL_0__13760_ gnd vdd FILL
XFILL_0__10972_ gnd vdd FILL
XFILL_5__11712_ gnd vdd FILL
XFILL_3_BUFX2_insert371 gnd vdd FILL
XFILL_4__13141_ gnd vdd FILL
X_15955_ _15949_/Y _15955_/B gnd _15955_/Y vdd NAND2X1
XFILL_2__14320_ gnd vdd FILL
X_11078_ _12250_/Y gnd _11078_/Y vdd INVX2
XFILL_5__15480_ gnd vdd FILL
XFILL_3_BUFX2_insert382 gnd vdd FILL
XFILL_3_BUFX2_insert393 gnd vdd FILL
XFILL_2__11532_ gnd vdd FILL
XFILL_3__13871_ gnd vdd FILL
XFILL_0__12711_ gnd vdd FILL
XFILL_1__10173_ gnd vdd FILL
X_10029_ _9993_/A _6957_/B gnd _10030_/C vdd NAND2X1
XFILL_0__13691_ gnd vdd FILL
X_14906_ _14906_/A _14905_/Y gnd _14907_/A vdd NAND2X1
XFILL_5__14431_ gnd vdd FILL
XFILL_2__8125_ gnd vdd FILL
XFILL_5__11643_ gnd vdd FILL
XFILL_3__15610_ gnd vdd FILL
XFILL_2__14251_ gnd vdd FILL
XFILL_4__10284_ gnd vdd FILL
X_15886_ _7658_/Q gnd _15886_/Y vdd INVX1
XFILL_0__15430_ gnd vdd FILL
XFILL_2__11463_ gnd vdd FILL
XFILL_0__12642_ gnd vdd FILL
XFILL_1__14981_ gnd vdd FILL
XFILL_5__9923_ gnd vdd FILL
XSFILL99480x69050 gnd vdd FILL
X_14837_ _14836_/Y _14567_/D gnd _14838_/C vdd NOR2X1
XFILL_4__12023_ gnd vdd FILL
XFILL_5__14362_ gnd vdd FILL
XSFILL99400x3050 gnd vdd FILL
XSFILL74120x67050 gnd vdd FILL
XFILL_2__8056_ gnd vdd FILL
XFILL_3__15541_ gnd vdd FILL
XFILL_2__10414_ gnd vdd FILL
XFILL_5__11574_ gnd vdd FILL
XFILL_2__14182_ gnd vdd FILL
XFILL_3__12753_ gnd vdd FILL
XFILL_1__13932_ gnd vdd FILL
XFILL_0__15361_ gnd vdd FILL
XFILL_5__16101_ gnd vdd FILL
XFILL_2__11394_ gnd vdd FILL
XFILL_5__13313_ gnd vdd FILL
XFILL_0__12573_ gnd vdd FILL
XFILL_5__9854_ gnd vdd FILL
XFILL_0__7071_ gnd vdd FILL
XFILL_5__10525_ gnd vdd FILL
XFILL_2__13133_ gnd vdd FILL
X_14768_ _14725_/A _14768_/B _14768_/C _14768_/D gnd _14772_/A vdd OAI22X1
XFILL_3__11704_ gnd vdd FILL
XFILL_5__14293_ gnd vdd FILL
XFILL_3__15472_ gnd vdd FILL
XFILL_0__14312_ gnd vdd FILL
XFILL_1__13863_ gnd vdd FILL
XFILL_0__11524_ gnd vdd FILL
XFILL_5__16032_ gnd vdd FILL
XFILL_0__15292_ gnd vdd FILL
XFILL_5__13244_ gnd vdd FILL
XFILL_5__9785_ gnd vdd FILL
X_13719_ _7173_/A _13434_/B _13883_/B _9435_/Q gnd _13719_/Y vdd AOI22X1
XSFILL53960x25050 gnd vdd FILL
XFILL_5__6997_ gnd vdd FILL
XFILL_3__14423_ gnd vdd FILL
XFILL_3__7820_ gnd vdd FILL
XFILL_4_CLKBUF1_insert150 gnd vdd FILL
X_14699_ _7748_/A gnd _14700_/B vdd INVX1
XFILL_3__11635_ gnd vdd FILL
XFILL_4__13974_ gnd vdd FILL
XFILL_1__15602_ gnd vdd FILL
XFILL_2__10276_ gnd vdd FILL
XFILL_0__14243_ gnd vdd FILL
XFILL_4_CLKBUF1_insert161 gnd vdd FILL
XFILL_1__13794_ gnd vdd FILL
XFILL_5__8736_ gnd vdd FILL
XFILL_4_CLKBUF1_insert172 gnd vdd FILL
XFILL_0__11455_ gnd vdd FILL
X_16438_ _16438_/Q _7261_/CLK _8669_/R vdd _16386_/Y gnd vdd DFFSR
XFILL_4__15713_ gnd vdd FILL
XSFILL13800x7050 gnd vdd FILL
XFILL_2__12015_ gnd vdd FILL
XFILL_4_CLKBUF1_insert183 gnd vdd FILL
XFILL_4_CLKBUF1_insert194 gnd vdd FILL
XFILL_1__15533_ gnd vdd FILL
XFILL_3__14354_ gnd vdd FILL
XFILL_5__10387_ gnd vdd FILL
XFILL_3__11566_ gnd vdd FILL
XFILL_0__10406_ gnd vdd FILL
XFILL_1__12745_ gnd vdd FILL
XSFILL18760x50 gnd vdd FILL
XFILL_2__8958_ gnd vdd FILL
XFILL_3__7751_ gnd vdd FILL
XFILL_0_BUFX2_insert250 gnd vdd FILL
XFILL_0__14174_ gnd vdd FILL
X_8320_ _8321_/B _9344_/B gnd _8320_/Y vdd NAND2X1
XFILL_5__12126_ gnd vdd FILL
XFILL_0_BUFX2_insert261 gnd vdd FILL
XFILL_0__11386_ gnd vdd FILL
XFILL_3__13305_ gnd vdd FILL
X_16369_ _14262_/A gnd _16369_/Y vdd INVX1
XFILL_0__7973_ gnd vdd FILL
XFILL_4__15644_ gnd vdd FILL
XFILL_3__10517_ gnd vdd FILL
XFILL_0_BUFX2_insert272 gnd vdd FILL
XFILL_0_BUFX2_insert283 gnd vdd FILL
XFILL_4__12856_ gnd vdd FILL
XFILL_0__13125_ gnd vdd FILL
XFILL_3__7682_ gnd vdd FILL
XFILL_0_BUFX2_insert294 gnd vdd FILL
XFILL_1__15464_ gnd vdd FILL
XFILL_3__11497_ gnd vdd FILL
XFILL_3__14285_ gnd vdd FILL
XFILL_2__8889_ gnd vdd FILL
XFILL_5__7618_ gnd vdd FILL
X_8251_ _8301_/Q gnd _8251_/Y vdd INVX1
XFILL_0__6924_ gnd vdd FILL
XFILL_3__16024_ gnd vdd FILL
XFILL_5__12057_ gnd vdd FILL
XFILL_5__8598_ gnd vdd FILL
XFILL_4__11807_ gnd vdd FILL
XFILL_3__13236_ gnd vdd FILL
XSFILL43880x77050 gnd vdd FILL
XFILL_3__9421_ gnd vdd FILL
XFILL_3__10448_ gnd vdd FILL
XFILL_4__15575_ gnd vdd FILL
XFILL_1__14415_ gnd vdd FILL
XFILL_4__12787_ gnd vdd FILL
XFILL_1__11627_ gnd vdd FILL
XFILL_1__15395_ gnd vdd FILL
XFILL_0__10268_ gnd vdd FILL
XFILL_2__13966_ gnd vdd FILL
XFILL_6__13347_ gnd vdd FILL
X_7202_ _7202_/A _7202_/B _7201_/Y gnd _7268_/D vdd OAI21X1
XFILL_5__7549_ gnd vdd FILL
XFILL_6__16135_ gnd vdd FILL
XFILL_5__11008_ gnd vdd FILL
XFILL_4__14526_ gnd vdd FILL
XFILL_0__6855_ gnd vdd FILL
XFILL_0__9643_ gnd vdd FILL
XFILL_2_BUFX2_insert10 gnd vdd FILL
XFILL_2__15705_ gnd vdd FILL
XFILL_3__13167_ gnd vdd FILL
X_8182_ _8278_/Q gnd _8182_/Y vdd INVX1
XFILL_4__11738_ gnd vdd FILL
XFILL_3__10379_ gnd vdd FILL
XFILL_3__9352_ gnd vdd FILL
XFILL_0__12007_ gnd vdd FILL
XFILL_1__14346_ gnd vdd FILL
XFILL_2__12917_ gnd vdd FILL
XSFILL48920x14050 gnd vdd FILL
XFILL_2_BUFX2_insert21 gnd vdd FILL
XFILL_1__11558_ gnd vdd FILL
XSFILL74200x47050 gnd vdd FILL
XFILL_2__13897_ gnd vdd FILL
XFILL_2_BUFX2_insert32 gnd vdd FILL
X_7133_ _7133_/Q _7147_/CLK _7133_/R vdd _7133_/D gnd vdd DFFSR
XFILL_2_BUFX2_insert43 gnd vdd FILL
XFILL_5__15816_ gnd vdd FILL
XFILL_4__14457_ gnd vdd FILL
XFILL_3__12118_ gnd vdd FILL
XFILL_2_BUFX2_insert54 gnd vdd FILL
XFILL_1__10509_ gnd vdd FILL
XFILL_2__15636_ gnd vdd FILL
XFILL_3__13098_ gnd vdd FILL
XFILL_2_BUFX2_insert65 gnd vdd FILL
XFILL_4__11669_ gnd vdd FILL
XFILL_2__12848_ gnd vdd FILL
XFILL_5__9219_ gnd vdd FILL
XFILL_3__9283_ gnd vdd FILL
XFILL_1__14277_ gnd vdd FILL
XFILL_2_BUFX2_insert76 gnd vdd FILL
XFILL_6__12229_ gnd vdd FILL
XFILL_1__11489_ gnd vdd FILL
XFILL_0__8525_ gnd vdd FILL
XFILL_4__13408_ gnd vdd FILL
XFILL_2_BUFX2_insert87 gnd vdd FILL
XSFILL49000x23050 gnd vdd FILL
XFILL_1__16016_ gnd vdd FILL
XFILL_2_BUFX2_insert98 gnd vdd FILL
XFILL_3__12049_ gnd vdd FILL
X_7064_ _7064_/A _8088_/B gnd _7065_/C vdd NAND2X1
XFILL_5__15747_ gnd vdd FILL
XFILL_5__12959_ gnd vdd FILL
XFILL_1__13228_ gnd vdd FILL
XFILL_4__14388_ gnd vdd FILL
XFILL_3__8234_ gnd vdd FILL
XFILL_2__12779_ gnd vdd FILL
XFILL_2__15567_ gnd vdd FILL
XFILL_0__13958_ gnd vdd FILL
XFILL_0__8456_ gnd vdd FILL
XSFILL109560x34050 gnd vdd FILL
XFILL_4__16127_ gnd vdd FILL
XFILL_4__13339_ gnd vdd FILL
XFILL_5__15678_ gnd vdd FILL
XFILL_2__14518_ gnd vdd FILL
XFILL_1__13159_ gnd vdd FILL
XFILL_0__12909_ gnd vdd FILL
XSFILL38840x66050 gnd vdd FILL
XFILL_2__15498_ gnd vdd FILL
XFILL112360x73050 gnd vdd FILL
XFILL_0__13889_ gnd vdd FILL
XFILL_3__7116_ gnd vdd FILL
XFILL_1__7180_ gnd vdd FILL
XFILL_5__14629_ gnd vdd FILL
XFILL_3__15808_ gnd vdd FILL
XFILL_0__8387_ gnd vdd FILL
XFILL_4__16058_ gnd vdd FILL
XSFILL54120x14050 gnd vdd FILL
XFILL_0__15628_ gnd vdd FILL
XFILL_3__8096_ gnd vdd FILL
XFILL_2__14449_ gnd vdd FILL
XFILL_4__15009_ gnd vdd FILL
XFILL_0__7338_ gnd vdd FILL
XFILL_3__15739_ gnd vdd FILL
X_7966_ _7955_/B _9246_/B gnd _7966_/Y vdd NAND2X1
XFILL_3__7047_ gnd vdd FILL
XFILL_0__15559_ gnd vdd FILL
X_9705_ _9647_/A _9705_/CLK _7649_/R vdd _9705_/D gnd vdd DFFSR
X_6917_ _6917_/A gnd _6919_/A vdd INVX1
XFILL_2__16119_ gnd vdd FILL
X_7897_ _7807_/A _8921_/CLK _9049_/R vdd _7897_/D gnd vdd DFFSR
XSFILL84920x50 gnd vdd FILL
XFILL_0__9008_ gnd vdd FILL
XFILL_4__7860_ gnd vdd FILL
X_9636_ _9615_/A _8868_/B gnd _9637_/C vdd NAND2X1
XSFILL18760x33050 gnd vdd FILL
XSFILL8600x43050 gnd vdd FILL
X_6848_ _6848_/A gnd memoryAddress[10] vdd BUFX2
XSFILL44040x66050 gnd vdd FILL
XFILL_3__8998_ gnd vdd FILL
XFILL_5_BUFX2_insert400 gnd vdd FILL
XFILL_5_BUFX2_insert411 gnd vdd FILL
X_9567_ _9567_/Q _9194_/CLK _9460_/R vdd _9491_/Y gnd vdd DFFSR
XFILL_4__9530_ gnd vdd FILL
XFILL_5_BUFX2_insert422 gnd vdd FILL
XFILL_3__7949_ gnd vdd FILL
XFILL_5_BUFX2_insert433 gnd vdd FILL
XFILL_5_BUFX2_insert444 gnd vdd FILL
X_8518_ _8518_/A _8460_/A _8518_/C gnd _8560_/D vdd OAI21X1
XFILL_1__9752_ gnd vdd FILL
XFILL_5_BUFX2_insert455 gnd vdd FILL
XSFILL23880x24050 gnd vdd FILL
XFILL_5_BUFX2_insert466 gnd vdd FILL
X_9498_ _9570_/Q gnd _9500_/A vdd INVX1
XFILL_1__6964_ gnd vdd FILL
XFILL_5_BUFX2_insert477 gnd vdd FILL
X_10380_ _10423_/B _9100_/B gnd _10381_/C vdd NAND2X1
XFILL_1__8703_ gnd vdd FILL
XFILL_5_BUFX2_insert488 gnd vdd FILL
X_8449_ _8447_/Y _8508_/A _8449_/C gnd _8537_/D vdd OAI21X1
XFILL_5_BUFX2_insert499 gnd vdd FILL
XSFILL38920x46050 gnd vdd FILL
XFILL_1__9683_ gnd vdd FILL
XFILL_1__6895_ gnd vdd FILL
XFILL_3__9619_ gnd vdd FILL
XFILL112440x53050 gnd vdd FILL
XSFILL64200x79050 gnd vdd FILL
XFILL_4__9392_ gnd vdd FILL
XFILL_1__8634_ gnd vdd FILL
XFILL_4__8343_ gnd vdd FILL
X_12050_ _12047_/Y _12050_/B _12049_/Y gnd _12050_/Y vdd NAND3X1
XSFILL39000x55050 gnd vdd FILL
X_11001_ _11013_/B gnd _11002_/B vdd INVX1
XFILL_4__8274_ gnd vdd FILL
XFILL_1__8496_ gnd vdd FILL
XFILL_4__7225_ gnd vdd FILL
XSFILL18840x13050 gnd vdd FILL
XSFILL94280x74050 gnd vdd FILL
XFILL_1__7447_ gnd vdd FILL
XFILL_2_BUFX2_insert301 gnd vdd FILL
XFILL_2_BUFX2_insert312 gnd vdd FILL
X_15740_ _15739_/Y _15740_/B _15740_/C gnd _15746_/B vdd NAND3X1
XFILL_2_BUFX2_insert323 gnd vdd FILL
XSFILL69080x50050 gnd vdd FILL
X_12952_ _12952_/A vdd gnd _12953_/C vdd NAND2X1
XFILL_2_BUFX2_insert334 gnd vdd FILL
XSFILL99320x11050 gnd vdd FILL
XFILL_2_BUFX2_insert345 gnd vdd FILL
XFILL_1__7378_ gnd vdd FILL
XFILL_2_BUFX2_insert356 gnd vdd FILL
XFILL_4__7087_ gnd vdd FILL
X_11903_ _11900_/A _12454_/A gnd _11903_/Y vdd NAND2X1
XFILL_2_BUFX2_insert367 gnd vdd FILL
X_15671_ _10531_/A gnd _15672_/D vdd INVX1
XFILL_2_BUFX2_insert378 gnd vdd FILL
XFILL_1__9117_ gnd vdd FILL
XFILL_2_BUFX2_insert389 gnd vdd FILL
XSFILL48760x49050 gnd vdd FILL
X_12883_ _12176_/B gnd _12883_/Y vdd INVX1
XFILL_5__6920_ gnd vdd FILL
XSFILL23800x2050 gnd vdd FILL
X_14622_ _9454_/Q gnd _14622_/Y vdd INVX1
X_11834_ _11834_/A _11834_/B gnd _11841_/B vdd NAND2X1
XFILL_2__9930_ gnd vdd FILL
XSFILL49640x77050 gnd vdd FILL
XFILL_5__10310_ gnd vdd FILL
XFILL_5__6851_ gnd vdd FILL
X_14553_ _10683_/A gnd _14553_/Y vdd INVX1
X_11765_ _11383_/A _11732_/B _11846_/C _11254_/Y gnd _11765_/Y vdd AOI22X1
XFILL_5__11290_ gnd vdd FILL
XFILL_2__10130_ gnd vdd FILL
XBUFX2_insert300 _12414_/Y gnd _9532_/B vdd BUFX2
XSFILL89240x63050 gnd vdd FILL
XFILL_2__9861_ gnd vdd FILL
XBUFX2_insert311 _11222_/Y gnd _11573_/C vdd BUFX2
XBUFX2_insert322 _13345_/Y gnd _9917_/B vdd BUFX2
X_10716_ _10716_/Q _7662_/CLK _9454_/R vdd _10634_/Y gnd vdd DFFSR
X_13504_ _13503_/Y _13489_/Y gnd _13504_/Y vdd NOR2X1
XFILL_4__7989_ gnd vdd FILL
XFILL_5__10241_ gnd vdd FILL
XFILL_3__11420_ gnd vdd FILL
XBUFX2_insert333 _12405_/Y gnd _9011_/B vdd BUFX2
X_14484_ _8811_/Q gnd _14484_/Y vdd INVX1
XBUFX2_insert344 _12396_/Y gnd _8874_/B vdd BUFX2
X_11696_ _11046_/Y _11676_/B _11835_/C gnd _11696_/Y vdd AOI21X1
XFILL_4__10971_ gnd vdd FILL
XFILL_2__10061_ gnd vdd FILL
XSFILL3720x66050 gnd vdd FILL
XFILL_2__9792_ gnd vdd FILL
XFILL_4__9728_ gnd vdd FILL
XBUFX2_insert355 _13306_/Y gnd _7970_/B vdd BUFX2
XFILL_5__8521_ gnd vdd FILL
XFILL_0__11240_ gnd vdd FILL
X_16223_ _15169_/A _14860_/Y _16222_/Y _16002_/A gnd _16226_/B vdd OAI22X1
XFILL_1__10791_ gnd vdd FILL
XBUFX2_insert366 _13487_/Y gnd _14909_/C vdd BUFX2
XFILL_4__12710_ gnd vdd FILL
XFILL_5_CLKBUF1_insert201 gnd vdd FILL
X_13435_ _13423_/A _13404_/B _13718_/B gnd _13435_/Y vdd NAND3X1
X_10647_ _10647_/A gnd _10649_/A vdd INVX1
XBUFX2_insert377 _12211_/Y gnd _12239_/C vdd BUFX2
XFILL_5__10172_ gnd vdd FILL
XBUFX2_insert388 _13331_/Y gnd _9101_/B vdd BUFX2
XFILL_5_CLKBUF1_insert212 gnd vdd FILL
XFILL_3__11351_ gnd vdd FILL
XFILL_5_CLKBUF1_insert223 gnd vdd FILL
XSFILL28920x78050 gnd vdd FILL
XFILL_2__8743_ gnd vdd FILL
XFILL_1__12530_ gnd vdd FILL
XBUFX2_insert399 _13293_/Y gnd _7570_/A vdd BUFX2
XFILL_4__13690_ gnd vdd FILL
XSFILL94360x54050 gnd vdd FILL
XFILL_0__11171_ gnd vdd FILL
XFILL_4__9659_ gnd vdd FILL
XFILL_5__8452_ gnd vdd FILL
XFILL_3__10302_ gnd vdd FILL
X_13366_ _12808_/Q gnd _13371_/B vdd INVX1
X_16154_ _14748_/Y _15940_/B _15802_/D _14784_/Y gnd _16156_/A vdd OAI22X1
XFILL_4__12641_ gnd vdd FILL
XFILL_5__14980_ gnd vdd FILL
XFILL_3__14070_ gnd vdd FILL
X_10578_ _10578_/A _10548_/B _10577_/Y gnd _10578_/Y vdd OAI21X1
XFILL_2__13820_ gnd vdd FILL
XFILL_0__10122_ gnd vdd FILL
XFILL_3__11282_ gnd vdd FILL
XFILL_1__12461_ gnd vdd FILL
XFILL_6__10413_ gnd vdd FILL
XSFILL69160x30050 gnd vdd FILL
X_15105_ _9815_/Q gnd _15106_/B vdd INVX1
XFILL_3__13021_ gnd vdd FILL
XFILL_5__8383_ gnd vdd FILL
XFILL_5__13931_ gnd vdd FILL
X_12317_ _6895_/A _12237_/B _12269_/C _12308_/B gnd _12318_/C vdd AOI22X1
X_13297_ _13297_/A _13296_/Y _13297_/C gnd _13297_/Y vdd NOR3X1
XFILL_1__14200_ gnd vdd FILL
XFILL_4__15360_ gnd vdd FILL
XFILL_3__10233_ gnd vdd FILL
X_16085_ _16085_/A _16085_/B _16085_/C gnd _16086_/B vdd NAND3X1
XFILL_4__12572_ gnd vdd FILL
XFILL_2__7625_ gnd vdd FILL
XFILL_1__11412_ gnd vdd FILL
XFILL_1__15180_ gnd vdd FILL
XFILL_2__10963_ gnd vdd FILL
XFILL_2__13751_ gnd vdd FILL
XFILL_0__14930_ gnd vdd FILL
XFILL_0__10053_ gnd vdd FILL
XFILL_1__12392_ gnd vdd FILL
XFILL_5__7334_ gnd vdd FILL
X_15036_ _15036_/A _12767_/A gnd _15037_/C vdd NOR2X1
X_12248_ _12248_/A _12719_/A _12248_/C gnd _12250_/B vdd NAND3X1
XSFILL48840x29050 gnd vdd FILL
XFILL_4__14311_ gnd vdd FILL
XFILL_5__13862_ gnd vdd FILL
XFILL_4__11523_ gnd vdd FILL
XFILL_2__12702_ gnd vdd FILL
XFILL_1__14131_ gnd vdd FILL
XFILL_3__10164_ gnd vdd FILL
XFILL_4__15291_ gnd vdd FILL
XFILL_2__13682_ gnd vdd FILL
XFILL_2__7556_ gnd vdd FILL
XFILL_1__11343_ gnd vdd FILL
XFILL_0__14861_ gnd vdd FILL
XFILL_2__10894_ gnd vdd FILL
XFILL_5__15601_ gnd vdd FILL
XSFILL74280x21050 gnd vdd FILL
XFILL_4__14242_ gnd vdd FILL
X_12179_ _12179_/A _12886_/A gnd _12180_/C vdd NAND2X1
XFILL_2__12633_ gnd vdd FILL
XFILL_5__13793_ gnd vdd FILL
XFILL_4__11454_ gnd vdd FILL
XFILL_2__15421_ gnd vdd FILL
XFILL_0__13812_ gnd vdd FILL
XFILL_2__7487_ gnd vdd FILL
XFILL_1__14062_ gnd vdd FILL
XFILL_5__9004_ gnd vdd FILL
XFILL_3__14972_ gnd vdd FILL
XFILL_6__12014_ gnd vdd FILL
XFILL_0__8310_ gnd vdd FILL
XFILL_1__11274_ gnd vdd FILL
XFILL_0__14792_ gnd vdd FILL
XFILL_5__15532_ gnd vdd FILL
XFILL_5__7196_ gnd vdd FILL
XSFILL59080x82050 gnd vdd FILL
XFILL_5__12744_ gnd vdd FILL
XFILL_4__10405_ gnd vdd FILL
XSFILL89320x43050 gnd vdd FILL
XFILL_0__9290_ gnd vdd FILL
XFILL_4__14173_ gnd vdd FILL
XFILL_2__9226_ gnd vdd FILL
XFILL_3__13923_ gnd vdd FILL
XFILL_1__13013_ gnd vdd FILL
XFILL_2__15352_ gnd vdd FILL
XFILL_4__11385_ gnd vdd FILL
XFILL_0__13743_ gnd vdd FILL
XSFILL109480x49050 gnd vdd FILL
XFILL_0__10955_ gnd vdd FILL
XFILL_0__8241_ gnd vdd FILL
XFILL_4__13124_ gnd vdd FILL
X_15938_ _8760_/A _15821_/B _15937_/Y gnd _15942_/C vdd AOI21X1
XFILL_5__15463_ gnd vdd FILL
XFILL_2__14303_ gnd vdd FILL
XFILL_2__11515_ gnd vdd FILL
XFILL_3__13854_ gnd vdd FILL
XFILL_2__9157_ gnd vdd FILL
XFILL_2__15283_ gnd vdd FILL
XFILL_2__12495_ gnd vdd FILL
XFILL_1__10156_ gnd vdd FILL
XSFILL54040x29050 gnd vdd FILL
XFILL_0__13674_ gnd vdd FILL
XFILL_5__14414_ gnd vdd FILL
X_7820_ _7887_/B _7948_/B gnd _7821_/C vdd NAND2X1
XFILL_6__6960_ gnd vdd FILL
XFILL_0__10886_ gnd vdd FILL
XFILL_5__11626_ gnd vdd FILL
XFILL_5__15394_ gnd vdd FILL
XFILL_2__14234_ gnd vdd FILL
X_15869_ _15632_/A _15869_/B _15869_/C gnd _15871_/A vdd OAI21X1
XFILL_2__8108_ gnd vdd FILL
XFILL_2__9088_ gnd vdd FILL
XFILL_0__15413_ gnd vdd FILL
XFILL_4__10267_ gnd vdd FILL
XFILL_2__11446_ gnd vdd FILL
XFILL_2_BUFX2_insert890 gnd vdd FILL
XFILL_0__12625_ gnd vdd FILL
XFILL_3__13785_ gnd vdd FILL
XSFILL68600x44050 gnd vdd FILL
XFILL_5__9906_ gnd vdd FILL
XFILL_0__16393_ gnd vdd FILL
XFILL_0__7123_ gnd vdd FILL
XFILL_1__14964_ gnd vdd FILL
XFILL_3__10997_ gnd vdd FILL
XFILL_4__12006_ gnd vdd FILL
XFILL_5__14345_ gnd vdd FILL
XFILL_3__15524_ gnd vdd FILL
XFILL_5__11557_ gnd vdd FILL
X_7751_ _7751_/A gnd _7753_/A vdd INVX1
XFILL_3__12736_ gnd vdd FILL
XFILL_2__14165_ gnd vdd FILL
XSFILL69240x10050 gnd vdd FILL
XFILL_0__15344_ gnd vdd FILL
XFILL_1__13915_ gnd vdd FILL
XFILL_2__11377_ gnd vdd FILL
XFILL_1__14895_ gnd vdd FILL
XFILL_0__7054_ gnd vdd FILL
XFILL_5__10508_ gnd vdd FILL
XFILL_2__13116_ gnd vdd FILL
XFILL_5__14276_ gnd vdd FILL
X_7682_ _7682_/A gnd _7682_/Y vdd INVX1
XFILL_4_BUFX2_insert0 gnd vdd FILL
XFILL_3__15455_ gnd vdd FILL
XFILL_5__11488_ gnd vdd FILL
XFILL_1__13846_ gnd vdd FILL
XSFILL18680x48050 gnd vdd FILL
XFILL_3__8852_ gnd vdd FILL
XFILL_0__11507_ gnd vdd FILL
XFILL_2__14096_ gnd vdd FILL
XFILL_5__16015_ gnd vdd FILL
XFILL_0__15275_ gnd vdd FILL
XFILL_5__9768_ gnd vdd FILL
XFILL_5__13227_ gnd vdd FILL
X_9421_ _9459_/Q gnd _9421_/Y vdd INVX1
XFILL_0__12487_ gnd vdd FILL
XSFILL58280x34050 gnd vdd FILL
XFILL_5__10439_ gnd vdd FILL
XFILL_3__14406_ gnd vdd FILL
XFILL_3__7803_ gnd vdd FILL
XFILL_4__13957_ gnd vdd FILL
XFILL_3__11618_ gnd vdd FILL
XFILL_3__15386_ gnd vdd FILL
XFILL_0__14226_ gnd vdd FILL
XFILL_2__10259_ gnd vdd FILL
XFILL_5__8719_ gnd vdd FILL
XFILL_3__8783_ gnd vdd FILL
XFILL_3__12598_ gnd vdd FILL
XFILL_1__13777_ gnd vdd FILL
XFILL_0__11438_ gnd vdd FILL
XFILL_1__10989_ gnd vdd FILL
X_9352_ _9352_/A gnd _9354_/A vdd INVX1
XFILL_4__12908_ gnd vdd FILL
XFILL_5__13158_ gnd vdd FILL
XSFILL49000x18050 gnd vdd FILL
XFILL_3__14337_ gnd vdd FILL
XFILL_1__12728_ gnd vdd FILL
XFILL_3__7734_ gnd vdd FILL
XFILL_1__15516_ gnd vdd FILL
XFILL_3__11549_ gnd vdd FILL
XFILL_4__13888_ gnd vdd FILL
XFILL_0__14157_ gnd vdd FILL
XFILL_5__12109_ gnd vdd FILL
X_8303_ _8303_/Q _7651_/CLK _7011_/R vdd _8303_/D gnd vdd DFFSR
XFILL_0__11369_ gnd vdd FILL
XFILL_4__15627_ gnd vdd FILL
XSFILL109560x29050 gnd vdd FILL
XFILL_4_BUFX2_insert407 gnd vdd FILL
XFILL_5__13089_ gnd vdd FILL
X_9283_ _9281_/Y _9282_/A _9283_/C gnd _9283_/Y vdd OAI21X1
XFILL_0__7956_ gnd vdd FILL
XFILL_4__12839_ gnd vdd FILL
XFILL_0__13108_ gnd vdd FILL
XFILL_3__14268_ gnd vdd FILL
XFILL_4_BUFX2_insert418 gnd vdd FILL
XFILL_1__12659_ gnd vdd FILL
XFILL_1__15447_ gnd vdd FILL
XFILL111880x61050 gnd vdd FILL
XFILL_2__14998_ gnd vdd FILL
XFILL_4_BUFX2_insert429 gnd vdd FILL
XFILL_0__14088_ gnd vdd FILL
XFILL112360x68050 gnd vdd FILL
XFILL_3__16007_ gnd vdd FILL
XFILL_0__6907_ gnd vdd FILL
X_8234_ _8237_/A _7594_/B gnd _8235_/C vdd NAND2X1
XFILL_3__13219_ gnd vdd FILL
XFILL_3__9404_ gnd vdd FILL
XFILL_4__15558_ gnd vdd FILL
XFILL_0__7887_ gnd vdd FILL
XSFILL109160x31050 gnd vdd FILL
XFILL_3__14199_ gnd vdd FILL
XFILL_1__15378_ gnd vdd FILL
XFILL_0__13039_ gnd vdd FILL
XFILL_2__13949_ gnd vdd FILL
XFILL_3__7596_ gnd vdd FILL
XFILL_4__14509_ gnd vdd FILL
XFILL_0__9626_ gnd vdd FILL
X_8165_ _8165_/Q _8165_/CLK _8165_/R vdd _8101_/Y gnd vdd DFFSR
XFILL_0__6838_ gnd vdd FILL
XSFILL79080x13050 gnd vdd FILL
XFILL_3__9335_ gnd vdd FILL
XFILL_4__15489_ gnd vdd FILL
XFILL_1__14329_ gnd vdd FILL
X_7116_ _7116_/A _7055_/A _7116_/C gnd _7154_/D vdd OAI21X1
XSFILL79320x75050 gnd vdd FILL
XFILL_1__8350_ gnd vdd FILL
XFILL_0__9557_ gnd vdd FILL
XFILL_2__15619_ gnd vdd FILL
X_8096_ _8096_/A gnd _8098_/A vdd INVX1
XFILL_3__9266_ gnd vdd FILL
XFILL_1__7301_ gnd vdd FILL
XFILL_0__8508_ gnd vdd FILL
XSFILL18760x28050 gnd vdd FILL
X_7047_ _7045_/Y _7067_/A _7046_/Y gnd _7131_/D vdd OAI21X1
XFILL_0__9488_ gnd vdd FILL
XFILL_3__8217_ gnd vdd FILL
XSFILL8600x38050 gnd vdd FILL
XFILL_1__7232_ gnd vdd FILL
XFILL_0__8439_ gnd vdd FILL
XFILL_3__8148_ gnd vdd FILL
XFILL_1__7163_ gnd vdd FILL
XFILL_3__8079_ gnd vdd FILL
X_8998_ _9062_/Q gnd _8998_/Y vdd INVX1
XFILL_1_BUFX2_insert308 gnd vdd FILL
XFILL_4__8961_ gnd vdd FILL
XFILL_1_BUFX2_insert319 gnd vdd FILL
X_7949_ _7947_/Y _7948_/A _7948_/Y gnd _8029_/D vdd OAI21X1
XFILL_1__7094_ gnd vdd FILL
XFILL112440x48050 gnd vdd FILL
XFILL_4__8892_ gnd vdd FILL
XSFILL23720x83050 gnd vdd FILL
XFILL_4__7843_ gnd vdd FILL
X_11550_ _11550_/A _11637_/B _11550_/C gnd _11551_/A vdd AOI21X1
XFILL_6__8759_ gnd vdd FILL
X_9619_ _9617_/Y _9652_/B _9619_/C gnd _9695_/D vdd OAI21X1
X_10501_ _10501_/A gnd _10503_/A vdd INVX1
XFILL_1__9804_ gnd vdd FILL
XFILL_5_BUFX2_insert230 gnd vdd FILL
X_11481_ _11415_/C _11480_/Y _11461_/C gnd _11481_/Y vdd NAND3X1
XFILL_5_BUFX2_insert241 gnd vdd FILL
XSFILL3720x9050 gnd vdd FILL
XFILL_4__9513_ gnd vdd FILL
X_13220_ _13220_/A gnd _13266_/A vdd INVX2
XFILL_1__7996_ gnd vdd FILL
XFILL_5_BUFX2_insert252 gnd vdd FILL
X_10432_ _10432_/A _10405_/B _10432_/C gnd _10432_/Y vdd OAI21X1
XFILL_5_BUFX2_insert263 gnd vdd FILL
XSFILL114600x64050 gnd vdd FILL
XFILL_5_BUFX2_insert274 gnd vdd FILL
XFILL_5_BUFX2_insert285 gnd vdd FILL
XFILL_1__9735_ gnd vdd FILL
XFILL_1__6947_ gnd vdd FILL
XFILL_5_BUFX2_insert296 gnd vdd FILL
X_13151_ _11959_/A gnd _13151_/Y vdd INVX1
X_10363_ _10363_/A _10363_/B _10362_/Y gnd _10363_/Y vdd OAI21X1
XFILL_4_BUFX2_insert930 gnd vdd FILL
XFILL_1__9666_ gnd vdd FILL
XFILL_4_BUFX2_insert941 gnd vdd FILL
X_12102_ _12102_/A _12102_/B _12102_/C gnd _13164_/B vdd NAND3X1
XFILL_1__6878_ gnd vdd FILL
XFILL_4_BUFX2_insert952 gnd vdd FILL
XFILL_4_BUFX2_insert963 gnd vdd FILL
XFILL_4__9375_ gnd vdd FILL
X_13082_ _11890_/A gnd _13082_/Y vdd INVX1
XFILL_1__8617_ gnd vdd FILL
X_10294_ _10294_/A _7222_/B gnd _10295_/C vdd NAND2X1
XFILL_4_BUFX2_insert974 gnd vdd FILL
XFILL_2__8390_ gnd vdd FILL
XFILL_4_BUFX2_insert985 gnd vdd FILL
XFILL_4_BUFX2_insert996 gnd vdd FILL
XFILL_1__9597_ gnd vdd FILL
XFILL_4__8326_ gnd vdd FILL
X_12033_ _12473_/B _12025_/B _12025_/C gnd gnd _12033_/Y vdd AOI22X1
XFILL_2__7341_ gnd vdd FILL
XFILL_5__7050_ gnd vdd FILL
XFILL_4__8257_ gnd vdd FILL
XFILL_5__10790_ gnd vdd FILL
XSFILL89240x58050 gnd vdd FILL
XFILL_4__7208_ gnd vdd FILL
XFILL_1__8479_ gnd vdd FILL
XSFILL18760x9050 gnd vdd FILL
XFILL112120x30050 gnd vdd FILL
XFILL_4__8188_ gnd vdd FILL
XFILL_4__11170_ gnd vdd FILL
XFILL_2__9011_ gnd vdd FILL
XFILL_3__10920_ gnd vdd FILL
X_13984_ _9751_/A gnd _13985_/A vdd INVX1
XFILL_1__10010_ gnd vdd FILL
X_15723_ _9766_/A gnd _15724_/D vdd INVX1
XFILL_4__10121_ gnd vdd FILL
XFILL_5__12460_ gnd vdd FILL
X_12935_ _12871_/A _7532_/CLK _8816_/R vdd _12935_/D gnd vdd DFFSR
XFILL_2__11300_ gnd vdd FILL
XFILL_2__12280_ gnd vdd FILL
XSFILL94360x49050 gnd vdd FILL
XSFILL43720x14050 gnd vdd FILL
XFILL_5__7952_ gnd vdd FILL
XFILL_0__10671_ gnd vdd FILL
XFILL_5__11411_ gnd vdd FILL
X_15654_ _15654_/A _15169_/D gnd _15658_/A vdd NOR2X1
XFILL_4__10052_ gnd vdd FILL
XFILL_5__12391_ gnd vdd FILL
X_12866_ vdd _12866_/B gnd _12867_/C vdd NAND2X1
XFILL_1_BUFX2_insert820 gnd vdd FILL
XFILL_2__11231_ gnd vdd FILL
XFILL_0__12410_ gnd vdd FILL
XFILL_1_BUFX2_insert831 gnd vdd FILL
XFILL_3__10782_ gnd vdd FILL
XFILL_3__13570_ gnd vdd FILL
XFILL_1__11961_ gnd vdd FILL
XFILL_5__6903_ gnd vdd FILL
XFILL_1_BUFX2_insert842 gnd vdd FILL
XFILL_1_BUFX2_insert853 gnd vdd FILL
X_14605_ _8430_/Q _13848_/B _13592_/A _8254_/A gnd _14607_/A vdd AOI22X1
XFILL_5__14130_ gnd vdd FILL
XFILL_0__13390_ gnd vdd FILL
XSFILL69160x25050 gnd vdd FILL
XFILL_5__7883_ gnd vdd FILL
XFILL_5__11342_ gnd vdd FILL
X_11817_ _11005_/Y _11816_/Y _11835_/C gnd _11818_/C vdd AOI21X1
XFILL_4__14860_ gnd vdd FILL
XFILL_1_BUFX2_insert864 gnd vdd FILL
XFILL_3__12521_ gnd vdd FILL
XFILL_2__9913_ gnd vdd FILL
XFILL_1__13700_ gnd vdd FILL
X_15585_ _15585_/A _15585_/B _15582_/Y gnd _15586_/A vdd NAND3X1
XFILL_1__10912_ gnd vdd FILL
X_12797_ _12713_/A _7005_/CLK _12799_/R vdd _12797_/D gnd vdd DFFSR
XFILL_1_BUFX2_insert875 gnd vdd FILL
XFILL_2__11162_ gnd vdd FILL
XFILL_1_BUFX2_insert886 gnd vdd FILL
XFILL_0__12341_ gnd vdd FILL
XFILL_1__14680_ gnd vdd FILL
XFILL_5__9622_ gnd vdd FILL
XFILL_1_BUFX2_insert897 gnd vdd FILL
XFILL_1__11892_ gnd vdd FILL
XSFILL7960x66050 gnd vdd FILL
XFILL_4__13811_ gnd vdd FILL
XFILL_5__14061_ gnd vdd FILL
X_14536_ _14536_/A _14536_/B gnd _14537_/C vdd NOR2X1
XFILL_2__10113_ gnd vdd FILL
XFILL_3__15240_ gnd vdd FILL
XSFILL104360x34050 gnd vdd FILL
XFILL_5__11273_ gnd vdd FILL
X_11748_ _11748_/A _11270_/Y _11682_/B gnd _11748_/Y vdd OAI21X1
XFILL_1__13631_ gnd vdd FILL
XFILL_3__12452_ gnd vdd FILL
XFILL_4__14791_ gnd vdd FILL
XFILL_2__15970_ gnd vdd FILL
XFILL_0__15060_ gnd vdd FILL
XFILL_2__11093_ gnd vdd FILL
XFILL_0__12272_ gnd vdd FILL
XFILL_5__9553_ gnd vdd FILL
XFILL_5__13012_ gnd vdd FILL
XSFILL74280x16050 gnd vdd FILL
X_14467_ _14466_/Y _14467_/B gnd _14467_/Y vdd NOR2X1
XFILL_4__13742_ gnd vdd FILL
XFILL_3__11403_ gnd vdd FILL
XFILL_4__10954_ gnd vdd FILL
XFILL_2__10044_ gnd vdd FILL
XFILL_3__15171_ gnd vdd FILL
XFILL_3__12383_ gnd vdd FILL
XFILL_0__14011_ gnd vdd FILL
XFILL_2__14921_ gnd vdd FILL
XSFILL79320x2050 gnd vdd FILL
X_11679_ _11045_/Y _11678_/A _11835_/C gnd _11679_/Y vdd AOI21X1
XFILL_1__16350_ gnd vdd FILL
XFILL_5__8504_ gnd vdd FILL
XFILL_2__9775_ gnd vdd FILL
XFILL_1__13562_ gnd vdd FILL
XFILL_0__11223_ gnd vdd FILL
X_16206_ _15922_/C _14871_/Y _15972_/C _14836_/Y gnd _16209_/B vdd OAI22X1
XFILL_2__6987_ gnd vdd FILL
XFILL_1__10774_ gnd vdd FILL
XFILL_5__9484_ gnd vdd FILL
XFILL_0__7810_ gnd vdd FILL
XSFILL105240x62050 gnd vdd FILL
X_13418_ _13418_/A _13377_/Y gnd _13418_/Y vdd NAND2X1
XSFILL59080x77050 gnd vdd FILL
XSFILL89320x38050 gnd vdd FILL
XFILL_5__10155_ gnd vdd FILL
XFILL_3__14122_ gnd vdd FILL
XFILL_1__12513_ gnd vdd FILL
XFILL_1__15301_ gnd vdd FILL
XFILL_4__13673_ gnd vdd FILL
X_14398_ _10671_/A _14868_/A _14214_/C _15846_/A gnd _14400_/A vdd AOI22X1
XFILL_2__8726_ gnd vdd FILL
XFILL112200x10050 gnd vdd FILL
XFILL_3__11334_ gnd vdd FILL
XFILL_2__14852_ gnd vdd FILL
XFILL_4__10885_ gnd vdd FILL
XFILL_1__16281_ gnd vdd FILL
XSFILL99480x82050 gnd vdd FILL
XFILL_0__11154_ gnd vdd FILL
XFILL_1__13493_ gnd vdd FILL
XFILL_4__15412_ gnd vdd FILL
X_16137_ _16137_/A _15025_/B _16137_/C _16135_/Y gnd _16137_/Y vdd OAI22X1
XFILL_0__7741_ gnd vdd FILL
X_13349_ _13341_/Y gnd _13350_/C vdd INVX1
XFILL_4__12624_ gnd vdd FILL
XFILL_2__13803_ gnd vdd FILL
XFILL_1__15232_ gnd vdd FILL
XFILL_3__14053_ gnd vdd FILL
XFILL_5__14963_ gnd vdd FILL
XFILL_4__16392_ gnd vdd FILL
XFILL_3__11265_ gnd vdd FILL
XFILL_3__7450_ gnd vdd FILL
XFILL_1__12444_ gnd vdd FILL
XFILL_0__10105_ gnd vdd FILL
XFILL_2__8657_ gnd vdd FILL
XFILL_2__11995_ gnd vdd FILL
XFILL_0__15962_ gnd vdd FILL
XFILL_0__11085_ gnd vdd FILL
XFILL_2__14783_ gnd vdd FILL
XFILL_5__8366_ gnd vdd FILL
XFILL_4__15343_ gnd vdd FILL
XFILL_0__7672_ gnd vdd FILL
XSFILL79800x8050 gnd vdd FILL
X_16068_ _10305_/A _15863_/A gnd _16075_/A vdd NAND2X1
XFILL_5__13914_ gnd vdd FILL
XFILL_3__13004_ gnd vdd FILL
XSFILL53800x79050 gnd vdd FILL
XFILL_2__7608_ gnd vdd FILL
XSFILL94440x29050 gnd vdd FILL
XFILL_5__14894_ gnd vdd FILL
XFILL_3__7381_ gnd vdd FILL
XFILL_1__15163_ gnd vdd FILL
XFILL_2__13734_ gnd vdd FILL
XFILL_3__11196_ gnd vdd FILL
XFILL_2__8588_ gnd vdd FILL
XFILL_2__10946_ gnd vdd FILL
XFILL_6__13115_ gnd vdd FILL
XFILL_1__12375_ gnd vdd FILL
XFILL_0__10036_ gnd vdd FILL
XFILL_5__7317_ gnd vdd FILL
XFILL_0__14913_ gnd vdd FILL
XFILL_0__15893_ gnd vdd FILL
X_15019_ _15313_/B _16037_/B _14981_/Y gnd _15019_/Y vdd NAND3X1
XFILL_0__9411_ gnd vdd FILL
XFILL_4__11506_ gnd vdd FILL
XFILL_5__13845_ gnd vdd FILL
XFILL_3__9120_ gnd vdd FILL
XFILL_3__10147_ gnd vdd FILL
XFILL_1__14114_ gnd vdd FILL
XFILL_4__15274_ gnd vdd FILL
XFILL_4__12486_ gnd vdd FILL
XFILL_1__11326_ gnd vdd FILL
XFILL_0__14844_ gnd vdd FILL
XFILL_2__13665_ gnd vdd FILL
XFILL_2__10877_ gnd vdd FILL
XFILL_1__15094_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1075 gnd vdd FILL
XFILL_5__7248_ gnd vdd FILL
XFILL_4__14225_ gnd vdd FILL
XFILL_0__9342_ gnd vdd FILL
XFILL_2__15404_ gnd vdd FILL
XFILL_5__13776_ gnd vdd FILL
X_9970_ _9970_/Q _8562_/CLK _7270_/R vdd _9970_/D gnd vdd DFFSR
XFILL_4__11437_ gnd vdd FILL
XFILL_2__12616_ gnd vdd FILL
XFILL_1__14045_ gnd vdd FILL
XFILL_5__10988_ gnd vdd FILL
XFILL_3__14955_ gnd vdd FILL
XFILL_2__16384_ gnd vdd FILL
XFILL_1__11257_ gnd vdd FILL
XFILL_2__13596_ gnd vdd FILL
XSFILL104440x14050 gnd vdd FILL
XFILL_0__14775_ gnd vdd FILL
X_8921_ _8831_/A _8921_/CLK _8942_/R vdd _8833_/Y gnd vdd DFFSR
XFILL_5__7179_ gnd vdd FILL
XFILL_5__12727_ gnd vdd FILL
XFILL_0__11987_ gnd vdd FILL
XFILL_0__9273_ gnd vdd FILL
XFILL_5__15515_ gnd vdd FILL
XFILL_4__14156_ gnd vdd FILL
XFILL_3__8002_ gnd vdd FILL
XFILL_3__13906_ gnd vdd FILL
XFILL_2__9209_ gnd vdd FILL
XFILL_2__15335_ gnd vdd FILL
XSFILL8680x12050 gnd vdd FILL
XFILL_4__11368_ gnd vdd FILL
XFILL_0__13726_ gnd vdd FILL
XFILL_3__14886_ gnd vdd FILL
XFILL_0__10938_ gnd vdd FILL
XFILL_0__8224_ gnd vdd FILL
XFILL_1__11188_ gnd vdd FILL
XFILL_4__13107_ gnd vdd FILL
XFILL_5__12658_ gnd vdd FILL
XFILL_4__10319_ gnd vdd FILL
X_8852_ _8928_/Q gnd _8854_/A vdd INVX1
XFILL_5__15446_ gnd vdd FILL
XFILL_3__13837_ gnd vdd FILL
XFILL_4__14087_ gnd vdd FILL
XFILL_2__12478_ gnd vdd FILL
XFILL_1__10139_ gnd vdd FILL
XFILL_4__11299_ gnd vdd FILL
XFILL_2__15266_ gnd vdd FILL
XFILL_0__13657_ gnd vdd FILL
XFILL_6__9731_ gnd vdd FILL
XSFILL89400x18050 gnd vdd FILL
XFILL_1__15996_ gnd vdd FILL
X_7803_ _7803_/A _7814_/A _7802_/Y gnd _7895_/D vdd OAI21X1
XFILL_5__11609_ gnd vdd FILL
XFILL_5__15377_ gnd vdd FILL
XFILL_4__13038_ gnd vdd FILL
XFILL_5__12589_ gnd vdd FILL
XFILL_2__14217_ gnd vdd FILL
X_8783_ _8783_/A _8765_/B _8782_/Y gnd _8819_/D vdd OAI21X1
XFILL_2__11429_ gnd vdd FILL
XFILL_0__12608_ gnd vdd FILL
XFILL_3__13768_ gnd vdd FILL
XFILL_2__15197_ gnd vdd FILL
XSFILL74200x60050 gnd vdd FILL
XFILL_1__14947_ gnd vdd FILL
XFILL_0__16376_ gnd vdd FILL
XFILL_0__7106_ gnd vdd FILL
XFILL_0__13588_ gnd vdd FILL
XFILL_5__14328_ gnd vdd FILL
X_7734_ _7759_/B _7990_/B gnd _7734_/Y vdd NAND2X1
XFILL_3__15507_ gnd vdd FILL
XFILL_0__8086_ gnd vdd FILL
XSFILL89000x20050 gnd vdd FILL
XFILL_3__12719_ gnd vdd FILL
XFILL_6__13879_ gnd vdd FILL
XFILL_3__8904_ gnd vdd FILL
XFILL_2__14148_ gnd vdd FILL
XFILL_0__15327_ gnd vdd FILL
XFILL_3__9884_ gnd vdd FILL
XFILL_3__13699_ gnd vdd FILL
XFILL_1__14878_ gnd vdd FILL
XFILL_6__15618_ gnd vdd FILL
XFILL_0__7037_ gnd vdd FILL
XSFILL13640x13050 gnd vdd FILL
XFILL_5__14259_ gnd vdd FILL
X_7665_ _7623_/A _9077_/CLK _7665_/R vdd _7665_/D gnd vdd DFFSR
XFILL_3__15438_ gnd vdd FILL
XFILL_3__8835_ gnd vdd FILL
XFILL_4__14989_ gnd vdd FILL
XFILL_2__14079_ gnd vdd FILL
XFILL_1__13829_ gnd vdd FILL
XFILL_0__15258_ gnd vdd FILL
XFILL_5_BUFX2_insert80 gnd vdd FILL
X_9404_ _9356_/A _8764_/B gnd _9405_/C vdd NAND2X1
XFILL_5_BUFX2_insert91 gnd vdd FILL
XFILL_1__7850_ gnd vdd FILL
XSFILL104920x4050 gnd vdd FILL
XFILL_3__15369_ gnd vdd FILL
XFILL_0__14209_ gnd vdd FILL
X_7596_ _7656_/Q gnd _7596_/Y vdd INVX1
XFILL_3__8766_ gnd vdd FILL
XFILL_0__15189_ gnd vdd FILL
X_9335_ _8823_/A _9420_/B gnd _9335_/Y vdd NAND2X1
XFILL_6__8475_ gnd vdd FILL
XFILL_3__7717_ gnd vdd FILL
XFILL_0__8988_ gnd vdd FILL
XSFILL114520x79050 gnd vdd FILL
XFILL_6__7426_ gnd vdd FILL
XFILL_4__7490_ gnd vdd FILL
XFILL_3__8697_ gnd vdd FILL
XFILL_4_BUFX2_insert226 gnd vdd FILL
XFILL_1__9520_ gnd vdd FILL
XFILL_0__7939_ gnd vdd FILL
X_9266_ _9266_/A gnd _9268_/A vdd INVX1
XFILL_4_BUFX2_insert237 gnd vdd FILL
XSFILL33800x26050 gnd vdd FILL
XFILL_4_BUFX2_insert248 gnd vdd FILL
XSFILL43960x70050 gnd vdd FILL
XFILL_4_BUFX2_insert259 gnd vdd FILL
X_8217_ _8217_/A _8216_/A _8217_/C gnd _8289_/D vdd OAI21X1
X_9197_ _9197_/Q _8051_/CLK _8038_/R vdd _9149_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert904 gnd vdd FILL
XFILL_4__9160_ gnd vdd FILL
XFILL_3__7579_ gnd vdd FILL
XFILL_3_BUFX2_insert915 gnd vdd FILL
XFILL_0__9609_ gnd vdd FILL
XFILL_1__8402_ gnd vdd FILL
X_8148_ _8098_/B _7508_/B gnd _8149_/C vdd NAND2X1
XFILL_3_BUFX2_insert926 gnd vdd FILL
XFILL_1__9382_ gnd vdd FILL
XFILL_3_BUFX2_insert937 gnd vdd FILL
XFILL_4__8111_ gnd vdd FILL
XFILL_3_BUFX2_insert948 gnd vdd FILL
XFILL111960x36050 gnd vdd FILL
XFILL_4__9091_ gnd vdd FILL
XFILL_3_BUFX2_insert959 gnd vdd FILL
XFILL_6__9027_ gnd vdd FILL
XFILL_1__8333_ gnd vdd FILL
X_8079_ _8079_/A _8207_/B gnd _8080_/C vdd NAND2X1
XSFILL23720x78050 gnd vdd FILL
XFILL_3__9249_ gnd vdd FILL
XFILL_1__8264_ gnd vdd FILL
X_10981_ _10987_/Q gnd _10983_/A vdd INVX1
XFILL_1__7215_ gnd vdd FILL
XFILL_1__8195_ gnd vdd FILL
XFILL_3_BUFX2_insert1009 gnd vdd FILL
X_12720_ _12762_/A memoryOutData[8] gnd _12721_/C vdd NAND2X1
XFILL_1_BUFX2_insert105 gnd vdd FILL
XFILL_4__9993_ gnd vdd FILL
X_12651_ _12428_/B gnd _12651_/Y vdd INVX1
XFILL_1__7077_ gnd vdd FILL
XFILL_0_CLKBUF1_insert220 gnd vdd FILL
XFILL_0_BUFX2_insert805 gnd vdd FILL
XFILL_4__8875_ gnd vdd FILL
X_11602_ _11602_/A gnd _11604_/B vdd INVX1
X_15370_ _15370_/A _15369_/Y gnd _15370_/Y vdd NOR2X1
X_12582_ _12668_/Q gnd _12582_/Y vdd INVX1
XFILL_0_BUFX2_insert816 gnd vdd FILL
XFILL_2__6910_ gnd vdd FILL
XFILL_0_BUFX2_insert827 gnd vdd FILL
XFILL_0_BUFX2_insert838 gnd vdd FILL
XFILL_1_BUFX2_insert1002 gnd vdd FILL
XFILL_4__7826_ gnd vdd FILL
XFILL_2__7890_ gnd vdd FILL
X_14321_ _14317_/Y _14321_/B gnd _14321_/Y vdd NOR2X1
XFILL_0_BUFX2_insert849 gnd vdd FILL
XFILL_1_BUFX2_insert1013 gnd vdd FILL
X_11533_ _11533_/A _11533_/B _11294_/Y gnd _11534_/A vdd AOI21X1
XFILL_1_BUFX2_insert1024 gnd vdd FILL
XFILL_1_BUFX2_insert1035 gnd vdd FILL
XFILL_2__6841_ gnd vdd FILL
XFILL_1_BUFX2_insert1046 gnd vdd FILL
XFILL_4__7757_ gnd vdd FILL
XFILL_1_BUFX2_insert1057 gnd vdd FILL
X_14252_ _10406_/A _14389_/B _14572_/C _14252_/D gnd _14253_/B vdd AOI22X1
X_11464_ _11191_/A _11480_/C _11480_/A gnd _11464_/Y vdd AOI21X1
XSFILL23800x58050 gnd vdd FILL
XFILL_1_BUFX2_insert1068 gnd vdd FILL
XFILL_1__7979_ gnd vdd FILL
X_13203_ _11971_/A _13175_/CLK _13199_/R vdd _13203_/D gnd vdd DFFSR
X_10415_ _15822_/B gnd _10415_/Y vdd INVX1
XFILL112120x25050 gnd vdd FILL
XFILL_4__7688_ gnd vdd FILL
XFILL_2__8511_ gnd vdd FILL
X_14183_ _7459_/A gnd _14184_/A vdd INVX1
XFILL_1__9718_ gnd vdd FILL
X_11395_ _11395_/A _11054_/A _11394_/Y gnd _11395_/Y vdd OAI21X1
XFILL_4__10670_ gnd vdd FILL
XFILL_5__8220_ gnd vdd FILL
XFILL_4__9427_ gnd vdd FILL
XSFILL64040x10050 gnd vdd FILL
XFILL_2__9491_ gnd vdd FILL
XFILL_1__10490_ gnd vdd FILL
X_13134_ _13134_/A _13134_/B gnd _13135_/C vdd NAND2X1
X_10346_ _15863_/B _9834_/CLK _7793_/R vdd _10292_/Y gnd vdd DFFSR
XFILL_5__11960_ gnd vdd FILL
XFILL_4_BUFX2_insert760 gnd vdd FILL
XFILL_3__11050_ gnd vdd FILL
XFILL_3_CLKBUF1_insert1081 gnd vdd FILL
XFILL_4_BUFX2_insert771 gnd vdd FILL
XFILL_1__9649_ gnd vdd FILL
XFILL_2__10800_ gnd vdd FILL
XFILL_2__8442_ gnd vdd FILL
XFILL_4_BUFX2_insert782 gnd vdd FILL
XFILL_2__11780_ gnd vdd FILL
XFILL_4__9358_ gnd vdd FILL
XFILL_6_CLKBUF1_insert137 gnd vdd FILL
XFILL_5__10911_ gnd vdd FILL
XFILL_4_BUFX2_insert793 gnd vdd FILL
X_13065_ _6888_/A _8169_/CLK _7408_/R vdd _13007_/Y gnd vdd DFFSR
XFILL_3__10001_ gnd vdd FILL
X_10277_ _10277_/A _10304_/B _10276_/Y gnd _10277_/Y vdd OAI21X1
XFILL_4__12340_ gnd vdd FILL
XFILL_5__11891_ gnd vdd FILL
XFILL_2__8373_ gnd vdd FILL
XFILL_5__7102_ gnd vdd FILL
XFILL_0__11910_ gnd vdd FILL
XFILL_1__12160_ gnd vdd FILL
X_12016_ _12084_/A _12710_/A _12084_/C gnd _12018_/B vdd NAND3X1
XFILL_5__13630_ gnd vdd FILL
XFILL_0__12890_ gnd vdd FILL
XFILL_4__9289_ gnd vdd FILL
XFILL_5__8082_ gnd vdd FILL
XSFILL69240x50 gnd vdd FILL
XFILL_2__7324_ gnd vdd FILL
XFILL_4__12271_ gnd vdd FILL
XFILL_1__11111_ gnd vdd FILL
XFILL_2__10662_ gnd vdd FILL
XFILL_2__13450_ gnd vdd FILL
XFILL_1__12091_ gnd vdd FILL
XFILL_5__7033_ gnd vdd FILL
XFILL_0__11841_ gnd vdd FILL
XFILL_4__14010_ gnd vdd FILL
XFILL_5__13561_ gnd vdd FILL
XFILL_4__11222_ gnd vdd FILL
XFILL_2__12401_ gnd vdd FILL
XFILL_3__14740_ gnd vdd FILL
XFILL_5__10773_ gnd vdd FILL
XFILL_3__11952_ gnd vdd FILL
XFILL_2__13381_ gnd vdd FILL
XFILL_1__11042_ gnd vdd FILL
XFILL_0__14560_ gnd vdd FILL
XFILL_5__12512_ gnd vdd FILL
XFILL_5__15300_ gnd vdd FILL
XFILL_0__11772_ gnd vdd FILL
XFILL_6__14851_ gnd vdd FILL
XFILL_5__16280_ gnd vdd FILL
XFILL_3__10903_ gnd vdd FILL
XFILL_2__12332_ gnd vdd FILL
XFILL_4__11153_ gnd vdd FILL
XFILL_5__13492_ gnd vdd FILL
X_13967_ _10720_/Q gnd _13969_/B vdd INVX1
XFILL_2__15120_ gnd vdd FILL
XFILL_2__7186_ gnd vdd FILL
XFILL_3__14671_ gnd vdd FILL
XFILL_0__13511_ gnd vdd FILL
XFILL_3__11883_ gnd vdd FILL
XFILL_1__15850_ gnd vdd FILL
XFILL_0__14491_ gnd vdd FILL
XFILL_6__13802_ gnd vdd FILL
X_15706_ _15697_/Y _15706_/B gnd _15732_/A vdd NOR2X1
XFILL_5__15231_ gnd vdd FILL
XFILL_3__16410_ gnd vdd FILL
XFILL_5__8984_ gnd vdd FILL
XFILL_4__10104_ gnd vdd FILL
XFILL_5__12443_ gnd vdd FILL
X_12918_ _12916_/Y vdd _12918_/C gnd _12918_/Y vdd OAI21X1
XFILL_3__13622_ gnd vdd FILL
XFILL_0__16230_ gnd vdd FILL
XFILL_1__14801_ gnd vdd FILL
XFILL_2__15051_ gnd vdd FILL
XFILL_4__15961_ gnd vdd FILL
XFILL_2__12263_ gnd vdd FILL
XFILL_4__11084_ gnd vdd FILL
X_13898_ _9361_/A _13883_/B _14868_/A _15439_/A gnd _13907_/A vdd AOI22X1
XFILL_3__10834_ gnd vdd FILL
XFILL_0__13442_ gnd vdd FILL
XFILL_5__7935_ gnd vdd FILL
XFILL_1__12993_ gnd vdd FILL
XFILL_1__15781_ gnd vdd FILL
XFILL_0__10654_ gnd vdd FILL
X_15637_ _15637_/A _15342_/B _15637_/C gnd _15637_/Y vdd OAI21X1
XFILL_5__15162_ gnd vdd FILL
XSFILL74120x75050 gnd vdd FILL
XFILL_3__16341_ gnd vdd FILL
X_12849_ _12847_/Y vdd _12849_/C gnd _12927_/D vdd OAI21X1
XFILL_2__14002_ gnd vdd FILL
XFILL_5__12374_ gnd vdd FILL
XFILL_1_BUFX2_insert650 gnd vdd FILL
XFILL_4__10035_ gnd vdd FILL
XFILL_4__14912_ gnd vdd FILL
XFILL_2__11214_ gnd vdd FILL
XFILL_4__15892_ gnd vdd FILL
XFILL_1_BUFX2_insert661 gnd vdd FILL
XFILL_3__13553_ gnd vdd FILL
XFILL_3__6950_ gnd vdd FILL
XFILL_3__10765_ gnd vdd FILL
XFILL_1_BUFX2_insert672 gnd vdd FILL
XFILL_1__11944_ gnd vdd FILL
XFILL_1__14732_ gnd vdd FILL
XFILL_2__12194_ gnd vdd FILL
XFILL_0__16161_ gnd vdd FILL
XFILL_0__13373_ gnd vdd FILL
XFILL_5__14113_ gnd vdd FILL
XFILL_1_BUFX2_insert683 gnd vdd FILL
XFILL_5__7866_ gnd vdd FILL
XFILL_5__11325_ gnd vdd FILL
XFILL_4__14843_ gnd vdd FILL
XFILL_3__12504_ gnd vdd FILL
XFILL_6__13664_ gnd vdd FILL
XFILL_1_BUFX2_insert694 gnd vdd FILL
X_15568_ _15568_/A _15313_/B _15568_/C gnd _15570_/C vdd NOR3X1
XFILL_5__15093_ gnd vdd FILL
XFILL_2__11145_ gnd vdd FILL
XFILL_0__15112_ gnd vdd FILL
XFILL_3__16272_ gnd vdd FILL
XFILL_3__13484_ gnd vdd FILL
XFILL_0__12324_ gnd vdd FILL
XFILL_5__9605_ gnd vdd FILL
XFILL_1__11875_ gnd vdd FILL
XFILL_6__15403_ gnd vdd FILL
XFILL_0__16092_ gnd vdd FILL
XFILL_3__6881_ gnd vdd FILL
XFILL_1__14663_ gnd vdd FILL
XFILL_3__10696_ gnd vdd FILL
XFILL_0__8911_ gnd vdd FILL
X_14519_ _14519_/A _14518_/Y gnd _14526_/C vdd NOR2X1
XFILL_5__14044_ gnd vdd FILL
XFILL_3__15223_ gnd vdd FILL
X_7450_ _7522_/Q gnd _7450_/Y vdd INVX1
XFILL_5__11256_ gnd vdd FILL
XFILL_0__9891_ gnd vdd FILL
X_15499_ _13991_/Y _16213_/B _15980_/C _13990_/Y gnd _15500_/B vdd OAI22X1
XFILL_3__8620_ gnd vdd FILL
XFILL_3__12435_ gnd vdd FILL
XFILL_1__16402_ gnd vdd FILL
XFILL_4__14774_ gnd vdd FILL
XFILL_1__13614_ gnd vdd FILL
XFILL_1__10826_ gnd vdd FILL
XFILL_4__11986_ gnd vdd FILL
XFILL_0__15043_ gnd vdd FILL
XFILL_2__15953_ gnd vdd FILL
XFILL_2__11076_ gnd vdd FILL
XFILL_1__14594_ gnd vdd FILL
XFILL_5__9536_ gnd vdd FILL
XFILL_0__12255_ gnd vdd FILL
XFILL_0__8842_ gnd vdd FILL
XFILL_4__13725_ gnd vdd FILL
XFILL_4__10937_ gnd vdd FILL
X_7381_ _7381_/A _7369_/B _7381_/C gnd _7381_/Y vdd OAI21X1
XFILL_3__15154_ gnd vdd FILL
XFILL_5__11187_ gnd vdd FILL
XFILL_2__14904_ gnd vdd FILL
XFILL_2__10027_ gnd vdd FILL
XFILL_3__12366_ gnd vdd FILL
XFILL_1__16333_ gnd vdd FILL
XFILL_2__9758_ gnd vdd FILL
XFILL_1__13545_ gnd vdd FILL
XFILL_0__11206_ gnd vdd FILL
XFILL_1__10757_ gnd vdd FILL
XFILL_2__15884_ gnd vdd FILL
X_9120_ _9188_/Q gnd _9120_/Y vdd INVX1
XFILL_0__12186_ gnd vdd FILL
XFILL_5__9467_ gnd vdd FILL
XFILL_5__10138_ gnd vdd FILL
XFILL_6__15265_ gnd vdd FILL
XFILL_3__14105_ gnd vdd FILL
XFILL_3__7502_ gnd vdd FILL
XFILL_4__13656_ gnd vdd FILL
XFILL_0__8773_ gnd vdd FILL
XFILL_3__11317_ gnd vdd FILL
XFILL_2__8709_ gnd vdd FILL
XFILL_2__14835_ gnd vdd FILL
XFILL_5__15995_ gnd vdd FILL
XFILL_3__15085_ gnd vdd FILL
XFILL_3__8482_ gnd vdd FILL
XFILL_1__13476_ gnd vdd FILL
XFILL_0__11137_ gnd vdd FILL
XFILL_1__16264_ gnd vdd FILL
XFILL_3__12297_ gnd vdd FILL
XFILL_1__10688_ gnd vdd FILL
XFILL_6__14216_ gnd vdd FILL
XFILL_6__8191_ gnd vdd FILL
XFILL_5__9398_ gnd vdd FILL
XFILL_4__12607_ gnd vdd FILL
XFILL_0__7724_ gnd vdd FILL
X_9051_ _9051_/Q _8151_/CLK _9048_/R vdd _9051_/D gnd vdd DFFSR
XFILL_3__14036_ gnd vdd FILL
XFILL_5__10069_ gnd vdd FILL
XFILL_5__14946_ gnd vdd FILL
XFILL_4__16375_ gnd vdd FILL
XSFILL89960x9050 gnd vdd FILL
XFILL_4__13587_ gnd vdd FILL
XFILL_1__15215_ gnd vdd FILL
XFILL_1__12427_ gnd vdd FILL
XFILL_3__7433_ gnd vdd FILL
XFILL_3__11248_ gnd vdd FILL
XFILL_1__16195_ gnd vdd FILL
XFILL_4__10799_ gnd vdd FILL
XFILL_2__14766_ gnd vdd FILL
XFILL_0__15945_ gnd vdd FILL
XFILL_2__11978_ gnd vdd FILL
XFILL_0__11068_ gnd vdd FILL
XFILL_5__8349_ gnd vdd FILL
X_8002_ _7955_/B _6978_/B gnd _8002_/Y vdd NAND2X1
XFILL_4__15326_ gnd vdd FILL
XFILL_6__11359_ gnd vdd FILL
XFILL_5__14877_ gnd vdd FILL
XSFILL18680x61050 gnd vdd FILL
XFILL_2__13717_ gnd vdd FILL
XFILL_3__11179_ gnd vdd FILL
XFILL_1__15146_ gnd vdd FILL
XSFILL48920x22050 gnd vdd FILL
XFILL_0__10019_ gnd vdd FILL
XFILL_2__10929_ gnd vdd FILL
XSFILL19160x68050 gnd vdd FILL
XFILL_1__12358_ gnd vdd FILL
XFILL_3__7364_ gnd vdd FILL
XSFILL74200x55050 gnd vdd FILL
XFILL_2__14697_ gnd vdd FILL
XFILL_6__14078_ gnd vdd FILL
XFILL_0__15876_ gnd vdd FILL
XFILL_5__13828_ gnd vdd FILL
XFILL_3__9103_ gnd vdd FILL
XFILL_4__15257_ gnd vdd FILL
XFILL_0__7586_ gnd vdd FILL
XFILL_4__12469_ gnd vdd FILL
XFILL_1__11309_ gnd vdd FILL
XFILL_3__15987_ gnd vdd FILL
XFILL_2__13648_ gnd vdd FILL
XFILL_1__15077_ gnd vdd FILL
XFILL_3__7295_ gnd vdd FILL
XFILL_0__14827_ gnd vdd FILL
XFILL_1__12289_ gnd vdd FILL
XFILL_4__14208_ gnd vdd FILL
XSFILL49000x31050 gnd vdd FILL
XFILL_3__9034_ gnd vdd FILL
XFILL_4__15188_ gnd vdd FILL
XFILL_5__13759_ gnd vdd FILL
X_9953_ _9879_/A _9953_/CLK _9441_/R vdd _9953_/D gnd vdd DFFSR
XFILL_1__14028_ gnd vdd FILL
XFILL_3__14938_ gnd vdd FILL
XFILL_2__16367_ gnd vdd FILL
XFILL_2__13579_ gnd vdd FILL
XFILL_0__14758_ gnd vdd FILL
XSFILL109560x42050 gnd vdd FILL
XFILL_0__9256_ gnd vdd FILL
XFILL_4__14139_ gnd vdd FILL
X_8904_ _8859_/A _7496_/B gnd _8905_/C vdd NAND2X1
XFILL_2__15318_ gnd vdd FILL
XFILL_3__14869_ gnd vdd FILL
X_9884_ _9884_/A _9865_/A _9883_/Y gnd _9884_/Y vdd OAI21X1
XFILL_0__13709_ gnd vdd FILL
XSFILL38840x74050 gnd vdd FILL
XFILL_2__16298_ gnd vdd FILL
XFILL_0__8207_ gnd vdd FILL
XFILL112360x81050 gnd vdd FILL
XFILL_0__14689_ gnd vdd FILL
XFILL_5__15429_ gnd vdd FILL
XSFILL54120x22050 gnd vdd FILL
X_8835_ _8845_/B _9347_/B gnd _8835_/Y vdd NAND2X1
XFILL_2__15249_ gnd vdd FILL
XFILL_4__6990_ gnd vdd FILL
XFILL_1__15979_ gnd vdd FILL
XFILL_0__8138_ gnd vdd FILL
XFILL_6_BUFX2_insert822 gnd vdd FILL
X_8766_ _8814_/Q gnd _8766_/Y vdd INVX1
XFILL_6_BUFX2_insert833 gnd vdd FILL
XFILL_3__9936_ gnd vdd FILL
XFILL_0__16359_ gnd vdd FILL
XSFILL43960x65050 gnd vdd FILL
X_7717_ _7715_/Y _7690_/B _7716_/Y gnd _7781_/D vdd OAI21X1
XFILL_0__8069_ gnd vdd FILL
XFILL_1__8951_ gnd vdd FILL
X_8697_ _8791_/Q gnd _8699_/A vdd INVX1
XFILL_3__9867_ gnd vdd FILL
XFILL_6_BUFX2_insert899 gnd vdd FILL
XFILL_4__8660_ gnd vdd FILL
XSFILL18760x41050 gnd vdd FILL
XSFILL8600x51050 gnd vdd FILL
X_7648_ _7572_/A _7791_/CLK _7648_/R vdd _7574_/Y gnd vdd DFFSR
XFILL_4__7611_ gnd vdd FILL
XSFILL44040x74050 gnd vdd FILL
XFILL_1__8882_ gnd vdd FILL
XFILL_4__8591_ gnd vdd FILL
XFILL_3__9798_ gnd vdd FILL
XFILL_1__7833_ gnd vdd FILL
X_7579_ _7562_/B _7579_/B gnd _7579_/Y vdd NAND2X1
XSFILL63880x16050 gnd vdd FILL
XFILL_4__7542_ gnd vdd FILL
XFILL_3__8749_ gnd vdd FILL
X_9318_ _9318_/Q _7411_/CLK _8929_/R vdd _9318_/D gnd vdd DFFSR
XFILL_1__7764_ gnd vdd FILL
X_10200_ _13572_/A _8152_/CLK _9944_/R vdd _10110_/Y gnd vdd DFFSR
XFILL_4__7473_ gnd vdd FILL
XFILL_1__9503_ gnd vdd FILL
X_11180_ _12314_/Y gnd _11180_/Y vdd INVX1
X_9249_ _9228_/A _9889_/B gnd _9249_/Y vdd NAND2X1
XFILL_4__9212_ gnd vdd FILL
XFILL_1__7695_ gnd vdd FILL
XFILL112440x61050 gnd vdd FILL
X_10131_ _10129_/Y _10193_/A _10131_/C gnd _10207_/D vdd OAI21X1
XFILL_3_BUFX2_insert701 gnd vdd FILL
XFILL_3_BUFX2_insert712 gnd vdd FILL
XFILL_3_BUFX2_insert723 gnd vdd FILL
XFILL_4__9143_ gnd vdd FILL
XFILL_3_BUFX2_insert734 gnd vdd FILL
X_10062_ _9985_/B _8526_/B gnd _10063_/C vdd NAND2X1
XSFILL39000x63050 gnd vdd FILL
XFILL_3_BUFX2_insert745 gnd vdd FILL
XFILL_3_BUFX2_insert756 gnd vdd FILL
XFILL_3_BUFX2_insert767 gnd vdd FILL
XFILL_1__9365_ gnd vdd FILL
XFILL_3_BUFX2_insert778 gnd vdd FILL
XFILL_3_BUFX2_insert789 gnd vdd FILL
X_14870_ _10061_/A gnd _14870_/Y vdd INVX1
XFILL_1__8316_ gnd vdd FILL
XFILL_1__9296_ gnd vdd FILL
XSFILL18840x21050 gnd vdd FILL
XSFILL94280x82050 gnd vdd FILL
X_13821_ _13820_/Y _14045_/A _14200_/C _13821_/D gnd _13825_/A vdd OAI22X1
XFILL_2__7040_ gnd vdd FILL
XFILL_1__8247_ gnd vdd FILL
X_13752_ _15300_/A _14389_/B _14868_/D _9180_/Q gnd _13760_/B vdd AOI22X1
X_10964_ _10964_/A _10963_/Y _10964_/C gnd _10979_/B vdd NAND3X1
X_12703_ _12703_/A _10944_/C _12703_/C gnd _12793_/D vdd OAI21X1
XFILL_4__9976_ gnd vdd FILL
X_13683_ _15246_/A _14344_/B _13818_/A _7298_/A gnd _13683_/Y vdd AOI22X1
X_10895_ _10895_/A _10894_/Y _10891_/Y gnd _10896_/A vdd OAI21X1
XFILL_5__7720_ gnd vdd FILL
XFILL_2__8991_ gnd vdd FILL
X_15422_ _9745_/A gnd _15423_/B vdd INVX1
X_12634_ vdd memoryOutData[22] gnd _12635_/C vdd NAND2X1
XFILL_0_BUFX2_insert602 gnd vdd FILL
XFILL_3__10550_ gnd vdd FILL
XFILL_0_BUFX2_insert613 gnd vdd FILL
XFILL_2__7942_ gnd vdd FILL
XFILL_0_BUFX2_insert624 gnd vdd FILL
XFILL_0__10370_ gnd vdd FILL
XFILL_4__8858_ gnd vdd FILL
XFILL_5__11110_ gnd vdd FILL
XFILL_0_BUFX2_insert635 gnd vdd FILL
X_15353_ _15353_/A _15351_/Y gnd _15353_/Y vdd NOR2X1
XFILL_0_BUFX2_insert646 gnd vdd FILL
XFILL_5__12090_ gnd vdd FILL
X_12565_ _12107_/B _13180_/CLK _13180_/R vdd _12565_/D gnd vdd DFFSR
XFILL_4__11840_ gnd vdd FILL
XSFILL89240x71050 gnd vdd FILL
XSFILL53880x48050 gnd vdd FILL
XFILL_0_BUFX2_insert657 gnd vdd FILL
XFILL_4__7809_ gnd vdd FILL
XFILL_0_BUFX2_insert668 gnd vdd FILL
XFILL_1__11660_ gnd vdd FILL
XFILL_2__7873_ gnd vdd FILL
XSFILL3480x12050 gnd vdd FILL
XFILL_0_BUFX2_insert679 gnd vdd FILL
X_14304_ _14643_/C _14302_/Y _14640_/C _15760_/B gnd _14305_/B vdd OAI22X1
X_11516_ _11516_/A gnd _12512_/B vdd INVX1
XFILL_5__7582_ gnd vdd FILL
XFILL_5__11041_ gnd vdd FILL
XFILL_4__8789_ gnd vdd FILL
XFILL_2__9612_ gnd vdd FILL
XFILL_3__12220_ gnd vdd FILL
X_15284_ _15284_/A _15284_/B gnd _15285_/B vdd NOR2X1
X_12496_ _12496_/A gnd _12496_/Y vdd INVX1
XFILL_4__11771_ gnd vdd FILL
XSFILL3720x74050 gnd vdd FILL
XFILL_0__12040_ gnd vdd FILL
XSFILL28680x24050 gnd vdd FILL
XFILL_6__12331_ gnd vdd FILL
XFILL_1__11591_ gnd vdd FILL
X_14235_ _9958_/Q gnd _14237_/D vdd INVX1
XSFILL84200x18050 gnd vdd FILL
XFILL_4__13510_ gnd vdd FILL
X_11447_ _11241_/Y _11447_/B _11447_/C gnd _11447_/Y vdd AOI21X1
XFILL_1__13330_ gnd vdd FILL
XFILL_4__14490_ gnd vdd FILL
XFILL_2__11901_ gnd vdd FILL
XFILL_3__12151_ gnd vdd FILL
XFILL_2__9543_ gnd vdd FILL
XSFILL94360x62050 gnd vdd FILL
XFILL_1__10542_ gnd vdd FILL
XFILL_5__9252_ gnd vdd FILL
XFILL_2__12881_ gnd vdd FILL
XSFILL68520x72050 gnd vdd FILL
XFILL_5__14800_ gnd vdd FILL
XFILL_6__15050_ gnd vdd FILL
X_14166_ _8608_/A gnd _15611_/B vdd INVX1
XFILL_4__13441_ gnd vdd FILL
XFILL_3__11102_ gnd vdd FILL
X_11378_ _11021_/Y _11027_/B gnd _11379_/C vdd NOR2X1
XFILL_2__14620_ gnd vdd FILL
XFILL_3__12082_ gnd vdd FILL
XFILL_5__15780_ gnd vdd FILL
XFILL_4__10653_ gnd vdd FILL
XFILL_5__12992_ gnd vdd FILL
XFILL_2__9474_ gnd vdd FILL
XFILL_1__13261_ gnd vdd FILL
XFILL_5__8203_ gnd vdd FILL
XFILL_2__11832_ gnd vdd FILL
XFILL_6__14001_ gnd vdd FILL
X_10329_ _10239_/A _7129_/CLK _8542_/R vdd _10329_/D gnd vdd DFFSR
XFILL_0__13991_ gnd vdd FILL
X_13117_ _13117_/A _13108_/B _13117_/C gnd _13187_/D vdd OAI21X1
XFILL_3__15910_ gnd vdd FILL
XFILL_5__11943_ gnd vdd FILL
XFILL_1__15000_ gnd vdd FILL
XFILL_5__14731_ gnd vdd FILL
XFILL_4_BUFX2_insert590 gnd vdd FILL
XFILL_6__12193_ gnd vdd FILL
XFILL_4__16160_ gnd vdd FILL
XFILL_3__11033_ gnd vdd FILL
XFILL_4__13372_ gnd vdd FILL
XFILL_1__12212_ gnd vdd FILL
X_14097_ _13865_/C _7709_/A _7581_/A _14290_/C gnd _14106_/B vdd AOI22X1
XFILL_2__14551_ gnd vdd FILL
XFILL_0__15730_ gnd vdd FILL
XFILL_5__8134_ gnd vdd FILL
XFILL_2__11763_ gnd vdd FILL
XFILL_0__7440_ gnd vdd FILL
XFILL_6__11144_ gnd vdd FILL
XFILL_4__15111_ gnd vdd FILL
XFILL_4__12323_ gnd vdd FILL
X_13048_ _6871_/A _8180_/CLK _7391_/R vdd _13048_/D gnd vdd DFFSR
XFILL_5__11874_ gnd vdd FILL
XFILL_4__16091_ gnd vdd FILL
XFILL_3__15841_ gnd vdd FILL
XSFILL99400x6050 gnd vdd FILL
XFILL_5__14662_ gnd vdd FILL
XFILL_2__13502_ gnd vdd FILL
XFILL_2__8356_ gnd vdd FILL
XFILL_1__12143_ gnd vdd FILL
XFILL_2__14482_ gnd vdd FILL
XFILL_0__15661_ gnd vdd FILL
XFILL_2__11694_ gnd vdd FILL
XFILL_5__8065_ gnd vdd FILL
XFILL_0__12873_ gnd vdd FILL
XFILL_5__16401_ gnd vdd FILL
XFILL_5__13613_ gnd vdd FILL
XFILL_0__7371_ gnd vdd FILL
XFILL_4__15042_ gnd vdd FILL
XFILL_5__10825_ gnd vdd FILL
XFILL_5__14593_ gnd vdd FILL
XFILL_2__7307_ gnd vdd FILL
XFILL_2__16221_ gnd vdd FILL
XFILL_4__12254_ gnd vdd FILL
XFILL_0__14612_ gnd vdd FILL
XFILL_3__7080_ gnd vdd FILL
XFILL_2__13433_ gnd vdd FILL
XFILL_3__15772_ gnd vdd FILL
XFILL_2__10645_ gnd vdd FILL
XFILL_1__12074_ gnd vdd FILL
XFILL_3__12984_ gnd vdd FILL
XFILL_0__11824_ gnd vdd FILL
XFILL_0__9110_ gnd vdd FILL
XFILL_0__15592_ gnd vdd FILL
XFILL_6__10026_ gnd vdd FILL
XFILL_5__16332_ gnd vdd FILL
XSFILL89320x51050 gnd vdd FILL
XFILL_4__11205_ gnd vdd FILL
XFILL_5__13544_ gnd vdd FILL
X_6950_ _7014_/Q gnd _6950_/Y vdd INVX1
XFILL_5__10756_ gnd vdd FILL
XFILL_3__14723_ gnd vdd FILL
XFILL_1__15902_ gnd vdd FILL
XFILL_4__12185_ gnd vdd FILL
XFILL_2__7238_ gnd vdd FILL
XFILL_3__11935_ gnd vdd FILL
X_14999_ _14999_/A gnd _16293_/A vdd INVX4
XFILL_1__11025_ gnd vdd FILL
XFILL_2__16152_ gnd vdd FILL
XFILL_2__13364_ gnd vdd FILL
XSFILL109480x57050 gnd vdd FILL
XFILL_0__14543_ gnd vdd FILL
XFILL_2__10576_ gnd vdd FILL
XFILL_0__11755_ gnd vdd FILL
XFILL_0__9041_ gnd vdd FILL
XFILL_5__13475_ gnd vdd FILL
XFILL_5__16263_ gnd vdd FILL
XFILL_4__11136_ gnd vdd FILL
XFILL_2__15103_ gnd vdd FILL
XFILL_5__10687_ gnd vdd FILL
X_6881_ _6881_/A gnd memoryWriteData[11] vdd BUFX2
XFILL_2__12315_ gnd vdd FILL
XFILL_3__14654_ gnd vdd FILL
XFILL_2__13295_ gnd vdd FILL
XFILL_2__7169_ gnd vdd FILL
XSFILL54040x37050 gnd vdd FILL
XFILL_1__15833_ gnd vdd FILL
XFILL_3__11866_ gnd vdd FILL
XFILL_2__16083_ gnd vdd FILL
XFILL_0__10706_ gnd vdd FILL
XFILL_0__14474_ gnd vdd FILL
XFILL_5__15214_ gnd vdd FILL
X_8620_ _8620_/A gnd _8620_/Y vdd INVX1
XFILL_5__12426_ gnd vdd FILL
XFILL_5__8967_ gnd vdd FILL
XFILL_0__11686_ gnd vdd FILL
XFILL_3__13605_ gnd vdd FILL
XFILL_5__16194_ gnd vdd FILL
XSFILL94440x42050 gnd vdd FILL
XFILL_0__16213_ gnd vdd FILL
XFILL_4__15944_ gnd vdd FILL
XFILL_2__15034_ gnd vdd FILL
XFILL_2__12246_ gnd vdd FILL
XFILL_3__10817_ gnd vdd FILL
XFILL_4__11067_ gnd vdd FILL
XFILL_3__14585_ gnd vdd FILL
XFILL_0__13425_ gnd vdd FILL
XFILL_0__10637_ gnd vdd FILL
XFILL_3__7982_ gnd vdd FILL
XFILL_1__15764_ gnd vdd FILL
XFILL_3__11797_ gnd vdd FILL
XFILL_1__12976_ gnd vdd FILL
XFILL_5__15145_ gnd vdd FILL
XFILL_4__10018_ gnd vdd FILL
XFILL_5__12357_ gnd vdd FILL
XFILL_1_BUFX2_insert480 gnd vdd FILL
XFILL_3__16324_ gnd vdd FILL
X_8551_ _8551_/Q _8551_/CLK _9064_/R vdd _8551_/D gnd vdd DFFSR
XFILL_5__8898_ gnd vdd FILL
XFILL_3__13536_ gnd vdd FILL
XFILL_3__9721_ gnd vdd FILL
XFILL_1_BUFX2_insert491 gnd vdd FILL
XFILL_1__14715_ gnd vdd FILL
XFILL_3__6933_ gnd vdd FILL
XFILL_3__10748_ gnd vdd FILL
XFILL_2__12177_ gnd vdd FILL
XFILL_4__15875_ gnd vdd FILL
XFILL_0__16144_ gnd vdd FILL
XFILL_0__13356_ gnd vdd FILL
XFILL_1__11927_ gnd vdd FILL
X_7502_ _7503_/B _7502_/B gnd _7502_/Y vdd NAND2X1
XFILL_1__15695_ gnd vdd FILL
XFILL_5_BUFX2_insert807 gnd vdd FILL
XFILL_5__7849_ gnd vdd FILL
XFILL_5__11308_ gnd vdd FILL
XFILL_0__10568_ gnd vdd FILL
XFILL_5__15076_ gnd vdd FILL
XFILL_5_BUFX2_insert818 gnd vdd FILL
XFILL_4__14826_ gnd vdd FILL
X_8482_ _8480_/Y _8460_/A _8482_/C gnd _8548_/D vdd OAI21X1
XFILL_5_BUFX2_insert829 gnd vdd FILL
XFILL_5__12288_ gnd vdd FILL
XFILL_2__11128_ gnd vdd FILL
XFILL_3__16255_ gnd vdd FILL
XSFILL18680x56050 gnd vdd FILL
XFILL_3__13467_ gnd vdd FILL
XBUFX2_insert1004 _12399_/Y gnd _6957_/B vdd BUFX2
XFILL_0__12307_ gnd vdd FILL
XFILL_3__9652_ gnd vdd FILL
XFILL_3__10679_ gnd vdd FILL
XFILL_1__14646_ gnd vdd FILL
XFILL_3__6864_ gnd vdd FILL
XBUFX2_insert1015 _15054_/Y gnd _16314_/A vdd BUFX2
XFILL_0__16075_ gnd vdd FILL
XFILL_1__11858_ gnd vdd FILL
XFILL_0__13287_ gnd vdd FILL
XBUFX2_insert1026 _13340_/Y gnd _9625_/B vdd BUFX2
XFILL_5__14027_ gnd vdd FILL
XFILL_3__15206_ gnd vdd FILL
X_7433_ _7460_/A _9993_/B gnd _7433_/Y vdd NAND2X1
XFILL_0__10499_ gnd vdd FILL
XFILL_5__11239_ gnd vdd FILL
XBUFX2_insert1037 _12390_/Y gnd _7972_/B vdd BUFX2
XFILL_3__12418_ gnd vdd FILL
XFILL_3__8603_ gnd vdd FILL
XFILL_0__9874_ gnd vdd FILL
XFILL_4__14757_ gnd vdd FILL
XBUFX2_insert1048 _12806_/Q gnd _11885_/B vdd BUFX2
XFILL_3__16186_ gnd vdd FILL
XFILL_0__15026_ gnd vdd FILL
XFILL_2__15936_ gnd vdd FILL
XFILL_4__11969_ gnd vdd FILL
XFILL_2__11059_ gnd vdd FILL
XFILL_3__13398_ gnd vdd FILL
XBUFX2_insert1059 _15051_/Y gnd _15995_/C vdd BUFX2
XFILL_1__10809_ gnd vdd FILL
XFILL_5__9519_ gnd vdd FILL
XFILL_0__12238_ gnd vdd FILL
XFILL_1__14577_ gnd vdd FILL
XFILL_1__11789_ gnd vdd FILL
XFILL_0__8825_ gnd vdd FILL
XSFILL49000x26050 gnd vdd FILL
XSFILL74600x71050 gnd vdd FILL
X_7364_ _7364_/A gnd _7366_/A vdd INVX1
XFILL_4__13708_ gnd vdd FILL
XFILL_3__15137_ gnd vdd FILL
XFILL_3__12349_ gnd vdd FILL
XFILL_1__16316_ gnd vdd FILL
XFILL_4__14688_ gnd vdd FILL
XSFILL59160x70050 gnd vdd FILL
XSFILL89400x31050 gnd vdd FILL
XFILL_2__15867_ gnd vdd FILL
XFILL_1__13528_ gnd vdd FILL
X_9103_ _9163_/A _7439_/B gnd _9104_/C vdd NAND2X1
XFILL_0__12169_ gnd vdd FILL
XFILL_4__13639_ gnd vdd FILL
XSFILL109560x37050 gnd vdd FILL
XFILL_0__8756_ gnd vdd FILL
X_7295_ _7295_/A gnd _7297_/A vdd INVX1
XFILL_5__15978_ gnd vdd FILL
XFILL_2__14818_ gnd vdd FILL
XFILL_3__15068_ gnd vdd FILL
XSFILL64680x59050 gnd vdd FILL
XFILL_1__13459_ gnd vdd FILL
XFILL_3__8465_ gnd vdd FILL
XFILL_1__16247_ gnd vdd FILL
XFILL_2__15798_ gnd vdd FILL
X_9034_ _9034_/A gnd _9036_/A vdd INVX1
XFILL_0__7707_ gnd vdd FILL
XFILL112360x76050 gnd vdd FILL
XFILL_3__14019_ gnd vdd FILL
XFILL_1__7480_ gnd vdd FILL
XFILL_5__14929_ gnd vdd FILL
XFILL_3__7416_ gnd vdd FILL
XFILL_4__16358_ gnd vdd FILL
XFILL_2__14749_ gnd vdd FILL
XFILL_0__15928_ gnd vdd FILL
XFILL_3__8396_ gnd vdd FILL
XFILL_1__16178_ gnd vdd FILL
XFILL_6__7125_ gnd vdd FILL
XFILL_4__15309_ gnd vdd FILL
XSFILL79080x21050 gnd vdd FILL
XFILL_4__16289_ gnd vdd FILL
XFILL_1__15129_ gnd vdd FILL
XFILL_3__7347_ gnd vdd FILL
XFILL_0__15859_ gnd vdd FILL
XFILL_1__9150_ gnd vdd FILL
XFILL_2_BUFX2_insert708 gnd vdd FILL
XFILL_2_BUFX2_insert719 gnd vdd FILL
XFILL_0__7569_ gnd vdd FILL
XFILL_1__8101_ gnd vdd FILL
XSFILL18760x36050 gnd vdd FILL
XSFILL8600x46050 gnd vdd FILL
XFILL_3__9017_ gnd vdd FILL
XFILL_1__9081_ gnd vdd FILL
X_9936_ _9936_/A gnd _9936_/Y vdd INVX1
XSFILL44040x69050 gnd vdd FILL
XSFILL84440x74050 gnd vdd FILL
XFILL_0__9239_ gnd vdd FILL
X_9867_ _9949_/Q gnd _9869_/A vdd INVX1
XFILL_6__7958_ gnd vdd FILL
X_8818_ _8778_/A _8818_/CLK _7270_/R vdd _8818_/D gnd vdd DFFSR
XSFILL23880x27050 gnd vdd FILL
XFILL_4__9761_ gnd vdd FILL
X_9798_ _9798_/A _9798_/B _9797_/Y gnd _9798_/Y vdd OAI21X1
XFILL_4__6973_ gnd vdd FILL
XFILL_6__6909_ gnd vdd FILL
XBUFX2_insert707 _12816_/Q gnd _15036_/A vdd BUFX2
X_10680_ _14504_/A gnd _10680_/Y vdd INVX1
XBUFX2_insert718 _13418_/Y gnd _14160_/B vdd BUFX2
XFILL_1__9983_ gnd vdd FILL
XFILL_3__9919_ gnd vdd FILL
XFILL_4__8712_ gnd vdd FILL
XSFILL38920x49050 gnd vdd FILL
XBUFX2_insert729 _12411_/Y gnd _9657_/B vdd BUFX2
X_8749_ _8695_/B _6957_/B gnd _8750_/C vdd NAND2X1
XFILL112440x56050 gnd vdd FILL
XFILL_6_BUFX2_insert674 gnd vdd FILL
XFILL112360x1050 gnd vdd FILL
XFILL_4__8643_ gnd vdd FILL
X_12350_ _12380_/A _12573_/A gnd _12351_/C vdd NAND2X1
XFILL_1__8865_ gnd vdd FILL
XFILL_1_CLKBUF1_insert112 gnd vdd FILL
XFILL_1_CLKBUF1_insert123 gnd vdd FILL
X_11301_ _11138_/Y _11614_/A gnd _11301_/Y vdd NOR2X1
XFILL_4__8574_ gnd vdd FILL
X_12281_ _6886_/A _12277_/B _12309_/C _11882_/B gnd _12282_/C vdd AOI22X1
XFILL_1_CLKBUF1_insert134 gnd vdd FILL
XFILL_1__7816_ gnd vdd FILL
XFILL_1_CLKBUF1_insert145 gnd vdd FILL
XFILL_1_CLKBUF1_insert156 gnd vdd FILL
XSFILL74040x3050 gnd vdd FILL
X_14020_ _14868_/A _10647_/A _15509_/D _13621_/B gnd _14022_/A vdd AOI22X1
XFILL_1_CLKBUF1_insert167 gnd vdd FILL
X_11232_ _12226_/Y _11013_/B gnd _11376_/A vdd AND2X2
XSFILL114600x72050 gnd vdd FILL
XFILL_1_CLKBUF1_insert178 gnd vdd FILL
XSFILL94280x77050 gnd vdd FILL
XSFILL44120x49050 gnd vdd FILL
XFILL_1_CLKBUF1_insert189 gnd vdd FILL
XFILL_1__7747_ gnd vdd FILL
XFILL_4__7456_ gnd vdd FILL
X_11163_ _11102_/Y _12310_/Y _11162_/Y gnd _11163_/Y vdd OAI21X1
XSFILL69080x53050 gnd vdd FILL
XSFILL99320x14050 gnd vdd FILL
XFILL_1__7678_ gnd vdd FILL
X_10114_ _10114_/A gnd _10114_/Y vdd INVX1
XFILL_3_BUFX2_insert520 gnd vdd FILL
XFILL_3_BUFX2_insert531 gnd vdd FILL
X_15971_ _10861_/Q gnd _15972_/A vdd INVX1
XFILL_3_BUFX2_insert542 gnd vdd FILL
XFILL_1__9417_ gnd vdd FILL
X_11094_ _12278_/Y _11094_/B gnd _11094_/Y vdd NOR2X1
XFILL_2__8210_ gnd vdd FILL
XFILL_3_BUFX2_insert553 gnd vdd FILL
XSFILL73560x78050 gnd vdd FILL
XFILL_4__9126_ gnd vdd FILL
XSFILL23800x5050 gnd vdd FILL
XFILL_3_BUFX2_insert564 gnd vdd FILL
X_10045_ _10045_/A _9985_/B _10045_/C gnd _10093_/D vdd OAI21X1
XFILL_3_BUFX2_insert575 gnd vdd FILL
X_14922_ _8052_/Q gnd _14923_/D vdd INVX1
XFILL_3_BUFX2_insert586 gnd vdd FILL
XFILL_2__8141_ gnd vdd FILL
XFILL_1__9348_ gnd vdd FILL
XFILL_3_BUFX2_insert597 gnd vdd FILL
X_14853_ _14852_/Y _13860_/B _14203_/B _14853_/D gnd _14857_/B vdd OAI22X1
XFILL_2__10430_ gnd vdd FILL
XFILL_5__11590_ gnd vdd FILL
XFILL_1__9279_ gnd vdd FILL
XSFILL89240x66050 gnd vdd FILL
XFILL_2__8072_ gnd vdd FILL
XFILL_4__8008_ gnd vdd FILL
XFILL_5__9870_ gnd vdd FILL
X_13804_ _13804_/A _13800_/Y _13804_/C gnd _13804_/Y vdd NOR3X1
XFILL_5__10541_ gnd vdd FILL
XSFILL49240x82050 gnd vdd FILL
XFILL_3__11720_ gnd vdd FILL
XFILL_6_BUFX2_insert24 gnd vdd FILL
X_14784_ _8049_/Q gnd _14784_/Y vdd INVX1
XFILL_6_BUFX2_insert35 gnd vdd FILL
X_11996_ _12012_/A _12695_/A _11996_/C gnd _11998_/B vdd NAND3X1
XFILL_2__10361_ gnd vdd FILL
XSFILL3720x69050 gnd vdd FILL
XFILL_0__11540_ gnd vdd FILL
XSFILL28680x19050 gnd vdd FILL
XFILL_5__13260_ gnd vdd FILL
XFILL_2__12100_ gnd vdd FILL
X_13735_ _7301_/A _14353_/A _13864_/B _8667_/Q gnd _13737_/A vdd AOI22X1
X_10947_ _12773_/A _12818_/Q gnd _10948_/B vdd NOR2X1
XFILL_2__13080_ gnd vdd FILL
XFILL_4__13990_ gnd vdd FILL
XFILL_3__11651_ gnd vdd FILL
XFILL_1__12830_ gnd vdd FILL
XFILL_2__10292_ gnd vdd FILL
XFILL_5__12211_ gnd vdd FILL
XFILL_0__11471_ gnd vdd FILL
XFILL_5__8752_ gnd vdd FILL
X_13666_ _14868_/A _15235_/A _15237_/A _14877_/D gnd _13666_/Y vdd AOI22X1
XFILL_2__12031_ gnd vdd FILL
XFILL_0__13210_ gnd vdd FILL
X_10878_ _10963_/A _10877_/Y gnd _10878_/Y vdd NAND2X1
XFILL_3__14370_ gnd vdd FILL
XFILL_0__10422_ gnd vdd FILL
XFILL_1__12761_ gnd vdd FILL
XFILL_2__8974_ gnd vdd FILL
XFILL_5__7703_ gnd vdd FILL
XFILL_3__11582_ gnd vdd FILL
XFILL_0__14190_ gnd vdd FILL
X_15405_ _15405_/A _15405_/B gnd _15412_/A vdd NOR2X1
XFILL_0_BUFX2_insert410 gnd vdd FILL
XSFILL69160x33050 gnd vdd FILL
X_12617_ _12615_/Y vdd _12617_/C gnd _12679_/D vdd OAI21X1
XFILL_0_BUFX2_insert421 gnd vdd FILL
XFILL_5__12142_ gnd vdd FILL
XFILL_3__13321_ gnd vdd FILL
X_16385_ gnd gnd gnd _16385_/Y vdd NAND2X1
XFILL_4__15660_ gnd vdd FILL
XFILL_0_BUFX2_insert432 gnd vdd FILL
X_13597_ _8831_/A gnd _13597_/Y vdd INVX1
XFILL_3__10533_ gnd vdd FILL
XFILL_1__14500_ gnd vdd FILL
XFILL_4__12872_ gnd vdd FILL
XFILL_0_BUFX2_insert443 gnd vdd FILL
XFILL_1__11712_ gnd vdd FILL
XFILL_0_BUFX2_insert454 gnd vdd FILL
XFILL_0__13141_ gnd vdd FILL
XFILL_1__15480_ gnd vdd FILL
XFILL_5__7634_ gnd vdd FILL
XFILL_4__14611_ gnd vdd FILL
X_15336_ _15336_/A _15335_/Y _15336_/C gnd _15337_/B vdd NAND3X1
XFILL_0_BUFX2_insert465 gnd vdd FILL
XFILL_3__16040_ gnd vdd FILL
XSFILL73640x58050 gnd vdd FILL
XFILL_5__12073_ gnd vdd FILL
XFILL_0__6940_ gnd vdd FILL
X_12548_ _12382_/A _12537_/CLK _12536_/R vdd _12548_/D gnd vdd DFFSR
XFILL_0_BUFX2_insert476 gnd vdd FILL
XFILL_4__11823_ gnd vdd FILL
XFILL_3__13252_ gnd vdd FILL
XFILL_0_BUFX2_insert487 gnd vdd FILL
XFILL_4__15591_ gnd vdd FILL
XFILL_2__7856_ gnd vdd FILL
XFILL_0_BUFX2_insert498 gnd vdd FILL
XFILL_1__11643_ gnd vdd FILL
XFILL_1__14431_ gnd vdd FILL
XFILL_2__13982_ gnd vdd FILL
XFILL_5__7565_ gnd vdd FILL
XFILL_5__15901_ gnd vdd FILL
XFILL_0__10284_ gnd vdd FILL
XFILL_5__11024_ gnd vdd FILL
XSFILL74280x24050 gnd vdd FILL
XFILL_3__12203_ gnd vdd FILL
XFILL_4__14542_ gnd vdd FILL
X_15267_ _7173_/A _15177_/B _16014_/C _8283_/Q gnd _15273_/B vdd AOI22X1
XFILL_2__15721_ gnd vdd FILL
XFILL_4__11754_ gnd vdd FILL
X_12479_ vdd _12041_/A gnd _12479_/Y vdd NAND2X1
XFILL_0__6871_ gnd vdd FILL
XFILL_0__12023_ gnd vdd FILL
XFILL_3__10395_ gnd vdd FILL
XFILL_1__14362_ gnd vdd FILL
XFILL_1__11574_ gnd vdd FILL
X_14218_ _8422_/Q gnd _14218_/Y vdd INVX1
XFILL_0__8610_ gnd vdd FILL
XSFILL89320x46050 gnd vdd FILL
XFILL_5__7496_ gnd vdd FILL
XFILL_5__15832_ gnd vdd FILL
XFILL_4__10705_ gnd vdd FILL
XFILL_1__13313_ gnd vdd FILL
XFILL_2__9526_ gnd vdd FILL
XFILL_4__14473_ gnd vdd FILL
X_15198_ _9945_/Q gnd _15198_/Y vdd INVX1
XFILL_3__12134_ gnd vdd FILL
XFILL_0__9590_ gnd vdd FILL
XFILL_1__16101_ gnd vdd FILL
XFILL_2__15652_ gnd vdd FILL
XFILL_4__11685_ gnd vdd FILL
XFILL_1__10525_ gnd vdd FILL
XFILL_5__9235_ gnd vdd FILL
XFILL_2__12864_ gnd vdd FILL
XFILL_1__14293_ gnd vdd FILL
XFILL_4__16212_ gnd vdd FILL
X_14149_ _14149_/A _13824_/B _14575_/C _14149_/D gnd _14153_/B vdd OAI22X1
XFILL_4__13424_ gnd vdd FILL
XCLKBUF1_insert111 CLKBUF1_insert220/A gnd _8680_/CLK vdd CLKBUF1
XFILL_4__10636_ gnd vdd FILL
XFILL_2__14603_ gnd vdd FILL
X_7080_ _7078_/Y _7100_/A _7080_/C gnd _7142_/D vdd OAI21X1
XCLKBUF1_insert122 CLKBUF1_insert206/A gnd _9060_/CLK vdd CLKBUF1
XFILL_5__15763_ gnd vdd FILL
XFILL_1__13244_ gnd vdd FILL
XFILL_3__8250_ gnd vdd FILL
XFILL_1__16032_ gnd vdd FILL
XFILL_5__12975_ gnd vdd FILL
XCLKBUF1_insert133 CLKBUF1_insert216/A gnd _9436_/CLK vdd CLKBUF1
XFILL_3__12065_ gnd vdd FILL
XFILL_2__11815_ gnd vdd FILL
XFILL_2__15583_ gnd vdd FILL
XCLKBUF1_insert144 CLKBUF1_insert192/A gnd _8306_/CLK vdd CLKBUF1
XFILL_5__9166_ gnd vdd FILL
XFILL_0__13974_ gnd vdd FILL
XFILL_5__14714_ gnd vdd FILL
XFILL_4__16143_ gnd vdd FILL
XCLKBUF1_insert155 CLKBUF1_insert182/A gnd _6999_/CLK vdd CLKBUF1
XFILL_4__13355_ gnd vdd FILL
XCLKBUF1_insert166 CLKBUF1_insert206/A gnd _8541_/CLK vdd CLKBUF1
XFILL_0__8472_ gnd vdd FILL
XFILL_3__7201_ gnd vdd FILL
XFILL_5__11926_ gnd vdd FILL
XFILL_3__11016_ gnd vdd FILL
XFILL_5__15694_ gnd vdd FILL
XFILL_2__14534_ gnd vdd FILL
XCLKBUF1_insert177 CLKBUF1_insert220/A gnd _9589_/CLK vdd CLKBUF1
XFILL_4__10567_ gnd vdd FILL
XFILL_5__8117_ gnd vdd FILL
XFILL_0__15713_ gnd vdd FILL
XFILL_2__9388_ gnd vdd FILL
XFILL_2__11746_ gnd vdd FILL
XCLKBUF1_insert188 CLKBUF1_insert187/A gnd _12667_/CLK vdd CLKBUF1
XFILL_1__10387_ gnd vdd FILL
XFILL_0__7423_ gnd vdd FILL
XCLKBUF1_insert199 CLKBUF1_insert206/A gnd _9050_/CLK vdd CLKBUF1
XFILL_5__9097_ gnd vdd FILL
XFILL_4__12306_ gnd vdd FILL
XFILL_5__14645_ gnd vdd FILL
XFILL_4__16074_ gnd vdd FILL
XFILL_4__13286_ gnd vdd FILL
XFILL_1__12126_ gnd vdd FILL
XFILL_3__15824_ gnd vdd FILL
XFILL_2__8339_ gnd vdd FILL
XSFILL69240x13050 gnd vdd FILL
XFILL_5__11857_ gnd vdd FILL
XFILL_2__14465_ gnd vdd FILL
XFILL_4__10498_ gnd vdd FILL
XFILL_0__15644_ gnd vdd FILL
XFILL_0__12856_ gnd vdd FILL
XFILL_2__11677_ gnd vdd FILL
XFILL_4__15025_ gnd vdd FILL
XFILL_6__15935_ gnd vdd FILL
XFILL_2__16204_ gnd vdd FILL
XFILL_0__7354_ gnd vdd FILL
XFILL_5__10808_ gnd vdd FILL
XFILL_4__12237_ gnd vdd FILL
XFILL_5__14576_ gnd vdd FILL
XFILL_2__13416_ gnd vdd FILL
X_7982_ _7982_/A _7972_/A _7982_/C gnd _8040_/D vdd OAI21X1
XFILL_5__11788_ gnd vdd FILL
XFILL_3__15755_ gnd vdd FILL
XFILL_2__10628_ gnd vdd FILL
XFILL_3__7063_ gnd vdd FILL
XFILL_1__12057_ gnd vdd FILL
XFILL_0__11807_ gnd vdd FILL
XFILL_3__12967_ gnd vdd FILL
XFILL_2__14396_ gnd vdd FILL
XFILL_0__15575_ gnd vdd FILL
XSFILL104440x22050 gnd vdd FILL
XFILL_0__12787_ gnd vdd FILL
XFILL_5__16315_ gnd vdd FILL
XFILL_5__13527_ gnd vdd FILL
XFILL_3__14706_ gnd vdd FILL
X_6933_ _6985_/B _6933_/B gnd _6934_/C vdd NAND2X1
X_9721_ _9815_/Q gnd _9721_/Y vdd INVX1
XFILL_3__11918_ gnd vdd FILL
XFILL_4__12168_ gnd vdd FILL
XFILL_2__16135_ gnd vdd FILL
XFILL_1__11008_ gnd vdd FILL
XFILL_2__13347_ gnd vdd FILL
XFILL_3__15686_ gnd vdd FILL
XSFILL8680x20050 gnd vdd FILL
XFILL_2__10559_ gnd vdd FILL
XFILL_0__14526_ gnd vdd FILL
XFILL_0__11738_ gnd vdd FILL
XFILL_3__12898_ gnd vdd FILL
XFILL_0__9024_ gnd vdd FILL
XFILL_4__11119_ gnd vdd FILL
XFILL_5__9999_ gnd vdd FILL
XFILL_5__16246_ gnd vdd FILL
XFILL_3__14637_ gnd vdd FILL
X_6864_ _6864_/A gnd memoryAddress[26] vdd BUFX2
XFILL_5__13458_ gnd vdd FILL
XFILL_6__15797_ gnd vdd FILL
XSFILL34360x20050 gnd vdd FILL
X_9652_ _9650_/Y _9652_/B _9651_/Y gnd _9652_/Y vdd OAI21X1
XFILL_4__12099_ gnd vdd FILL
XFILL_1__15816_ gnd vdd FILL
XFILL_2__16066_ gnd vdd FILL
XFILL_3__11849_ gnd vdd FILL
XFILL_2__13278_ gnd vdd FILL
XFILL_0__14457_ gnd vdd FILL
XSFILL59160x65050 gnd vdd FILL
XFILL_0__11669_ gnd vdd FILL
XFILL_5__12409_ gnd vdd FILL
X_8603_ _8567_/B _8091_/B gnd _8604_/C vdd NAND2X1
XFILL_6__14748_ gnd vdd FILL
XFILL_4__15927_ gnd vdd FILL
XFILL_5__16177_ gnd vdd FILL
XFILL_5__13389_ gnd vdd FILL
XFILL_2__15017_ gnd vdd FILL
X_9583_ _9583_/Q _9568_/CLK _8431_/R vdd _9583_/D gnd vdd DFFSR
XFILL_3__14568_ gnd vdd FILL
XFILL_0__13408_ gnd vdd FILL
XFILL_2__12229_ gnd vdd FILL
XFILL_1__15747_ gnd vdd FILL
XFILL_3__7965_ gnd vdd FILL
XFILL_0__14388_ gnd vdd FILL
XFILL_1__12959_ gnd vdd FILL
XFILL111880x64050 gnd vdd FILL
XFILL_5_BUFX2_insert604 gnd vdd FILL
X_8534_ _8438_/A _8818_/CLK _8278_/R vdd _8534_/D gnd vdd DFFSR
XFILL_3__16307_ gnd vdd FILL
XFILL_5__15128_ gnd vdd FILL
XFILL_6__7674_ gnd vdd FILL
XFILL_5_BUFX2_insert615 gnd vdd FILL
XFILL_3__13519_ gnd vdd FILL
XFILL_3__6916_ gnd vdd FILL
XFILL_1__6980_ gnd vdd FILL
XFILL_4__15858_ gnd vdd FILL
XFILL_0__13339_ gnd vdd FILL
XFILL_3__14499_ gnd vdd FILL
XFILL_5_BUFX2_insert626 gnd vdd FILL
XFILL_0__16127_ gnd vdd FILL
XFILL_1__15678_ gnd vdd FILL
XFILL_5_BUFX2_insert637 gnd vdd FILL
XSFILL13640x21050 gnd vdd FILL
XFILL_5_BUFX2_insert648 gnd vdd FILL
XFILL_0__9926_ gnd vdd FILL
XFILL_3__16238_ gnd vdd FILL
XFILL_4__14809_ gnd vdd FILL
XFILL_5__15059_ gnd vdd FILL
XFILL_5_BUFX2_insert659 gnd vdd FILL
X_8465_ _8465_/A gnd _8465_/Y vdd INVX1
XSFILL79080x16050 gnd vdd FILL
XFILL_3__9635_ gnd vdd FILL
XFILL_1__14629_ gnd vdd FILL
XFILL_3__6847_ gnd vdd FILL
XFILL_4__15789_ gnd vdd FILL
XFILL_0__16058_ gnd vdd FILL
XSFILL79320x78050 gnd vdd FILL
X_7416_ _7416_/A _7416_/B _7415_/Y gnd _7416_/Y vdd OAI21X1
XFILL_0__9857_ gnd vdd FILL
XFILL_1__8650_ gnd vdd FILL
XFILL_2__15919_ gnd vdd FILL
X_8396_ _8394_/Y _8321_/B _8395_/Y gnd _8434_/D vdd OAI21X1
XFILL_3__16169_ gnd vdd FILL
XFILL_0__15009_ gnd vdd FILL
XFILL_6__9275_ gnd vdd FILL
XFILL_1__7601_ gnd vdd FILL
X_7347_ _7354_/B _9779_/B gnd _7347_/Y vdd NAND2X1
XFILL_0__9788_ gnd vdd FILL
XFILL_4__7310_ gnd vdd FILL
XFILL_3__8517_ gnd vdd FILL
XFILL_1__8581_ gnd vdd FILL
XFILL_3__9497_ gnd vdd FILL
XFILL_6__8226_ gnd vdd FILL
XFILL_2_CLKBUF1_insert207 gnd vdd FILL
XFILL_2_CLKBUF1_insert218 gnd vdd FILL
XFILL_0__8739_ gnd vdd FILL
XSFILL33800x34050 gnd vdd FILL
X_7278_ _7230_/A _8046_/CLK _9061_/R vdd _7278_/D gnd vdd DFFSR
XSFILL58600x79050 gnd vdd FILL
XFILL_3__8448_ gnd vdd FILL
XFILL_4__7241_ gnd vdd FILL
X_9017_ _9017_/A _9017_/B gnd _9018_/C vdd NAND2X1
XFILL_1__7463_ gnd vdd FILL
XFILL_3__8379_ gnd vdd FILL
XFILL_4__7172_ gnd vdd FILL
XFILL_2_BUFX2_insert505 gnd vdd FILL
XFILL111960x44050 gnd vdd FILL
XFILL_2_BUFX2_insert516 gnd vdd FILL
XFILL_2_BUFX2_insert527 gnd vdd FILL
XFILL_2_BUFX2_insert538 gnd vdd FILL
XFILL_1__9133_ gnd vdd FILL
XSFILL109240x14050 gnd vdd FILL
XFILL_2_BUFX2_insert549 gnd vdd FILL
XSFILL88680x74050 gnd vdd FILL
XFILL112040x53050 gnd vdd FILL
X_11850_ _11841_/B _12440_/A _11840_/Y gnd _11850_/Y vdd NOR3X1
X_9919_ _9920_/B _7359_/B gnd _9920_/C vdd NAND2X1
X_10801_ _10801_/A _10822_/B _10801_/C gnd _10857_/D vdd OAI21X1
XFILL_1__8015_ gnd vdd FILL
X_11781_ _11769_/A _11776_/A gnd _11781_/Y vdd AND2X2
XFILL_4__9813_ gnd vdd FILL
XFILL_6_BUFX2_insert1068 gnd vdd FILL
X_13520_ _8663_/Q gnd _13520_/Y vdd INVX1
X_10732_ _14504_/A _7020_/CLK _9964_/R vdd _10732_/D gnd vdd DFFSR
XBUFX2_insert504 BUFX2_insert494/A gnd _7648_/R vdd BUFX2
XBUFX2_insert515 BUFX2_insert559/A gnd _7262_/R vdd BUFX2
XFILL_4__9744_ gnd vdd FILL
XFILL_4__6956_ gnd vdd FILL
XBUFX2_insert526 BUFX2_insert496/A gnd _9048_/R vdd BUFX2
X_13451_ _13451_/A _13439_/Y _13451_/C gnd _13451_/Y vdd NAND3X1
XBUFX2_insert537 BUFX2_insert524/A gnd _7011_/R vdd BUFX2
XBUFX2_insert548 BUFX2_insert570/A gnd _7258_/R vdd BUFX2
X_10663_ _10700_/B _9895_/B gnd _10664_/C vdd NAND2X1
XBUFX2_insert559 BUFX2_insert559/A gnd _8025_/R vdd BUFX2
XFILL_4__9675_ gnd vdd FILL
X_12402_ _12400_/Y _12359_/A _12402_/C gnd _12402_/Y vdd OAI21X1
X_16170_ _16036_/A _16170_/B _15322_/A _14813_/Y gnd _16171_/B vdd OAI22X1
XFILL_4__6887_ gnd vdd FILL
XSFILL29080x64050 gnd vdd FILL
X_13382_ _13680_/B gnd _14389_/B vdd INVX8
X_10594_ _15545_/A _7778_/CLK _8418_/R vdd _10594_/D gnd vdd DFFSR
XFILL_2__7710_ gnd vdd FILL
XFILL_1__8917_ gnd vdd FILL
XFILL111960x3050 gnd vdd FILL
XFILL_4__8626_ gnd vdd FILL
XFILL_1__9897_ gnd vdd FILL
X_15121_ _13517_/A _15795_/B _15121_/C gnd _15124_/A vdd OAI21X1
X_12333_ _6899_/A _12301_/B _12301_/C _12313_/D gnd _12334_/C vdd AOI22X1
XFILL_4_BUFX2_insert1050 gnd vdd FILL
XFILL_4_BUFX2_insert1061 gnd vdd FILL
XFILL_1__8848_ gnd vdd FILL
XFILL_4_BUFX2_insert1072 gnd vdd FILL
XFILL_5__7350_ gnd vdd FILL
X_15052_ _16035_/B _16148_/C gnd _15052_/Y vdd NAND2X1
XSFILL23800x66050 gnd vdd FILL
X_12264_ _12272_/A _11876_/B _12272_/C gnd _12266_/B vdd NAND3X1
XFILL_3__10180_ gnd vdd FILL
XFILL_1__8779_ gnd vdd FILL
XFILL_4__7508_ gnd vdd FILL
XFILL_2__7572_ gnd vdd FILL
X_14003_ _14002_/Y _14862_/C gnd _14004_/C vdd NOR2X1
XFILL112120x33050 gnd vdd FILL
XFILL_4__8488_ gnd vdd FILL
X_11215_ _10882_/Y _11214_/Y gnd _11215_/Y vdd NOR2X1
X_12195_ _12195_/A _12201_/B _12195_/C gnd _12195_/Y vdd OAI21X1
XSFILL113800x19050 gnd vdd FILL
XFILL_1__10310_ gnd vdd FILL
XFILL_4__11470_ gnd vdd FILL
XFILL_5__9020_ gnd vdd FILL
XFILL_4__7439_ gnd vdd FILL
XFILL_1__11290_ gnd vdd FILL
XFILL_4__10421_ gnd vdd FILL
XFILL_5__12760_ gnd vdd FILL
X_11146_ _11582_/C _11146_/B gnd _11403_/A vdd NOR2X1
XFILL_2__9242_ gnd vdd FILL
XSFILL79880x3050 gnd vdd FILL
XFILL_2__11600_ gnd vdd FILL
XFILL_1__10241_ gnd vdd FILL
XFILL_2__12580_ gnd vdd FILL
XFILL_3_BUFX2_insert350 gnd vdd FILL
XFILL_0__10971_ gnd vdd FILL
XSFILL33960x6050 gnd vdd FILL
XFILL_3_BUFX2_insert361 gnd vdd FILL
XFILL_3_BUFX2_insert372 gnd vdd FILL
XFILL_4__13140_ gnd vdd FILL
X_15954_ _15954_/A _15954_/B gnd _15955_/B vdd NOR2X1
XFILL_5__11711_ gnd vdd FILL
X_11077_ _12254_/Y _11076_/Y gnd _11081_/C vdd NOR2X1
XFILL_3_BUFX2_insert383 gnd vdd FILL
XFILL_3__13870_ gnd vdd FILL
XFILL_0__12710_ gnd vdd FILL
XFILL_2__11531_ gnd vdd FILL
XFILL_4__9109_ gnd vdd FILL
XFILL_2__9173_ gnd vdd FILL
XFILL_1__10172_ gnd vdd FILL
XFILL_3_BUFX2_insert394 gnd vdd FILL
X_10028_ _15797_/A gnd _10028_/Y vdd INVX1
XSFILL69160x28050 gnd vdd FILL
XFILL_0__13690_ gnd vdd FILL
X_14905_ _14904_/Y _14901_/Y gnd _14905_/Y vdd NOR2X1
XFILL_5__11642_ gnd vdd FILL
XFILL_5__14430_ gnd vdd FILL
XFILL_2__8124_ gnd vdd FILL
XFILL_6__13981_ gnd vdd FILL
X_15885_ _14414_/D gnd _15885_/Y vdd INVX1
XFILL_2__14250_ gnd vdd FILL
XFILL_4__10283_ gnd vdd FILL
XFILL_2__11462_ gnd vdd FILL
XFILL_0__12641_ gnd vdd FILL
XFILL_6__15720_ gnd vdd FILL
XFILL_1__14980_ gnd vdd FILL
XSFILL84200x31050 gnd vdd FILL
XFILL_5__9922_ gnd vdd FILL
X_14836_ _8141_/A gnd _14836_/Y vdd INVX1
XFILL_4__12022_ gnd vdd FILL
XFILL_3__15540_ gnd vdd FILL
XFILL_5__14361_ gnd vdd FILL
XFILL_5__11573_ gnd vdd FILL
XFILL_3__12752_ gnd vdd FILL
XFILL_2__8055_ gnd vdd FILL
XSFILL104360x37050 gnd vdd FILL
XFILL_2__10413_ gnd vdd FILL
XFILL_0__15360_ gnd vdd FILL
XFILL_2__14181_ gnd vdd FILL
XFILL_2__11393_ gnd vdd FILL
XFILL_1__13931_ gnd vdd FILL
XFILL_0__12572_ gnd vdd FILL
XFILL_5__16100_ gnd vdd FILL
XFILL_5__9853_ gnd vdd FILL
XFILL_5__13312_ gnd vdd FILL
XFILL_5__10524_ gnd vdd FILL
XFILL_0__7070_ gnd vdd FILL
XFILL_3__11703_ gnd vdd FILL
XSFILL74280x19050 gnd vdd FILL
X_14767_ _8817_/Q gnd _14768_/B vdd INVX1
XFILL_5__14292_ gnd vdd FILL
XFILL_2__13132_ gnd vdd FILL
X_11979_ _11979_/A _11969_/A _11978_/Y gnd _6868_/A vdd OAI21X1
XFILL_0__14311_ gnd vdd FILL
XFILL_3__15471_ gnd vdd FILL
XFILL_0__11523_ gnd vdd FILL
XSFILL79320x5050 gnd vdd FILL
XFILL_1__13862_ gnd vdd FILL
XFILL_0__15291_ gnd vdd FILL
XFILL_5__13243_ gnd vdd FILL
XFILL_5__16031_ gnd vdd FILL
X_13718_ _13718_/A _13718_/B gnd _13883_/B vdd AND2X2
XFILL_5__9784_ gnd vdd FILL
XFILL_6__11814_ gnd vdd FILL
XFILL_5__6996_ gnd vdd FILL
XFILL_6__15582_ gnd vdd FILL
XFILL_3__14422_ gnd vdd FILL
XFILL_4_CLKBUF1_insert140 gnd vdd FILL
X_14698_ _8132_/A gnd _16098_/C vdd INVX1
XFILL_3__11634_ gnd vdd FILL
XFILL_1__15601_ gnd vdd FILL
XFILL112200x13050 gnd vdd FILL
XFILL_2__10275_ gnd vdd FILL
XFILL_0__14242_ gnd vdd FILL
XFILL_4__13973_ gnd vdd FILL
XFILL_0__11454_ gnd vdd FILL
XFILL_5__8735_ gnd vdd FILL
XFILL_4_CLKBUF1_insert151 gnd vdd FILL
XFILL_1__13793_ gnd vdd FILL
XFILL_6__14533_ gnd vdd FILL
XFILL_4_CLKBUF1_insert162 gnd vdd FILL
X_16437_ _14418_/A _7527_/CLK _8935_/R vdd _16437_/D gnd vdd DFFSR
XSFILL74120x83050 gnd vdd FILL
XFILL_4_CLKBUF1_insert173 gnd vdd FILL
XFILL_4__15712_ gnd vdd FILL
X_13649_ _9818_/Q gnd _13649_/Y vdd INVX1
XFILL_5__13174_ gnd vdd FILL
XFILL_2__12014_ gnd vdd FILL
XFILL_4_CLKBUF1_insert184 gnd vdd FILL
XFILL_3__14353_ gnd vdd FILL
XFILL_5__10386_ gnd vdd FILL
XFILL_4_CLKBUF1_insert195 gnd vdd FILL
XFILL_0__10405_ gnd vdd FILL
XFILL_1__15532_ gnd vdd FILL
XFILL_2__8957_ gnd vdd FILL
XFILL_3__11565_ gnd vdd FILL
XFILL_3__7750_ gnd vdd FILL
XFILL_1__12744_ gnd vdd FILL
XFILL_0__14173_ gnd vdd FILL
XFILL_0_BUFX2_insert240 gnd vdd FILL
XFILL_5__12125_ gnd vdd FILL
XFILL_0__11385_ gnd vdd FILL
XFILL_0_BUFX2_insert251 gnd vdd FILL
XFILL_3__13304_ gnd vdd FILL
XFILL_0_BUFX2_insert262 gnd vdd FILL
X_16368_ _16368_/A gnd _16368_/C gnd _16368_/Y vdd OAI21X1
XFILL_0_BUFX2_insert273 gnd vdd FILL
XFILL_0__7972_ gnd vdd FILL
XFILL_4__15643_ gnd vdd FILL
XSFILL13560x36050 gnd vdd FILL
XFILL_6__11676_ gnd vdd FILL
XFILL_4__12855_ gnd vdd FILL
XFILL_3__10516_ gnd vdd FILL
XFILL_0__13124_ gnd vdd FILL
XFILL_3__14284_ gnd vdd FILL
XFILL_3__7681_ gnd vdd FILL
XFILL_2__8888_ gnd vdd FILL
XFILL_0_BUFX2_insert284 gnd vdd FILL
XFILL_5__7617_ gnd vdd FILL
XFILL_1__15463_ gnd vdd FILL
XFILL_3__11496_ gnd vdd FILL
XFILL_0_BUFX2_insert295 gnd vdd FILL
X_15319_ _9864_/A gnd _15321_/D vdd INVX1
XSFILL53960x41050 gnd vdd FILL
X_8250_ _8250_/A _8249_/A _8250_/C gnd _8250_/Y vdd OAI21X1
XFILL_0__6923_ gnd vdd FILL
XFILL_3__16023_ gnd vdd FILL
XFILL_5__12056_ gnd vdd FILL
XFILL_5__8597_ gnd vdd FILL
XFILL_4__11806_ gnd vdd FILL
XFILL_3__13235_ gnd vdd FILL
XFILL_3__9420_ gnd vdd FILL
XFILL_6__14395_ gnd vdd FILL
X_16299_ _15045_/D _14961_/Y _16299_/C gnd _16302_/A vdd OAI21X1
XFILL_4__12786_ gnd vdd FILL
XFILL_3__10447_ gnd vdd FILL
XFILL_2__7839_ gnd vdd FILL
XFILL_4__15574_ gnd vdd FILL
XFILL_1__14414_ gnd vdd FILL
XSFILL94840x53050 gnd vdd FILL
XFILL_1__11626_ gnd vdd FILL
XFILL_2__13965_ gnd vdd FILL
XFILL_1__15394_ gnd vdd FILL
X_7201_ _7202_/B _7713_/B gnd _7201_/Y vdd NAND2X1
XFILL_0__10267_ gnd vdd FILL
XFILL_5__7548_ gnd vdd FILL
XFILL_5__11007_ gnd vdd FILL
XFILL_0__9642_ gnd vdd FILL
XFILL_6__10558_ gnd vdd FILL
XFILL_2__15704_ gnd vdd FILL
XFILL_0__6854_ gnd vdd FILL
XFILL_4__14525_ gnd vdd FILL
X_8181_ _8147_/A _7010_/CLK _7413_/R vdd _8149_/Y gnd vdd DFFSR
XFILL_4__11737_ gnd vdd FILL
XFILL_3__13166_ gnd vdd FILL
XFILL_0__12006_ gnd vdd FILL
XFILL_2__12916_ gnd vdd FILL
XFILL_3__9351_ gnd vdd FILL
XFILL_2_BUFX2_insert11 gnd vdd FILL
XFILL_3__10378_ gnd vdd FILL
XFILL_1__14345_ gnd vdd FILL
XFILL_1__11557_ gnd vdd FILL
XFILL_2__13896_ gnd vdd FILL
XFILL_2_BUFX2_insert22 gnd vdd FILL
XFILL_5__7479_ gnd vdd FILL
X_7132_ _7048_/A _7534_/CLK _8156_/R vdd _7050_/Y gnd vdd DFFSR
XFILL_5__15815_ gnd vdd FILL
XFILL_2_BUFX2_insert33 gnd vdd FILL
XFILL_2__9509_ gnd vdd FILL
XFILL_4__14456_ gnd vdd FILL
XFILL_3__12117_ gnd vdd FILL
XFILL_1__10508_ gnd vdd FILL
XFILL_2__15635_ gnd vdd FILL
XFILL_2_BUFX2_insert44 gnd vdd FILL
XFILL_4__11668_ gnd vdd FILL
XFILL_2_BUFX2_insert55 gnd vdd FILL
XFILL_5__9218_ gnd vdd FILL
XFILL_2__12847_ gnd vdd FILL
XFILL_3__13097_ gnd vdd FILL
XFILL_3__9282_ gnd vdd FILL
XSFILL8680x15050 gnd vdd FILL
XFILL_2_BUFX2_insert66 gnd vdd FILL
XFILL_1__11488_ gnd vdd FILL
XFILL_1__14276_ gnd vdd FILL
XFILL_4__13407_ gnd vdd FILL
XFILL_2_BUFX2_insert77 gnd vdd FILL
XFILL_0__8524_ gnd vdd FILL
XFILL_2_BUFX2_insert88 gnd vdd FILL
X_7063_ _7137_/Q gnd _7065_/A vdd INVX1
XFILL_5__15746_ gnd vdd FILL
XFILL_4__10619_ gnd vdd FILL
XFILL_1__16015_ gnd vdd FILL
XFILL_3__12048_ gnd vdd FILL
XFILL_4__14387_ gnd vdd FILL
XFILL_5__12958_ gnd vdd FILL
XFILL_3__8233_ gnd vdd FILL
XFILL_1__13227_ gnd vdd FILL
XFILL_2__15566_ gnd vdd FILL
XFILL_2_BUFX2_insert99 gnd vdd FILL
XFILL_1__10439_ gnd vdd FILL
XFILL_4__11599_ gnd vdd FILL
XFILL_5__9149_ gnd vdd FILL
XFILL_2__12778_ gnd vdd FILL
XFILL_0__13957_ gnd vdd FILL
XFILL_4__13338_ gnd vdd FILL
XFILL_5__11909_ gnd vdd FILL
XFILL_4__16126_ gnd vdd FILL
XFILL_0__8455_ gnd vdd FILL
XFILL_5__15677_ gnd vdd FILL
XFILL_2__14517_ gnd vdd FILL
XSFILL48920x30050 gnd vdd FILL
XFILL_1__13158_ gnd vdd FILL
XFILL_5__12889_ gnd vdd FILL
XFILL_2__11729_ gnd vdd FILL
XSFILL74200x63050 gnd vdd FILL
XFILL_0__12908_ gnd vdd FILL
XFILL_2__15497_ gnd vdd FILL
XFILL_5__14628_ gnd vdd FILL
XFILL_0__13888_ gnd vdd FILL
XFILL_4__16057_ gnd vdd FILL
XFILL_3__7115_ gnd vdd FILL
XFILL_4__13269_ gnd vdd FILL
XFILL_1__12109_ gnd vdd FILL
XFILL_3__15807_ gnd vdd FILL
XFILL_0__8386_ gnd vdd FILL
XFILL_2__14448_ gnd vdd FILL
XFILL_1__13089_ gnd vdd FILL
XFILL_0__15627_ gnd vdd FILL
XFILL_3__13999_ gnd vdd FILL
XFILL_3__8095_ gnd vdd FILL
XFILL_4__15008_ gnd vdd FILL
XFILL_0__12839_ gnd vdd FILL
XSFILL13640x16050 gnd vdd FILL
XFILL_6__8913_ gnd vdd FILL
XFILL_0__7337_ gnd vdd FILL
XFILL_5__14559_ gnd vdd FILL
XFILL_3__15738_ gnd vdd FILL
X_7965_ _8035_/Q gnd _7967_/A vdd INVX1
XFILL_3__7046_ gnd vdd FILL
XFILL_2__14379_ gnd vdd FILL
XFILL_0__15558_ gnd vdd FILL
XSFILL109560x50050 gnd vdd FILL
X_9704_ _9644_/A _7400_/CLK _9704_/R vdd _9704_/D gnd vdd DFFSR
X_6916_ _6916_/A _6967_/B _6915_/Y gnd _7002_/D vdd OAI21X1
XFILL_2__16118_ gnd vdd FILL
XFILL_3__15669_ gnd vdd FILL
XSFILL38840x82050 gnd vdd FILL
XFILL_0__14509_ gnd vdd FILL
X_7896_ _7804_/A _8792_/CLK _7896_/R vdd _7806_/Y gnd vdd DFFSR
XFILL_0__9007_ gnd vdd FILL
XFILL_5__16229_ gnd vdd FILL
XSFILL54120x30050 gnd vdd FILL
XFILL_0__15489_ gnd vdd FILL
X_9635_ _9701_/Q gnd _9635_/Y vdd INVX1
XFILL_0__7199_ gnd vdd FILL
X_6847_ _6847_/A gnd memoryAddress[9] vdd BUFX2
XFILL_2__16049_ gnd vdd FILL
XFILL_3__8997_ gnd vdd FILL
XSFILL33800x29050 gnd vdd FILL
X_9566_ _9566_/Q _7790_/CLK _9566_/R vdd _9566_/D gnd vdd DFFSR
XFILL_5_BUFX2_insert401 gnd vdd FILL
XFILL_3__7948_ gnd vdd FILL
XFILL_5_BUFX2_insert412 gnd vdd FILL
XSFILL43960x73050 gnd vdd FILL
XFILL_5_BUFX2_insert423 gnd vdd FILL
XFILL_5_BUFX2_insert434 gnd vdd FILL
XFILL_1__9751_ gnd vdd FILL
X_8517_ _8460_/A _9413_/B gnd _8518_/C vdd NAND2X1
XSFILL28760x7050 gnd vdd FILL
XFILL_5_BUFX2_insert445 gnd vdd FILL
XFILL_1__6963_ gnd vdd FILL
X_9497_ _9495_/Y _9533_/B _9497_/C gnd _9497_/Y vdd OAI21X1
XFILL_5_BUFX2_insert456 gnd vdd FILL
XFILL_5_BUFX2_insert467 gnd vdd FILL
XFILL_3__7879_ gnd vdd FILL
XFILL_0__9909_ gnd vdd FILL
XFILL_5_BUFX2_insert478 gnd vdd FILL
XFILL_1__8702_ gnd vdd FILL
XFILL_5_BUFX2_insert489 gnd vdd FILL
XSFILL44040x82050 gnd vdd FILL
X_8448_ _8508_/A _9344_/B gnd _8449_/C vdd NAND2X1
XFILL_3__9618_ gnd vdd FILL
XFILL_1__9682_ gnd vdd FILL
XFILL_1__6894_ gnd vdd FILL
XFILL_4__9391_ gnd vdd FILL
XFILL_1__8633_ gnd vdd FILL
X_8379_ _8379_/A gnd _8381_/A vdd INVX1
XFILL_3__9549_ gnd vdd FILL
XFILL_4__8342_ gnd vdd FILL
XSFILL43960x1050 gnd vdd FILL
XFILL112040x48050 gnd vdd FILL
X_11000_ _12230_/Y _10999_/Y gnd _11006_/C vdd NOR2X1
XFILL_4__8273_ gnd vdd FILL
XFILL_4__7224_ gnd vdd FILL
XFILL_1__8495_ gnd vdd FILL
XSFILL79000x55050 gnd vdd FILL
XFILL_1__7446_ gnd vdd FILL
XFILL_2_BUFX2_insert302 gnd vdd FILL
XSFILL39000x71050 gnd vdd FILL
XFILL_2_BUFX2_insert313 gnd vdd FILL
XFILL_2_BUFX2_insert324 gnd vdd FILL
X_12951_ _6870_/A gnd _12951_/Y vdd INVX1
XFILL_2_BUFX2_insert335 gnd vdd FILL
XFILL_1__7377_ gnd vdd FILL
XFILL_2_BUFX2_insert346 gnd vdd FILL
XFILL_2_BUFX2_insert357 gnd vdd FILL
X_11902_ _13180_/Q gnd _11902_/Y vdd INVX1
XFILL_4__7086_ gnd vdd FILL
XFILL_2_BUFX2_insert368 gnd vdd FILL
X_15670_ _10853_/Q gnd _15670_/Y vdd INVX1
XFILL_1__9116_ gnd vdd FILL
X_12882_ _12880_/Y vdd _12882_/C gnd _12938_/D vdd OAI21X1
XFILL_2_BUFX2_insert379 gnd vdd FILL
X_14621_ _14211_/A _14620_/Y _13587_/C _14619_/Y gnd _14625_/A vdd OAI22X1
X_11833_ _11374_/Y _11848_/A _11846_/C _11011_/Y gnd _11834_/A vdd AOI22X1
XFILL_5__6850_ gnd vdd FILL
X_14552_ _14551_/Y _13876_/B _13876_/C _14550_/Y gnd _14552_/Y vdd OAI22X1
X_11764_ _11764_/A _11245_/Y _11018_/Y _11764_/D gnd _11772_/A vdd AOI22X1
XFILL_2__9860_ gnd vdd FILL
XBUFX2_insert301 _12414_/Y gnd _8636_/B vdd BUFX2
XBUFX2_insert312 _11222_/Y gnd _11495_/C vdd BUFX2
X_13503_ _13493_/Y _13503_/B _13503_/C gnd _13503_/Y vdd NAND3X1
XFILL_5__10240_ gnd vdd FILL
XFILL112120x28050 gnd vdd FILL
X_10715_ _13702_/A _8792_/CLK _7896_/R vdd _10715_/D gnd vdd DFFSR
XFILL_4__7988_ gnd vdd FILL
X_14483_ _14483_/A _14482_/Y _14483_/C gnd _14483_/Y vdd NAND3X1
XBUFX2_insert323 _13345_/Y gnd _9902_/B vdd BUFX2
XFILL_4__10970_ gnd vdd FILL
XFILL_2__10060_ gnd vdd FILL
XBUFX2_insert334 _13494_/Y gnd _13848_/B vdd BUFX2
X_11695_ _11065_/Y _11681_/B _11764_/A _11046_/Y gnd _11695_/Y vdd AOI22X1
XFILL_2__9791_ gnd vdd FILL
XFILL_5__8520_ gnd vdd FILL
XFILL_6_BUFX2_insert290 gnd vdd FILL
XBUFX2_insert345 _12396_/Y gnd _9258_/B vdd BUFX2
XSFILL64040x13050 gnd vdd FILL
XFILL_4__9727_ gnd vdd FILL
X_16222_ _9203_/Q gnd _16222_/Y vdd INVX1
XBUFX2_insert356 _13306_/Y gnd _7972_/A vdd BUFX2
XFILL_1__10790_ gnd vdd FILL
XFILL_4__6939_ gnd vdd FILL
X_13434_ _7158_/A _13434_/B _13434_/C gnd _13451_/A vdd AOI21X1
XBUFX2_insert367 _13487_/Y gnd _14344_/C vdd BUFX2
XFILL_5__10171_ gnd vdd FILL
XSFILL89640x77050 gnd vdd FILL
XFILL_5_CLKBUF1_insert202 gnd vdd FILL
X_10646_ _10646_/A _10681_/A _10645_/Y gnd _10646_/Y vdd OAI21X1
XFILL_2__8742_ gnd vdd FILL
XBUFX2_insert378 _12211_/Y gnd _12319_/C vdd BUFX2
XFILL_3__11350_ gnd vdd FILL
XBUFX2_insert389 _12387_/Y gnd _9633_/B vdd BUFX2
XFILL_5_CLKBUF1_insert213 gnd vdd FILL
XFILL_5_CLKBUF1_insert224 gnd vdd FILL
XFILL_5__8451_ gnd vdd FILL
XFILL_4__9658_ gnd vdd FILL
XFILL_0__11170_ gnd vdd FILL
X_16153_ _16153_/A _16152_/Y gnd _16163_/A vdd NAND2X1
X_13365_ _13326_/A _13365_/B gnd _13365_/Y vdd NOR2X1
XFILL_4__12640_ gnd vdd FILL
XFILL_3__10301_ gnd vdd FILL
XFILL_6__11461_ gnd vdd FILL
X_10577_ _10548_/B _8273_/B gnd _10577_/Y vdd NAND2X1
XFILL_0__10121_ gnd vdd FILL
XFILL_1__12460_ gnd vdd FILL
XFILL_4__8609_ gnd vdd FILL
XFILL_3__11281_ gnd vdd FILL
XFILL_5_BUFX2_insert990 gnd vdd FILL
X_15104_ _16141_/A _13496_/Y _16141_/C gnd _15104_/Y vdd NOR3X1
XFILL_5__8382_ gnd vdd FILL
X_12316_ _12224_/A _12308_/B _12224_/C gnd _12318_/B vdd NAND3X1
XFILL_3__13020_ gnd vdd FILL
XFILL_6__14180_ gnd vdd FILL
X_16084_ _16084_/A _16084_/B gnd _16085_/B vdd NOR2X1
XFILL_5__13930_ gnd vdd FILL
X_13296_ _13295_/Y _13290_/Y gnd _13296_/Y vdd NAND2X1
XFILL_4__12571_ gnd vdd FILL
XFILL_3__10232_ gnd vdd FILL
XFILL_2__7624_ gnd vdd FILL
XFILL_1__11411_ gnd vdd FILL
XSFILL68920x78050 gnd vdd FILL
XFILL_2__13750_ gnd vdd FILL
XFILL_2__10962_ gnd vdd FILL
XFILL_5__7333_ gnd vdd FILL
XFILL_1__12391_ gnd vdd FILL
XFILL_0__10052_ gnd vdd FILL
X_15035_ _15064_/A _15035_/B _15035_/C gnd _15035_/Y vdd OAI21X1
XFILL_4__14310_ gnd vdd FILL
XSFILL84200x26050 gnd vdd FILL
X_12247_ _12255_/A gnd _12255_/C gnd _12247_/Y vdd NAND3X1
XFILL_4__11522_ gnd vdd FILL
XFILL_2__12701_ gnd vdd FILL
XFILL_5__13861_ gnd vdd FILL
XFILL_4__15290_ gnd vdd FILL
XSFILL94360x70050 gnd vdd FILL
XFILL_2__7555_ gnd vdd FILL
XFILL_1__14130_ gnd vdd FILL
XFILL_3__10163_ gnd vdd FILL
XFILL_1__11342_ gnd vdd FILL
XFILL_2__13681_ gnd vdd FILL
XFILL_0__14860_ gnd vdd FILL
XFILL_2__10893_ gnd vdd FILL
XFILL_5__15600_ gnd vdd FILL
XFILL_4__14241_ gnd vdd FILL
XFILL_6__10274_ gnd vdd FILL
X_12178_ _13196_/Q gnd _12178_/Y vdd INVX1
XFILL_4__11453_ gnd vdd FILL
XFILL_2__15420_ gnd vdd FILL
XFILL_2__12632_ gnd vdd FILL
XFILL_5__13792_ gnd vdd FILL
XFILL_1__14061_ gnd vdd FILL
XFILL_3__14971_ gnd vdd FILL
XFILL_5__9003_ gnd vdd FILL
XFILL_0__13811_ gnd vdd FILL
XFILL_2__7486_ gnd vdd FILL
XFILL_1__11273_ gnd vdd FILL
XFILL_0__14791_ gnd vdd FILL
XFILL_4__10404_ gnd vdd FILL
XFILL_5__15531_ gnd vdd FILL
XFILL_5__7195_ gnd vdd FILL
X_11129_ _11590_/A _11591_/C gnd _11129_/Y vdd NAND2X1
XFILL_5__12743_ gnd vdd FILL
XFILL_4__14172_ gnd vdd FILL
XFILL_2__9225_ gnd vdd FILL
XFILL_3__13922_ gnd vdd FILL
XFILL_1__13012_ gnd vdd FILL
XFILL_2__15351_ gnd vdd FILL
XFILL_4__11384_ gnd vdd FILL
XFILL_0__10954_ gnd vdd FILL
XFILL_0__13742_ gnd vdd FILL
XFILL_4__13123_ gnd vdd FILL
XFILL_0__8240_ gnd vdd FILL
X_15937_ _15322_/A _14524_/A _15937_/C _15322_/D gnd _15937_/Y vdd OAI22X1
XFILL_5__15462_ gnd vdd FILL
XFILL_2__14302_ gnd vdd FILL
XFILL_3__13853_ gnd vdd FILL
XSFILL34680x51050 gnd vdd FILL
XFILL_2__9156_ gnd vdd FILL
XFILL_2__11514_ gnd vdd FILL
XFILL_1__10155_ gnd vdd FILL
XFILL_2__15282_ gnd vdd FILL
XFILL_0__13673_ gnd vdd FILL
XFILL_2__12494_ gnd vdd FILL
XFILL_0__10885_ gnd vdd FILL
XFILL_5__14413_ gnd vdd FILL
X_15868_ _7402_/Q _15631_/B _15945_/C gnd _15869_/C vdd NAND3X1
XFILL_5__11625_ gnd vdd FILL
XFILL_2__8107_ gnd vdd FILL
XFILL_5__15393_ gnd vdd FILL
XFILL_2__14233_ gnd vdd FILL
XFILL_4__10266_ gnd vdd FILL
XFILL_2__9087_ gnd vdd FILL
XFILL_0__15412_ gnd vdd FILL
XFILL_0__12624_ gnd vdd FILL
XFILL_3__13784_ gnd vdd FILL
XFILL_2_BUFX2_insert880 gnd vdd FILL
XFILL_2__11445_ gnd vdd FILL
XFILL_5__9905_ gnd vdd FILL
XFILL_1__14963_ gnd vdd FILL
XFILL_3__10996_ gnd vdd FILL
XFILL_2_BUFX2_insert891 gnd vdd FILL
X_14819_ _14815_/Y _14818_/Y gnd _14819_/Y vdd NOR2X1
XFILL_4__12005_ gnd vdd FILL
XFILL_0__16392_ gnd vdd FILL
XFILL_0__7122_ gnd vdd FILL
XFILL_3__15523_ gnd vdd FILL
XSFILL53960x36050 gnd vdd FILL
XFILL_5__14344_ gnd vdd FILL
XFILL_5__11556_ gnd vdd FILL
XFILL_3__12735_ gnd vdd FILL
X_15799_ _15795_/Y _15799_/B gnd _15799_/Y vdd NOR2X1
X_7750_ _7750_/A _7729_/B _7749_/Y gnd _7750_/Y vdd OAI21X1
XFILL_2__14164_ gnd vdd FILL
XFILL_4__10197_ gnd vdd FILL
XFILL_1__13914_ gnd vdd FILL
XFILL_0__15343_ gnd vdd FILL
XFILL_2__11376_ gnd vdd FILL
XFILL_5__10507_ gnd vdd FILL
XFILL_0__7053_ gnd vdd FILL
XFILL_1__14894_ gnd vdd FILL
XFILL_6__12846_ gnd vdd FILL
X_7681_ _7681_/A _7744_/B _7680_/Y gnd _7769_/D vdd OAI21X1
XFILL_2__13115_ gnd vdd FILL
XFILL_5__11487_ gnd vdd FILL
XFILL_3__15454_ gnd vdd FILL
XFILL_5__14275_ gnd vdd FILL
XSFILL54040x45050 gnd vdd FILL
XFILL_3__8851_ gnd vdd FILL
XFILL_0__11506_ gnd vdd FILL
XFILL_1__13845_ gnd vdd FILL
XFILL_4_BUFX2_insert1 gnd vdd FILL
XFILL_2__14095_ gnd vdd FILL
XFILL_0__15274_ gnd vdd FILL
XFILL_5__16014_ gnd vdd FILL
XFILL_0__12486_ gnd vdd FILL
XFILL_5__9767_ gnd vdd FILL
XFILL_5__13226_ gnd vdd FILL
X_9420_ _9418_/Y _9420_/B _9420_/C gnd _9458_/D vdd OAI21X1
XSFILL94440x50050 gnd vdd FILL
XFILL_5__10438_ gnd vdd FILL
XFILL_3__14405_ gnd vdd FILL
XFILL_5__6979_ gnd vdd FILL
XFILL_3__7802_ gnd vdd FILL
XFILL_3__11617_ gnd vdd FILL
XFILL_3__15385_ gnd vdd FILL
XFILL_0__14225_ gnd vdd FILL
XFILL_2__13046_ gnd vdd FILL
XFILL_2__10258_ gnd vdd FILL
XFILL_4__13956_ gnd vdd FILL
XFILL_3__8782_ gnd vdd FILL
XFILL_3__12597_ gnd vdd FILL
XFILL_0__11437_ gnd vdd FILL
XFILL_2__9989_ gnd vdd FILL
XFILL_5__8718_ gnd vdd FILL
XFILL_1__13776_ gnd vdd FILL
XFILL_5__13157_ gnd vdd FILL
XFILL_1__10988_ gnd vdd FILL
XFILL_5__10369_ gnd vdd FILL
XFILL_4__12907_ gnd vdd FILL
XFILL_3__14336_ gnd vdd FILL
X_9351_ _9351_/A _9339_/B _9351_/C gnd _9351_/Y vdd OAI21X1
XFILL_3__7733_ gnd vdd FILL
XFILL_1__15515_ gnd vdd FILL
XFILL_3__11548_ gnd vdd FILL
XFILL_2__10189_ gnd vdd FILL
XFILL_1__12727_ gnd vdd FILL
XFILL_4__13887_ gnd vdd FILL
XFILL_0__14156_ gnd vdd FILL
XBUFX2_insert890 _12369_/Y gnd _8719_/B vdd BUFX2
XFILL_5__8649_ gnd vdd FILL
XFILL_0__11368_ gnd vdd FILL
X_8302_ _8254_/A _7790_/CLK _9566_/R vdd _8302_/D gnd vdd DFFSR
XFILL_5__12108_ gnd vdd FILL
XFILL_6__14447_ gnd vdd FILL
XFILL_5__13088_ gnd vdd FILL
XFILL_4__15626_ gnd vdd FILL
X_9282_ _9282_/A _9282_/B gnd _9283_/C vdd NAND2X1
XFILL_0__7955_ gnd vdd FILL
XFILL_0__13107_ gnd vdd FILL
XFILL_4__12838_ gnd vdd FILL
XFILL_3__14267_ gnd vdd FILL
XSFILL48920x25050 gnd vdd FILL
XFILL_0__10319_ gnd vdd FILL
XFILL_4_BUFX2_insert408 gnd vdd FILL
XSFILL18680x64050 gnd vdd FILL
XFILL_1__15446_ gnd vdd FILL
XFILL_3__11479_ gnd vdd FILL
XFILL_1__12658_ gnd vdd FILL
XFILL_2__14997_ gnd vdd FILL
XFILL_4_BUFX2_insert419 gnd vdd FILL
XFILL_0__14087_ gnd vdd FILL
XFILL_3__16006_ gnd vdd FILL
XFILL_6__7373_ gnd vdd FILL
XFILL_5__12039_ gnd vdd FILL
XFILL_0__6906_ gnd vdd FILL
XFILL_0__11299_ gnd vdd FILL
X_8233_ _8233_/A gnd _8233_/Y vdd INVX1
XFILL_3__13218_ gnd vdd FILL
XFILL_3__9403_ gnd vdd FILL
XFILL_0__7886_ gnd vdd FILL
XFILL_4__12769_ gnd vdd FILL
XFILL_4__15557_ gnd vdd FILL
XFILL_3__14198_ gnd vdd FILL
XFILL_0__13038_ gnd vdd FILL
XFILL_1__11609_ gnd vdd FILL
XFILL_2__13948_ gnd vdd FILL
XFILL_1__15377_ gnd vdd FILL
XFILL_3__7595_ gnd vdd FILL
XFILL_1__12589_ gnd vdd FILL
XFILL_0__9625_ gnd vdd FILL
XSFILL49000x34050 gnd vdd FILL
XFILL_0__6837_ gnd vdd FILL
X_8164_ _8096_/A _7268_/CLK _8688_/R vdd _8098_/Y gnd vdd DFFSR
XFILL_4__14508_ gnd vdd FILL
XFILL_3__13149_ gnd vdd FILL
XFILL_3__9334_ gnd vdd FILL
XFILL_1__14328_ gnd vdd FILL
XFILL_4__15488_ gnd vdd FILL
XFILL_2__13879_ gnd vdd FILL
XFILL_6__9043_ gnd vdd FILL
X_7115_ _7055_/A _7499_/B gnd _7116_/C vdd NAND2X1
XFILL_6__16048_ gnd vdd FILL
XSFILL109560x45050 gnd vdd FILL
XFILL_0__9556_ gnd vdd FILL
XFILL_2__15618_ gnd vdd FILL
X_8095_ _8095_/A _8082_/A _8095_/C gnd _8163_/D vdd OAI21X1
XFILL_4__14439_ gnd vdd FILL
XFILL_3__9265_ gnd vdd FILL
XFILL_1__14259_ gnd vdd FILL
XFILL_0__8507_ gnd vdd FILL
XFILL_1__7300_ gnd vdd FILL
XSFILL79480x27050 gnd vdd FILL
XFILL_5__15729_ gnd vdd FILL
XFILL_0__14989_ gnd vdd FILL
X_7046_ _7067_/A _9094_/B gnd _7046_/Y vdd NAND2X1
XSFILL54120x25050 gnd vdd FILL
XFILL_0__9487_ gnd vdd FILL
XFILL_3__8216_ gnd vdd FILL
XFILL_2__15549_ gnd vdd FILL
XSFILL39480x43050 gnd vdd FILL
XFILL_1__7231_ gnd vdd FILL
XFILL_0__8438_ gnd vdd FILL
XFILL_4__16109_ gnd vdd FILL
XFILL_3__8147_ gnd vdd FILL
XSFILL43960x68050 gnd vdd FILL
XFILL_0__8369_ gnd vdd FILL
XFILL_1__7162_ gnd vdd FILL
XSFILL83560x54050 gnd vdd FILL
XFILL_4__8960_ gnd vdd FILL
XFILL_3__8078_ gnd vdd FILL
X_8997_ _8997_/A _8996_/A _8997_/C gnd _8997_/Y vdd OAI21X1
XFILL_1_BUFX2_insert309 gnd vdd FILL
XSFILL18760x44050 gnd vdd FILL
XFILL_1__7093_ gnd vdd FILL
X_7948_ _7948_/A _7948_/B gnd _7948_/Y vdd NAND2X1
XSFILL8600x54050 gnd vdd FILL
XSFILL44040x77050 gnd vdd FILL
XFILL_4__8891_ gnd vdd FILL
XFILL_4__7842_ gnd vdd FILL
X_7879_ _7921_/Q gnd _7881_/A vdd INVX1
X_9618_ _9652_/B _8466_/B gnd _9619_/C vdd NAND2X1
XSFILL23880x35050 gnd vdd FILL
X_10500_ _10500_/A _10500_/B _10499_/Y gnd _10500_/Y vdd OAI21X1
XFILL_1__9803_ gnd vdd FILL
X_11480_ _11480_/A _11191_/A _11480_/C gnd _11480_/Y vdd NAND3X1
X_9549_ _9587_/Q gnd _9551_/A vdd INVX1
XFILL_4__9512_ gnd vdd FILL
XSFILL38920x57050 gnd vdd FILL
XFILL_5_BUFX2_insert231 gnd vdd FILL
XFILL_1__7995_ gnd vdd FILL
XFILL_5_BUFX2_insert242 gnd vdd FILL
XFILL112440x64050 gnd vdd FILL
XFILL_5_BUFX2_insert253 gnd vdd FILL
X_10431_ _10405_/B _8511_/B gnd _10432_/C vdd NAND2X1
XFILL_5_BUFX2_insert264 gnd vdd FILL
XFILL_1__9734_ gnd vdd FILL
XFILL_1__6946_ gnd vdd FILL
XFILL_5_BUFX2_insert275 gnd vdd FILL
XFILL_5_BUFX2_insert286 gnd vdd FILL
XFILL_5_BUFX2_insert297 gnd vdd FILL
XSFILL39000x66050 gnd vdd FILL
X_13150_ _13150_/A _13149_/A _13150_/C gnd _13150_/Y vdd OAI21X1
XFILL_4_BUFX2_insert920 gnd vdd FILL
X_10362_ _10363_/B _6906_/B gnd _10362_/Y vdd NAND2X1
XFILL_1__9665_ gnd vdd FILL
XFILL_4_BUFX2_insert931 gnd vdd FILL
XFILL_1__6877_ gnd vdd FILL
XSFILL114200x59050 gnd vdd FILL
X_12101_ _12101_/A _12073_/B _12073_/C gnd gnd _12102_/C vdd AOI22X1
XFILL_4_BUFX2_insert942 gnd vdd FILL
XFILL_4__9374_ gnd vdd FILL
XFILL_4_BUFX2_insert953 gnd vdd FILL
X_10293_ _10293_/A gnd _10295_/A vdd INVX1
XFILL_1__8616_ gnd vdd FILL
X_13081_ _13081_/A _13153_/B _13080_/Y gnd _13175_/D vdd OAI21X1
XFILL_4_BUFX2_insert964 gnd vdd FILL
XFILL_4_BUFX2_insert975 gnd vdd FILL
XFILL_4_BUFX2_insert986 gnd vdd FILL
XFILL_1__9596_ gnd vdd FILL
XFILL_4__8325_ gnd vdd FILL
XSFILL18840x24050 gnd vdd FILL
XSFILL69480x59050 gnd vdd FILL
X_12032_ _12028_/A _12800_/Q _12024_/C gnd _12032_/Y vdd NAND3X1
XFILL_4_BUFX2_insert997 gnd vdd FILL
XSFILL114600x80050 gnd vdd FILL
XFILL_2__7340_ gnd vdd FILL
XFILL_4__8256_ gnd vdd FILL
XFILL_4__7207_ gnd vdd FILL
XFILL_1__8478_ gnd vdd FILL
XFILL_4__8187_ gnd vdd FILL
XFILL_2__9010_ gnd vdd FILL
XFILL_2_BUFX2_insert110 gnd vdd FILL
X_13983_ _13983_/A gnd _13985_/D vdd INVX1
XFILL_1__7429_ gnd vdd FILL
X_15722_ _14252_/D gnd _15724_/A vdd INVX1
XFILL_4__10120_ gnd vdd FILL
X_12934_ _12934_/Q _9060_/CLK _7140_/R vdd _12934_/D gnd vdd DFFSR
XFILL_5__7951_ gnd vdd FILL
XFILL_0__10670_ gnd vdd FILL
XFILL_4__7069_ gnd vdd FILL
XFILL_5__11410_ gnd vdd FILL
X_15653_ _9123_/A gnd _15654_/A vdd INVX1
XFILL_6__10961_ gnd vdd FILL
XFILL_5__12390_ gnd vdd FILL
X_12865_ _12865_/A gnd _12865_/Y vdd INVX1
XFILL_4__10051_ gnd vdd FILL
XFILL_1_BUFX2_insert810 gnd vdd FILL
XFILL_1_BUFX2_insert821 gnd vdd FILL
XFILL_2__11230_ gnd vdd FILL
XFILL_5__6902_ gnd vdd FILL
XFILL_3__10781_ gnd vdd FILL
X_14604_ _14604_/A _14600_/Y gnd _14604_/Y vdd NOR2X1
XFILL_1__11960_ gnd vdd FILL
XFILL_1_BUFX2_insert832 gnd vdd FILL
XFILL_5__7882_ gnd vdd FILL
XFILL_1_BUFX2_insert843 gnd vdd FILL
X_11816_ _11015_/A _11240_/Y _11376_/A gnd _11816_/Y vdd AOI21X1
XFILL_5__11341_ gnd vdd FILL
XFILL_1_BUFX2_insert854 gnd vdd FILL
XFILL_3__12520_ gnd vdd FILL
XSFILL99960x7050 gnd vdd FILL
X_15584_ _8349_/A _15978_/B _16212_/A _8675_/Q gnd _15585_/B vdd AOI22X1
X_12796_ _12710_/A _12538_/CLK _12795_/R vdd _12796_/D gnd vdd DFFSR
XFILL_2__9912_ gnd vdd FILL
XFILL_2__11161_ gnd vdd FILL
XFILL_1_BUFX2_insert865 gnd vdd FILL
XSFILL3720x77050 gnd vdd FILL
XFILL_1__10911_ gnd vdd FILL
XFILL_1_BUFX2_insert876 gnd vdd FILL
XFILL_0__12340_ gnd vdd FILL
XFILL_5__9621_ gnd vdd FILL
XFILL_1_BUFX2_insert887 gnd vdd FILL
XFILL_5__14060_ gnd vdd FILL
X_14535_ _14535_/A _14045_/A _13868_/B _14533_/Y gnd _14536_/A vdd OAI22X1
XFILL_1__11891_ gnd vdd FILL
XFILL_2__10112_ gnd vdd FILL
XFILL_4__13810_ gnd vdd FILL
XFILL_1_BUFX2_insert898 gnd vdd FILL
XFILL_5__11272_ gnd vdd FILL
X_11747_ _11745_/Y _11366_/B _11746_/Y gnd _11749_/C vdd OAI21X1
XFILL_3__12451_ gnd vdd FILL
XFILL_1__13630_ gnd vdd FILL
XFILL_2__11092_ gnd vdd FILL
XFILL_4__14790_ gnd vdd FILL
XSFILL94360x65050 gnd vdd FILL
XSFILL44200x37050 gnd vdd FILL
XFILL_0__12271_ gnd vdd FILL
XFILL_5__9552_ gnd vdd FILL
XFILL_5__13011_ gnd vdd FILL
X_14466_ _14465_/Y _14865_/B _14466_/C _14464_/Y gnd _14466_/Y vdd OAI22X1
XFILL_3__11402_ gnd vdd FILL
XFILL_4__10953_ gnd vdd FILL
XFILL_2__10043_ gnd vdd FILL
XFILL_3__15170_ gnd vdd FILL
XFILL_4__13741_ gnd vdd FILL
XFILL_0__14010_ gnd vdd FILL
X_11678_ _11678_/A _11045_/Y gnd _11678_/Y vdd OR2X2
XFILL_2__14920_ gnd vdd FILL
XFILL_5__8503_ gnd vdd FILL
XFILL_3__12382_ gnd vdd FILL
XFILL_2__9774_ gnd vdd FILL
XFILL_0__11222_ gnd vdd FILL
X_16205_ _15978_/C _8525_/A _8269_/A _16014_/C gnd _16210_/B vdd AOI22X1
XFILL_2__6986_ gnd vdd FILL
XFILL_1__13561_ gnd vdd FILL
XFILL_1__10773_ gnd vdd FILL
XFILL_5__9483_ gnd vdd FILL
X_13417_ _7894_/Q gnd _13417_/Y vdd INVX1
XFILL_5__10154_ gnd vdd FILL
X_10629_ _13702_/A gnd _10629_/Y vdd INVX1
XFILL_3__14121_ gnd vdd FILL
XFILL_1__15300_ gnd vdd FILL
XFILL_4__13672_ gnd vdd FILL
X_14397_ _14393_/Y _14397_/B gnd _14400_/C vdd NOR2X1
XFILL_2__8725_ gnd vdd FILL
XFILL_3__11333_ gnd vdd FILL
XFILL_2__14851_ gnd vdd FILL
XFILL_1__12512_ gnd vdd FILL
XFILL_4__10884_ gnd vdd FILL
XFILL_0__11153_ gnd vdd FILL
XFILL_1__16280_ gnd vdd FILL
XFILL_6__14232_ gnd vdd FILL
XFILL_1__13492_ gnd vdd FILL
X_16136_ _8433_/Q gnd _16137_/A vdd INVX1
XFILL_0__7740_ gnd vdd FILL
XFILL_4__12623_ gnd vdd FILL
X_13348_ _13347_/Y _13226_/B gnd _13348_/Y vdd OR2X2
XFILL_4__15411_ gnd vdd FILL
XFILL_2__13802_ gnd vdd FILL
XSFILL104360x50050 gnd vdd FILL
XFILL_3__14052_ gnd vdd FILL
XFILL_5__14962_ gnd vdd FILL
XSFILL99400x9050 gnd vdd FILL
XFILL_1__15231_ gnd vdd FILL
XFILL_0__10104_ gnd vdd FILL
XFILL_4__16391_ gnd vdd FILL
XFILL_3__11264_ gnd vdd FILL
XFILL_2__8656_ gnd vdd FILL
XFILL_1__12443_ gnd vdd FILL
XFILL_2__14782_ gnd vdd FILL
XFILL_0__15961_ gnd vdd FILL
XFILL_2__11994_ gnd vdd FILL
XFILL_5__8365_ gnd vdd FILL
XFILL_0__11084_ gnd vdd FILL
XFILL_3__13003_ gnd vdd FILL
X_16067_ _16066_/Y _16059_/Y gnd _16087_/B vdd NOR2X1
XFILL_5__13913_ gnd vdd FILL
X_13279_ _13297_/A _13279_/B gnd _13280_/B vdd OR2X2
XFILL_2__7607_ gnd vdd FILL
XFILL_4__15342_ gnd vdd FILL
XFILL_0__7671_ gnd vdd FILL
XFILL_2__13733_ gnd vdd FILL
XFILL_5__14893_ gnd vdd FILL
XFILL_2__8587_ gnd vdd FILL
XFILL_2__10945_ gnd vdd FILL
XFILL_1__12374_ gnd vdd FILL
XFILL_3__7380_ gnd vdd FILL
XFILL_0__10035_ gnd vdd FILL
XFILL_1__15162_ gnd vdd FILL
XFILL_5__7316_ gnd vdd FILL
XFILL_3__11195_ gnd vdd FILL
XFILL_0__14912_ gnd vdd FILL
X_15018_ _7286_/A gnd _15022_/A vdd INVX1
XFILL_0__9410_ gnd vdd FILL
XFILL_0__15892_ gnd vdd FILL
XSFILL89320x54050 gnd vdd FILL
XFILL_4__11505_ gnd vdd FILL
XFILL_5__13844_ gnd vdd FILL
XFILL_6__14094_ gnd vdd FILL
XFILL_4__15273_ gnd vdd FILL
XFILL_4__12485_ gnd vdd FILL
XFILL_3__10146_ gnd vdd FILL
XFILL_1__14113_ gnd vdd FILL
XFILL_1__11325_ gnd vdd FILL
XFILL_2__13664_ gnd vdd FILL
XFILL_0__14843_ gnd vdd FILL
XFILL_5__7247_ gnd vdd FILL
XFILL_2__10876_ gnd vdd FILL
XFILL_1__15093_ gnd vdd FILL
XFILL_4__14224_ gnd vdd FILL
XFILL_0__9341_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1076 gnd vdd FILL
XFILL_2__15403_ gnd vdd FILL
XFILL_4__11436_ gnd vdd FILL
XFILL_2__12615_ gnd vdd FILL
XFILL_5__13775_ gnd vdd FILL
XFILL_2__16383_ gnd vdd FILL
XFILL_1__14044_ gnd vdd FILL
XFILL_3__14954_ gnd vdd FILL
XFILL_2__7469_ gnd vdd FILL
XFILL_1__11256_ gnd vdd FILL
XFILL_2__13595_ gnd vdd FILL
XFILL_5__7178_ gnd vdd FILL
XFILL_0__11986_ gnd vdd FILL
XFILL_5__15514_ gnd vdd FILL
XFILL_0__14774_ gnd vdd FILL
XFILL_5__12726_ gnd vdd FILL
XFILL_4__14155_ gnd vdd FILL
XFILL_2__9208_ gnd vdd FILL
XFILL_0__9272_ gnd vdd FILL
X_8920_ _8828_/A _7640_/CLK _7000_/R vdd _8830_/Y gnd vdd DFFSR
XFILL_3__8001_ gnd vdd FILL
XFILL_2__15334_ gnd vdd FILL
XFILL_3__13905_ gnd vdd FILL
XFILL_4__11367_ gnd vdd FILL
XFILL_3__14885_ gnd vdd FILL
XFILL_0__10937_ gnd vdd FILL
XFILL_1__11187_ gnd vdd FILL
XFILL_0__13725_ gnd vdd FILL
XFILL_4__13106_ gnd vdd FILL
XFILL_0__8223_ gnd vdd FILL
XFILL_4__10318_ gnd vdd FILL
XFILL_5__15445_ gnd vdd FILL
XFILL_5__12657_ gnd vdd FILL
XFILL_3__13836_ gnd vdd FILL
X_8851_ _8851_/A _8854_/B _8850_/Y gnd _8927_/D vdd OAI21X1
XFILL_4__14086_ gnd vdd FILL
XFILL_2__9139_ gnd vdd FILL
XFILL_1__10138_ gnd vdd FILL
XFILL_4__11298_ gnd vdd FILL
XFILL_2__15265_ gnd vdd FILL
XFILL_2__12477_ gnd vdd FILL
XFILL_1__15995_ gnd vdd FILL
XFILL_0__13656_ gnd vdd FILL
XFILL_4__13037_ gnd vdd FILL
XFILL_5__11608_ gnd vdd FILL
X_7802_ _7814_/A _6906_/B gnd _7802_/Y vdd NAND2X1
XFILL_4__10249_ gnd vdd FILL
XFILL_5__15376_ gnd vdd FILL
XFILL_2__14216_ gnd vdd FILL
XFILL_5__12588_ gnd vdd FILL
XFILL_3__13767_ gnd vdd FILL
X_8782_ _8765_/B _8526_/B gnd _8782_/Y vdd NAND2X1
XFILL_2__11428_ gnd vdd FILL
XFILL_3__10979_ gnd vdd FILL
XFILL_2__15196_ gnd vdd FILL
XFILL_0__12607_ gnd vdd FILL
XSFILL18680x59050 gnd vdd FILL
XFILL_1__10069_ gnd vdd FILL
XFILL_1__14946_ gnd vdd FILL
XFILL_0__13587_ gnd vdd FILL
XSFILL104440x30050 gnd vdd FILL
XFILL_0__16375_ gnd vdd FILL
XFILL_0__7105_ gnd vdd FILL
XFILL_6__6873_ gnd vdd FILL
XFILL_0__10799_ gnd vdd FILL
XFILL_5__14327_ gnd vdd FILL
X_7733_ _7787_/Q gnd _7735_/A vdd INVX1
XFILL_3__12718_ gnd vdd FILL
XFILL_3__15506_ gnd vdd FILL
XFILL_5__11539_ gnd vdd FILL
XFILL_0__8085_ gnd vdd FILL
XSFILL33720x62050 gnd vdd FILL
XFILL_2__14147_ gnd vdd FILL
XFILL_3__8903_ gnd vdd FILL
XFILL_0__15326_ gnd vdd FILL
XFILL_3__9883_ gnd vdd FILL
XFILL_3__13698_ gnd vdd FILL
XFILL_2__11359_ gnd vdd FILL
XFILL_1__14877_ gnd vdd FILL
XSFILL49000x29050 gnd vdd FILL
XFILL_0__7036_ gnd vdd FILL
XFILL_5__14258_ gnd vdd FILL
XFILL_3__12649_ gnd vdd FILL
XFILL_3__8834_ gnd vdd FILL
X_7664_ _7620_/A _7664_/CLK _7649_/R vdd _7622_/Y gnd vdd DFFSR
XFILL_3__15437_ gnd vdd FILL
XFILL_1__13828_ gnd vdd FILL
XFILL_4__14988_ gnd vdd FILL
XSFILL89400x34050 gnd vdd FILL
XFILL_2__14078_ gnd vdd FILL
XSFILL59160x73050 gnd vdd FILL
XFILL_0__15257_ gnd vdd FILL
XFILL_5_BUFX2_insert70 gnd vdd FILL
XFILL_0__12469_ gnd vdd FILL
XFILL_5__13209_ gnd vdd FILL
X_9403_ _9453_/Q gnd _9403_/Y vdd INVX1
XFILL_5_BUFX2_insert81 gnd vdd FILL
XFILL_5_BUFX2_insert92 gnd vdd FILL
XFILL_3__15368_ gnd vdd FILL
XFILL_5__14189_ gnd vdd FILL
XFILL_2__13029_ gnd vdd FILL
X_7595_ _7595_/A _7598_/B _7594_/Y gnd _7655_/D vdd OAI21X1
XFILL_4__13939_ gnd vdd FILL
XFILL_3__8765_ gnd vdd FILL
XFILL_0__14208_ gnd vdd FILL
XFILL_0__15188_ gnd vdd FILL
XFILL_1__13759_ gnd vdd FILL
X_9334_ _9334_/A gnd _9336_/A vdd INVX1
XFILL_3__14319_ gnd vdd FILL
XFILL_3__7716_ gnd vdd FILL
XFILL_0__8987_ gnd vdd FILL
XFILL_3__15299_ gnd vdd FILL
XFILL_0__14139_ gnd vdd FILL
XFILL_3__8696_ gnd vdd FILL
XFILL_0__7938_ gnd vdd FILL
XFILL_4__15609_ gnd vdd FILL
XFILL_4_BUFX2_insert227 gnd vdd FILL
X_9265_ _9263_/Y _9240_/A _9265_/C gnd _9265_/Y vdd OAI21X1
XFILL_1__15429_ gnd vdd FILL
XFILL_4_BUFX2_insert238 gnd vdd FILL
XFILL_4_BUFX2_insert249 gnd vdd FILL
X_8216_ _8216_/A _8600_/B gnd _8217_/C vdd NAND2X1
XFILL_0__7869_ gnd vdd FILL
X_9196_ _9144_/A _9958_/CLK _9580_/R vdd _9196_/D gnd vdd DFFSR
XSFILL83560x49050 gnd vdd FILL
XFILL_3__7578_ gnd vdd FILL
XFILL_3_BUFX2_insert905 gnd vdd FILL
XFILL_0__9608_ gnd vdd FILL
XFILL_1__8401_ gnd vdd FILL
XFILL_3_BUFX2_insert916 gnd vdd FILL
XFILL_1__9381_ gnd vdd FILL
XFILL_4__8110_ gnd vdd FILL
XSFILL18760x39050 gnd vdd FILL
X_8147_ _8147_/A gnd _8149_/A vdd INVX1
XFILL_3_BUFX2_insert927 gnd vdd FILL
XSFILL8600x49050 gnd vdd FILL
XFILL_3_BUFX2_insert938 gnd vdd FILL
XSFILL104520x10050 gnd vdd FILL
XFILL_4__9090_ gnd vdd FILL
XFILL_3_BUFX2_insert949 gnd vdd FILL
XFILL_1__8332_ gnd vdd FILL
XSFILL33800x42050 gnd vdd FILL
XFILL_0__9539_ gnd vdd FILL
X_8078_ _8158_/Q gnd _8078_/Y vdd INVX1
XFILL_3__9248_ gnd vdd FILL
X_7029_ _7029_/Q _9958_/CLK _8053_/R vdd _6997_/Y gnd vdd DFFSR
XFILL_1__8263_ gnd vdd FILL
XFILL_1__7214_ gnd vdd FILL
X_10980_ _10980_/A vdd _10980_/C gnd _10986_/D vdd OAI21X1
XFILL_1__8194_ gnd vdd FILL
XFILL111960x52050 gnd vdd FILL
XFILL112440x59050 gnd vdd FILL
XFILL_4__9992_ gnd vdd FILL
XFILL_1_BUFX2_insert106 gnd vdd FILL
X_12650_ _12648_/Y vdd _12649_/Y gnd _12690_/D vdd OAI21X1
XFILL112040x61050 gnd vdd FILL
XFILL_1__7076_ gnd vdd FILL
XSFILL24360x60050 gnd vdd FILL
XFILL_0_CLKBUF1_insert210 gnd vdd FILL
X_11601_ _11630_/B _11139_/Y _11406_/Y gnd _11602_/A vdd OAI21X1
XFILL_4__8874_ gnd vdd FILL
XFILL_0_CLKBUF1_insert221 gnd vdd FILL
X_12581_ _12579_/Y vdd _12580_/Y gnd _12667_/D vdd OAI21X1
XFILL_0_BUFX2_insert806 gnd vdd FILL
XFILL_0_BUFX2_insert817 gnd vdd FILL
XFILL_0_BUFX2_insert828 gnd vdd FILL
XFILL_4__7825_ gnd vdd FILL
X_14320_ _14211_/A _14320_/B _14320_/C _14318_/Y gnd _14321_/B vdd OAI22X1
XFILL_1_BUFX2_insert1003 gnd vdd FILL
XFILL_0_BUFX2_insert839 gnd vdd FILL
X_11532_ _11431_/Y _11616_/B _11550_/A gnd _11533_/B vdd OAI21X1
XSFILL18840x19050 gnd vdd FILL
XFILL_1_BUFX2_insert1014 gnd vdd FILL
XFILL_1_BUFX2_insert1025 gnd vdd FILL
XFILL_2__6840_ gnd vdd FILL
XFILL_1_BUFX2_insert1036 gnd vdd FILL
XFILL_4__7756_ gnd vdd FILL
X_14251_ _9766_/A _14213_/A _14180_/C _10534_/A gnd _14253_/A vdd AOI22X1
XFILL_1_BUFX2_insert1047 gnd vdd FILL
XFILL_1_BUFX2_insert1058 gnd vdd FILL
X_11463_ _11185_/A _11185_/B _11463_/C gnd _11480_/C vdd OAI21X1
XSFILL99320x17050 gnd vdd FILL
XFILL_1_BUFX2_insert1069 gnd vdd FILL
XFILL_1__7978_ gnd vdd FILL
X_13202_ _13202_/Q _13180_/CLK _13180_/R vdd _13202_/D gnd vdd DFFSR
X_10414_ _10414_/A _10395_/A _10413_/Y gnd _10472_/D vdd OAI21X1
XFILL_4__7687_ gnd vdd FILL
X_14182_ _14182_/A _14182_/B _14179_/Y gnd _14195_/B vdd NAND3X1
XFILL_2__8510_ gnd vdd FILL
X_11394_ _11085_/C gnd _11394_/Y vdd INVX1
XFILL_1__6929_ gnd vdd FILL
XFILL_2__9490_ gnd vdd FILL
XFILL_4__9426_ gnd vdd FILL
X_13133_ _13133_/A gnd _13135_/A vdd INVX1
XSFILL23800x8050 gnd vdd FILL
XFILL_4_BUFX2_insert750 gnd vdd FILL
X_10345_ _14359_/D _9705_/CLK _7649_/R vdd _10345_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert761 gnd vdd FILL
XFILL_1__9648_ gnd vdd FILL
XFILL_2__8441_ gnd vdd FILL
XFILL_6_CLKBUF1_insert116 gnd vdd FILL
XFILL_4__9357_ gnd vdd FILL
XFILL_6_CLKBUF1_insert127 gnd vdd FILL
XFILL_4_BUFX2_insert772 gnd vdd FILL
XFILL_3_CLKBUF1_insert1082 gnd vdd FILL
XFILL_4_BUFX2_insert783 gnd vdd FILL
XFILL_5__10910_ gnd vdd FILL
XFILL_4_BUFX2_insert794 gnd vdd FILL
XFILL_3__10000_ gnd vdd FILL
X_13064_ _6887_/A _8169_/CLK _8937_/R vdd _13064_/D gnd vdd DFFSR
XSFILL23800x74050 gnd vdd FILL
X_10276_ _10304_/B _9380_/B gnd _10276_/Y vdd NAND2X1
XFILL_5__7101_ gnd vdd FILL
XFILL_5__11890_ gnd vdd FILL
XFILL_2__8372_ gnd vdd FILL
XSFILL89240x69050 gnd vdd FILL
X_12015_ _11999_/A _12364_/A _11999_/C gnd _12018_/A vdd NAND3X1
XFILL_4__9288_ gnd vdd FILL
XFILL_5__8081_ gnd vdd FILL
XSFILL24440x40050 gnd vdd FILL
XFILL_2__7323_ gnd vdd FILL
XFILL_4__12270_ gnd vdd FILL
XFILL_1__11110_ gnd vdd FILL
XFILL_2__10661_ gnd vdd FILL
XFILL_5__7032_ gnd vdd FILL
XFILL_1__12090_ gnd vdd FILL
XFILL_0__11840_ gnd vdd FILL
XFILL_4__8239_ gnd vdd FILL
XFILL_4__11221_ gnd vdd FILL
XFILL_2__12400_ gnd vdd FILL
XFILL_5__13560_ gnd vdd FILL
XFILL_5__10772_ gnd vdd FILL
XFILL_3__11951_ gnd vdd FILL
XFILL_1__11041_ gnd vdd FILL
XFILL_2__13380_ gnd vdd FILL
XFILL_0__11771_ gnd vdd FILL
XFILL_5__12511_ gnd vdd FILL
XFILL_3__10902_ gnd vdd FILL
XFILL_4__11152_ gnd vdd FILL
X_13966_ _13966_/A _13879_/B _13479_/C _15458_/A gnd _13966_/Y vdd OAI22X1
XFILL_2__12331_ gnd vdd FILL
XFILL_3__14670_ gnd vdd FILL
XFILL_5__13491_ gnd vdd FILL
XFILL_3__11882_ gnd vdd FILL
XFILL_2__7185_ gnd vdd FILL
XFILL_0__13510_ gnd vdd FILL
XSFILL115320x21050 gnd vdd FILL
XFILL_0__14490_ gnd vdd FILL
X_15705_ _15705_/A _15705_/B _15705_/C gnd _15706_/B vdd NAND3X1
XFILL_5__15230_ gnd vdd FILL
XSFILL69160x36050 gnd vdd FILL
X_12917_ vdd _12917_/B gnd _12918_/C vdd NAND2X1
XFILL_4__10103_ gnd vdd FILL
XFILL_3__13621_ gnd vdd FILL
XFILL_5__8983_ gnd vdd FILL
XFILL_5__12442_ gnd vdd FILL
XSFILL3640x1050 gnd vdd FILL
XFILL_1__14800_ gnd vdd FILL
XFILL_2__15050_ gnd vdd FILL
XFILL_4__15960_ gnd vdd FILL
XFILL_6__11993_ gnd vdd FILL
XFILL_4__11083_ gnd vdd FILL
X_13897_ _13895_/Y _13897_/B _13897_/C gnd _13908_/B vdd NAND3X1
XFILL_3__10833_ gnd vdd FILL
XFILL_0__13441_ gnd vdd FILL
XFILL_2__12262_ gnd vdd FILL
XFILL_1__15780_ gnd vdd FILL
XFILL_0__10653_ gnd vdd FILL
XFILL_5__7934_ gnd vdd FILL
XFILL_1__12992_ gnd vdd FILL
XFILL_3__16340_ gnd vdd FILL
X_12848_ vdd _12848_/B gnd _12849_/C vdd NAND2X1
X_15636_ _9376_/A _15636_/B _15995_/C gnd _15637_/C vdd NAND3X1
XFILL_2__14001_ gnd vdd FILL
XFILL_5__12373_ gnd vdd FILL
XFILL_1_BUFX2_insert640 gnd vdd FILL
XFILL_4__10034_ gnd vdd FILL
XFILL_5__15161_ gnd vdd FILL
XFILL_4__14911_ gnd vdd FILL
XFILL_1_BUFX2_insert651 gnd vdd FILL
XSFILL104360x45050 gnd vdd FILL
XFILL_3__13552_ gnd vdd FILL
XFILL_2__11213_ gnd vdd FILL
XFILL_3__10764_ gnd vdd FILL
XFILL_1__14731_ gnd vdd FILL
XFILL_4__15891_ gnd vdd FILL
XFILL_0__13372_ gnd vdd FILL
XFILL_1__11943_ gnd vdd FILL
XFILL_2__12193_ gnd vdd FILL
XFILL_1_BUFX2_insert662 gnd vdd FILL
XFILL_0__16160_ gnd vdd FILL
XFILL_5__7865_ gnd vdd FILL
XFILL_1_BUFX2_insert673 gnd vdd FILL
XFILL_5__14112_ gnd vdd FILL
XFILL_3__12503_ gnd vdd FILL
XFILL_1_BUFX2_insert684 gnd vdd FILL
X_15567_ _12813_/Q _14980_/Y _14982_/Y gnd _15568_/C vdd NAND3X1
XSFILL74280x27050 gnd vdd FILL
XFILL_5__11324_ gnd vdd FILL
X_12779_ _12779_/A gnd _12779_/Y vdd INVX1
XFILL_1_BUFX2_insert695 gnd vdd FILL
XFILL_4__14842_ gnd vdd FILL
XFILL_5__15092_ gnd vdd FILL
XFILL_3__16271_ gnd vdd FILL
XFILL_0__12323_ gnd vdd FILL
XFILL_2__11144_ gnd vdd FILL
XFILL_0__15111_ gnd vdd FILL
XFILL_3__13483_ gnd vdd FILL
XFILL_5__9604_ gnd vdd FILL
XFILL_0__16091_ gnd vdd FILL
XFILL_3__6880_ gnd vdd FILL
XFILL_1__14662_ gnd vdd FILL
XFILL_3__10695_ gnd vdd FILL
XFILL_0__8910_ gnd vdd FILL
XFILL_1__11874_ gnd vdd FILL
XFILL_6__12614_ gnd vdd FILL
X_14518_ _14518_/A _13803_/A _14865_/C _14518_/D gnd _14518_/Y vdd OAI22X1
XFILL_3__15222_ gnd vdd FILL
XFILL_5__14043_ gnd vdd FILL
XFILL_5__11255_ gnd vdd FILL
XFILL_3__12434_ gnd vdd FILL
XFILL_0__9890_ gnd vdd FILL
X_15498_ _15922_/C _15498_/B _15351_/D _15498_/D gnd _15500_/A vdd OAI22X1
XSFILL89320x49050 gnd vdd FILL
XFILL_1__16401_ gnd vdd FILL
XFILL112200x21050 gnd vdd FILL
XFILL_1__13613_ gnd vdd FILL
XFILL_4__11985_ gnd vdd FILL
XFILL_0__15042_ gnd vdd FILL
XFILL_2__15952_ gnd vdd FILL
XFILL_4__14773_ gnd vdd FILL
XFILL_0__12254_ gnd vdd FILL
XFILL_2__11075_ gnd vdd FILL
XFILL_1__10825_ gnd vdd FILL
XFILL_1__14593_ gnd vdd FILL
XFILL_5__9535_ gnd vdd FILL
XFILL_0__8841_ gnd vdd FILL
X_14449_ _14449_/A _14448_/Y gnd _14450_/A vdd NOR2X1
X_7380_ _7369_/B _7380_/B gnd _7381_/C vdd NAND2X1
XFILL_3__15153_ gnd vdd FILL
XFILL_5__11186_ gnd vdd FILL
XFILL_4__13724_ gnd vdd FILL
XFILL_3__12365_ gnd vdd FILL
XFILL_4__10936_ gnd vdd FILL
XFILL_1__16332_ gnd vdd FILL
XFILL_2__9757_ gnd vdd FILL
XFILL_0__11205_ gnd vdd FILL
XFILL_2__14903_ gnd vdd FILL
XFILL_2__10026_ gnd vdd FILL
XFILL_2__6969_ gnd vdd FILL
XFILL_1__13544_ gnd vdd FILL
XFILL_2__15883_ gnd vdd FILL
XFILL_0__12185_ gnd vdd FILL
XFILL_1__10756_ gnd vdd FILL
XFILL_5__9466_ gnd vdd FILL
XFILL_5__10137_ gnd vdd FILL
XFILL_3__14104_ gnd vdd FILL
XFILL_3__7501_ gnd vdd FILL
XFILL_0__8772_ gnd vdd FILL
XFILL_3__11316_ gnd vdd FILL
XSFILL18680x1050 gnd vdd FILL
XFILL_5__15994_ gnd vdd FILL
XFILL_2__8708_ gnd vdd FILL
XFILL_4__13655_ gnd vdd FILL
XFILL_2__14834_ gnd vdd FILL
XSFILL13560x44050 gnd vdd FILL
XFILL_3__15084_ gnd vdd FILL
XFILL_3__8481_ gnd vdd FILL
XFILL_1__16263_ gnd vdd FILL
XFILL_3__12296_ gnd vdd FILL
XFILL_0__11136_ gnd vdd FILL
XFILL_1__10687_ gnd vdd FILL
XFILL_1__13475_ gnd vdd FILL
X_16119_ _8560_/Q gnd _16119_/Y vdd INVX1
XFILL_5__9397_ gnd vdd FILL
X_9050_ _8962_/A _9050_/CLK _9050_/R vdd _8964_/Y gnd vdd DFFSR
XFILL_0__7723_ gnd vdd FILL
XFILL_4__12606_ gnd vdd FILL
XFILL_3__14035_ gnd vdd FILL
XFILL_5__10068_ gnd vdd FILL
XFILL_5__14945_ gnd vdd FILL
XFILL_2__8639_ gnd vdd FILL
XFILL_1__15214_ gnd vdd FILL
XFILL_3__7432_ gnd vdd FILL
XFILL_4__16374_ gnd vdd FILL
XFILL_3__11247_ gnd vdd FILL
XFILL_4__13586_ gnd vdd FILL
XFILL_1__12426_ gnd vdd FILL
XFILL_4__10798_ gnd vdd FILL
XSFILL69240x16050 gnd vdd FILL
XFILL_2__14765_ gnd vdd FILL
XFILL_1__16194_ gnd vdd FILL
XFILL_0__15944_ gnd vdd FILL
XFILL_5__8348_ gnd vdd FILL
XFILL_2__11977_ gnd vdd FILL
XFILL_0__11067_ gnd vdd FILL
X_8001_ _8001_/A gnd _8001_/Y vdd INVX1
XFILL_4__15325_ gnd vdd FILL
XFILL_5__14876_ gnd vdd FILL
XFILL_2__13716_ gnd vdd FILL
XFILL_2__10928_ gnd vdd FILL
XFILL_0__10018_ gnd vdd FILL
XFILL_3__7363_ gnd vdd FILL
XFILL_3__11178_ gnd vdd FILL
XFILL_1__15145_ gnd vdd FILL
XFILL_1__12357_ gnd vdd FILL
XFILL_2__14696_ gnd vdd FILL
XFILL_0__15875_ gnd vdd FILL
XFILL_3__9102_ gnd vdd FILL
XFILL_5__13827_ gnd vdd FILL
XFILL_4__15256_ gnd vdd FILL
XFILL_0__7585_ gnd vdd FILL
XFILL_4__12468_ gnd vdd FILL
XFILL_3__10129_ gnd vdd FILL
XFILL_2__13647_ gnd vdd FILL
XFILL_1__11308_ gnd vdd FILL
XSFILL8680x23050 gnd vdd FILL
XFILL_0__14826_ gnd vdd FILL
XFILL_3__15986_ gnd vdd FILL
XFILL_1__15076_ gnd vdd FILL
XFILL_3__7294_ gnd vdd FILL
XFILL_1__12288_ gnd vdd FILL
XFILL_4__14207_ gnd vdd FILL
XFILL_4__11419_ gnd vdd FILL
XFILL_5__13758_ gnd vdd FILL
X_9952_ _9952_/Q _9568_/CLK _8431_/R vdd _9952_/D gnd vdd DFFSR
XFILL_3__9033_ gnd vdd FILL
XFILL_4__15187_ gnd vdd FILL
XFILL_4__12399_ gnd vdd FILL
XFILL_1__14027_ gnd vdd FILL
XFILL_3__14937_ gnd vdd FILL
XFILL_2__16366_ gnd vdd FILL
XFILL_2__13578_ gnd vdd FILL
XFILL_1__11239_ gnd vdd FILL
XSFILL59160x68050 gnd vdd FILL
XFILL_0__14757_ gnd vdd FILL
XFILL_5__12709_ gnd vdd FILL
XFILL_0__9255_ gnd vdd FILL
XFILL_0__11969_ gnd vdd FILL
X_8903_ _8945_/Q gnd _8903_/Y vdd INVX1
XFILL_2__15317_ gnd vdd FILL
XFILL_4__14138_ gnd vdd FILL
X_9883_ _9865_/A _9371_/B gnd _9883_/Y vdd NAND2X1
XFILL_2__12529_ gnd vdd FILL
XFILL_5__13689_ gnd vdd FILL
XFILL_3__14868_ gnd vdd FILL
XSFILL49400x45050 gnd vdd FILL
XFILL_2__16297_ gnd vdd FILL
XFILL_0__13708_ gnd vdd FILL
XFILL_0__8206_ gnd vdd FILL
XFILL_5__15428_ gnd vdd FILL
XFILL_0__14688_ gnd vdd FILL
X_8834_ _8834_/A gnd _8836_/A vdd INVX1
XFILL_6__14979_ gnd vdd FILL
XFILL_4__14069_ gnd vdd FILL
XFILL_3__13819_ gnd vdd FILL
XFILL_2__15248_ gnd vdd FILL
XSFILL108680x30050 gnd vdd FILL
XFILL_1__15978_ gnd vdd FILL
XFILL_0__13639_ gnd vdd FILL
XFILL_3__14799_ gnd vdd FILL
XSFILL37960x62050 gnd vdd FILL
XFILL_0__8137_ gnd vdd FILL
XFILL_6_BUFX2_insert812 gnd vdd FILL
XFILL_5__15359_ gnd vdd FILL
X_8765_ _8765_/A _8765_/B _8764_/Y gnd _8765_/Y vdd OAI21X1
XFILL_3__9935_ gnd vdd FILL
XFILL_2__15179_ gnd vdd FILL
XFILL_1__14929_ gnd vdd FILL
XFILL_0__16358_ gnd vdd FILL
XFILL_1__8950_ gnd vdd FILL
X_7716_ _7690_/B _8228_/B gnd _7716_/Y vdd NAND2X1
XFILL_0__8068_ gnd vdd FILL
XFILL_0__15309_ gnd vdd FILL
X_8696_ _8694_/Y _8695_/B _8696_/C gnd _8696_/Y vdd OAI21X1
XFILL_3__9866_ gnd vdd FILL
XFILL_6_BUFX2_insert889 gnd vdd FILL
XFILL_0__16289_ gnd vdd FILL
XFILL_4__7610_ gnd vdd FILL
X_7647_ _7647_/Q _7647_/CLK _7775_/R vdd _7647_/D gnd vdd DFFSR
XFILL_1__8881_ gnd vdd FILL
XFILL_4__8590_ gnd vdd FILL
XFILL_3__9797_ gnd vdd FILL
XFILL_6__8526_ gnd vdd FILL
XFILL_1__7832_ gnd vdd FILL
XSFILL33800x37050 gnd vdd FILL
X_7578_ _7578_/A gnd _7578_/Y vdd INVX1
XFILL_3__8748_ gnd vdd FILL
XSFILL43960x81050 gnd vdd FILL
X_9317_ _9317_/Q _8537_/CLK _9054_/R vdd _9253_/Y gnd vdd DFFSR
XFILL_1__7763_ gnd vdd FILL
XFILL_4__7472_ gnd vdd FILL
XFILL_1__9502_ gnd vdd FILL
X_9248_ _9248_/A gnd _9250_/A vdd INVX1
XFILL_4__9211_ gnd vdd FILL
XFILL_1__7694_ gnd vdd FILL
X_10130_ _10193_/A _7954_/B gnd _10131_/C vdd NAND2X1
XFILL_3_BUFX2_insert702 gnd vdd FILL
XFILL_4__9142_ gnd vdd FILL
XFILL_3_BUFX2_insert713 gnd vdd FILL
X_9179_ _9179_/Q _8151_/CLK _9944_/R vdd _9095_/Y gnd vdd DFFSR
XFILL_3_BUFX2_insert724 gnd vdd FILL
X_10061_ _10061_/A gnd _10061_/Y vdd INVX1
XFILL_3_BUFX2_insert735 gnd vdd FILL
XFILL_3_BUFX2_insert746 gnd vdd FILL
XFILL112040x56050 gnd vdd FILL
XFILL_3_BUFX2_insert757 gnd vdd FILL
XFILL_1__9364_ gnd vdd FILL
XFILL_3_BUFX2_insert768 gnd vdd FILL
XFILL_3_BUFX2_insert779 gnd vdd FILL
XSFILL64760x60050 gnd vdd FILL
XFILL_1__8315_ gnd vdd FILL
XSFILL38920x70050 gnd vdd FILL
XFILL_1__9295_ gnd vdd FILL
X_13820_ _7261_/Q gnd _13820_/Y vdd INVX1
XFILL_1_BUFX2_insert90 gnd vdd FILL
XSFILL2760x82050 gnd vdd FILL
XFILL_1__8246_ gnd vdd FILL
X_13751_ _9820_/Q _13751_/B _13751_/C _9864_/A gnd _13751_/Y vdd AOI22X1
X_10963_ _10963_/A _10924_/Y gnd _10963_/Y vdd NOR2X1
X_12702_ _10944_/C memoryOutData[2] gnd _12703_/C vdd NAND2X1
XFILL_4__9975_ gnd vdd FILL
X_13682_ _14878_/C _13682_/B _9986_/A _14214_/C gnd _13684_/A vdd AOI22X1
X_10894_ _12704_/A _10894_/B _10881_/A gnd _10894_/Y vdd NOR3X1
XFILL111960x6050 gnd vdd FILL
XFILL_2__8990_ gnd vdd FILL
X_15421_ _15416_/Y _15421_/B _15421_/C gnd _15426_/C vdd NOR3X1
X_12633_ _12633_/A gnd _12635_/A vdd INVX1
XFILL_0_BUFX2_insert603 gnd vdd FILL
XFILL_2__7941_ gnd vdd FILL
XFILL_1__7059_ gnd vdd FILL
XFILL_0_BUFX2_insert614 gnd vdd FILL
X_15352_ _13811_/Y _16213_/B _16208_/B _13802_/Y gnd _15353_/A vdd OAI22X1
XFILL_0_BUFX2_insert625 gnd vdd FILL
XFILL_4__8857_ gnd vdd FILL
XSFILL63960x12050 gnd vdd FILL
XFILL_0_BUFX2_insert636 gnd vdd FILL
X_12564_ _12430_/A _13175_/CLK _12536_/R vdd _12564_/D gnd vdd DFFSR
XSFILL23800x69050 gnd vdd FILL
XFILL_0_BUFX2_insert647 gnd vdd FILL
XSFILL33480x3050 gnd vdd FILL
XFILL_2__7872_ gnd vdd FILL
XFILL_4__7808_ gnd vdd FILL
XFILL_0_BUFX2_insert658 gnd vdd FILL
X_14303_ _7527_/Q gnd _15760_/B vdd INVX1
XFILL_0_BUFX2_insert669 gnd vdd FILL
XFILL112120x36050 gnd vdd FILL
XFILL_5__7581_ gnd vdd FILL
X_11515_ _11507_/Y _11514_/Y gnd _11516_/A vdd NOR2X1
XFILL_5__11040_ gnd vdd FILL
XFILL_2__9611_ gnd vdd FILL
X_15283_ _16306_/A _13725_/D _15558_/D _15283_/D gnd _15284_/B vdd OAI22X1
XFILL_4__8788_ gnd vdd FILL
X_12495_ _12493_/Y vdd _12494_/Y gnd _12495_/Y vdd OAI21X1
XFILL_4__11770_ gnd vdd FILL
XSFILL64040x21050 gnd vdd FILL
XFILL_1__11590_ gnd vdd FILL
XFILL_4__7739_ gnd vdd FILL
X_14234_ _14234_/A _14233_/Y gnd _14234_/Y vdd NOR2X1
X_11446_ _11446_/A _11445_/Y gnd _11447_/C vdd NAND2X1
XFILL_2__11900_ gnd vdd FILL
XFILL_2__9542_ gnd vdd FILL
XFILL_3__12150_ gnd vdd FILL
XFILL_1__10541_ gnd vdd FILL
XFILL_5__9251_ gnd vdd FILL
XFILL_2__12880_ gnd vdd FILL
X_14165_ _8992_/A gnd _15646_/C vdd INVX1
XFILL_3__11101_ gnd vdd FILL
XSFILL33960x9050 gnd vdd FILL
XFILL_4__13440_ gnd vdd FILL
XFILL_4__10652_ gnd vdd FILL
X_11377_ _11839_/A _11377_/B _11376_/Y gnd _11377_/Y vdd AOI21X1
XFILL_2__9473_ gnd vdd FILL
XFILL_3__12081_ gnd vdd FILL
XFILL_5__8202_ gnd vdd FILL
XFILL_5__12991_ gnd vdd FILL
XFILL_2__11831_ gnd vdd FILL
XFILL_1__13260_ gnd vdd FILL
XFILL_4__9409_ gnd vdd FILL
X_13116_ _13108_/B _13116_/B gnd _13117_/C vdd NAND2X1
XFILL_0__13990_ gnd vdd FILL
XFILL_5__14730_ gnd vdd FILL
X_10328_ _13537_/A _8663_/CLK _8664_/R vdd _10238_/Y gnd vdd DFFSR
XFILL_4_BUFX2_insert580 gnd vdd FILL
XSFILL13880x80050 gnd vdd FILL
XFILL_4__13371_ gnd vdd FILL
XFILL_5__11942_ gnd vdd FILL
X_14096_ _14095_/Y _14096_/B gnd _14122_/B vdd NOR2X1
XFILL_3__11032_ gnd vdd FILL
XFILL_2__14550_ gnd vdd FILL
XFILL_4_BUFX2_insert591 gnd vdd FILL
XFILL_1__12211_ gnd vdd FILL
XFILL_5__8133_ gnd vdd FILL
XFILL_2__11762_ gnd vdd FILL
XSFILL84200x34050 gnd vdd FILL
X_13047_ _6870_/A _8176_/CLK _8176_/R vdd _13047_/D gnd vdd DFFSR
XFILL_4__12322_ gnd vdd FILL
XFILL_4__15110_ gnd vdd FILL
XFILL_4__16090_ gnd vdd FILL
X_10259_ _10259_/A _10264_/A _10258_/Y gnd _10335_/D vdd OAI21X1
XFILL_5__14661_ gnd vdd FILL
XFILL_2__13501_ gnd vdd FILL
XFILL_5__11873_ gnd vdd FILL
XFILL_2__8355_ gnd vdd FILL
XFILL_3__15840_ gnd vdd FILL
XFILL_2__14481_ gnd vdd FILL
XFILL_1__12142_ gnd vdd FILL
XFILL_5__8064_ gnd vdd FILL
XFILL_0__15660_ gnd vdd FILL
XFILL_5__16400_ gnd vdd FILL
XFILL_2__11693_ gnd vdd FILL
XFILL_5__13612_ gnd vdd FILL
XFILL_0__12872_ gnd vdd FILL
XSFILL59000x10050 gnd vdd FILL
XFILL_0__7370_ gnd vdd FILL
XFILL_2__16220_ gnd vdd FILL
XFILL_2__7306_ gnd vdd FILL
XFILL_4__15041_ gnd vdd FILL
XFILL_6__15951_ gnd vdd FILL
XFILL_4__12253_ gnd vdd FILL
XFILL_5__10824_ gnd vdd FILL
XFILL_5__14592_ gnd vdd FILL
XFILL_2__13432_ gnd vdd FILL
XFILL_0__14611_ gnd vdd FILL
XFILL_1__12073_ gnd vdd FILL
XFILL_3__15771_ gnd vdd FILL
XFILL_3__12983_ gnd vdd FILL
XFILL_2__10644_ gnd vdd FILL
XFILL_0__11823_ gnd vdd FILL
XFILL_5__16331_ gnd vdd FILL
XFILL_0__15591_ gnd vdd FILL
XFILL_4__11204_ gnd vdd FILL
XFILL_6__14902_ gnd vdd FILL
XFILL_5__13543_ gnd vdd FILL
XFILL_1__15901_ gnd vdd FILL
XFILL_3__11934_ gnd vdd FILL
XFILL_4__12184_ gnd vdd FILL
XFILL_2__7237_ gnd vdd FILL
XFILL_5__10755_ gnd vdd FILL
XFILL_3__14722_ gnd vdd FILL
XFILL_1__11024_ gnd vdd FILL
XFILL_2__16151_ gnd vdd FILL
XFILL_2__13363_ gnd vdd FILL
X_14998_ _14989_/A _16037_/B _15024_/C gnd _14998_/Y vdd NAND3X1
XFILL112200x16050 gnd vdd FILL
XFILL_2__10575_ gnd vdd FILL
XFILL_0__14542_ gnd vdd FILL
XFILL_0__11754_ gnd vdd FILL
XFILL_0__9040_ gnd vdd FILL
XFILL_4__11135_ gnd vdd FILL
XFILL_2__15102_ gnd vdd FILL
XFILL_5__16262_ gnd vdd FILL
XFILL_5__13474_ gnd vdd FILL
XFILL_2__12314_ gnd vdd FILL
X_13949_ _13949_/A _13948_/Y gnd _13952_/C vdd NOR2X1
XFILL_5__10686_ gnd vdd FILL
XFILL_2__7168_ gnd vdd FILL
XFILL_1__15832_ gnd vdd FILL
XFILL_3__11865_ gnd vdd FILL
X_6880_ _6880_/A gnd memoryWriteData[10] vdd BUFX2
XFILL_3__14653_ gnd vdd FILL
XFILL_2__16082_ gnd vdd FILL
XFILL_2__13294_ gnd vdd FILL
XFILL_0__10705_ gnd vdd FILL
XFILL_0__14473_ gnd vdd FILL
XFILL_5__15213_ gnd vdd FILL
XFILL_0__11685_ gnd vdd FILL
XFILL_5__12425_ gnd vdd FILL
XFILL_5__8966_ gnd vdd FILL
XFILL_6__14764_ gnd vdd FILL
XFILL_3__10816_ gnd vdd FILL
XFILL_3__13604_ gnd vdd FILL
XFILL_5__16193_ gnd vdd FILL
XFILL_2__15033_ gnd vdd FILL
XFILL_4__15943_ gnd vdd FILL
XFILL_4__11066_ gnd vdd FILL
XFILL_0__16212_ gnd vdd FILL
XFILL_3__14584_ gnd vdd FILL
XFILL_2__12245_ gnd vdd FILL
XFILL_2__7099_ gnd vdd FILL
XFILL_0__10636_ gnd vdd FILL
XFILL_0__13424_ gnd vdd FILL
XFILL_3__7981_ gnd vdd FILL
XFILL_1__15763_ gnd vdd FILL
XFILL_3__11796_ gnd vdd FILL
XFILL_1__12975_ gnd vdd FILL
XFILL_6__13715_ gnd vdd FILL
XFILL_4__10017_ gnd vdd FILL
X_15619_ _8736_/A _15821_/B gnd _15619_/Y vdd NAND2X1
XSFILL53960x44050 gnd vdd FILL
XFILL_1_BUFX2_insert470 gnd vdd FILL
XFILL_5__15144_ gnd vdd FILL
X_8550_ _8550_/Q _7282_/CLK _9054_/R vdd _8488_/Y gnd vdd DFFSR
XFILL_5__12356_ gnd vdd FILL
XFILL_3__16323_ gnd vdd FILL
XFILL_3__13535_ gnd vdd FILL
XFILL_5__8897_ gnd vdd FILL
XSFILL109480x73050 gnd vdd FILL
XFILL_3__9720_ gnd vdd FILL
XFILL_1_BUFX2_insert481 gnd vdd FILL
XFILL_1__14714_ gnd vdd FILL
XFILL_3__6932_ gnd vdd FILL
XFILL_3__10747_ gnd vdd FILL
XFILL_4__15874_ gnd vdd FILL
XFILL_1__11926_ gnd vdd FILL
XFILL_0__16143_ gnd vdd FILL
XFILL_2__12176_ gnd vdd FILL
XFILL_1_BUFX2_insert492 gnd vdd FILL
XFILL_0__13355_ gnd vdd FILL
XFILL_1__15694_ gnd vdd FILL
XSFILL13160x41050 gnd vdd FILL
XFILL_0__10567_ gnd vdd FILL
XFILL_5__7848_ gnd vdd FILL
X_7501_ _7539_/Q gnd _7503_/A vdd INVX1
XFILL_5_BUFX2_insert808 gnd vdd FILL
XFILL_5__11307_ gnd vdd FILL
XFILL_4__14825_ gnd vdd FILL
XFILL_5__15075_ gnd vdd FILL
XFILL_5_BUFX2_insert819 gnd vdd FILL
XFILL_3__13466_ gnd vdd FILL
X_8481_ _8460_/A _7329_/B gnd _8482_/C vdd NAND2X1
XFILL_5__12287_ gnd vdd FILL
XFILL_2__11127_ gnd vdd FILL
XFILL_3__16254_ gnd vdd FILL
XFILL_3__9651_ gnd vdd FILL
XFILL_3__10678_ gnd vdd FILL
XFILL_1__14645_ gnd vdd FILL
XFILL_3__6863_ gnd vdd FILL
XFILL_0__12306_ gnd vdd FILL
XFILL_0__13286_ gnd vdd FILL
XBUFX2_insert1005 _10928_/Y gnd _12272_/A vdd BUFX2
XFILL_0__16074_ gnd vdd FILL
XSFILL103960x13050 gnd vdd FILL
XFILL_1__11857_ gnd vdd FILL
XBUFX2_insert1016 _15054_/Y gnd _15169_/A vdd BUFX2
XFILL_6__16365_ gnd vdd FILL
XFILL_0__10498_ gnd vdd FILL
XFILL_5__14026_ gnd vdd FILL
XFILL_3__12417_ gnd vdd FILL
XFILL_3__15205_ gnd vdd FILL
X_7432_ _7432_/A gnd _7434_/A vdd INVX1
XFILL_0__9873_ gnd vdd FILL
XFILL_6__13577_ gnd vdd FILL
XBUFX2_insert1027 _13333_/Y gnd _9238_/B vdd BUFX2
XFILL_5__11238_ gnd vdd FILL
XBUFX2_insert1038 _12390_/Y gnd _8868_/B vdd BUFX2
XFILL_3__16185_ gnd vdd FILL
XFILL_3__8602_ gnd vdd FILL
XFILL_4__14756_ gnd vdd FILL
XFILL_2__9809_ gnd vdd FILL
XFILL_3__13397_ gnd vdd FILL
XFILL_0__15025_ gnd vdd FILL
XFILL_2__15935_ gnd vdd FILL
XFILL_4__11968_ gnd vdd FILL
XFILL_1__10808_ gnd vdd FILL
XFILL_0__12237_ gnd vdd FILL
XFILL_2__11058_ gnd vdd FILL
XSFILL8680x18050 gnd vdd FILL
XFILL_1__14576_ gnd vdd FILL
XFILL_6__15316_ gnd vdd FILL
XFILL_5__9518_ gnd vdd FILL
XBUFX2_insert1049 _12806_/Q gnd _12308_/B vdd BUFX2
XFILL_0__8824_ gnd vdd FILL
XFILL_6__9291_ gnd vdd FILL
XFILL_1__11788_ gnd vdd FILL
XFILL_3__15136_ gnd vdd FILL
XFILL_4__13707_ gnd vdd FILL
XFILL_5__11169_ gnd vdd FILL
XFILL_4__10919_ gnd vdd FILL
XFILL_2__10009_ gnd vdd FILL
XFILL_3__8533_ gnd vdd FILL
XFILL_3__12348_ gnd vdd FILL
XFILL_1__16315_ gnd vdd FILL
X_7363_ _7361_/Y _7354_/B _7363_/C gnd _7407_/D vdd OAI21X1
XSFILL33880x11050 gnd vdd FILL
XFILL_1__13527_ gnd vdd FILL
XFILL_4__14687_ gnd vdd FILL
XFILL_4__11899_ gnd vdd FILL
XFILL_0__12168_ gnd vdd FILL
XFILL_6__8242_ gnd vdd FILL
XFILL_2__15866_ gnd vdd FILL
X_9102_ _9102_/A gnd _9104_/A vdd INVX1
XFILL_6__12459_ gnd vdd FILL
XFILL_0__8755_ gnd vdd FILL
XFILL_5__15977_ gnd vdd FILL
XFILL_4__13638_ gnd vdd FILL
XFILL_3__15067_ gnd vdd FILL
X_7294_ _7292_/Y _7323_/A _7293_/Y gnd _7384_/D vdd OAI21X1
XFILL_3__8464_ gnd vdd FILL
XFILL_2__14817_ gnd vdd FILL
XFILL_3__12279_ gnd vdd FILL
XFILL_0__11119_ gnd vdd FILL
XFILL_1__16246_ gnd vdd FILL
XFILL_1__13458_ gnd vdd FILL
XFILL_2__15797_ gnd vdd FILL
XSFILL74200x66050 gnd vdd FILL
XFILL_0__12099_ gnd vdd FILL
XFILL_0__7706_ gnd vdd FILL
XFILL_6__15178_ gnd vdd FILL
XFILL_3__14018_ gnd vdd FILL
X_9033_ _9033_/A _9044_/A _9033_/C gnd _9073_/D vdd OAI21X1
XFILL_5__14928_ gnd vdd FILL
XFILL_3__7415_ gnd vdd FILL
XFILL_4__16357_ gnd vdd FILL
XFILL_1__12409_ gnd vdd FILL
XFILL_4__13569_ gnd vdd FILL
XFILL_2__14748_ gnd vdd FILL
XFILL_0__15927_ gnd vdd FILL
XFILL_3__8395_ gnd vdd FILL
XFILL_1__16177_ gnd vdd FILL
XFILL_6__14129_ gnd vdd FILL
XFILL_1__13389_ gnd vdd FILL
XFILL_4__15308_ gnd vdd FILL
XFILL_0__7637_ gnd vdd FILL
XSFILL13640x19050 gnd vdd FILL
XFILL_5__14859_ gnd vdd FILL
XFILL_4__16288_ gnd vdd FILL
XFILL_1__15128_ gnd vdd FILL
XFILL_3__7346_ gnd vdd FILL
XFILL_2__14679_ gnd vdd FILL
XFILL_0__15858_ gnd vdd FILL
XFILL_0__7568_ gnd vdd FILL
XFILL_4__15239_ gnd vdd FILL
XFILL_2_BUFX2_insert709 gnd vdd FILL
XFILL_3__15969_ gnd vdd FILL
XFILL_0__14809_ gnd vdd FILL
XFILL_1__15059_ gnd vdd FILL
XFILL_1__8100_ gnd vdd FILL
XFILL_0__15789_ gnd vdd FILL
X_9935_ _9933_/Y _9917_/B _9935_/C gnd _9971_/D vdd OAI21X1
XFILL_1__9080_ gnd vdd FILL
XFILL_3__9016_ gnd vdd FILL
XSFILL54120x33050 gnd vdd FILL
XFILL_0__7499_ gnd vdd FILL
XFILL_2__16349_ gnd vdd FILL
XFILL_0__9238_ gnd vdd FILL
X_9866_ _9864_/Y _9865_/A _9866_/C gnd _9948_/D vdd OAI21X1
X_8817_ _8817_/Q _9834_/CLK _7793_/R vdd _8817_/D gnd vdd DFFSR
XFILL_0__9169_ gnd vdd FILL
X_9797_ _9798_/B _9797_/B gnd _9797_/Y vdd NAND2X1
XFILL_4__6972_ gnd vdd FILL
XFILL_4__9760_ gnd vdd FILL
XSFILL8600x62050 gnd vdd FILL
XBUFX2_insert708 _12816_/Q gnd _12770_/A vdd BUFX2
X_8748_ _8808_/Q gnd _8748_/Y vdd INVX1
XFILL_1__9982_ gnd vdd FILL
XFILL_3__9918_ gnd vdd FILL
XBUFX2_insert719 _13418_/Y gnd _13420_/B vdd BUFX2
XFILL_4__8711_ gnd vdd FILL
XFILL_6_BUFX2_insert664 gnd vdd FILL
XFILL_6__9627_ gnd vdd FILL
X_8679_ _8617_/A _8679_/CLK _9959_/R vdd _8679_/D gnd vdd DFFSR
XFILL_3__9849_ gnd vdd FILL
XFILL_4__8642_ gnd vdd FILL
XFILL_1__8864_ gnd vdd FILL
XFILL_1_CLKBUF1_insert113 gnd vdd FILL
XFILL_4__8573_ gnd vdd FILL
X_11300_ _11300_/A _11620_/B gnd _11614_/A vdd NAND2X1
XFILL_1_CLKBUF1_insert124 gnd vdd FILL
X_12280_ _12272_/A _11885_/B _12272_/C gnd _12282_/B vdd NAND3X1
XFILL_1__7815_ gnd vdd FILL
XFILL_1_CLKBUF1_insert135 gnd vdd FILL
XSFILL38920x65050 gnd vdd FILL
XFILL_1_CLKBUF1_insert146 gnd vdd FILL
XFILL_1_CLKBUF1_insert157 gnd vdd FILL
XFILL112440x72050 gnd vdd FILL
XFILL_1_CLKBUF1_insert168 gnd vdd FILL
X_11231_ _10997_/B gnd _11231_/Y vdd INVX1
XFILL_1_CLKBUF1_insert179 gnd vdd FILL
XSFILL79000x58050 gnd vdd FILL
XFILL_1__7746_ gnd vdd FILL
XFILL_4__7455_ gnd vdd FILL
XSFILL39000x74050 gnd vdd FILL
X_11162_ _11529_/A _11105_/Y _11527_/B gnd _11162_/Y vdd OAI21X1
XSFILL89320x3050 gnd vdd FILL
XFILL_1__7677_ gnd vdd FILL
XFILL_3_BUFX2_insert510 gnd vdd FILL
X_10113_ _10111_/Y _10191_/B _10113_/C gnd _10113_/Y vdd OAI21X1
XFILL_3_BUFX2_insert521 gnd vdd FILL
XFILL_3_BUFX2_insert532 gnd vdd FILL
XFILL_1__9416_ gnd vdd FILL
X_15970_ _10427_/A _15175_/B _15383_/A _7611_/A gnd _15976_/B vdd AOI22X1
X_11093_ _12162_/Y gnd _11094_/B vdd INVX1
XFILL_4__9125_ gnd vdd FILL
XFILL_3_BUFX2_insert543 gnd vdd FILL
XFILL_3_BUFX2_insert554 gnd vdd FILL
XFILL_3_BUFX2_insert565 gnd vdd FILL
XSFILL18840x32050 gnd vdd FILL
X_10044_ _9985_/B _9532_/B gnd _10045_/C vdd NAND2X1
X_14921_ _9040_/A gnd _16263_/A vdd INVX1
XFILL_3_BUFX2_insert576 gnd vdd FILL
XSFILL44120x65050 gnd vdd FILL
XFILL_1__9347_ gnd vdd FILL
XFILL_2__8140_ gnd vdd FILL
XFILL_3_BUFX2_insert587 gnd vdd FILL
XFILL_3_BUFX2_insert598 gnd vdd FILL
XSFILL99320x30050 gnd vdd FILL
XSFILL89800x9050 gnd vdd FILL
X_14852_ _8909_/A gnd _14852_/Y vdd INVX1
XFILL_1__9278_ gnd vdd FILL
XFILL_2__8071_ gnd vdd FILL
XFILL_4__8007_ gnd vdd FILL
X_13803_ _13803_/A _13801_/Y _14567_/A _13802_/Y gnd _13804_/C vdd OAI22X1
XFILL_1__8229_ gnd vdd FILL
XFILL_5__10540_ gnd vdd FILL
X_14783_ _7921_/Q _13865_/B _13865_/C _7751_/A gnd _14783_/Y vdd AOI22X1
X_11995_ _12007_/A _12349_/A _12059_/C gnd _11998_/A vdd NAND3X1
XFILL_6_BUFX2_insert14 gnd vdd FILL
XFILL_2__10360_ gnd vdd FILL
XSFILL64040x16050 gnd vdd FILL
XFILL_6__11830_ gnd vdd FILL
X_13734_ _13733_/Y _13730_/Y gnd _13737_/C vdd NOR2X1
X_10946_ _10944_/A _10944_/B gnd _10946_/Y vdd NAND2X1
XFILL_3__11650_ gnd vdd FILL
XFILL_0__11470_ gnd vdd FILL
XFILL_2__10291_ gnd vdd FILL
XFILL_5__12210_ gnd vdd FILL
XFILL_5__8751_ gnd vdd FILL
X_13665_ _13865_/C _7682_/A _7554_/A _13848_/C gnd _13665_/Y vdd AOI22X1
XFILL_2__12030_ gnd vdd FILL
X_10877_ _12111_/A gnd _10877_/Y vdd INVX1
XFILL_0__10421_ gnd vdd FILL
XSFILL89240x82050 gnd vdd FILL
XFILL_2__8973_ gnd vdd FILL
XFILL_3__11581_ gnd vdd FILL
XFILL_4__8909_ gnd vdd FILL
XFILL_1__12760_ gnd vdd FILL
XFILL_5__7702_ gnd vdd FILL
XFILL_6__13500_ gnd vdd FILL
XFILL_0_BUFX2_insert400 gnd vdd FILL
X_12616_ vdd memoryOutData[16] gnd _12617_/C vdd NAND2X1
X_15404_ _15404_/A _15683_/B _15683_/C _15403_/Y gnd _15405_/A vdd OAI22X1
XFILL_0_BUFX2_insert411 gnd vdd FILL
XFILL_3__13320_ gnd vdd FILL
X_16384_ _16438_/Q gnd _16386_/A vdd INVX1
XFILL_4__9889_ gnd vdd FILL
XFILL_5__12141_ gnd vdd FILL
XSFILL113800x40050 gnd vdd FILL
XFILL_0_BUFX2_insert422 gnd vdd FILL
X_13596_ _9983_/A gnd _13596_/Y vdd INVX1
XFILL_3__10532_ gnd vdd FILL
XFILL_0_BUFX2_insert433 gnd vdd FILL
XFILL_0__13140_ gnd vdd FILL
XFILL_4__12871_ gnd vdd FILL
XFILL_1__11711_ gnd vdd FILL
XFILL_0_BUFX2_insert444 gnd vdd FILL
X_15335_ _15335_/A _15334_/Y gnd _15335_/Y vdd NOR2X1
XFILL_0_BUFX2_insert455 gnd vdd FILL
XFILL_5__7633_ gnd vdd FILL
XFILL_0_BUFX2_insert466 gnd vdd FILL
XFILL_4__14610_ gnd vdd FILL
XFILL_5__12072_ gnd vdd FILL
X_12547_ _12035_/B _13184_/CLK _8033_/R vdd _12477_/Y gnd vdd DFFSR
XSFILL84200x29050 gnd vdd FILL
XFILL_3__13251_ gnd vdd FILL
XFILL_4__11822_ gnd vdd FILL
XFILL_0_BUFX2_insert477 gnd vdd FILL
XFILL_2__7855_ gnd vdd FILL
XFILL_4__15590_ gnd vdd FILL
XFILL_1__14430_ gnd vdd FILL
XSFILL94360x73050 gnd vdd FILL
XFILL_2__13981_ gnd vdd FILL
XFILL_0_BUFX2_insert488 gnd vdd FILL
XFILL_1__11642_ gnd vdd FILL
XFILL_5__7564_ gnd vdd FILL
XFILL_5__15900_ gnd vdd FILL
XFILL_0__10283_ gnd vdd FILL
XFILL_5__11023_ gnd vdd FILL
XFILL_0_BUFX2_insert499 gnd vdd FILL
XFILL_6__16150_ gnd vdd FILL
XFILL_6__13362_ gnd vdd FILL
XFILL_3__12202_ gnd vdd FILL
X_15266_ _7771_/Q _15969_/C gnd _15273_/A vdd NAND2X1
XFILL_4__14541_ gnd vdd FILL
X_12478_ _12382_/A gnd _12480_/A vdd INVX1
XFILL_0__6870_ gnd vdd FILL
XFILL_2__15720_ gnd vdd FILL
XFILL_0__12022_ gnd vdd FILL
XFILL_4__11753_ gnd vdd FILL
XFILL_3__10394_ gnd vdd FILL
XFILL_1__14361_ gnd vdd FILL
XSFILL99400x10050 gnd vdd FILL
XFILL_6__15101_ gnd vdd FILL
X_14217_ _14217_/A _14217_/B _14265_/C gnd _12997_/B vdd AOI21X1
XFILL_1__11573_ gnd vdd FILL
XFILL_5__7495_ gnd vdd FILL
XFILL_5__15831_ gnd vdd FILL
X_11429_ _11429_/A _11242_/Y _11251_/Y gnd _11431_/B vdd OAI21X1
X_15197_ _13616_/Y _15197_/B _15197_/C _13600_/Y gnd _15201_/A vdd OAI22X1
XFILL_3__12133_ gnd vdd FILL
XFILL_1__16100_ gnd vdd FILL
XFILL_4__10704_ gnd vdd FILL
XFILL_1__13312_ gnd vdd FILL
XFILL_2__9525_ gnd vdd FILL
XFILL_4__14472_ gnd vdd FILL
XFILL_2__15651_ gnd vdd FILL
XFILL_4__11684_ gnd vdd FILL
XFILL_1__10524_ gnd vdd FILL
XFILL_2__12863_ gnd vdd FILL
XFILL_5__9234_ gnd vdd FILL
XFILL_1__14292_ gnd vdd FILL
XFILL_4__16211_ gnd vdd FILL
X_14148_ _9572_/Q gnd _14149_/D vdd INVX1
XFILL_6__12244_ gnd vdd FILL
XFILL_4__10635_ gnd vdd FILL
XFILL_2__14602_ gnd vdd FILL
XFILL_4__13423_ gnd vdd FILL
XFILL_5__15762_ gnd vdd FILL
XFILL_1__16031_ gnd vdd FILL
XFILL_5__12974_ gnd vdd FILL
XCLKBUF1_insert112 CLKBUF1_insert216/A gnd _7406_/CLK vdd CLKBUF1
XFILL_3__12064_ gnd vdd FILL
XFILL_2__11814_ gnd vdd FILL
XFILL_1__13243_ gnd vdd FILL
XCLKBUF1_insert123 CLKBUF1_insert220/A gnd _7778_/CLK vdd CLKBUF1
XFILL_2__15582_ gnd vdd FILL
XFILL_5__9165_ gnd vdd FILL
XCLKBUF1_insert134 CLKBUF1_insert169/A gnd _8297_/CLK vdd CLKBUF1
XFILL_5__14713_ gnd vdd FILL
XSFILL74280x40050 gnd vdd FILL
XCLKBUF1_insert145 CLKBUF1_insert150/A gnd _9953_/CLK vdd CLKBUF1
XFILL_0__13973_ gnd vdd FILL
XFILL_0__8471_ gnd vdd FILL
XFILL_3__7200_ gnd vdd FILL
XFILL_5__11925_ gnd vdd FILL
XFILL_4__16142_ gnd vdd FILL
X_14079_ _7523_/Q gnd _15589_/B vdd INVX1
XFILL_3__11015_ gnd vdd FILL
XFILL_4__13354_ gnd vdd FILL
XCLKBUF1_insert156 CLKBUF1_insert218/A gnd _7261_/CLK vdd CLKBUF1
XFILL_2__14533_ gnd vdd FILL
XFILL_5__15693_ gnd vdd FILL
XFILL_4__10566_ gnd vdd FILL
XFILL_0__15712_ gnd vdd FILL
XFILL_5__8116_ gnd vdd FILL
XFILL_2__9387_ gnd vdd FILL
XCLKBUF1_insert167 CLKBUF1_insert182/A gnd _9077_/CLK vdd CLKBUF1
XFILL_2__11745_ gnd vdd FILL
XCLKBUF1_insert178 CLKBUF1_insert220/A gnd _8562_/CLK vdd CLKBUF1
XFILL_1__13174_ gnd vdd FILL
XFILL_1__10386_ gnd vdd FILL
XFILL_5__9096_ gnd vdd FILL
XCLKBUF1_insert189 CLKBUF1_insert182/A gnd _7515_/CLK vdd CLKBUF1
XFILL_0__7422_ gnd vdd FILL
XFILL_5__14644_ gnd vdd FILL
XSFILL89320x62050 gnd vdd FILL
XSFILL53960x39050 gnd vdd FILL
XFILL_4__12305_ gnd vdd FILL
XFILL_4__13285_ gnd vdd FILL
XFILL_3__15823_ gnd vdd FILL
XFILL_2__8338_ gnd vdd FILL
XFILL_5__11856_ gnd vdd FILL
XFILL_4__16073_ gnd vdd FILL
XFILL_4__10497_ gnd vdd FILL
XFILL_2__14464_ gnd vdd FILL
XFILL_1__12125_ gnd vdd FILL
XFILL_0__15643_ gnd vdd FILL
XFILL_2__11676_ gnd vdd FILL
XFILL_0__12855_ gnd vdd FILL
XFILL_5__10807_ gnd vdd FILL
XFILL_2__16203_ gnd vdd FILL
XFILL_4__15024_ gnd vdd FILL
XFILL_0__7353_ gnd vdd FILL
XFILL_4__12236_ gnd vdd FILL
XFILL_6__11057_ gnd vdd FILL
XFILL_5__14575_ gnd vdd FILL
XFILL_2__13415_ gnd vdd FILL
XSFILL28760x15050 gnd vdd FILL
XFILL_2__8269_ gnd vdd FILL
XFILL_2__10627_ gnd vdd FILL
X_7981_ _7972_/A _9517_/B gnd _7982_/C vdd NAND2X1
XFILL_5__11787_ gnd vdd FILL
XFILL_3__7062_ gnd vdd FILL
XFILL_3__15754_ gnd vdd FILL
XFILL_1__12056_ gnd vdd FILL
XFILL_2__14395_ gnd vdd FILL
XFILL_0__11806_ gnd vdd FILL
XFILL_3__12966_ gnd vdd FILL
XSFILL109080x70050 gnd vdd FILL
XFILL_5__16314_ gnd vdd FILL
XFILL_0__15574_ gnd vdd FILL
XFILL_0__12786_ gnd vdd FILL
X_9720_ _9718_/Y _9737_/A _9720_/C gnd _9814_/D vdd OAI21X1
XFILL_5__13526_ gnd vdd FILL
XFILL_3__14705_ gnd vdd FILL
XFILL_4__12167_ gnd vdd FILL
X_6932_ _7008_/Q gnd _6932_/Y vdd INVX1
XFILL_2__16134_ gnd vdd FILL
XFILL_2__13346_ gnd vdd FILL
XFILL_3__11917_ gnd vdd FILL
XFILL_1__11007_ gnd vdd FILL
XFILL_2__10558_ gnd vdd FILL
XFILL_3__15685_ gnd vdd FILL
XFILL_3__12897_ gnd vdd FILL
XFILL_0__14525_ gnd vdd FILL
XFILL_0__9023_ gnd vdd FILL
XFILL_0__11737_ gnd vdd FILL
XFILL_4__11118_ gnd vdd FILL
XFILL_5__16245_ gnd vdd FILL
XFILL_5__13457_ gnd vdd FILL
XFILL_5__9998_ gnd vdd FILL
X_9651_ _9652_/B _9779_/B gnd _9651_/Y vdd NAND2X1
XFILL_3__14636_ gnd vdd FILL
X_6863_ _6863_/A gnd memoryAddress[25] vdd BUFX2
XFILL_4__12098_ gnd vdd FILL
XFILL_5__10669_ gnd vdd FILL
XFILL_1__15815_ gnd vdd FILL
XFILL_2__16065_ gnd vdd FILL
XFILL_3__11848_ gnd vdd FILL
XFILL_2__13277_ gnd vdd FILL
XFILL_0__14456_ gnd vdd FILL
XFILL_2__10489_ gnd vdd FILL
XFILL_5__12408_ gnd vdd FILL
X_8602_ _8602_/A gnd _8604_/A vdd INVX1
XFILL_0__11668_ gnd vdd FILL
XFILL_4__15926_ gnd vdd FILL
XFILL_5__16176_ gnd vdd FILL
XFILL_2__15016_ gnd vdd FILL
XFILL_4__11049_ gnd vdd FILL
X_9582_ _9534_/A _8165_/CLK _9046_/R vdd _9582_/D gnd vdd DFFSR
XFILL_5__13388_ gnd vdd FILL
XFILL_2__12228_ gnd vdd FILL
XFILL_3__14567_ gnd vdd FILL
XFILL_0__13407_ gnd vdd FILL
XFILL_1__15746_ gnd vdd FILL
XFILL_3__11779_ gnd vdd FILL
XFILL_3__7964_ gnd vdd FILL
XFILL_0__10619_ gnd vdd FILL
XFILL_1__12958_ gnd vdd FILL
XFILL_0__14387_ gnd vdd FILL
XFILL_0__11599_ gnd vdd FILL
XFILL_5__15127_ gnd vdd FILL
X_8533_ _8533_/A _8440_/B _8532_/Y gnd _8533_/Y vdd OAI21X1
XFILL_5__12339_ gnd vdd FILL
XFILL_3__16306_ gnd vdd FILL
XFILL_5_BUFX2_insert605 gnd vdd FILL
XFILL_3__13518_ gnd vdd FILL
XFILL_4__15857_ gnd vdd FILL
XFILL_3__14498_ gnd vdd FILL
XFILL_1__11909_ gnd vdd FILL
XFILL_3__6915_ gnd vdd FILL
XFILL_5_BUFX2_insert616 gnd vdd FILL
XFILL_2__12159_ gnd vdd FILL
XFILL_0__16126_ gnd vdd FILL
XFILL_0__13338_ gnd vdd FILL
XFILL_1__15677_ gnd vdd FILL
XFILL_5_BUFX2_insert627 gnd vdd FILL
XFILL_1__12889_ gnd vdd FILL
XFILL_5_BUFX2_insert638 gnd vdd FILL
XFILL_4__14808_ gnd vdd FILL
XFILL_5__15058_ gnd vdd FILL
XFILL_0__9925_ gnd vdd FILL
XSFILL49000x37050 gnd vdd FILL
X_8464_ _8464_/A _8508_/A _8464_/C gnd _8542_/D vdd OAI21X1
XFILL_3__16237_ gnd vdd FILL
XFILL_5_BUFX2_insert649 gnd vdd FILL
XFILL_1__14628_ gnd vdd FILL
XFILL_3__9634_ gnd vdd FILL
XFILL_3__6846_ gnd vdd FILL
XFILL_3__13449_ gnd vdd FILL
XFILL_4__15788_ gnd vdd FILL
XSFILL59160x81050 gnd vdd FILL
XSFILL89400x42050 gnd vdd FILL
XFILL_0__16057_ gnd vdd FILL
XFILL_0__13269_ gnd vdd FILL
XFILL_6__9343_ gnd vdd FILL
XFILL_5__14009_ gnd vdd FILL
X_7415_ _8951_/A _7416_/B gnd _7415_/Y vdd NAND2X1
XSFILL109560x48050 gnd vdd FILL
XFILL_0__9856_ gnd vdd FILL
XFILL_4__14739_ gnd vdd FILL
XFILL_2__15918_ gnd vdd FILL
X_8395_ _8321_/B _7883_/B gnd _8395_/Y vdd NAND2X1
XFILL_3__16168_ gnd vdd FILL
XFILL_0__15008_ gnd vdd FILL
XFILL_1__14559_ gnd vdd FILL
XFILL_1__7600_ gnd vdd FILL
XFILL_0__9787_ gnd vdd FILL
XFILL_1__8580_ gnd vdd FILL
XFILL_3__15119_ gnd vdd FILL
X_7346_ _7402_/Q gnd _7346_/Y vdd INVX1
XFILL_3__8516_ gnd vdd FILL
XFILL_3__16099_ gnd vdd FILL
XFILL_3__9496_ gnd vdd FILL
XFILL_2__15849_ gnd vdd FILL
XFILL_4__16409_ gnd vdd FILL
XFILL_0__8738_ gnd vdd FILL
XFILL_2_CLKBUF1_insert208 gnd vdd FILL
XFILL_3__8447_ gnd vdd FILL
X_7277_ _7277_/Q _8429_/CLK _7533_/R vdd _7229_/Y gnd vdd DFFSR
XFILL_1__16229_ gnd vdd FILL
XFILL_2_CLKBUF1_insert219 gnd vdd FILL
XFILL_4__7240_ gnd vdd FILL
XSFILL13720x2050 gnd vdd FILL
X_9016_ _9016_/A gnd _9016_/Y vdd INVX1
XFILL_1__7462_ gnd vdd FILL
XFILL_3__8378_ gnd vdd FILL
XFILL_4__7171_ gnd vdd FILL
XFILL_6__8087_ gnd vdd FILL
XSFILL18760x47050 gnd vdd FILL
XFILL_3__7329_ gnd vdd FILL
XFILL_2_BUFX2_insert506 gnd vdd FILL
XFILL_2_BUFX2_insert517 gnd vdd FILL
XFILL_6__7038_ gnd vdd FILL
XFILL_2_BUFX2_insert528 gnd vdd FILL
XFILL_1__9132_ gnd vdd FILL
XFILL_2_BUFX2_insert539 gnd vdd FILL
X_9918_ _9918_/A gnd _9918_/Y vdd INVX1
X_10800_ _10822_/B _9008_/B gnd _10801_/C vdd NAND2X1
XFILL_1__8014_ gnd vdd FILL
X_11780_ _11779_/Y _11778_/Y gnd _11784_/A vdd NOR2X1
X_9849_ _9849_/A gnd _9851_/A vdd INVX1
XFILL_6_BUFX2_insert1047 gnd vdd FILL
XFILL_4__9812_ gnd vdd FILL
XFILL112440x67050 gnd vdd FILL
XFILL_6_BUFX2_insert1058 gnd vdd FILL
X_10731_ _10677_/A _9195_/CLK _8051_/R vdd _10731_/D gnd vdd DFFSR
XBUFX2_insert505 BUFX2_insert607/A gnd _8418_/R vdd BUFX2
XFILL_4__9743_ gnd vdd FILL
XBUFX2_insert516 BUFX2_insert556/A gnd _8053_/R vdd BUFX2
X_13450_ _13449_/Y _13450_/B gnd _13451_/C vdd NOR2X1
XSFILL79160x12050 gnd vdd FILL
XFILL_4__6955_ gnd vdd FILL
XSFILL39000x69050 gnd vdd FILL
X_10662_ _15704_/B gnd _10664_/A vdd INVX1
XBUFX2_insert527 BUFX2_insert494/A gnd _7523_/R vdd BUFX2
XBUFX2_insert538 BUFX2_insert556/A gnd _7276_/R vdd BUFX2
XBUFX2_insert549 BUFX2_insert559/A gnd _9062_/R vdd BUFX2
X_12401_ _12359_/A _12624_/A gnd _12402_/C vdd NAND2X1
XFILL_4__9674_ gnd vdd FILL
XFILL_4__6886_ gnd vdd FILL
X_13381_ _13381_/A _13381_/B _13398_/A gnd _13381_/Y vdd NAND3X1
X_10593_ _13983_/A _7268_/CLK _8688_/R vdd _10521_/Y gnd vdd DFFSR
XFILL_1__8916_ gnd vdd FILL
XFILL_1__9896_ gnd vdd FILL
XFILL_4__8625_ gnd vdd FILL
X_15120_ _9431_/Q _15794_/B _15764_/C gnd _15121_/C vdd NAND3X1
X_12332_ _12312_/A _12340_/B _12312_/C gnd _12332_/Y vdd NAND3X1
XFILL_4_BUFX2_insert1040 gnd vdd FILL
XFILL_4_BUFX2_insert1051 gnd vdd FILL
XFILL_1__8847_ gnd vdd FILL
XFILL_4_BUFX2_insert1062 gnd vdd FILL
XFILL_4_BUFX2_insert1073 gnd vdd FILL
XFILL_4_BUFX2_insert1084 gnd vdd FILL
X_15051_ _12813_/Q _12812_/Q _14989_/A gnd _15051_/Y vdd NOR3X1
X_12263_ _12239_/A gnd _12239_/C gnd _12263_/Y vdd NAND3X1
XSFILL69080x64050 gnd vdd FILL
XFILL_1__8778_ gnd vdd FILL
XFILL_2__7571_ gnd vdd FILL
X_14002_ _9057_/Q gnd _14002_/Y vdd INVX1
XFILL_4__7507_ gnd vdd FILL
XFILL_4__8487_ gnd vdd FILL
X_11214_ _10889_/Y gnd _11214_/Y vdd INVX2
X_12194_ _12150_/B _12901_/A gnd _12195_/C vdd NAND2X1
XFILL_1__7729_ gnd vdd FILL
XSFILL99480x4050 gnd vdd FILL
XFILL_4__7438_ gnd vdd FILL
XFILL_4__10420_ gnd vdd FILL
X_11145_ _11591_/A _11126_/A gnd _11146_/B vdd NOR2X1
XSFILL53560x7050 gnd vdd FILL
XFILL_2__9241_ gnd vdd FILL
XFILL_1__10240_ gnd vdd FILL
XFILL_3_BUFX2_insert340 gnd vdd FILL
XFILL_4__7369_ gnd vdd FILL
XFILL_3_BUFX2_insert351 gnd vdd FILL
XFILL_0__10970_ gnd vdd FILL
XFILL_5__11710_ gnd vdd FILL
XSFILL23800x82050 gnd vdd FILL
X_15953_ _15953_/A _15953_/B _15521_/C _14509_/A gnd _15954_/B vdd OAI22X1
XFILL_3_BUFX2_insert362 gnd vdd FILL
X_11076_ _12144_/Y gnd _11076_/Y vdd INVX1
XFILL_3_BUFX2_insert373 gnd vdd FILL
XFILL_2__11530_ gnd vdd FILL
XFILL_2__9172_ gnd vdd FILL
XFILL_1__10171_ gnd vdd FILL
XFILL_3_BUFX2_insert384 gnd vdd FILL
XFILL_4__9108_ gnd vdd FILL
XFILL_3_BUFX2_insert395 gnd vdd FILL
X_14904_ _14904_/A _14697_/B _14752_/C _16254_/C gnd _14904_/Y vdd OAI22X1
X_10027_ _10025_/Y _9979_/B _10027_/C gnd _10027_/Y vdd OAI21X1
XFILL_2__8123_ gnd vdd FILL
XFILL_5__11641_ gnd vdd FILL
XFILL_4__10282_ gnd vdd FILL
X_15884_ _16089_/B _15884_/B _15883_/Y _15848_/A gnd _15884_/Y vdd OAI22X1
XFILL_2__11461_ gnd vdd FILL
XFILL_4__9039_ gnd vdd FILL
XFILL_0__12640_ gnd vdd FILL
XFILL_5__9921_ gnd vdd FILL
XFILL_4__12021_ gnd vdd FILL
X_14835_ _7245_/A _13619_/B _14626_/A _7411_/Q gnd _14846_/A vdd AOI22X1
XFILL_5__14360_ gnd vdd FILL
XFILL_3__12751_ gnd vdd FILL
XFILL_2__10412_ gnd vdd FILL
XFILL_5__11572_ gnd vdd FILL
XFILL_2__8054_ gnd vdd FILL
XFILL_2__14180_ gnd vdd FILL
XFILL_1__13930_ gnd vdd FILL
XFILL_2__11392_ gnd vdd FILL
XFILL_5__13311_ gnd vdd FILL
XFILL_0__12571_ gnd vdd FILL
XFILL_5__9852_ gnd vdd FILL
XFILL_5__10523_ gnd vdd FILL
XFILL_3__11702_ gnd vdd FILL
XFILL_6__12862_ gnd vdd FILL
XFILL_2__13131_ gnd vdd FILL
X_11978_ _11969_/A _12107_/B gnd _11978_/Y vdd NAND2X1
X_14766_ _9671_/A gnd _14768_/C vdd INVX1
XFILL_5__14291_ gnd vdd FILL
XFILL_0__14310_ gnd vdd FILL
XFILL_3__15470_ gnd vdd FILL
XFILL_1__13861_ gnd vdd FILL
XFILL_0__11522_ gnd vdd FILL
XFILL_5__16030_ gnd vdd FILL
XFILL_0__15290_ gnd vdd FILL
XFILL_5__9783_ gnd vdd FILL
XFILL_5__13242_ gnd vdd FILL
X_10929_ _10929_/A _10938_/B gnd _10936_/B vdd NOR2X1
X_13717_ _7813_/A _13865_/B _13717_/C gnd _13717_/Y vdd AOI21X1
XFILL_5__6995_ gnd vdd FILL
X_14697_ _16099_/A _14697_/B _14697_/C _16090_/A gnd _14701_/A vdd OAI22X1
XFILL_3__14421_ gnd vdd FILL
XFILL_3__11633_ gnd vdd FILL
XFILL_1__15600_ gnd vdd FILL
XFILL_4_CLKBUF1_insert130 gnd vdd FILL
XFILL_4__13972_ gnd vdd FILL
XFILL_0__14241_ gnd vdd FILL
XFILL_4_CLKBUF1_insert141 gnd vdd FILL
XFILL_2__10274_ gnd vdd FILL
XFILL_0__11453_ gnd vdd FILL
XFILL_1__13792_ gnd vdd FILL
XFILL_4_CLKBUF1_insert152 gnd vdd FILL
XFILL_5__8734_ gnd vdd FILL
XFILL_4__15711_ gnd vdd FILL
X_16436_ _15826_/A _9953_/CLK _7649_/R vdd _16380_/Y gnd vdd DFFSR
XFILL_4_CLKBUF1_insert163 gnd vdd FILL
X_13648_ _13648_/A _13647_/Y _13648_/C gnd _13664_/B vdd NAND3X1
XFILL_2__12013_ gnd vdd FILL
XFILL_5__13173_ gnd vdd FILL
XFILL_3__14352_ gnd vdd FILL
XFILL_5__10385_ gnd vdd FILL
XFILL_0__10404_ gnd vdd FILL
XFILL_1__15531_ gnd vdd FILL
XFILL_3__11564_ gnd vdd FILL
XFILL_4_CLKBUF1_insert174 gnd vdd FILL
XFILL_1__12743_ gnd vdd FILL
XFILL_4_CLKBUF1_insert185 gnd vdd FILL
XFILL_2__8956_ gnd vdd FILL
XFILL_0_BUFX2_insert230 gnd vdd FILL
XFILL_4_CLKBUF1_insert196 gnd vdd FILL
XFILL_0__14172_ gnd vdd FILL
XFILL_0_BUFX2_insert241 gnd vdd FILL
XFILL_0__11384_ gnd vdd FILL
XFILL_5__12124_ gnd vdd FILL
XSFILL74280x35050 gnd vdd FILL
XFILL_3__13303_ gnd vdd FILL
X_16367_ gnd gnd gnd _16368_/C vdd NAND2X1
XFILL_0__7971_ gnd vdd FILL
XFILL_4__15642_ gnd vdd FILL
XFILL_0_BUFX2_insert252 gnd vdd FILL
X_13579_ _13865_/C _7768_/Q _7128_/Q _14344_/C gnd _13582_/A vdd AOI22X1
XFILL_3__10515_ gnd vdd FILL
XFILL_4__12854_ gnd vdd FILL
XFILL_0_BUFX2_insert263 gnd vdd FILL
XFILL_3__14283_ gnd vdd FILL
XFILL_3__7680_ gnd vdd FILL
XFILL_0_BUFX2_insert274 gnd vdd FILL
XFILL_0__13123_ gnd vdd FILL
XFILL_3__11495_ gnd vdd FILL
XFILL_1__15462_ gnd vdd FILL
XFILL_2__8887_ gnd vdd FILL
XFILL_5__7616_ gnd vdd FILL
XFILL_0_BUFX2_insert285 gnd vdd FILL
XFILL_0_BUFX2_insert296 gnd vdd FILL
XFILL_0__6922_ gnd vdd FILL
X_15318_ _15318_/A _15317_/Y _15318_/C gnd _15318_/Y vdd NOR3X1
XFILL_6__10626_ gnd vdd FILL
XFILL_3__13234_ gnd vdd FILL
XFILL_3__16022_ gnd vdd FILL
XSFILL89320x57050 gnd vdd FILL
XFILL_5__12055_ gnd vdd FILL
X_16298_ _7413_/Q _15789_/B _15794_/B gnd _16299_/C vdd NAND3X1
XFILL_5__8596_ gnd vdd FILL
XSFILL49080x11050 gnd vdd FILL
XFILL_4__11805_ gnd vdd FILL
XFILL_3__10446_ gnd vdd FILL
XFILL_4__15573_ gnd vdd FILL
XFILL_1__14413_ gnd vdd FILL
XFILL_4__12785_ gnd vdd FILL
XFILL_2__7838_ gnd vdd FILL
XFILL_1__11625_ gnd vdd FILL
XFILL_2__13964_ gnd vdd FILL
XFILL_1__15393_ gnd vdd FILL
XFILL_0__10266_ gnd vdd FILL
X_7200_ _7268_/Q gnd _7202_/A vdd INVX1
XFILL_5__7547_ gnd vdd FILL
XFILL_5__11006_ gnd vdd FILL
XFILL_0__9641_ gnd vdd FILL
XFILL_0__6853_ gnd vdd FILL
X_15249_ _13675_/Y _15981_/B _15922_/C _15248_/Y gnd _15249_/Y vdd OAI22X1
XFILL_4__14524_ gnd vdd FILL
XFILL_2__15703_ gnd vdd FILL
XFILL_3__13165_ gnd vdd FILL
XFILL_2__12915_ gnd vdd FILL
XFILL_4__11736_ gnd vdd FILL
XFILL_3__9350_ gnd vdd FILL
X_8180_ _8180_/Q _8180_/CLK _8937_/R vdd _8180_/D gnd vdd DFFSR
XFILL_3__10377_ gnd vdd FILL
XFILL_0__12005_ gnd vdd FILL
XFILL_1__14344_ gnd vdd FILL
XFILL_2__13895_ gnd vdd FILL
XFILL_1__11556_ gnd vdd FILL
XFILL_5__7478_ gnd vdd FILL
XFILL_2_BUFX2_insert12 gnd vdd FILL
XFILL_0__10197_ gnd vdd FILL
XFILL_3__12116_ gnd vdd FILL
XFILL_5__15814_ gnd vdd FILL
XFILL112200x1050 gnd vdd FILL
X_7131_ _7045_/A _8663_/CLK _7131_/R vdd _7131_/D gnd vdd DFFSR
XFILL_2_BUFX2_insert23 gnd vdd FILL
XFILL_2__9508_ gnd vdd FILL
XFILL_4__14455_ gnd vdd FILL
XFILL_2_BUFX2_insert34 gnd vdd FILL
XSFILL94440x48050 gnd vdd FILL
XFILL_1__10507_ gnd vdd FILL
XFILL_2__12846_ gnd vdd FILL
XSFILL14040x59050 gnd vdd FILL
XFILL_2__15634_ gnd vdd FILL
XFILL_3__13096_ gnd vdd FILL
XFILL_2_BUFX2_insert45 gnd vdd FILL
XFILL_3__9281_ gnd vdd FILL
XFILL_4__11667_ gnd vdd FILL
XFILL_5__9217_ gnd vdd FILL
XFILL_2_BUFX2_insert56 gnd vdd FILL
XFILL_1__14275_ gnd vdd FILL
XFILL_0__8523_ gnd vdd FILL
XFILL_1__11487_ gnd vdd FILL
XFILL_4__13406_ gnd vdd FILL
XFILL_2_BUFX2_insert67 gnd vdd FILL
X_7062_ _7060_/Y _7124_/A _7061_/Y gnd _7136_/D vdd OAI21X1
XFILL_5__15745_ gnd vdd FILL
XFILL_1__16014_ gnd vdd FILL
XFILL_3__8232_ gnd vdd FILL
XFILL_2_BUFX2_insert78 gnd vdd FILL
XFILL_3__12047_ gnd vdd FILL
XFILL_4__10618_ gnd vdd FILL
XFILL_5__12957_ gnd vdd FILL
XFILL_1__13226_ gnd vdd FILL
XFILL_2_BUFX2_insert89 gnd vdd FILL
XFILL_2__15565_ gnd vdd FILL
XFILL_4__14386_ gnd vdd FILL
XSFILL69240x24050 gnd vdd FILL
XFILL_2__12777_ gnd vdd FILL
XFILL_1__10438_ gnd vdd FILL
XFILL_4__11598_ gnd vdd FILL
XFILL_5__9148_ gnd vdd FILL
XFILL_0__13956_ gnd vdd FILL
XFILL_5__11908_ gnd vdd FILL
XFILL_4__16125_ gnd vdd FILL
XFILL_0__8454_ gnd vdd FILL
XFILL_4__13337_ gnd vdd FILL
XFILL_5__15676_ gnd vdd FILL
XFILL_4__10549_ gnd vdd FILL
XFILL_5__12888_ gnd vdd FILL
XFILL_2__14516_ gnd vdd FILL
XFILL_2__11728_ gnd vdd FILL
XFILL_1__13157_ gnd vdd FILL
XFILL_0__12907_ gnd vdd FILL
XFILL_2__15496_ gnd vdd FILL
XFILL_1__10369_ gnd vdd FILL
XSFILL104440x33050 gnd vdd FILL
XFILL_0__13887_ gnd vdd FILL
XFILL_5__14627_ gnd vdd FILL
XFILL_5__9079_ gnd vdd FILL
XFILL_3__7114_ gnd vdd FILL
XFILL_3__15806_ gnd vdd FILL
XFILL_0__8385_ gnd vdd FILL
XFILL_4__16056_ gnd vdd FILL
XFILL_5__11839_ gnd vdd FILL
XFILL_4__13268_ gnd vdd FILL
XFILL_1__12108_ gnd vdd FILL
XSFILL8680x31050 gnd vdd FILL
XFILL_2__14447_ gnd vdd FILL
XSFILL33720x65050 gnd vdd FILL
XFILL_0__15626_ gnd vdd FILL
XFILL_2__11659_ gnd vdd FILL
XFILL_3__8094_ gnd vdd FILL
XSFILL74360x15050 gnd vdd FILL
XFILL_1__13088_ gnd vdd FILL
XFILL_3__13998_ gnd vdd FILL
XFILL_0__12838_ gnd vdd FILL
XFILL_0__7336_ gnd vdd FILL
XFILL_4__15007_ gnd vdd FILL
XFILL_5__14558_ gnd vdd FILL
XFILL_4__12219_ gnd vdd FILL
X_7964_ _7964_/A _7972_/A _7963_/Y gnd _7964_/Y vdd OAI21X1
XFILL_3__15737_ gnd vdd FILL
XFILL_3__7045_ gnd vdd FILL
XFILL_1__12039_ gnd vdd FILL
XFILL_2__14378_ gnd vdd FILL
XFILL_0__15557_ gnd vdd FILL
XSFILL89400x37050 gnd vdd FILL
XFILL_0__12769_ gnd vdd FILL
XFILL_5__13509_ gnd vdd FILL
X_9703_ _9641_/A _7527_/CLK _8935_/R vdd _9703_/D gnd vdd DFFSR
X_6915_ _6967_/B _8195_/B gnd _6915_/Y vdd NAND2X1
XFILL_6__15848_ gnd vdd FILL
XFILL_2__13329_ gnd vdd FILL
XFILL_5__14489_ gnd vdd FILL
XFILL_2__16117_ gnd vdd FILL
XFILL_3__15668_ gnd vdd FILL
XFILL_0__14508_ gnd vdd FILL
X_7895_ _7895_/Q _6999_/CLK _7000_/R vdd _7895_/D gnd vdd DFFSR
XFILL_0__9006_ gnd vdd FILL
XFILL111880x75050 gnd vdd FILL
XFILL_5__16228_ gnd vdd FILL
XFILL_0__15488_ gnd vdd FILL
X_9634_ _9632_/Y _9613_/B _9633_/Y gnd _9700_/D vdd OAI21X1
XFILL_6__8774_ gnd vdd FILL
XFILL_3__14619_ gnd vdd FILL
X_6846_ _6846_/A gnd memoryAddress[8] vdd BUFX2
XFILL_0__7198_ gnd vdd FILL
XFILL_2__16048_ gnd vdd FILL
XFILL_3__15599_ gnd vdd FILL
XFILL_0__14439_ gnd vdd FILL
XFILL_3__8996_ gnd vdd FILL
XFILL_6__7725_ gnd vdd FILL
XSFILL13640x32050 gnd vdd FILL
XFILL_4__15909_ gnd vdd FILL
XFILL_5__16159_ gnd vdd FILL
X_9565_ _9565_/Q _9195_/CLK _8051_/R vdd _9485_/Y gnd vdd DFFSR
XFILL_5_BUFX2_insert402 gnd vdd FILL
XFILL_3__7947_ gnd vdd FILL
XFILL_1__15729_ gnd vdd FILL
XFILL_5_BUFX2_insert413 gnd vdd FILL
XFILL_5_BUFX2_insert424 gnd vdd FILL
X_8516_ _8560_/Q gnd _8518_/A vdd INVX1
XFILL_1__9750_ gnd vdd FILL
XFILL_1__6962_ gnd vdd FILL
XFILL_5_BUFX2_insert435 gnd vdd FILL
X_9496_ _9533_/B _8472_/B gnd _9497_/C vdd NAND2X1
XFILL_5_BUFX2_insert446 gnd vdd FILL
XFILL_0__16109_ gnd vdd FILL
XFILL_5_BUFX2_insert457 gnd vdd FILL
XFILL_3__7878_ gnd vdd FILL
XFILL_5_BUFX2_insert468 gnd vdd FILL
XFILL_0__9908_ gnd vdd FILL
XFILL_1__8701_ gnd vdd FILL
X_8447_ _8447_/A gnd _8447_/Y vdd INVX1
XFILL_5_BUFX2_insert479 gnd vdd FILL
XFILL_1__9681_ gnd vdd FILL
XFILL_1__6893_ gnd vdd FILL
XFILL_3__9617_ gnd vdd FILL
XFILL_4__9390_ gnd vdd FILL
XFILL_1__8632_ gnd vdd FILL
XSFILL33800x45050 gnd vdd FILL
X_8378_ _8378_/A _8360_/B _8377_/Y gnd _8428_/D vdd OAI21X1
XFILL_4__8341_ gnd vdd FILL
XFILL_3__9548_ gnd vdd FILL
X_7329_ _7308_/A _7329_/B gnd _7329_/Y vdd NAND2X1
XFILL_4__8272_ gnd vdd FILL
XFILL_3__9479_ gnd vdd FILL
XSFILL23880x3050 gnd vdd FILL
XFILL_4__7223_ gnd vdd FILL
XFILL_1__8494_ gnd vdd FILL
XFILL_1__7445_ gnd vdd FILL
XFILL112360x7050 gnd vdd FILL
XSFILL13720x12050 gnd vdd FILL
XFILL_2_BUFX2_insert303 gnd vdd FILL
X_12950_ _12950_/Q _7020_/CLK _8053_/R vdd _12918_/Y gnd vdd DFFSR
XFILL112040x64050 gnd vdd FILL
XFILL_2_BUFX2_insert314 gnd vdd FILL
XFILL_1__7376_ gnd vdd FILL
XFILL_2_BUFX2_insert325 gnd vdd FILL
XFILL_2_BUFX2_insert336 gnd vdd FILL
X_11901_ _11901_/A _11900_/A _11901_/C gnd _6842_/A vdd OAI21X1
XFILL_4__7085_ gnd vdd FILL
XFILL_2_BUFX2_insert347 gnd vdd FILL
XFILL_1__9115_ gnd vdd FILL
XFILL_2_BUFX2_insert358 gnd vdd FILL
X_12881_ vdd _12881_/B gnd _12882_/C vdd NAND2X1
XFILL_2_BUFX2_insert369 gnd vdd FILL
XSFILL69240x2050 gnd vdd FILL
X_14620_ _7790_/Q gnd _14620_/Y vdd INVX1
X_11832_ _11764_/A _11835_/A _11238_/Y _11223_/B gnd _11834_/B vdd AOI22X1
XSFILL114600x78050 gnd vdd FILL
X_14551_ _9197_/Q gnd _14551_/Y vdd INVX1
X_11763_ _11245_/Y _11758_/Y _11763_/C gnd _11763_/Y vdd AOI21X1
XBUFX2_insert302 _12414_/Y gnd _7868_/B vdd BUFX2
X_10714_ _15235_/A _9818_/CLK _9441_/R vdd _10714_/D gnd vdd DFFSR
X_13502_ _13498_/Y _13502_/B gnd _13503_/C vdd NOR2X1
X_14482_ _8939_/Q _14482_/B _13854_/B _9269_/A gnd _14482_/Y vdd AOI22X1
XBUFX2_insert313 _13454_/Y gnd _13857_/C vdd BUFX2
XFILL_4__7987_ gnd vdd FILL
XBUFX2_insert324 _13345_/Y gnd _9896_/B vdd BUFX2
X_11694_ _11066_/Y _11846_/C _11693_/Y gnd _11698_/A vdd OAI21X1
XFILL_6_BUFX2_insert280 gnd vdd FILL
XBUFX2_insert335 _13494_/Y gnd _13647_/B vdd BUFX2
XFILL_2__9790_ gnd vdd FILL
XFILL_4__9726_ gnd vdd FILL
XSFILL104280x68050 gnd vdd FILL
X_16221_ _15187_/A _14854_/Y _15187_/C gnd _16243_/B vdd NOR3X1
X_13433_ _13433_/A _14636_/C gnd _13434_/C vdd NOR2X1
XFILL_4__6938_ gnd vdd FILL
XBUFX2_insert346 _12396_/Y gnd _9898_/B vdd BUFX2
XBUFX2_insert357 _13306_/Y gnd _7997_/B vdd BUFX2
XFILL_5__10170_ gnd vdd FILL
X_10645_ _10681_/A _7061_/B gnd _10645_/Y vdd NAND2X1
XBUFX2_insert368 _13338_/Y gnd _9548_/B vdd BUFX2
XFILL_5_CLKBUF1_insert203 gnd vdd FILL
XFILL_2__8741_ gnd vdd FILL
XBUFX2_insert379 _12211_/Y gnd _12311_/C vdd BUFX2
XFILL_5_CLKBUF1_insert214 gnd vdd FILL
XFILL_5__8450_ gnd vdd FILL
XFILL_4__9657_ gnd vdd FILL
X_16152_ _16152_/A _16151_/Y gnd _16152_/Y vdd NOR2X1
X_13364_ _13361_/A _13363_/Y gnd _13364_/Y vdd NOR2X1
XFILL_3__10300_ gnd vdd FILL
XFILL_4__6869_ gnd vdd FILL
XSFILL23800x77050 gnd vdd FILL
X_10576_ _16246_/A gnd _10578_/A vdd INVX1
XFILL_0__10120_ gnd vdd FILL
XFILL_3__11280_ gnd vdd FILL
XFILL_4__8608_ gnd vdd FILL
XFILL_1__9879_ gnd vdd FILL
XFILL_5_BUFX2_insert980 gnd vdd FILL
XFILL_5__8381_ gnd vdd FILL
XFILL_5_BUFX2_insert991 gnd vdd FILL
XFILL112120x44050 gnd vdd FILL
X_12315_ _12227_/A gnd _12307_/C gnd _12318_/A vdd NAND3X1
X_15103_ _15103_/A _15094_/Y _15103_/C gnd _15127_/A vdd NOR3X1
XSFILL24440x43050 gnd vdd FILL
X_16083_ _15842_/A _16083_/B _16083_/C _16137_/C gnd _16084_/B vdd OAI22X1
X_13295_ _13295_/A _13294_/Y _13295_/C gnd _13295_/Y vdd OAI21X1
XSFILL48760x81050 gnd vdd FILL
XFILL_3__10231_ gnd vdd FILL
XFILL_2__7623_ gnd vdd FILL
XFILL_4__12570_ gnd vdd FILL
XFILL_1__11410_ gnd vdd FILL
XFILL_2__10961_ gnd vdd FILL
XFILL_5__7332_ gnd vdd FILL
XFILL_0__10051_ gnd vdd FILL
XFILL_1__12390_ gnd vdd FILL
X_15034_ _14981_/Y _15212_/B _15044_/C gnd _15035_/B vdd OAI21X1
XFILL_6__13130_ gnd vdd FILL
X_12246_ _12246_/A _12246_/B _12246_/C gnd _11384_/A vdd NAND3X1
XFILL_2__12700_ gnd vdd FILL
XFILL_5__13860_ gnd vdd FILL
XFILL_4__11521_ gnd vdd FILL
XFILL_2__7554_ gnd vdd FILL
XFILL_3__10162_ gnd vdd FILL
XFILL_2__13680_ gnd vdd FILL
XFILL_1__11341_ gnd vdd FILL
XFILL_2__10892_ gnd vdd FILL
XFILL_4__14240_ gnd vdd FILL
X_12177_ _12177_/A _12123_/B _12176_/Y gnd _12177_/Y vdd OAI21X1
XFILL_2__12631_ gnd vdd FILL
XFILL_5__13791_ gnd vdd FILL
XFILL_4__11452_ gnd vdd FILL
XFILL_2__7485_ gnd vdd FILL
XFILL_0__13810_ gnd vdd FILL
XFILL_1__14060_ gnd vdd FILL
XFILL_3__14970_ gnd vdd FILL
XFILL_5__9002_ gnd vdd FILL
XFILL_1__11272_ gnd vdd FILL
XFILL_5__15530_ gnd vdd FILL
XFILL_5__7194_ gnd vdd FILL
XSFILL69160x39050 gnd vdd FILL
X_11128_ _11591_/A gnd _11590_/A vdd INVX1
XFILL_0__14790_ gnd vdd FILL
XFILL_4__10403_ gnd vdd FILL
XFILL_5__12742_ gnd vdd FILL
XFILL_2__9224_ gnd vdd FILL
XFILL_2__15350_ gnd vdd FILL
XFILL_4__14171_ gnd vdd FILL
XSFILL3640x4050 gnd vdd FILL
XFILL_3__13921_ gnd vdd FILL
XFILL_4__11383_ gnd vdd FILL
XFILL_1__13011_ gnd vdd FILL
XFILL_0__13741_ gnd vdd FILL
XFILL_0__10953_ gnd vdd FILL
X_15936_ _15934_/Y _15936_/B _15936_/C gnd _15943_/A vdd NAND3X1
XFILL_4__13122_ gnd vdd FILL
XFILL_2__14301_ gnd vdd FILL
X_11059_ _12274_/Y _12159_/Y gnd _11059_/Y vdd AND2X2
XFILL_5__15461_ gnd vdd FILL
XFILL_2__9155_ gnd vdd FILL
XFILL_2__11513_ gnd vdd FILL
XFILL_3__13852_ gnd vdd FILL
XSFILL104360x48050 gnd vdd FILL
XFILL_2__15281_ gnd vdd FILL
XFILL_2__12493_ gnd vdd FILL
XFILL_1__10154_ gnd vdd FILL
XFILL_0__13672_ gnd vdd FILL
XFILL_5__14412_ gnd vdd FILL
XFILL_0__10884_ gnd vdd FILL
XFILL_5__11624_ gnd vdd FILL
XFILL_2__8106_ gnd vdd FILL
XFILL_2__14232_ gnd vdd FILL
XFILL_5__15392_ gnd vdd FILL
XFILL_4__10265_ gnd vdd FILL
X_15867_ _15550_/A _14418_/Y _15550_/C gnd _15890_/B vdd NOR3X1
XFILL_0__15411_ gnd vdd FILL
XFILL_2__9086_ gnd vdd FILL
XFILL_2__11444_ gnd vdd FILL
XFILL_0__12623_ gnd vdd FILL
XFILL_3__13783_ gnd vdd FILL
XFILL_5__9904_ gnd vdd FILL
XFILL_2_BUFX2_insert870 gnd vdd FILL
XFILL_1__14962_ gnd vdd FILL
XFILL_3__10995_ gnd vdd FILL
XFILL_0__16391_ gnd vdd FILL
XFILL_2_BUFX2_insert881 gnd vdd FILL
XFILL_0__7121_ gnd vdd FILL
XFILL_2_BUFX2_insert892 gnd vdd FILL
X_14818_ _16180_/B _13420_/B _13633_/C _14818_/D gnd _14818_/Y vdd OAI22X1
XFILL_4__12004_ gnd vdd FILL
XFILL_5__14343_ gnd vdd FILL
XFILL_3__15522_ gnd vdd FILL
XFILL_6__13894_ gnd vdd FILL
XFILL_5__11555_ gnd vdd FILL
XFILL_3__12734_ gnd vdd FILL
XFILL_2__14163_ gnd vdd FILL
X_15798_ _15796_/Y _15392_/B _16199_/C _15798_/D gnd _15799_/B vdd OAI22X1
XFILL_4__10196_ gnd vdd FILL
XFILL_1__13913_ gnd vdd FILL
XFILL_0__15342_ gnd vdd FILL
XFILL_2__11375_ gnd vdd FILL
XFILL_1__14893_ gnd vdd FILL
XFILL_0__7052_ gnd vdd FILL
XFILL_5__10506_ gnd vdd FILL
XFILL_6__15633_ gnd vdd FILL
XFILL_2__13114_ gnd vdd FILL
X_14749_ _14748_/Y _14934_/B _14697_/C _14747_/Y gnd _14753_/A vdd OAI22X1
XFILL_5__14274_ gnd vdd FILL
X_7680_ _7744_/B _8832_/B gnd _7680_/Y vdd NAND2X1
XFILL_5__11486_ gnd vdd FILL
XFILL_3__15453_ gnd vdd FILL
XFILL_1__13844_ gnd vdd FILL
XFILL_3__8850_ gnd vdd FILL
XFILL_0__11505_ gnd vdd FILL
XFILL_2__14094_ gnd vdd FILL
XFILL_5__16013_ gnd vdd FILL
XFILL_0__15273_ gnd vdd FILL
XFILL_5__9766_ gnd vdd FILL
XFILL_5__13225_ gnd vdd FILL
XFILL_0__12485_ gnd vdd FILL
XFILL_4_BUFX2_insert2 gnd vdd FILL
XFILL_5__10437_ gnd vdd FILL
XFILL_5__6978_ gnd vdd FILL
XFILL_3__14404_ gnd vdd FILL
XFILL_2__13045_ gnd vdd FILL
XFILL_3__11616_ gnd vdd FILL
XSFILL18680x4050 gnd vdd FILL
XFILL_3__7801_ gnd vdd FILL
XFILL_4__13955_ gnd vdd FILL
XFILL_3__15384_ gnd vdd FILL
XFILL_3__12596_ gnd vdd FILL
XFILL_0__14224_ gnd vdd FILL
XFILL_2__10257_ gnd vdd FILL
XFILL_3__8781_ gnd vdd FILL
XFILL_5__8717_ gnd vdd FILL
XFILL_2__9988_ gnd vdd FILL
XFILL_1__13775_ gnd vdd FILL
XFILL_0__11436_ gnd vdd FILL
XSFILL53960x52050 gnd vdd FILL
XFILL_6__11727_ gnd vdd FILL
X_16419_ _16419_/Q _8152_/CLK _9944_/R vdd _16329_/Y gnd vdd DFFSR
XFILL_5__13156_ gnd vdd FILL
XFILL_4__12906_ gnd vdd FILL
XFILL_6__8490_ gnd vdd FILL
XFILL_6__15495_ gnd vdd FILL
X_9350_ _9339_/B _7558_/B gnd _9351_/C vdd NAND2X1
XFILL_5__10368_ gnd vdd FILL
XFILL_1__15514_ gnd vdd FILL
XFILL_3__14335_ gnd vdd FILL
XFILL_3__11547_ gnd vdd FILL
XFILL_1__12726_ gnd vdd FILL
XFILL_4__13886_ gnd vdd FILL
XFILL_3__7732_ gnd vdd FILL
XSFILL69240x19050 gnd vdd FILL
XFILL_2__10188_ gnd vdd FILL
XFILL_0__14155_ gnd vdd FILL
XBUFX2_insert880 _12216_/Y gnd _12301_/C vdd BUFX2
X_8301_ _8301_/Q _8306_/CLK _7533_/R vdd _8253_/Y gnd vdd DFFSR
XFILL_5__12107_ gnd vdd FILL
XFILL_6__7441_ gnd vdd FILL
XFILL_5__8648_ gnd vdd FILL
XFILL_0__11367_ gnd vdd FILL
XBUFX2_insert891 _12369_/Y gnd _7439_/B vdd BUFX2
XFILL_4__15625_ gnd vdd FILL
XFILL_0__7954_ gnd vdd FILL
XFILL_4__12837_ gnd vdd FILL
XFILL_5__13087_ gnd vdd FILL
X_9281_ _9281_/A gnd _9281_/Y vdd INVX1
XFILL_5__10299_ gnd vdd FILL
XSFILL54040x61050 gnd vdd FILL
XFILL_0__13106_ gnd vdd FILL
XFILL_3__11478_ gnd vdd FILL
XFILL_1__15445_ gnd vdd FILL
XFILL_3__14266_ gnd vdd FILL
XFILL_1__12657_ gnd vdd FILL
XFILL_0__10318_ gnd vdd FILL
XFILL_4_BUFX2_insert409 gnd vdd FILL
XFILL_2__14996_ gnd vdd FILL
XSFILL104440x28050 gnd vdd FILL
XFILL_0__6905_ gnd vdd FILL
XFILL_0__11298_ gnd vdd FILL
XFILL_0__14086_ gnd vdd FILL
XFILL_3__16005_ gnd vdd FILL
XFILL_5__8579_ gnd vdd FILL
X_8232_ _8232_/A _8232_/B _8231_/Y gnd _8232_/Y vdd OAI21X1
XFILL_5__12038_ gnd vdd FILL
XFILL_0__7885_ gnd vdd FILL
XFILL_3__10429_ gnd vdd FILL
XFILL_3__13217_ gnd vdd FILL
XFILL_4__15556_ gnd vdd FILL
XFILL_3__9402_ gnd vdd FILL
XFILL_6__11589_ gnd vdd FILL
XFILL_4__12768_ gnd vdd FILL
XFILL_3__14197_ gnd vdd FILL
XFILL_1__11608_ gnd vdd FILL
XFILL_0__10249_ gnd vdd FILL
XFILL_1__15376_ gnd vdd FILL
XFILL_0__13037_ gnd vdd FILL
XFILL_3__7594_ gnd vdd FILL
XFILL_2__13947_ gnd vdd FILL
XFILL_1__12588_ gnd vdd FILL
XFILL_0__6836_ gnd vdd FILL
XFILL_0__9624_ gnd vdd FILL
XFILL_4__14507_ gnd vdd FILL
XFILL_3__13148_ gnd vdd FILL
XFILL_4__11719_ gnd vdd FILL
X_8163_ _8163_/Q _7791_/CLK _7648_/R vdd _8163_/D gnd vdd DFFSR
XFILL_1__14327_ gnd vdd FILL
XFILL_4__15487_ gnd vdd FILL
XFILL_4__12699_ gnd vdd FILL
XFILL_1__11539_ gnd vdd FILL
XFILL_2__13878_ gnd vdd FILL
X_7114_ _7114_/A gnd _7116_/A vdd INVX1
XFILL_0__9555_ gnd vdd FILL
XFILL111800x3050 gnd vdd FILL
XFILL_4__14438_ gnd vdd FILL
XSFILL18680x80050 gnd vdd FILL
XFILL_3__13079_ gnd vdd FILL
XFILL_2__15617_ gnd vdd FILL
XFILL_5__13989_ gnd vdd FILL
XSFILL48920x41050 gnd vdd FILL
XFILL_3__9264_ gnd vdd FILL
X_8094_ _8082_/A _9246_/B gnd _8095_/C vdd NAND2X1
XFILL_1__14258_ gnd vdd FILL
XFILL_2__12829_ gnd vdd FILL
XFILL_0__8506_ gnd vdd FILL
XFILL_0__14988_ gnd vdd FILL
XFILL_0__9486_ gnd vdd FILL
XFILL_5__15728_ gnd vdd FILL
XSFILL89800x53050 gnd vdd FILL
X_7045_ _7045_/A gnd _7045_/Y vdd INVX1
XFILL_1__13209_ gnd vdd FILL
XFILL_3__8215_ gnd vdd FILL
XFILL_4__14369_ gnd vdd FILL
XFILL_2__15548_ gnd vdd FILL
XFILL_1__14189_ gnd vdd FILL
XFILL_0__13939_ gnd vdd FILL
XFILL_1__7230_ gnd vdd FILL
XSFILL49000x50050 gnd vdd FILL
XFILL_4__16108_ gnd vdd FILL
XSFILL13640x27050 gnd vdd FILL
XFILL_5__15659_ gnd vdd FILL
XFILL_3__8146_ gnd vdd FILL
XFILL_2__15479_ gnd vdd FILL
XSFILL78840x77050 gnd vdd FILL
XSFILL109560x61050 gnd vdd FILL
XFILL_4__16039_ gnd vdd FILL
XFILL_0__8368_ gnd vdd FILL
XFILL_1__7161_ gnd vdd FILL
X_8996_ _8996_/A _8356_/B gnd _8997_/C vdd NAND2X1
XFILL_3__8077_ gnd vdd FILL
XFILL_0__15609_ gnd vdd FILL
XFILL_0__7319_ gnd vdd FILL
XSFILL54120x41050 gnd vdd FILL
XFILL_6__9875_ gnd vdd FILL
X_7947_ _7947_/A gnd _7947_/Y vdd INVX1
XFILL_1__7092_ gnd vdd FILL
XSFILL69720x20050 gnd vdd FILL
XFILL_4__8890_ gnd vdd FILL
XFILL_6__8826_ gnd vdd FILL
X_7878_ _7876_/Y _7878_/B _7878_/C gnd _7878_/Y vdd OAI21X1
XFILL_4__7841_ gnd vdd FILL
X_9617_ _9695_/Q gnd _9617_/Y vdd INVX1
XFILL_3__8979_ gnd vdd FILL
XFILL_1__9802_ gnd vdd FILL
X_9548_ _9546_/Y _9548_/B _9548_/C gnd _9586_/D vdd OAI21X1
XFILL_4__9511_ gnd vdd FILL
XFILL_1__7994_ gnd vdd FILL
XFILL_5_BUFX2_insert232 gnd vdd FILL
X_10430_ _10430_/A gnd _10432_/A vdd INVX1
XFILL_5_BUFX2_insert243 gnd vdd FILL
XFILL_5_BUFX2_insert254 gnd vdd FILL
XFILL_1__6945_ gnd vdd FILL
XFILL_5_BUFX2_insert265 gnd vdd FILL
XFILL_1__9733_ gnd vdd FILL
X_9479_ _9479_/A _9514_/A _9479_/C gnd _9479_/Y vdd OAI21X1
XFILL_5_BUFX2_insert276 gnd vdd FILL
XFILL_5_BUFX2_insert287 gnd vdd FILL
X_10361_ _13528_/A gnd _10363_/A vdd INVX1
XFILL_5_BUFX2_insert298 gnd vdd FILL
XFILL_4_BUFX2_insert910 gnd vdd FILL
XFILL112040x59050 gnd vdd FILL
XFILL_1__9664_ gnd vdd FILL
XFILL_4_BUFX2_insert921 gnd vdd FILL
XFILL_1__6876_ gnd vdd FILL
X_12100_ _12072_/A _11971_/A _12072_/C gnd _12102_/B vdd NAND3X1
XFILL_4_BUFX2_insert932 gnd vdd FILL
XFILL_4__9373_ gnd vdd FILL
XFILL_4_BUFX2_insert943 gnd vdd FILL
XFILL_4_BUFX2_insert954 gnd vdd FILL
X_13080_ _13080_/A _13153_/B gnd _13080_/Y vdd NAND2X1
XFILL_1__8615_ gnd vdd FILL
X_10292_ _10290_/Y _10325_/B _10292_/C gnd _10292_/Y vdd OAI21X1
XFILL_4_BUFX2_insert965 gnd vdd FILL
XSFILL38920x73050 gnd vdd FILL
XFILL_1__9595_ gnd vdd FILL
XFILL112440x80050 gnd vdd FILL
XFILL_4__8324_ gnd vdd FILL
XFILL_4_BUFX2_insert976 gnd vdd FILL
X_12031_ _12031_/A _12031_/B _12031_/C gnd _12034_/A vdd NAND3X1
XFILL_4_BUFX2_insert987 gnd vdd FILL
XFILL_4_BUFX2_insert998 gnd vdd FILL
XFILL_4__8255_ gnd vdd FILL
XSFILL39000x82050 gnd vdd FILL
XFILL_1__8477_ gnd vdd FILL
XFILL_4__7206_ gnd vdd FILL
XFILL_4__8186_ gnd vdd FILL
XFILL_1__7428_ gnd vdd FILL
XFILL_2_BUFX2_insert100 gnd vdd FILL
X_13982_ _15512_/B _14160_/B _14865_/C _15514_/B gnd _13982_/Y vdd OAI22X1
XSFILL18840x40050 gnd vdd FILL
X_15721_ _15410_/D _14228_/Y _15972_/C _14219_/Y gnd _15725_/B vdd OAI22X1
X_12933_ _12865_/A _8161_/CLK _8033_/R vdd _12933_/D gnd vdd DFFSR
XFILL_1__7359_ gnd vdd FILL
XFILL_4__7068_ gnd vdd FILL
XFILL_5__7950_ gnd vdd FILL
X_15652_ _15652_/A _9507_/A _9701_/Q _15652_/D gnd _15660_/A vdd AOI22X1
XFILL_1_BUFX2_insert800 gnd vdd FILL
XFILL_4__10050_ gnd vdd FILL
X_12864_ _12862_/Y vdd _12864_/C gnd _12864_/Y vdd OAI21X1
XFILL_1_BUFX2_insert811 gnd vdd FILL
XFILL_3__10780_ gnd vdd FILL
XFILL_5__6901_ gnd vdd FILL
XFILL_1_BUFX2_insert822 gnd vdd FILL
X_14603_ _14601_/Y _13860_/B _13857_/B _14602_/Y gnd _14604_/A vdd OAI22X1
XFILL_1_BUFX2_insert833 gnd vdd FILL
XFILL_1__9029_ gnd vdd FILL
X_11815_ _11815_/A _11815_/B gnd _11819_/B vdd NOR2X1
XFILL_1_BUFX2_insert844 gnd vdd FILL
XFILL_5__7881_ gnd vdd FILL
XFILL_5__11340_ gnd vdd FILL
XFILL_2__9911_ gnd vdd FILL
X_12795_ _12707_/A _12667_/CLK _12795_/R vdd _12795_/D gnd vdd DFFSR
X_15583_ _15583_/A _15357_/B _16294_/C _14077_/C gnd _15585_/A vdd AOI22X1
XSFILL109720x21050 gnd vdd FILL
XFILL_1__10910_ gnd vdd FILL
XFILL_1_BUFX2_insert855 gnd vdd FILL
XFILL_2__11160_ gnd vdd FILL
XFILL_1_BUFX2_insert866 gnd vdd FILL
XFILL_5__9620_ gnd vdd FILL
XSFILL64040x24050 gnd vdd FILL
XFILL_1_BUFX2_insert877 gnd vdd FILL
XFILL_1__11890_ gnd vdd FILL
X_14534_ _7276_/Q gnd _14535_/A vdd INVX1
XFILL_1_BUFX2_insert888 gnd vdd FILL
X_11746_ _11270_/Y _11732_/B gnd _11746_/Y vdd NAND2X1
XFILL_2__10111_ gnd vdd FILL
XFILL_3__12450_ gnd vdd FILL
XBUFX2_insert110 _10925_/Y gnd _11934_/B vdd BUFX2
XFILL_1_BUFX2_insert899 gnd vdd FILL
XFILL_5__11271_ gnd vdd FILL
XFILL_0__12270_ gnd vdd FILL
XFILL_2__11091_ gnd vdd FILL
XFILL_5__9551_ gnd vdd FILL
XFILL_5__13010_ gnd vdd FILL
XFILL_3__11401_ gnd vdd FILL
X_14465_ _8427_/Q gnd _14465_/Y vdd INVX1
XFILL_4__13740_ gnd vdd FILL
X_11677_ _11063_/Y _11064_/Y _11677_/C gnd _11678_/A vdd OAI21X1
XFILL_4__10952_ gnd vdd FILL
XFILL_3__12381_ gnd vdd FILL
XFILL_2__10042_ gnd vdd FILL
XFILL_5__8502_ gnd vdd FILL
XFILL_2__9773_ gnd vdd FILL
XFILL_1__13560_ gnd vdd FILL
XFILL_2__6985_ gnd vdd FILL
XFILL_0__11221_ gnd vdd FILL
X_16204_ _7885_/A _16204_/B _15390_/B _9843_/Q gnd _16210_/A vdd AOI22X1
XFILL_6__11512_ gnd vdd FILL
XFILL_1__10772_ gnd vdd FILL
XFILL_5__9482_ gnd vdd FILL
X_13416_ _16417_/Q gnd _13416_/Y vdd INVX1
X_10628_ _10626_/Y _10658_/B _10627_/Y gnd _10714_/D vdd OAI21X1
XFILL_6__15280_ gnd vdd FILL
XFILL_5__10153_ gnd vdd FILL
X_14396_ _14721_/A _15845_/B _14718_/B _14394_/Y gnd _14397_/B vdd OAI22X1
XFILL_3__14120_ gnd vdd FILL
XFILL_3__11332_ gnd vdd FILL
XSFILL43320x25050 gnd vdd FILL
XFILL_1__12511_ gnd vdd FILL
XFILL_4__13671_ gnd vdd FILL
XFILL_2__8724_ gnd vdd FILL
XFILL_2__14850_ gnd vdd FILL
XFILL_4__10883_ gnd vdd FILL
XFILL_0__11152_ gnd vdd FILL
XFILL_1__13491_ gnd vdd FILL
X_13347_ _13246_/A _13352_/B _13295_/C gnd _13347_/Y vdd AOI21X1
XFILL_4__15410_ gnd vdd FILL
XSFILL84200x37050 gnd vdd FILL
X_16135_ _8647_/A gnd _16135_/Y vdd INVX1
XFILL_4__12622_ gnd vdd FILL
X_10559_ _10511_/A _7231_/B gnd _10560_/C vdd NAND2X1
XFILL_3__14051_ gnd vdd FILL
XFILL_5__14961_ gnd vdd FILL
XFILL_4__16390_ gnd vdd FILL
XFILL_2__13801_ gnd vdd FILL
XFILL_1__15230_ gnd vdd FILL
XFILL_3__11263_ gnd vdd FILL
XFILL_0__10103_ gnd vdd FILL
XSFILL94360x81050 gnd vdd FILL
XFILL_2__8655_ gnd vdd FILL
XFILL_1__12442_ gnd vdd FILL
XFILL_0__15960_ gnd vdd FILL
XFILL_2__11993_ gnd vdd FILL
XFILL_0__11083_ gnd vdd FILL
XFILL_2__14781_ gnd vdd FILL
XFILL_5__8364_ gnd vdd FILL
XFILL_5__13912_ gnd vdd FILL
XFILL_3__13002_ gnd vdd FILL
X_13278_ _13285_/B _13278_/B gnd _13279_/B vdd NAND2X1
XFILL_4__15341_ gnd vdd FILL
XFILL_0__7670_ gnd vdd FILL
X_16066_ _16066_/A _16066_/B _16065_/Y gnd _16066_/Y vdd NAND3X1
XSFILL59000x13050 gnd vdd FILL
XFILL_6__11374_ gnd vdd FILL
XFILL_2__7606_ gnd vdd FILL
XFILL_5__14892_ gnd vdd FILL
XFILL_2__10944_ gnd vdd FILL
XFILL_2__13732_ gnd vdd FILL
XFILL_0__10034_ gnd vdd FILL
XFILL_1__15161_ gnd vdd FILL
XFILL_3__11194_ gnd vdd FILL
XFILL_0__14911_ gnd vdd FILL
XFILL_2__8586_ gnd vdd FILL
XFILL_1__12373_ gnd vdd FILL
XFILL_5__7315_ gnd vdd FILL
X_15017_ _7158_/A _15177_/B _16014_/C _8278_/Q gnd _15027_/B vdd AOI22X1
X_12229_ _6873_/A _12277_/B _12309_/C _12792_/Q gnd _12230_/C vdd AOI22X1
XFILL_6__10325_ gnd vdd FILL
XFILL_0__15891_ gnd vdd FILL
XFILL_5__13843_ gnd vdd FILL
XFILL_4__11504_ gnd vdd FILL
XFILL_3__10145_ gnd vdd FILL
XFILL_1__14112_ gnd vdd FILL
XFILL_4__15272_ gnd vdd FILL
XFILL_2__16451_ gnd vdd FILL
XFILL_2__13663_ gnd vdd FILL
XFILL_4__12484_ gnd vdd FILL
XFILL_1__11324_ gnd vdd FILL
XFILL112200x19050 gnd vdd FILL
XFILL_0__14842_ gnd vdd FILL
XFILL_2__10875_ gnd vdd FILL
XFILL_1__15092_ gnd vdd FILL
XFILL_5__7246_ gnd vdd FILL
XFILL_0__9340_ gnd vdd FILL
XFILL_4__14223_ gnd vdd FILL
XFILL_4_CLKBUF1_insert1077 gnd vdd FILL
XFILL_5__13774_ gnd vdd FILL
XFILL_2__15402_ gnd vdd FILL
XFILL_2__12614_ gnd vdd FILL
XFILL_4__11435_ gnd vdd FILL
XFILL_1__14043_ gnd vdd FILL
XFILL_2__7468_ gnd vdd FILL
XFILL_3__14953_ gnd vdd FILL
XFILL_2__16382_ gnd vdd FILL
XFILL_2__13594_ gnd vdd FILL
XFILL_1__11255_ gnd vdd FILL
XFILL_5__7177_ gnd vdd FILL
XFILL_5__15513_ gnd vdd FILL
XFILL_0__14773_ gnd vdd FILL
XFILL_5__12725_ gnd vdd FILL
XFILL_3__8000_ gnd vdd FILL
XFILL_0__9271_ gnd vdd FILL
XFILL_0__11985_ gnd vdd FILL
XFILL_4__14154_ gnd vdd FILL
XFILL_2__9207_ gnd vdd FILL
XFILL_3__13904_ gnd vdd FILL
XFILL_2__15333_ gnd vdd FILL
XFILL_4__11366_ gnd vdd FILL
XFILL_0__13724_ gnd vdd FILL
XFILL_3__14884_ gnd vdd FILL
XFILL_0__10936_ gnd vdd FILL
XFILL_0__8222_ gnd vdd FILL
XFILL_1__11186_ gnd vdd FILL
XSFILL89320x70050 gnd vdd FILL
X_15919_ _7275_/Q gnd _15920_/A vdd INVX1
XFILL_4__13105_ gnd vdd FILL
XSFILL53960x47050 gnd vdd FILL
XFILL_5__15444_ gnd vdd FILL
XFILL_5__12656_ gnd vdd FILL
XFILL_4__10317_ gnd vdd FILL
X_8850_ _8854_/B _9362_/B gnd _8850_/Y vdd NAND2X1
XSFILL3560x11050 gnd vdd FILL
XFILL_3__13835_ gnd vdd FILL
XFILL_2__9138_ gnd vdd FILL
XFILL_4__11297_ gnd vdd FILL
XFILL_2__15264_ gnd vdd FILL
XFILL_4__14085_ gnd vdd FILL
XSFILL109480x76050 gnd vdd FILL
XFILL_1__10137_ gnd vdd FILL
XFILL_2__12476_ gnd vdd FILL
XFILL_0__13655_ gnd vdd FILL
XFILL_1__15994_ gnd vdd FILL
XFILL_5__11607_ gnd vdd FILL
X_7801_ _7895_/Q gnd _7803_/A vdd INVX1
XFILL_4__10248_ gnd vdd FILL
XFILL_5__15375_ gnd vdd FILL
XFILL_2__14215_ gnd vdd FILL
XFILL_4__13036_ gnd vdd FILL
XSFILL28760x23050 gnd vdd FILL
XFILL_5__12587_ gnd vdd FILL
X_8781_ _8819_/Q gnd _8783_/A vdd INVX1
XFILL_2__11427_ gnd vdd FILL
XFILL_2__15195_ gnd vdd FILL
XFILL_0__12606_ gnd vdd FILL
XFILL_3__13766_ gnd vdd FILL
XSFILL54040x56050 gnd vdd FILL
XFILL_0__7104_ gnd vdd FILL
XFILL_3__10978_ gnd vdd FILL
XFILL_1__10068_ gnd vdd FILL
XFILL_1__14945_ gnd vdd FILL
XFILL_0__16374_ gnd vdd FILL
XFILL_0__13586_ gnd vdd FILL
XFILL_5__14326_ gnd vdd FILL
XFILL_3__15505_ gnd vdd FILL
X_7732_ _7730_/Y _7684_/B _7732_/C gnd _7786_/D vdd OAI21X1
XFILL_0__10798_ gnd vdd FILL
XFILL_5__11538_ gnd vdd FILL
XFILL_0__8084_ gnd vdd FILL
XFILL_3__12717_ gnd vdd FILL
XFILL_2__14146_ gnd vdd FILL
XFILL_3__8902_ gnd vdd FILL
XFILL_4__10179_ gnd vdd FILL
XFILL_0__15325_ gnd vdd FILL
XFILL_2__11358_ gnd vdd FILL
XFILL_1__14876_ gnd vdd FILL
XFILL_3__9882_ gnd vdd FILL
XFILL_3__13697_ gnd vdd FILL
XFILL_0__7035_ gnd vdd FILL
XFILL_5__14257_ gnd vdd FILL
XFILL_6__9591_ gnd vdd FILL
XFILL_2__10309_ gnd vdd FILL
X_7663_ _7663_/Q _7791_/CLK _7648_/R vdd _7663_/D gnd vdd DFFSR
XFILL_3__15436_ gnd vdd FILL
XFILL_5__11469_ gnd vdd FILL
XFILL_3__8833_ gnd vdd FILL
XFILL_3__12648_ gnd vdd FILL
XFILL_1__13827_ gnd vdd FILL
XFILL_4__14987_ gnd vdd FILL
XFILL_2__14077_ gnd vdd FILL
XFILL_0__15256_ gnd vdd FILL
XFILL_5_BUFX2_insert60 gnd vdd FILL
XFILL_2__11289_ gnd vdd FILL
XFILL_5__13208_ gnd vdd FILL
XFILL_0__12468_ gnd vdd FILL
X_9402_ _9400_/Y _9401_/A _9402_/C gnd _9452_/D vdd OAI21X1
XFILL_5_BUFX2_insert71 gnd vdd FILL
XFILL_5__9749_ gnd vdd FILL
XFILL_5__14188_ gnd vdd FILL
XFILL_5_BUFX2_insert82 gnd vdd FILL
XFILL_4__13938_ gnd vdd FILL
XFILL_2__13028_ gnd vdd FILL
XSFILL18680x75050 gnd vdd FILL
XFILL_3__15367_ gnd vdd FILL
XFILL_0__14207_ gnd vdd FILL
XFILL_5_BUFX2_insert93 gnd vdd FILL
XSFILL48920x36050 gnd vdd FILL
X_7594_ _7598_/B _7594_/B gnd _7594_/Y vdd NAND2X1
XFILL_3__12579_ gnd vdd FILL
XFILL_3__8764_ gnd vdd FILL
XFILL_1__13758_ gnd vdd FILL
XSFILL104440x7050 gnd vdd FILL
XFILL_0__11419_ gnd vdd FILL
XSFILL74200x69050 gnd vdd FILL
XFILL_0__15187_ gnd vdd FILL
XFILL_0__12399_ gnd vdd FILL
XFILL_5__13139_ gnd vdd FILL
X_9333_ _9333_/Q _7537_/CLK _7537_/R vdd _9333_/D gnd vdd DFFSR
XFILL_3__14318_ gnd vdd FILL
XFILL_4__13869_ gnd vdd FILL
XFILL_3__7715_ gnd vdd FILL
XFILL_1__12709_ gnd vdd FILL
XFILL_0__8986_ gnd vdd FILL
XFILL_3__15298_ gnd vdd FILL
XFILL_0__14138_ gnd vdd FILL
XFILL_3__8695_ gnd vdd FILL
XFILL_1__13689_ gnd vdd FILL
XSFILL49800x64050 gnd vdd FILL
XFILL_4__15608_ gnd vdd FILL
XFILL_0__7937_ gnd vdd FILL
X_9264_ _9240_/A _6960_/B gnd _9265_/C vdd NAND2X1
XFILL_4_BUFX2_insert228 gnd vdd FILL
XFILL_3__14249_ gnd vdd FILL
XFILL_1__15428_ gnd vdd FILL
XSFILL89400x50050 gnd vdd FILL
XFILL_2__14979_ gnd vdd FILL
XFILL_4_BUFX2_insert239 gnd vdd FILL
XFILL_0__14069_ gnd vdd FILL
X_8215_ _8215_/A gnd _8217_/A vdd INVX1
XSFILL109560x56050 gnd vdd FILL
XFILL_4__15539_ gnd vdd FILL
X_9195_ _9195_/Q _9195_/CLK _8051_/R vdd _9143_/Y gnd vdd DFFSR
XFILL_0__7868_ gnd vdd FILL
XFILL_1__15359_ gnd vdd FILL
XFILL_3__7577_ gnd vdd FILL
XFILL_3_BUFX2_insert906 gnd vdd FILL
XFILL_0__9607_ gnd vdd FILL
XFILL_1__8400_ gnd vdd FILL
XFILL_1__9380_ gnd vdd FILL
XFILL_6__7286_ gnd vdd FILL
XSFILL54120x36050 gnd vdd FILL
X_8146_ _8146_/A _8133_/A _8146_/C gnd _8180_/D vdd OAI21X1
XFILL_0__7799_ gnd vdd FILL
XFILL_3_BUFX2_insert917 gnd vdd FILL
XSFILL39480x54050 gnd vdd FILL
XFILL_3_BUFX2_insert928 gnd vdd FILL
XFILL_3_BUFX2_insert939 gnd vdd FILL
XFILL_1__8331_ gnd vdd FILL
XFILL_0__9538_ gnd vdd FILL
X_8077_ _8077_/A _8118_/A _8077_/C gnd _8157_/D vdd OAI21X1
XFILL_3__9247_ gnd vdd FILL
XSFILL43960x79050 gnd vdd FILL
XFILL_1__8262_ gnd vdd FILL
X_7028_ _6992_/A _8297_/CLK _7796_/R vdd _7028_/D gnd vdd DFFSR
XFILL_0__9469_ gnd vdd FILL
XFILL_1__7213_ gnd vdd FILL
XSFILL18760x55050 gnd vdd FILL
XFILL_1__8193_ gnd vdd FILL
XFILL_3__8129_ gnd vdd FILL
XFILL_4__9991_ gnd vdd FILL
XFILL_6__9927_ gnd vdd FILL
XFILL_1_BUFX2_insert107 gnd vdd FILL
X_8979_ _8979_/A _9011_/A _8979_/C gnd _9055_/D vdd OAI21X1
XSFILL43960x7050 gnd vdd FILL
XFILL_1__7075_ gnd vdd FILL
XSFILL33800x50 gnd vdd FILL
X_11600_ _11600_/A _11600_/B _11599_/Y gnd _12065_/A vdd NAND3X1
XFILL_0_CLKBUF1_insert200 gnd vdd FILL
XFILL_0_CLKBUF1_insert211 gnd vdd FILL
XFILL_4__8873_ gnd vdd FILL
X_12580_ vdd memoryOutData[4] gnd _12580_/Y vdd NAND2X1
XFILL_0_CLKBUF1_insert222 gnd vdd FILL
XSFILL38920x68050 gnd vdd FILL
XFILL_0_BUFX2_insert807 gnd vdd FILL
XFILL_4__7824_ gnd vdd FILL
XFILL112440x75050 gnd vdd FILL
XFILL_0_BUFX2_insert818 gnd vdd FILL
XFILL_0_BUFX2_insert829 gnd vdd FILL
X_11531_ _11531_/A _11846_/C _11530_/Y gnd _11531_/Y vdd AOI21X1
XFILL_1_BUFX2_insert1004 gnd vdd FILL
XFILL_1_BUFX2_insert1015 gnd vdd FILL
XFILL_1_BUFX2_insert1026 gnd vdd FILL
XFILL_1_BUFX2_insert1037 gnd vdd FILL
XFILL_4__7755_ gnd vdd FILL
X_14250_ _14250_/A _14250_/B gnd _14250_/Y vdd NOR2X1
XFILL_1_BUFX2_insert1048 gnd vdd FILL
X_11462_ _11184_/A gnd _11463_/C vdd INVX1
XFILL_1_BUFX2_insert1059 gnd vdd FILL
XSFILL89320x6050 gnd vdd FILL
X_13201_ _13157_/A _13201_/CLK _13201_/R vdd _13201_/D gnd vdd DFFSR
XFILL_1__7977_ gnd vdd FILL
X_10413_ _10395_/A _7853_/B gnd _10413_/Y vdd NAND2X1
X_14181_ _9317_/Q _13854_/B _13853_/B _8805_/Q gnd _14182_/B vdd AOI22X1
XFILL_4__7686_ gnd vdd FILL
X_11393_ _11393_/A gnd _11395_/A vdd INVX1
XFILL_1__6928_ gnd vdd FILL
XFILL_4__9425_ gnd vdd FILL
X_13132_ _13130_/Y _13173_/A _13132_/C gnd _13132_/Y vdd OAI21X1
XSFILL18840x35050 gnd vdd FILL
X_10344_ _10284_/A _7400_/CLK _9704_/R vdd _10344_/D gnd vdd DFFSR
XSFILL84280x11050 gnd vdd FILL
XFILL_4_BUFX2_insert740 gnd vdd FILL
XFILL_4_BUFX2_insert751 gnd vdd FILL
XFILL_2__8440_ gnd vdd FILL
XFILL_1__9647_ gnd vdd FILL
XFILL_1__6859_ gnd vdd FILL
XFILL_4_BUFX2_insert762 gnd vdd FILL
XFILL_4_BUFX2_insert773 gnd vdd FILL
XFILL_4__9356_ gnd vdd FILL
XFILL_3_CLKBUF1_insert1083 gnd vdd FILL
X_13063_ _6886_/A _8176_/CLK _8816_/R vdd _13063_/D gnd vdd DFFSR
X_10275_ _10341_/Q gnd _10277_/A vdd INVX1
XSFILL99320x33050 gnd vdd FILL
XFILL_4_BUFX2_insert784 gnd vdd FILL
XFILL_4_BUFX2_insert795 gnd vdd FILL
XFILL_2__8371_ gnd vdd FILL
XFILL_5__7100_ gnd vdd FILL
XFILL_5__8080_ gnd vdd FILL
X_12014_ _12014_/A _12012_/Y _12014_/C gnd _13098_/B vdd NAND3X1
XFILL_4__9287_ gnd vdd FILL
XFILL_2__7322_ gnd vdd FILL
XFILL_1__8529_ gnd vdd FILL
XFILL_2__10660_ gnd vdd FILL
XFILL_5__7031_ gnd vdd FILL
XFILL_4__8238_ gnd vdd FILL
XSFILL64040x19050 gnd vdd FILL
XFILL_6__10041_ gnd vdd FILL
XFILL_4__11220_ gnd vdd FILL
XFILL_5__10771_ gnd vdd FILL
XFILL_2__7253_ gnd vdd FILL
XFILL_3__11950_ gnd vdd FILL
XFILL_1__11040_ gnd vdd FILL
XFILL_5__12510_ gnd vdd FILL
XFILL_0__11770_ gnd vdd FILL
XFILL_4__11151_ gnd vdd FILL
XFILL_3__10901_ gnd vdd FILL
XFILL_5__13490_ gnd vdd FILL
XFILL_2__12330_ gnd vdd FILL
X_13965_ _8980_/A gnd _15458_/A vdd INVX1
XFILL_2__7184_ gnd vdd FILL
XFILL_3__11881_ gnd vdd FILL
X_15704_ _15916_/B _15704_/B _10534_/A _15356_/C gnd _15705_/B vdd AOI22X1
XFILL_4__10102_ gnd vdd FILL
XSFILL3480x26050 gnd vdd FILL
XFILL_5__12441_ gnd vdd FILL
X_12916_ _12950_/Q gnd _12916_/Y vdd INVX1
XFILL_5__8982_ gnd vdd FILL
XFILL_3__13620_ gnd vdd FILL
XFILL_4__11082_ gnd vdd FILL
XFILL_2__12261_ gnd vdd FILL
X_13896_ _7185_/A _14762_/B _14413_/A _8209_/A gnd _13897_/B vdd AOI22X1
XFILL_3__10832_ gnd vdd FILL
XFILL_0__13440_ gnd vdd FILL
XFILL_0__10652_ gnd vdd FILL
XFILL_5__7933_ gnd vdd FILL
XFILL_1__12991_ gnd vdd FILL
X_15635_ _9248_/A gnd _15637_/A vdd INVX1
XFILL_2__14000_ gnd vdd FILL
XFILL_4__10033_ gnd vdd FILL
XFILL_5__15160_ gnd vdd FILL
XFILL_4__14910_ gnd vdd FILL
XFILL_1_BUFX2_insert630 gnd vdd FILL
X_12847_ _12847_/A gnd _12847_/Y vdd INVX1
XFILL_5__12372_ gnd vdd FILL
XFILL_2__11212_ gnd vdd FILL
XFILL_3__10763_ gnd vdd FILL
XFILL_1__14730_ gnd vdd FILL
XFILL_3__13551_ gnd vdd FILL
XFILL_4__15890_ gnd vdd FILL
XFILL_1_BUFX2_insert641 gnd vdd FILL
XSFILL94360x76050 gnd vdd FILL
XFILL_1_BUFX2_insert652 gnd vdd FILL
XFILL_1__11942_ gnd vdd FILL
XFILL_2__12192_ gnd vdd FILL
XFILL_0__13371_ gnd vdd FILL
XFILL_1_BUFX2_insert663 gnd vdd FILL
XFILL_5__14111_ gnd vdd FILL
XFILL_5__7864_ gnd vdd FILL
XFILL_5__11323_ gnd vdd FILL
XFILL_4__14841_ gnd vdd FILL
XFILL_3__12502_ gnd vdd FILL
X_15566_ _15566_/A gnd _15568_/A vdd INVX1
XFILL_1_BUFX2_insert674 gnd vdd FILL
XFILL_6__10874_ gnd vdd FILL
XFILL_5__15091_ gnd vdd FILL
X_12778_ _12776_/Y _12777_/A _12778_/C gnd _12818_/D vdd OAI21X1
XFILL_1_BUFX2_insert685 gnd vdd FILL
XFILL_2__11143_ gnd vdd FILL
XFILL_0__15110_ gnd vdd FILL
XFILL_3__16270_ gnd vdd FILL
XFILL_5__9603_ gnd vdd FILL
XFILL_1_BUFX2_insert696 gnd vdd FILL
XFILL_3__10694_ gnd vdd FILL
XFILL_0__12322_ gnd vdd FILL
XFILL_1__14661_ gnd vdd FILL
XFILL_3__13482_ gnd vdd FILL
XFILL_1__11873_ gnd vdd FILL
XSFILL69160x52050 gnd vdd FILL
XFILL_0__16090_ gnd vdd FILL
XSFILL99400x13050 gnd vdd FILL
X_14517_ _7480_/A gnd _14518_/D vdd INVX1
XFILL_5__14042_ gnd vdd FILL
XFILL_3__15221_ gnd vdd FILL
X_11729_ _11078_/Y _11270_/B _11728_/Y gnd _11729_/Y vdd OAI21X1
XFILL_5__11254_ gnd vdd FILL
XFILL_1__13612_ gnd vdd FILL
XFILL_1__16400_ gnd vdd FILL
XFILL_3__12433_ gnd vdd FILL
X_15497_ _15496_/Y _15473_/Y _14791_/C gnd _12854_/B vdd AOI21X1
XFILL_4__14772_ gnd vdd FILL
XFILL_4__11984_ gnd vdd FILL
XFILL_0__15041_ gnd vdd FILL
XFILL_2__15951_ gnd vdd FILL
XFILL_2__11074_ gnd vdd FILL
XFILL_1__10824_ gnd vdd FILL
XFILL_1__14592_ gnd vdd FILL
XFILL_5__9534_ gnd vdd FILL
XFILL_0__12253_ gnd vdd FILL
XFILL_6__15332_ gnd vdd FILL
XFILL_0__8840_ gnd vdd FILL
XSFILL73640x77050 gnd vdd FILL
XSFILL104360x61050 gnd vdd FILL
XFILL_4__13723_ gnd vdd FILL
X_14448_ _14448_/A _14447_/Y _14445_/Y gnd _14448_/Y vdd NAND3X1
XFILL_4__10935_ gnd vdd FILL
XFILL_3__12364_ gnd vdd FILL
XFILL_1__16331_ gnd vdd FILL
XFILL_5__11185_ gnd vdd FILL
XFILL_3__15152_ gnd vdd FILL
XFILL_2__14902_ gnd vdd FILL
XFILL_2__10025_ gnd vdd FILL
XFILL_2__9756_ gnd vdd FILL
XFILL_0__11204_ gnd vdd FILL
XFILL_1__13543_ gnd vdd FILL
XFILL_1__10755_ gnd vdd FILL
XFILL_2__6968_ gnd vdd FILL
XFILL_2__15882_ gnd vdd FILL
XFILL_0__12184_ gnd vdd FILL
XFILL_5__9465_ gnd vdd FILL
XFILL_5__10136_ gnd vdd FILL
XFILL_3__14103_ gnd vdd FILL
XFILL_3__11315_ gnd vdd FILL
XFILL_0__8771_ gnd vdd FILL
XFILL_3__7500_ gnd vdd FILL
XFILL_2__8707_ gnd vdd FILL
XFILL_4__13654_ gnd vdd FILL
X_14379_ _14379_/A _14379_/B _14374_/Y gnd _14380_/B vdd NAND3X1
XFILL_5__15993_ gnd vdd FILL
XFILL_2__14833_ gnd vdd FILL
XFILL_3__15083_ gnd vdd FILL
XFILL_3__12295_ gnd vdd FILL
XFILL_1__16262_ gnd vdd FILL
XFILL_3__8480_ gnd vdd FILL
XFILL_1__13474_ gnd vdd FILL
XFILL_0__11135_ gnd vdd FILL
XFILL_1__10686_ gnd vdd FILL
X_16118_ _8688_/Q gnd _16118_/Y vdd INVX1
XFILL_2__6899_ gnd vdd FILL
XFILL_4__12605_ gnd vdd FILL
XFILL_5__9396_ gnd vdd FILL
XFILL_0__7722_ gnd vdd FILL
XFILL_1__15213_ gnd vdd FILL
XFILL_3__14034_ gnd vdd FILL
XFILL_5__10067_ gnd vdd FILL
XFILL_5__14944_ gnd vdd FILL
XFILL_3__11246_ gnd vdd FILL
XFILL_4__16373_ gnd vdd FILL
XFILL_2__8638_ gnd vdd FILL
XFILL_4__13585_ gnd vdd FILL
XFILL_1__12425_ gnd vdd FILL
XFILL_3__7431_ gnd vdd FILL
XFILL_2__11976_ gnd vdd FILL
XFILL_1__16193_ gnd vdd FILL
XFILL_0__15943_ gnd vdd FILL
XFILL_4__10797_ gnd vdd FILL
XFILL_0__11066_ gnd vdd FILL
XFILL_2__14764_ gnd vdd FILL
X_8000_ _7998_/Y _7937_/B _8000_/C gnd _8046_/D vdd OAI21X1
XFILL_6__14145_ gnd vdd FILL
XFILL_5__8347_ gnd vdd FILL
XFILL_4__15324_ gnd vdd FILL
X_16049_ _9455_/Q gnd _16049_/Y vdd INVX1
XFILL_5__14875_ gnd vdd FILL
XSFILL28760x18050 gnd vdd FILL
XFILL_2__10927_ gnd vdd FILL
XFILL_2__13715_ gnd vdd FILL
XFILL_3__7362_ gnd vdd FILL
XFILL_1__15144_ gnd vdd FILL
XFILL_3__11177_ gnd vdd FILL
XFILL_1__12356_ gnd vdd FILL
XFILL_0__10017_ gnd vdd FILL
XFILL_2__8569_ gnd vdd FILL
XFILL_2__14695_ gnd vdd FILL
XFILL_0__15874_ gnd vdd FILL
XFILL_3__9101_ gnd vdd FILL
XFILL_3__10128_ gnd vdd FILL
XFILL_5__13826_ gnd vdd FILL
XFILL_4__15255_ gnd vdd FILL
XSFILL94440x56050 gnd vdd FILL
XFILL_0__7584_ gnd vdd FILL
XSFILL43800x21050 gnd vdd FILL
XFILL_4__12467_ gnd vdd FILL
XFILL_1__11307_ gnd vdd FILL
XFILL_3__15985_ gnd vdd FILL
XFILL_2__13646_ gnd vdd FILL
XFILL_0__14825_ gnd vdd FILL
XFILL_1__15075_ gnd vdd FILL
XFILL_3__7293_ gnd vdd FILL
XSFILL28360x20050 gnd vdd FILL
XFILL_5__7229_ gnd vdd FILL
XFILL_1__12287_ gnd vdd FILL
XFILL_6__13027_ gnd vdd FILL
XFILL_4__14206_ gnd vdd FILL
XFILL_5__13757_ gnd vdd FILL
X_9951_ _9951_/Q _7274_/CLK _7274_/R vdd _9951_/D gnd vdd DFFSR
XFILL_4__11418_ gnd vdd FILL
XFILL_5__10969_ gnd vdd FILL
XFILL_4__15186_ gnd vdd FILL
XFILL_3__10059_ gnd vdd FILL
XFILL_1__14026_ gnd vdd FILL
XFILL_3__14936_ gnd vdd FILL
XSFILL69240x32050 gnd vdd FILL
XSFILL53960x2050 gnd vdd FILL
XFILL_3__9032_ gnd vdd FILL
XFILL_4__12398_ gnd vdd FILL
XFILL_2__16365_ gnd vdd FILL
XFILL_2__13577_ gnd vdd FILL
XFILL_1__11238_ gnd vdd FILL
XFILL_2__10789_ gnd vdd FILL
XFILL_0__14756_ gnd vdd FILL
XFILL_5__12708_ gnd vdd FILL
XFILL_0__9254_ gnd vdd FILL
XFILL_0__11968_ gnd vdd FILL
X_8902_ _8902_/A _8902_/B _8901_/Y gnd _8902_/Y vdd OAI21X1
XFILL_4__14137_ gnd vdd FILL
XFILL_2__15316_ gnd vdd FILL
X_9882_ _9954_/Q gnd _9884_/A vdd INVX1
XFILL_5__13688_ gnd vdd FILL
XFILL_4__11349_ gnd vdd FILL
XFILL_3__14867_ gnd vdd FILL
XFILL_2__12528_ gnd vdd FILL
XFILL_0__13707_ gnd vdd FILL
XFILL_0__10919_ gnd vdd FILL
XFILL_0__8205_ gnd vdd FILL
XSFILL104440x41050 gnd vdd FILL
XFILL_2__16296_ gnd vdd FILL
XFILL_1__11169_ gnd vdd FILL
XFILL_0__14687_ gnd vdd FILL
X_8833_ _8833_/A _8896_/B _8832_/Y gnd _8833_/Y vdd OAI21X1
XFILL_5__12639_ gnd vdd FILL
XFILL_6__7973_ gnd vdd FILL
XFILL_0__11899_ gnd vdd FILL
XFILL_5__15427_ gnd vdd FILL
XFILL_3__13818_ gnd vdd FILL
XFILL_4__14068_ gnd vdd FILL
XFILL_2__15247_ gnd vdd FILL
XFILL_2__12459_ gnd vdd FILL
XFILL_0__13638_ gnd vdd FILL
XFILL_3__14798_ gnd vdd FILL
XFILL_1__15977_ gnd vdd FILL
XFILL_6__6924_ gnd vdd FILL
XFILL_0__8136_ gnd vdd FILL
XFILL_5__15358_ gnd vdd FILL
XFILL_4__13019_ gnd vdd FILL
XFILL_6_BUFX2_insert802 gnd vdd FILL
X_8764_ _8765_/B _8764_/B gnd _8764_/Y vdd NAND2X1
XFILL_3__9934_ gnd vdd FILL
XFILL_2__15178_ gnd vdd FILL
XFILL_3__13749_ gnd vdd FILL
XSFILL89400x45050 gnd vdd FILL
XFILL_0__16357_ gnd vdd FILL
XFILL_1__14928_ gnd vdd FILL
XFILL_0__13569_ gnd vdd FILL
XFILL_5__14309_ gnd vdd FILL
XFILL_6__9643_ gnd vdd FILL
X_7715_ _7781_/Q gnd _7715_/Y vdd INVX1
XFILL_0__8067_ gnd vdd FILL
XSFILL99320x1050 gnd vdd FILL
XFILL_5__15289_ gnd vdd FILL
XFILL_0__15308_ gnd vdd FILL
XFILL_2__14129_ gnd vdd FILL
XFILL_6_BUFX2_insert868 gnd vdd FILL
X_8695_ _6903_/A _8695_/B gnd _8696_/C vdd NAND2X1
XFILL_3__9865_ gnd vdd FILL
XFILL_6_BUFX2_insert879 gnd vdd FILL
XFILL_1__14859_ gnd vdd FILL
XFILL_0__16288_ gnd vdd FILL
X_7646_ _7646_/Q _7902_/CLK _7150_/R vdd _7568_/Y gnd vdd DFFSR
XFILL_3__15419_ gnd vdd FILL
XFILL_1__8880_ gnd vdd FILL
XFILL_0__15239_ gnd vdd FILL
XFILL_3__16399_ gnd vdd FILL
XSFILL13640x40050 gnd vdd FILL
XFILL_3__9796_ gnd vdd FILL
XFILL_1__7831_ gnd vdd FILL
X_7577_ _7577_/A _7577_/B _7576_/Y gnd _7577_/Y vdd OAI21X1
XFILL_3__8747_ gnd vdd FILL
XSFILL13720x5050 gnd vdd FILL
XSFILL99800x7050 gnd vdd FILL
X_9316_ _9248_/A _9306_/CLK _9306_/R vdd _9316_/D gnd vdd DFFSR
XSFILL69320x12050 gnd vdd FILL
XFILL_0__8969_ gnd vdd FILL
XFILL_1__7762_ gnd vdd FILL
XFILL_4__7471_ gnd vdd FILL
XFILL_1__9501_ gnd vdd FILL
X_9247_ _9247_/A _9282_/A _9246_/Y gnd _9315_/D vdd OAI21X1
XFILL_1__7693_ gnd vdd FILL
XFILL_4__9210_ gnd vdd FILL
XSFILL104520x21050 gnd vdd FILL
XFILL_3__7629_ gnd vdd FILL
X_9178_ _9090_/A _9195_/CLK _9963_/R vdd _9178_/D gnd vdd DFFSR
XFILL_3_BUFX2_insert703 gnd vdd FILL
XFILL_4__9141_ gnd vdd FILL
XFILL_3_BUFX2_insert714 gnd vdd FILL
XFILL_3_BUFX2_insert725 gnd vdd FILL
X_10060_ _10058_/Y _9985_/B _10059_/Y gnd _10098_/D vdd OAI21X1
XFILL_3_BUFX2_insert736 gnd vdd FILL
X_8129_ _8129_/A gnd _8131_/A vdd INVX1
XFILL_3_BUFX2_insert747 gnd vdd FILL
XFILL_1__9363_ gnd vdd FILL
XFILL_3_BUFX2_insert758 gnd vdd FILL
XFILL_3_BUFX2_insert769 gnd vdd FILL
XFILL_1__8314_ gnd vdd FILL
XFILL_1__9294_ gnd vdd FILL
XFILL111960x63050 gnd vdd FILL
XFILL_1_BUFX2_insert80 gnd vdd FILL
XFILL_1__8245_ gnd vdd FILL
XFILL_1_BUFX2_insert91 gnd vdd FILL
XSFILL94600x16050 gnd vdd FILL
XSFILL13720x20050 gnd vdd FILL
X_10962_ _10936_/B _10962_/B gnd _10964_/C vdd NAND2X1
X_13750_ _13741_/Y _13750_/B _13750_/C gnd _13761_/A vdd NAND3X1
XSFILL24360x71050 gnd vdd FILL
XSFILL39160x31050 gnd vdd FILL
X_12701_ _12701_/A gnd _12703_/A vdd INVX1
XFILL_4__9974_ gnd vdd FILL
X_13681_ _13680_/Y _13681_/B gnd _13684_/C vdd NOR2X1
X_10893_ _12701_/A gnd _10894_/B vdd INVX1
X_15420_ _15419_/Y _15848_/A gnd _15421_/C vdd NOR2X1
X_12632_ _12632_/A vdd _12632_/C gnd _12684_/D vdd OAI21X1
XFILL_1__7058_ gnd vdd FILL
XFILL_2__7940_ gnd vdd FILL
XFILL_0_BUFX2_insert604 gnd vdd FILL
XFILL_4__8856_ gnd vdd FILL
XFILL_0_BUFX2_insert615 gnd vdd FILL
X_15351_ _15351_/A _13828_/Y _13813_/D _15351_/D gnd _15351_/Y vdd OAI22X1
X_12563_ _12427_/A _13175_/CLK _13199_/R vdd _12525_/Y gnd vdd DFFSR
XFILL_0_BUFX2_insert626 gnd vdd FILL
XSFILL99320x28050 gnd vdd FILL
XFILL_0_BUFX2_insert637 gnd vdd FILL
XFILL_2__7871_ gnd vdd FILL
XFILL_4__7807_ gnd vdd FILL
XFILL_0_BUFX2_insert648 gnd vdd FILL
XFILL_0_BUFX2_insert659 gnd vdd FILL
X_11514_ _11514_/A _11512_/Y _11514_/C gnd _11514_/Y vdd OAI21X1
X_14302_ _9063_/Q gnd _14302_/Y vdd INVX1
XFILL_5__7580_ gnd vdd FILL
XFILL_4__8787_ gnd vdd FILL
XFILL_2__9610_ gnd vdd FILL
X_12494_ vdd _12494_/B gnd _12494_/Y vdd NAND2X1
X_15282_ _13728_/Y _15795_/B _15282_/C gnd _15284_/A vdd OAI21X1
XFILL_4__7738_ gnd vdd FILL
X_14233_ _14555_/C _14232_/Y _14203_/C _14231_/Y gnd _14233_/Y vdd OAI22X1
X_11445_ _11034_/B _11444_/Y gnd _11445_/Y vdd NOR2X1
XFILL_2__9541_ gnd vdd FILL
XFILL_1__10540_ gnd vdd FILL
XFILL_5__9250_ gnd vdd FILL
X_14164_ _13467_/A _14164_/B _14865_/C _14164_/D gnd _14164_/Y vdd OAI22X1
XFILL_3__11100_ gnd vdd FILL
X_11376_ _11376_/A _11376_/B _11235_/Y _11236_/Y gnd _11376_/Y vdd OAI22X1
XFILL_3__12080_ gnd vdd FILL
XFILL_2__11830_ gnd vdd FILL
XFILL_4__10651_ gnd vdd FILL
XFILL_5__12990_ gnd vdd FILL
XFILL_2__9472_ gnd vdd FILL
XFILL_4__9408_ gnd vdd FILL
XFILL_5__8201_ gnd vdd FILL
XFILL112120x52050 gnd vdd FILL
XFILL_6__11211_ gnd vdd FILL
X_13115_ _12151_/A gnd _13117_/A vdd INVX1
X_10327_ _13497_/A _7515_/CLK _7665_/R vdd _10327_/D gnd vdd DFFSR
XFILL_4_BUFX2_insert570 gnd vdd FILL
XFILL_5__11941_ gnd vdd FILL
X_14095_ _14095_/A _14095_/B _14092_/Y gnd _14095_/Y vdd NAND3X1
XFILL_3__11031_ gnd vdd FILL
XFILL_4_BUFX2_insert581 gnd vdd FILL
XFILL_4__13370_ gnd vdd FILL
XFILL_1__12210_ gnd vdd FILL
XFILL_4_BUFX2_insert592 gnd vdd FILL
XFILL_2__11761_ gnd vdd FILL
XFILL_5__8132_ gnd vdd FILL
XFILL_4__9339_ gnd vdd FILL
X_13046_ _13044_/Y vdd _13045_/Y gnd _13078_/D vdd OAI21X1
XFILL_4__12321_ gnd vdd FILL
X_10258_ _10264_/A _7186_/B gnd _10258_/Y vdd NAND2X1
XFILL_5__14660_ gnd vdd FILL
XFILL_5__11872_ gnd vdd FILL
XFILL_2__13500_ gnd vdd FILL
XFILL_2__14480_ gnd vdd FILL
XFILL_2__8354_ gnd vdd FILL
XFILL_1__12141_ gnd vdd FILL
XFILL_2__11692_ gnd vdd FILL
XFILL_5__8063_ gnd vdd FILL
XFILL_5__13611_ gnd vdd FILL
XFILL_0__12871_ gnd vdd FILL
XFILL_4__15040_ gnd vdd FILL
XFILL_5__10823_ gnd vdd FILL
X_10189_ _10189_/A gnd _10189_/Y vdd INVX1
XFILL_5__14591_ gnd vdd FILL
XFILL_2__7305_ gnd vdd FILL
XFILL_2__13431_ gnd vdd FILL
XFILL_4__12252_ gnd vdd FILL
XFILL_0__14610_ gnd vdd FILL
XFILL_3__15770_ gnd vdd FILL
XFILL_2__10643_ gnd vdd FILL
XFILL_1__12072_ gnd vdd FILL
XFILL_3__12982_ gnd vdd FILL
XFILL_0__11822_ gnd vdd FILL
XFILL_5__16330_ gnd vdd FILL
XSFILL69160x47050 gnd vdd FILL
XFILL_0__15590_ gnd vdd FILL
XFILL_5__13542_ gnd vdd FILL
XFILL_4__11203_ gnd vdd FILL
XFILL_2__7236_ gnd vdd FILL
XFILL_5__10754_ gnd vdd FILL
XFILL_3__14721_ gnd vdd FILL
XFILL_2__13362_ gnd vdd FILL
XFILL_1__15900_ gnd vdd FILL
X_14997_ _12767_/A _12764_/A gnd _16037_/B vdd NOR2X1
XFILL_3__11933_ gnd vdd FILL
XFILL_4__12183_ gnd vdd FILL
XFILL_1__11023_ gnd vdd FILL
XFILL_2__16150_ gnd vdd FILL
XFILL_2__10574_ gnd vdd FILL
XFILL_0__14541_ gnd vdd FILL
XFILL_0__11753_ gnd vdd FILL
XFILL_5__16261_ gnd vdd FILL
XFILL_5__13473_ gnd vdd FILL
XFILL_2__12313_ gnd vdd FILL
XFILL_4__11134_ gnd vdd FILL
X_13948_ _15461_/A _14897_/D _13876_/C _13948_/D gnd _13948_/Y vdd OAI22X1
XFILL_2__15101_ gnd vdd FILL
XFILL_5__10685_ gnd vdd FILL
XFILL_2__7167_ gnd vdd FILL
XSFILL104360x56050 gnd vdd FILL
XFILL_3__14652_ gnd vdd FILL
XFILL_2__16081_ gnd vdd FILL
XFILL_2__13293_ gnd vdd FILL
XFILL_1__15831_ gnd vdd FILL
XFILL_3__11864_ gnd vdd FILL
XFILL_0__10704_ gnd vdd FILL
XFILL_0__14472_ gnd vdd FILL
XFILL_5__15212_ gnd vdd FILL
XFILL_5__12424_ gnd vdd FILL
XSFILL74280x38050 gnd vdd FILL
XFILL_5__8965_ gnd vdd FILL
XFILL_0__11684_ gnd vdd FILL
XFILL_3__13603_ gnd vdd FILL
XFILL_5__16192_ gnd vdd FILL
XFILL_2__15032_ gnd vdd FILL
XFILL_4__15942_ gnd vdd FILL
XFILL_3__10815_ gnd vdd FILL
X_13879_ _13879_/A _13879_/B _14456_/C _13877_/Y gnd _13880_/A vdd OAI22X1
XFILL_0__16211_ gnd vdd FILL
XFILL_2__12244_ gnd vdd FILL
XFILL_4__11065_ gnd vdd FILL
XFILL_3__14583_ gnd vdd FILL
XFILL_0__13423_ gnd vdd FILL
XFILL_2__7098_ gnd vdd FILL
XFILL_0__10635_ gnd vdd FILL
XFILL_1__12974_ gnd vdd FILL
XFILL_3__7980_ gnd vdd FILL
XFILL_1__15762_ gnd vdd FILL
XFILL_3__11795_ gnd vdd FILL
X_15618_ _15616_/Y _15618_/B _15618_/C gnd _15629_/A vdd NAND3X1
XFILL_5__15143_ gnd vdd FILL
XFILL_5__8896_ gnd vdd FILL
XFILL_4__10016_ gnd vdd FILL
XFILL_3__16322_ gnd vdd FILL
XFILL_1_BUFX2_insert460 gnd vdd FILL
XFILL_5__12355_ gnd vdd FILL
XSFILL49080x14050 gnd vdd FILL
XFILL_1_BUFX2_insert471 gnd vdd FILL
XFILL112200x32050 gnd vdd FILL
XFILL_4__15873_ gnd vdd FILL
XFILL_3__13534_ gnd vdd FILL
XFILL_1_BUFX2_insert482 gnd vdd FILL
XFILL_1__11925_ gnd vdd FILL
XFILL_2__12175_ gnd vdd FILL
XFILL_1__14713_ gnd vdd FILL
XFILL_0__16142_ gnd vdd FILL
XFILL_3__6931_ gnd vdd FILL
XFILL_3__10746_ gnd vdd FILL
XFILL_0__13354_ gnd vdd FILL
XFILL_1_BUFX2_insert493 gnd vdd FILL
XFILL_1__15693_ gnd vdd FILL
XFILL_5__7847_ gnd vdd FILL
X_7500_ _7498_/Y _7460_/A _7499_/Y gnd _7500_/Y vdd OAI21X1
XFILL_0__10566_ gnd vdd FILL
XFILL_5__11306_ gnd vdd FILL
XFILL_4__14824_ gnd vdd FILL
XFILL_5__15074_ gnd vdd FILL
X_15549_ _15549_/A _15549_/B gnd _15573_/A vdd NOR2X1
XFILL_0__9941_ gnd vdd FILL
XFILL_5_BUFX2_insert809 gnd vdd FILL
X_8480_ _8548_/Q gnd _8480_/Y vdd INVX1
XFILL_2__11126_ gnd vdd FILL
XFILL_3__16253_ gnd vdd FILL
XFILL_5__12286_ gnd vdd FILL
XFILL_1__14644_ gnd vdd FILL
XFILL_3__13465_ gnd vdd FILL
XFILL_0__12305_ gnd vdd FILL
XFILL_3__9650_ gnd vdd FILL
XFILL_3__10677_ gnd vdd FILL
XFILL_3__6862_ gnd vdd FILL
XFILL_1__11856_ gnd vdd FILL
XFILL_0__16073_ gnd vdd FILL
XFILL_0__13285_ gnd vdd FILL
XFILL_5__14025_ gnd vdd FILL
XBUFX2_insert1006 _10928_/Y gnd _12224_/A vdd BUFX2
XFILL_0__10497_ gnd vdd FILL
XFILL_3__15204_ gnd vdd FILL
X_7431_ _7429_/Y _7430_/A _7431_/C gnd _7515_/D vdd OAI21X1
XFILL_5__11237_ gnd vdd FILL
XFILL_0__9872_ gnd vdd FILL
XFILL_3__12416_ gnd vdd FILL
XFILL_3__8601_ gnd vdd FILL
XBUFX2_insert1017 _15054_/Y gnd _16089_/B vdd BUFX2
XFILL_4__14755_ gnd vdd FILL
XFILL_2__9808_ gnd vdd FILL
XFILL_1__10807_ gnd vdd FILL
XFILL_3__16184_ gnd vdd FILL
XFILL_4__11967_ gnd vdd FILL
XFILL_2__15934_ gnd vdd FILL
XFILL_0__15024_ gnd vdd FILL
XBUFX2_insert1028 _13333_/Y gnd _9208_/B vdd BUFX2
XFILL_2__11057_ gnd vdd FILL
XFILL_1__14575_ gnd vdd FILL
XBUFX2_insert1039 _12390_/Y gnd _8356_/B vdd BUFX2
XFILL_6__8310_ gnd vdd FILL
XFILL_3__13396_ gnd vdd FILL
XFILL_5__9517_ gnd vdd FILL
XFILL_0__12236_ gnd vdd FILL
XFILL_1__11787_ gnd vdd FILL
XFILL_0__8823_ gnd vdd FILL
XFILL_4__13706_ gnd vdd FILL
XFILL_4__10918_ gnd vdd FILL
XFILL_2__10008_ gnd vdd FILL
X_7362_ _7354_/B _7490_/B gnd _7363_/C vdd NAND2X1
XFILL_3__15135_ gnd vdd FILL
XFILL_5__11168_ gnd vdd FILL
XFILL_2__9739_ gnd vdd FILL
XFILL_3__12347_ gnd vdd FILL
XFILL_3__8532_ gnd vdd FILL
XFILL_1__16314_ gnd vdd FILL
XSFILL69240x27050 gnd vdd FILL
XFILL_4__14686_ gnd vdd FILL
XFILL_1__13526_ gnd vdd FILL
XFILL_4__11898_ gnd vdd FILL
XFILL_2__15865_ gnd vdd FILL
X_9101_ _9101_/A _9101_/B _9100_/Y gnd _9101_/Y vdd OAI21X1
XFILL_0__12167_ gnd vdd FILL
XFILL_5__10119_ gnd vdd FILL
XFILL_4__13637_ gnd vdd FILL
XFILL_0__8754_ gnd vdd FILL
XFILL_5__15976_ gnd vdd FILL
XFILL_3__15066_ gnd vdd FILL
XFILL_2__14816_ gnd vdd FILL
XFILL_5__11099_ gnd vdd FILL
X_7293_ _7323_/A _7293_/B gnd _7293_/Y vdd NAND2X1
XFILL_3__8463_ gnd vdd FILL
XFILL_1__13457_ gnd vdd FILL
XFILL_3__12278_ gnd vdd FILL
XFILL_0__11118_ gnd vdd FILL
XFILL_1__16245_ gnd vdd FILL
XFILL_2__15796_ gnd vdd FILL
XFILL_1__10669_ gnd vdd FILL
XFILL_5__9379_ gnd vdd FILL
XFILL_0__7705_ gnd vdd FILL
XFILL_0__12098_ gnd vdd FILL
XSFILL104440x36050 gnd vdd FILL
X_9032_ _9044_/A _7240_/B gnd _9033_/C vdd NAND2X1
XFILL_3__14017_ gnd vdd FILL
XFILL_4__16356_ gnd vdd FILL
XFILL_5__14927_ gnd vdd FILL
XFILL_1__12408_ gnd vdd FILL
XFILL_3__7414_ gnd vdd FILL
XFILL_4__13568_ gnd vdd FILL
XFILL_3__11229_ gnd vdd FILL
XFILL_1__16176_ gnd vdd FILL
XSFILL8680x34050 gnd vdd FILL
XFILL_2__14747_ gnd vdd FILL
XSFILL114520x50 gnd vdd FILL
XFILL_0__15926_ gnd vdd FILL
XFILL_2__11959_ gnd vdd FILL
XFILL_3__8394_ gnd vdd FILL
XFILL_1__13388_ gnd vdd FILL
XFILL_0__11049_ gnd vdd FILL
XFILL_4__15307_ gnd vdd FILL
XFILL_4__12519_ gnd vdd FILL
XFILL_0__7636_ gnd vdd FILL
XFILL_5__14858_ gnd vdd FILL
XFILL_4__16287_ gnd vdd FILL
XFILL_1__15127_ gnd vdd FILL
XFILL_1__12339_ gnd vdd FILL
XFILL_3__7345_ gnd vdd FILL
XFILL_4__13499_ gnd vdd FILL
XFILL_2__14678_ gnd vdd FILL
XFILL_0__15857_ gnd vdd FILL
XFILL_0__7567_ gnd vdd FILL
XFILL_5__13809_ gnd vdd FILL
XFILL_4__15238_ gnd vdd FILL
XFILL_2__13629_ gnd vdd FILL
XFILL_1__15058_ gnd vdd FILL
XFILL_3__15968_ gnd vdd FILL
XFILL_5__14789_ gnd vdd FILL
XFILL_0__14808_ gnd vdd FILL
XFILL_0__15788_ gnd vdd FILL
X_9934_ _9917_/B _7502_/B gnd _9935_/C vdd NAND2X1
XFILL_3__9015_ gnd vdd FILL
XFILL_4__15169_ gnd vdd FILL
XFILL_0__7498_ gnd vdd FILL
XFILL_1__14009_ gnd vdd FILL
XSFILL108680x41050 gnd vdd FILL
XFILL_3__14919_ gnd vdd FILL
XFILL_2__16348_ gnd vdd FILL
XFILL_3__15899_ gnd vdd FILL
XFILL_0__14739_ gnd vdd FILL
XSFILL13640x35050 gnd vdd FILL
XFILL_0__9237_ gnd vdd FILL
X_9865_ _9865_/A _9737_/B gnd _9866_/C vdd NAND2X1
XFILL_2__16279_ gnd vdd FILL
XFILL_0__9168_ gnd vdd FILL
X_8816_ _8772_/A _7532_/CLK _8816_/R vdd _8816_/D gnd vdd DFFSR
X_9796_ _9796_/A gnd _9798_/A vdd INVX1
XFILL_0__16409_ gnd vdd FILL
XFILL_4__6971_ gnd vdd FILL
XFILL_0__8119_ gnd vdd FILL
XFILL_0__9099_ gnd vdd FILL
XFILL_6_BUFX2_insert643 gnd vdd FILL
X_8747_ _8745_/Y _8695_/B _8747_/C gnd _8807_/D vdd OAI21X1
XFILL_3__9917_ gnd vdd FILL
XFILL_6_BUFX2_insert654 gnd vdd FILL
XBUFX2_insert709 _12816_/Q gnd _15000_/A vdd BUFX2
XFILL_4__8710_ gnd vdd FILL
XFILL_1__9981_ gnd vdd FILL
XSFILL104520x16050 gnd vdd FILL
XSFILL33800x48050 gnd vdd FILL
X_8678_ _8678_/Q _8306_/CLK _7533_/R vdd _8678_/D gnd vdd DFFSR
XFILL_3__9848_ gnd vdd FILL
XFILL_4__8641_ gnd vdd FILL
X_7629_ _7629_/A gnd _7631_/A vdd INVX1
XFILL_1__8863_ gnd vdd FILL
XFILL_4__8572_ gnd vdd FILL
XFILL_3__9779_ gnd vdd FILL
XFILL_1_CLKBUF1_insert114 gnd vdd FILL
XSFILL23880x6050 gnd vdd FILL
XFILL_6__9488_ gnd vdd FILL
XFILL_1__7814_ gnd vdd FILL
XFILL_1_CLKBUF1_insert125 gnd vdd FILL
XFILL_1_CLKBUF1_insert136 gnd vdd FILL
XFILL_1_CLKBUF1_insert147 gnd vdd FILL
XFILL111960x58050 gnd vdd FILL
X_11230_ _11229_/Y _11230_/B gnd _11230_/Y vdd NOR2X1
XFILL_1_CLKBUF1_insert158 gnd vdd FILL
XFILL_6__8439_ gnd vdd FILL
XFILL_1_CLKBUF1_insert169 gnd vdd FILL
XFILL_1__7745_ gnd vdd FILL
XSFILL13720x15050 gnd vdd FILL
XFILL_4__7454_ gnd vdd FILL
X_11161_ _12306_/Y _11160_/Y gnd _11527_/B vdd NOR2X1
XFILL112040x67050 gnd vdd FILL
XFILL_3_BUFX2_insert500 gnd vdd FILL
XFILL_1__7676_ gnd vdd FILL
X_10112_ _10191_/B _8832_/B gnd _10113_/C vdd NAND2X1
XFILL_3_BUFX2_insert511 gnd vdd FILL
XFILL_3_BUFX2_insert522 gnd vdd FILL
XFILL_1__9415_ gnd vdd FILL
X_11092_ _12274_/Y _11092_/B gnd _11092_/Y vdd NOR2X1
XSFILL38920x81050 gnd vdd FILL
XSFILL38120x62050 gnd vdd FILL
XFILL_3_BUFX2_insert533 gnd vdd FILL
XFILL_4__9124_ gnd vdd FILL
XFILL_3_BUFX2_insert544 gnd vdd FILL
XSFILL69240x5050 gnd vdd FILL
X_10043_ _10043_/A gnd _10045_/A vdd INVX1
XFILL_3_BUFX2_insert555 gnd vdd FILL
X_14920_ _16247_/A _14441_/B _14377_/B _14919_/Y gnd _14920_/Y vdd OAI22X1
XFILL_3_BUFX2_insert566 gnd vdd FILL
XFILL_1__9346_ gnd vdd FILL
XFILL_3_BUFX2_insert577 gnd vdd FILL
XFILL_3_BUFX2_insert588 gnd vdd FILL
XFILL_3_BUFX2_insert599 gnd vdd FILL
X_14851_ _9677_/A gnd _14853_/D vdd INVX1
XFILL_2__8070_ gnd vdd FILL
XFILL_1__9277_ gnd vdd FILL
XFILL_4__8006_ gnd vdd FILL
X_13802_ _8715_/A gnd _13802_/Y vdd INVX1
XFILL_1__8228_ gnd vdd FILL
X_14782_ _14781_/Y _14778_/Y gnd _14789_/C vdd NOR2X1
X_11994_ _11991_/Y _11994_/B _11994_/C gnd _13083_/B vdd NAND3X1
X_13733_ _13733_/A _14934_/B _14897_/D _13733_/D gnd _13733_/Y vdd OAI22X1
X_10945_ _10944_/Y _10945_/B _10945_/C gnd _10973_/A vdd NAND3X1
XFILL_2__10290_ gnd vdd FILL
XFILL_5__8750_ gnd vdd FILL
X_13664_ _13664_/A _13664_/B gnd _13686_/A vdd NOR2X1
XFILL_3__11580_ gnd vdd FILL
X_10876_ _12695_/A _12792_/Q gnd _10881_/A vdd NAND2X1
XFILL_2__8972_ gnd vdd FILL
XFILL_4__8908_ gnd vdd FILL
XFILL_0__10420_ gnd vdd FILL
XFILL_5__7701_ gnd vdd FILL
X_15403_ _7694_/A gnd _15403_/Y vdd INVX1
X_12615_ _12615_/A gnd _12615_/Y vdd INVX1
XFILL_0_BUFX2_insert401 gnd vdd FILL
XFILL_4__9888_ gnd vdd FILL
XFILL_5__12140_ gnd vdd FILL
X_16383_ _16381_/Y gnd _16382_/Y gnd _16437_/D vdd OAI21X1
XFILL_0_BUFX2_insert412 gnd vdd FILL
XFILL_6__11691_ gnd vdd FILL
XFILL_3__10531_ gnd vdd FILL
X_13595_ _13595_/A _13595_/B _13595_/C gnd _13611_/A vdd NAND3X1
XFILL_4__12870_ gnd vdd FILL
XFILL_1__11710_ gnd vdd FILL
XFILL_0_BUFX2_insert423 gnd vdd FILL
XFILL_0_BUFX2_insert434 gnd vdd FILL
XSFILL64040x32050 gnd vdd FILL
XFILL_0_BUFX2_insert445 gnd vdd FILL
XFILL_4__8839_ gnd vdd FILL
XFILL_5__7632_ gnd vdd FILL
X_15334_ _15687_/A _15334_/B _15334_/C _16018_/C gnd _15334_/Y vdd OAI22X1
XSFILL38200x42050 gnd vdd FILL
XFILL_5__12071_ gnd vdd FILL
XFILL_0_BUFX2_insert456 gnd vdd FILL
X_12546_ _12031_/B _9060_/CLK _9060_/R vdd _12474_/Y gnd vdd DFFSR
XFILL_4__11821_ gnd vdd FILL
XFILL_3__13250_ gnd vdd FILL
XFILL_0_BUFX2_insert467 gnd vdd FILL
XFILL_0_BUFX2_insert478 gnd vdd FILL
XFILL_2__7854_ gnd vdd FILL
XFILL_1__11641_ gnd vdd FILL
XFILL_2__13980_ gnd vdd FILL
XFILL_0_BUFX2_insert489 gnd vdd FILL
XFILL_0__10282_ gnd vdd FILL
XFILL_5__7563_ gnd vdd FILL
XFILL_5__11022_ gnd vdd FILL
XFILL_6__10573_ gnd vdd FILL
XFILL_4__14540_ gnd vdd FILL
XFILL_3__12201_ gnd vdd FILL
X_15265_ _15265_/A _15261_/Y _15265_/C gnd _15274_/B vdd NAND3X1
X_12477_ _12477_/A vdd _12476_/Y gnd _12477_/Y vdd OAI21X1
XFILL_4__11752_ gnd vdd FILL
XFILL_0__12021_ gnd vdd FILL
XFILL_3__10393_ gnd vdd FILL
XFILL_1__14360_ gnd vdd FILL
XFILL_1__11572_ gnd vdd FILL
X_14216_ _14216_/A _14216_/B gnd _14217_/A vdd NOR2X1
XFILL_4__10703_ gnd vdd FILL
XFILL_5__7494_ gnd vdd FILL
XFILL_5__15830_ gnd vdd FILL
X_11428_ _11809_/C _11005_/Y _11428_/C gnd _11429_/A vdd NOR3X1
XFILL_1__13311_ gnd vdd FILL
XFILL_4__14471_ gnd vdd FILL
X_15196_ _15196_/A _15196_/B gnd _15207_/A vdd NAND2X1
XFILL_2__9524_ gnd vdd FILL
XSFILL3640x7050 gnd vdd FILL
XFILL_3__12132_ gnd vdd FILL
XFILL_2__15650_ gnd vdd FILL
XFILL_1__10523_ gnd vdd FILL
XFILL_4__11683_ gnd vdd FILL
XFILL_1__14291_ gnd vdd FILL
XFILL_5__9233_ gnd vdd FILL
XFILL_2__12862_ gnd vdd FILL
XFILL_4__16210_ gnd vdd FILL
XSFILL84200x45050 gnd vdd FILL
X_14147_ _9700_/Q gnd _14149_/A vdd INVX1
XFILL_4__13422_ gnd vdd FILL
X_11359_ _11359_/A _11359_/B gnd _11359_/Y vdd AND2X2
XFILL_2__14601_ gnd vdd FILL
XFILL_1__16030_ gnd vdd FILL
XFILL_5__12973_ gnd vdd FILL
XFILL_4__10634_ gnd vdd FILL
XFILL_3__12063_ gnd vdd FILL
XFILL_5__15761_ gnd vdd FILL
XFILL_1__13242_ gnd vdd FILL
XCLKBUF1_insert113 CLKBUF1_insert182/A gnd _7791_/CLK vdd CLKBUF1
XFILL_2__11813_ gnd vdd FILL
XFILL_2__15581_ gnd vdd FILL
XFILL_5__9164_ gnd vdd FILL
XCLKBUF1_insert124 CLKBUF1_insert169/A gnd _8169_/CLK vdd CLKBUF1
XFILL_0__13972_ gnd vdd FILL
XFILL_5__11924_ gnd vdd FILL
XFILL_5__14712_ gnd vdd FILL
XCLKBUF1_insert135 CLKBUF1_insert193/A gnd _7016_/CLK vdd CLKBUF1
XFILL_0__8470_ gnd vdd FILL
XFILL_3__11014_ gnd vdd FILL
XSFILL59000x21050 gnd vdd FILL
XFILL_4__16141_ gnd vdd FILL
XFILL_4__13353_ gnd vdd FILL
XCLKBUF1_insert146 CLKBUF1_insert150/A gnd _7020_/CLK vdd CLKBUF1
X_14078_ _14078_/A gnd _14078_/Y vdd INVX1
XCLKBUF1_insert157 CLKBUF1_insert218/A gnd _8051_/CLK vdd CLKBUF1
XFILL_5__15692_ gnd vdd FILL
XFILL_2__14532_ gnd vdd FILL
XFILL_4__10565_ gnd vdd FILL
XCLKBUF1_insert168 CLKBUF1_insert216/A gnd _8926_/CLK vdd CLKBUF1
XFILL_0__15711_ gnd vdd FILL
XFILL_1__13173_ gnd vdd FILL
XFILL_2__9386_ gnd vdd FILL
XFILL_5__8115_ gnd vdd FILL
XFILL_2__11744_ gnd vdd FILL
XFILL_1__10385_ gnd vdd FILL
XFILL_0__7421_ gnd vdd FILL
XSFILL105240x79050 gnd vdd FILL
XCLKBUF1_insert179 CLKBUF1_insert187/A gnd _13175_/CLK vdd CLKBUF1
X_13029_ _6896_/A gnd _13029_/Y vdd INVX1
XFILL_4__12304_ gnd vdd FILL
XFILL_5__9095_ gnd vdd FILL
XFILL_5__14643_ gnd vdd FILL
XFILL_3__15822_ gnd vdd FILL
XFILL_4__16072_ gnd vdd FILL
XFILL_5__11855_ gnd vdd FILL
XFILL_4__13284_ gnd vdd FILL
XFILL_1__12124_ gnd vdd FILL
XFILL112200x27050 gnd vdd FILL
XFILL_2__8337_ gnd vdd FILL
XFILL_4__10496_ gnd vdd FILL
XFILL_2__14463_ gnd vdd FILL
XFILL_0__15642_ gnd vdd FILL
XFILL_2__11675_ gnd vdd FILL
XFILL_0__12854_ gnd vdd FILL
XFILL_5__10806_ gnd vdd FILL
XFILL_4__15023_ gnd vdd FILL
XFILL_0__7352_ gnd vdd FILL
XFILL_5__14574_ gnd vdd FILL
XFILL_2__16202_ gnd vdd FILL
XFILL_4__12235_ gnd vdd FILL
XSFILL64120x12050 gnd vdd FILL
XFILL_2__13414_ gnd vdd FILL
XFILL_2__10626_ gnd vdd FILL
X_7980_ _7980_/A gnd _7982_/A vdd INVX1
XFILL_3__7061_ gnd vdd FILL
XFILL_5__11786_ gnd vdd FILL
XFILL_3__15753_ gnd vdd FILL
XFILL_2__8268_ gnd vdd FILL
XFILL_3__12965_ gnd vdd FILL
XFILL_1__12055_ gnd vdd FILL
XFILL_0__11805_ gnd vdd FILL
XFILL_0__15573_ gnd vdd FILL
XFILL_2__14394_ gnd vdd FILL
XFILL_0__12785_ gnd vdd FILL
XFILL_5__16313_ gnd vdd FILL
XFILL_5__13525_ gnd vdd FILL
XFILL_3__14704_ gnd vdd FILL
XFILL_6__15864_ gnd vdd FILL
X_6931_ _6931_/A _6982_/B _6930_/Y gnd _7007_/D vdd OAI21X1
XFILL_3__11916_ gnd vdd FILL
XFILL_4__12166_ gnd vdd FILL
XSFILL18680x7050 gnd vdd FILL
XFILL_2__7219_ gnd vdd FILL
XFILL_1__11006_ gnd vdd FILL
XFILL_2__16133_ gnd vdd FILL
XFILL_2__13345_ gnd vdd FILL
XFILL_3__15684_ gnd vdd FILL
XFILL_2__10557_ gnd vdd FILL
XFILL_0__14524_ gnd vdd FILL
XFILL_3__12896_ gnd vdd FILL
XFILL_0__9022_ gnd vdd FILL
XFILL_0__11736_ gnd vdd FILL
XFILL_2__8199_ gnd vdd FILL
XSFILL53960x55050 gnd vdd FILL
XFILL_6__14815_ gnd vdd FILL
XFILL_5__9997_ gnd vdd FILL
XFILL_5__16244_ gnd vdd FILL
XFILL_5__13456_ gnd vdd FILL
XFILL_4__11117_ gnd vdd FILL
X_9650_ _9650_/A gnd _9650_/Y vdd INVX1
XFILL_3__14635_ gnd vdd FILL
X_6862_ _6862_/A gnd memoryAddress[24] vdd BUFX2
XFILL_5__10668_ gnd vdd FILL
XFILL_2__13276_ gnd vdd FILL
XFILL_4__12097_ gnd vdd FILL
XFILL_1__15814_ gnd vdd FILL
XFILL_2__16064_ gnd vdd FILL
XFILL_3__11847_ gnd vdd FILL
XFILL_0__14455_ gnd vdd FILL
XFILL_2__10488_ gnd vdd FILL
XFILL_5__12407_ gnd vdd FILL
X_8601_ _8601_/A _8609_/A _8600_/Y gnd _8673_/D vdd OAI21X1
XFILL_0__11667_ gnd vdd FILL
XFILL_5__16175_ gnd vdd FILL
XSFILL28760x31050 gnd vdd FILL
X_9581_ _9581_/Q _7021_/CLK _9062_/R vdd _9533_/Y gnd vdd DFFSR
XFILL_4__15925_ gnd vdd FILL
XFILL_5__13387_ gnd vdd FILL
XFILL_2__15015_ gnd vdd FILL
XFILL_2__12227_ gnd vdd FILL
XFILL_4__11048_ gnd vdd FILL
XFILL_3__14566_ gnd vdd FILL
XSFILL54040x64050 gnd vdd FILL
XFILL_0__13406_ gnd vdd FILL
XFILL_3__7963_ gnd vdd FILL
XFILL_0__10618_ gnd vdd FILL
XSFILL33880x1050 gnd vdd FILL
XFILL_3__11778_ gnd vdd FILL
XFILL_1__15745_ gnd vdd FILL
XFILL_0__14386_ gnd vdd FILL
XFILL_5__15126_ gnd vdd FILL
XFILL_1__12957_ gnd vdd FILL
X_8532_ _8440_/B _9556_/B gnd _8532_/Y vdd NAND2X1
XFILL_1_BUFX2_insert290 gnd vdd FILL
XFILL_3__16305_ gnd vdd FILL
XFILL_5__12338_ gnd vdd FILL
XFILL_0__11598_ gnd vdd FILL
XFILL_5__8879_ gnd vdd FILL
XSFILL14040x80050 gnd vdd FILL
XFILL_6__14677_ gnd vdd FILL
XFILL_3__13517_ gnd vdd FILL
XFILL_5_BUFX2_insert606 gnd vdd FILL
XFILL_3__6914_ gnd vdd FILL
XFILL_2__12158_ gnd vdd FILL
XFILL_0__16125_ gnd vdd FILL
XFILL_4__15856_ gnd vdd FILL
XFILL_0__13337_ gnd vdd FILL
XFILL_3__14497_ gnd vdd FILL
XFILL_1__11908_ gnd vdd FILL
XFILL_0__10549_ gnd vdd FILL
XFILL_1__15676_ gnd vdd FILL
XFILL_1__12888_ gnd vdd FILL
XFILL_5_BUFX2_insert617 gnd vdd FILL
XFILL_6__16416_ gnd vdd FILL
XFILL_6__13628_ gnd vdd FILL
XFILL_5_BUFX2_insert628 gnd vdd FILL
XFILL_5__15057_ gnd vdd FILL
XFILL_0__9924_ gnd vdd FILL
X_8463_ _8508_/A _7439_/B gnd _8464_/C vdd NAND2X1
XFILL_3__16236_ gnd vdd FILL
XFILL_4__14807_ gnd vdd FILL
XFILL_5_BUFX2_insert639 gnd vdd FILL
XFILL_5__12269_ gnd vdd FILL
XFILL_2__11109_ gnd vdd FILL
XFILL_3__9633_ gnd vdd FILL
XFILL_3__13448_ gnd vdd FILL
XFILL_4__15787_ gnd vdd FILL
XFILL_1__14627_ gnd vdd FILL
XFILL_3__6845_ gnd vdd FILL
XFILL_2__12089_ gnd vdd FILL
XFILL_4__12999_ gnd vdd FILL
XFILL_0__16056_ gnd vdd FILL
XFILL_1__11839_ gnd vdd FILL
XFILL_0__13268_ gnd vdd FILL
XFILL_5__14008_ gnd vdd FILL
X_7414_ _7510_/Q gnd _7416_/A vdd INVX1
XFILL_0_BUFX2_insert990 gnd vdd FILL
XFILL_0__9855_ gnd vdd FILL
XFILL_4__14738_ gnd vdd FILL
XFILL111800x6050 gnd vdd FILL
XSFILL18680x83050 gnd vdd FILL
XFILL_2__15917_ gnd vdd FILL
X_8394_ _8394_/A gnd _8394_/Y vdd INVX1
XFILL_3__16167_ gnd vdd FILL
XFILL_0__15007_ gnd vdd FILL
XSFILL48920x44050 gnd vdd FILL
XSFILL99560x79050 gnd vdd FILL
XFILL_3__13379_ gnd vdd FILL
XFILL_0__12219_ gnd vdd FILL
XFILL_1__14558_ gnd vdd FILL
X_7345_ _7345_/A _7366_/B _7344_/Y gnd _7345_/Y vdd OAI21X1
XFILL_3__15118_ gnd vdd FILL
XFILL_6__16278_ gnd vdd FILL
XFILL_0__9786_ gnd vdd FILL
XFILL_3__8515_ gnd vdd FILL
XFILL_4__14669_ gnd vdd FILL
XFILL_3__16098_ gnd vdd FILL
XFILL_2__15848_ gnd vdd FILL
XFILL_1__13509_ gnd vdd FILL
XFILL_1__14489_ gnd vdd FILL
XFILL_3__9495_ gnd vdd FILL
XFILL_6__15229_ gnd vdd FILL
XSFILL49000x53050 gnd vdd FILL
XSFILL33320x3050 gnd vdd FILL
XFILL_4__16408_ gnd vdd FILL
XFILL_0__8737_ gnd vdd FILL
XFILL_3__15049_ gnd vdd FILL
XFILL_5__15959_ gnd vdd FILL
X_7276_ _7276_/Q _9953_/CLK _7276_/R vdd _7226_/Y gnd vdd DFFSR
XFILL_1__16228_ gnd vdd FILL
XFILL_3__8446_ gnd vdd FILL
XFILL_2_CLKBUF1_insert209 gnd vdd FILL
XFILL_2__15779_ gnd vdd FILL
X_9015_ _9015_/A _9014_/A _9014_/Y gnd _9015_/Y vdd OAI21X1
XSFILL109560x64050 gnd vdd FILL
XFILL_1__7461_ gnd vdd FILL
XFILL_4__16339_ gnd vdd FILL
XFILL_4__7170_ gnd vdd FILL
XSFILL38040x77050 gnd vdd FILL
XFILL_3__8377_ gnd vdd FILL
XFILL_0__15909_ gnd vdd FILL
XSFILL28840x11050 gnd vdd FILL
XFILL_1__16159_ gnd vdd FILL
XSFILL54120x44050 gnd vdd FILL
XFILL_0__7619_ gnd vdd FILL
XFILL_3__7328_ gnd vdd FILL
XFILL_0__8599_ gnd vdd FILL
XSFILL33800x9050 gnd vdd FILL
XFILL_2_BUFX2_insert507 gnd vdd FILL
XFILL_2_BUFX2_insert518 gnd vdd FILL
XFILL_1__9131_ gnd vdd FILL
XFILL_2_BUFX2_insert529 gnd vdd FILL
X_9917_ _9915_/Y _9917_/B _9917_/C gnd _9917_/Y vdd OAI21X1
XFILL_1__8013_ gnd vdd FILL
XSFILL18760x63050 gnd vdd FILL
XSFILL8600x73050 gnd vdd FILL
XFILL_6_BUFX2_insert1037 gnd vdd FILL
X_9848_ _9848_/A _9865_/A _9847_/Y gnd _9942_/D vdd OAI21X1
XFILL_4__9811_ gnd vdd FILL
X_10730_ _14414_/D _7156_/CLK _7391_/R vdd _10730_/D gnd vdd DFFSR
XSFILL99240x61050 gnd vdd FILL
XFILL_4__9742_ gnd vdd FILL
X_9779_ _9785_/A _9779_/B gnd _9779_/Y vdd NAND2X1
XBUFX2_insert506 BUFX2_insert518/A gnd _9963_/R vdd BUFX2
XFILL_4__6954_ gnd vdd FILL
X_10661_ _10661_/A _10661_/B _10660_/Y gnd _10661_/Y vdd OAI21X1
XBUFX2_insert517 BUFX2_insert520/A gnd _9056_/R vdd BUFX2
XBUFX2_insert528 BUFX2_insert600/A gnd _13201_/R vdd BUFX2
XBUFX2_insert539 BUFX2_insert607/A gnd _8430_/R vdd BUFX2
XSFILL38680x14050 gnd vdd FILL
X_12400_ _12496_/A gnd _12400_/Y vdd INVX1
XFILL_4__9673_ gnd vdd FILL
XFILL_6_BUFX2_insert495 gnd vdd FILL
XFILL_4__6885_ gnd vdd FILL
X_13380_ _12808_/Q _12807_/Q gnd _13381_/B vdd NOR2X1
X_10592_ _10592_/Q _8433_/CLK _7921_/R vdd _10518_/Y gnd vdd DFFSR
XFILL_1__8915_ gnd vdd FILL
XSFILL38920x76050 gnd vdd FILL
XFILL_1__9895_ gnd vdd FILL
XFILL_4__8624_ gnd vdd FILL
XFILL112440x83050 gnd vdd FILL
X_12331_ _12327_/A gnd _12319_/C gnd _12331_/Y vdd NAND3X1
XFILL_4_BUFX2_insert1030 gnd vdd FILL
XFILL_4_BUFX2_insert1041 gnd vdd FILL
XFILL_1__8846_ gnd vdd FILL
XFILL_4_BUFX2_insert1052 gnd vdd FILL
XFILL_4_BUFX2_insert1063 gnd vdd FILL
X_15050_ _15000_/A _15061_/C _15044_/C gnd _15050_/Y vdd NAND3X1
X_12262_ _12259_/Y _12260_/Y _12262_/C gnd _12262_/Y vdd NAND3X1
XFILL_4_BUFX2_insert1085 gnd vdd FILL
XFILL_2__7570_ gnd vdd FILL
XFILL_4__7506_ gnd vdd FILL
XFILL_1__8777_ gnd vdd FILL
X_14001_ _9367_/A _13883_/B _14000_/Y gnd _14012_/A vdd AOI21X1
XSFILL84680x17050 gnd vdd FILL
X_11213_ _10993_/Y _12338_/Y _11212_/Y gnd _11220_/B vdd OAI21X1
XFILL_4__8486_ gnd vdd FILL
X_12193_ _13157_/A gnd _12195_/A vdd INVX1
XFILL_1__7728_ gnd vdd FILL
XFILL_4__7437_ gnd vdd FILL
XSFILL18840x43050 gnd vdd FILL
X_11144_ _11120_/Y _11130_/B gnd _11582_/C vdd NOR2X1
XSFILL44120x76050 gnd vdd FILL
XFILL_2__9240_ gnd vdd FILL
XFILL_3_BUFX2_insert330 gnd vdd FILL
XFILL_3_BUFX2_insert341 gnd vdd FILL
XFILL_4__7368_ gnd vdd FILL
X_15952_ _10552_/A gnd _15953_/B vdd INVX1
XSFILL99320x41050 gnd vdd FILL
X_11075_ _12254_/Y _12144_/Y gnd _11081_/A vdd XNOR2X1
XFILL_3_BUFX2_insert352 gnd vdd FILL
XFILL_3_BUFX2_insert363 gnd vdd FILL
XFILL_2__9171_ gnd vdd FILL
XFILL_4__9107_ gnd vdd FILL
XFILL_3_BUFX2_insert374 gnd vdd FILL
XFILL_1__10170_ gnd vdd FILL
XFILL_3_BUFX2_insert385 gnd vdd FILL
X_14903_ _8180_/Q gnd _16254_/C vdd INVX1
X_10026_ _9979_/B _9770_/B gnd _10027_/C vdd NAND2X1
XFILL_3_BUFX2_insert396 gnd vdd FILL
XFILL_4__7299_ gnd vdd FILL
XFILL_5__11640_ gnd vdd FILL
XFILL_2__8122_ gnd vdd FILL
X_15883_ _9194_/Q gnd _15883_/Y vdd INVX1
XFILL_4__10281_ gnd vdd FILL
XSFILL110200x12050 gnd vdd FILL
XFILL_2__11460_ gnd vdd FILL
XFILL_4__9038_ gnd vdd FILL
XFILL_5__9920_ gnd vdd FILL
XSFILL64040x27050 gnd vdd FILL
XFILL_4__12020_ gnd vdd FILL
X_14834_ _14834_/A _14833_/Y _15338_/C gnd _13036_/B vdd AOI21X1
XFILL_2__10411_ gnd vdd FILL
XFILL_5__11571_ gnd vdd FILL
XFILL_3__12750_ gnd vdd FILL
XFILL_2__11391_ gnd vdd FILL
XFILL_5__13310_ gnd vdd FILL
XFILL_0__12570_ gnd vdd FILL
XFILL_5__9851_ gnd vdd FILL
XFILL_5__10522_ gnd vdd FILL
XFILL_2__13130_ gnd vdd FILL
XFILL_5__14290_ gnd vdd FILL
XFILL_3__11701_ gnd vdd FILL
X_14765_ _14765_/A _14764_/Y gnd _14765_/Y vdd NOR2X1
X_11977_ _12108_/B gnd _11979_/A vdd INVX1
XFILL_0__11521_ gnd vdd FILL
XFILL_1__13860_ gnd vdd FILL
XFILL_6__14600_ gnd vdd FILL
XFILL_5__9782_ gnd vdd FILL
XFILL_5__13241_ gnd vdd FILL
X_13716_ _15286_/C _13461_/C gnd _13717_/C vdd NOR2X1
X_10928_ _10938_/A _10906_/A _10938_/B _10929_/A gnd _10928_/Y vdd OAI22X1
XFILL_5__10453_ gnd vdd FILL
XFILL_3__14420_ gnd vdd FILL
XFILL_5__6994_ gnd vdd FILL
XFILL_4_CLKBUF1_insert120 gnd vdd FILL
X_14696_ _8900_/A gnd _16099_/A vdd INVX1
XFILL_3__11632_ gnd vdd FILL
XFILL_4__13971_ gnd vdd FILL
XFILL_4_CLKBUF1_insert131 gnd vdd FILL
XFILL_0__14240_ gnd vdd FILL
XFILL_2__10273_ gnd vdd FILL
XFILL_1__13791_ gnd vdd FILL
XFILL_0__11452_ gnd vdd FILL
XFILL_5__8733_ gnd vdd FILL
XFILL_4_CLKBUF1_insert142 gnd vdd FILL
X_16435_ _15787_/A _7912_/CLK _7911_/R vdd _16435_/D gnd vdd DFFSR
XFILL_4__15710_ gnd vdd FILL
X_13647_ _8410_/Q _13647_/B _13864_/B _8666_/Q gnd _13647_/Y vdd AOI22X1
XFILL_2__12012_ gnd vdd FILL
XFILL_4_CLKBUF1_insert153 gnd vdd FILL
XFILL_5__13172_ gnd vdd FILL
XFILL_6__11743_ gnd vdd FILL
X_10859_ _10859_/Q _9963_/CLK _9963_/R vdd _10859_/D gnd vdd DFFSR
XFILL_5__10384_ gnd vdd FILL
XFILL_4_CLKBUF1_insert164 gnd vdd FILL
XFILL_3__14351_ gnd vdd FILL
XFILL_0__10403_ gnd vdd FILL
XFILL_1__12742_ gnd vdd FILL
XFILL_1__15530_ gnd vdd FILL
XFILL_2__8955_ gnd vdd FILL
XFILL_4_CLKBUF1_insert175 gnd vdd FILL
XFILL_3__11563_ gnd vdd FILL
XFILL_4_CLKBUF1_insert186 gnd vdd FILL
XSFILL44200x56050 gnd vdd FILL
XFILL_0__14171_ gnd vdd FILL
XFILL_0_BUFX2_insert231 gnd vdd FILL
XFILL_5__12123_ gnd vdd FILL
XFILL_0__11383_ gnd vdd FILL
XFILL_3__13302_ gnd vdd FILL
XFILL_6__14462_ gnd vdd FILL
XFILL_0_BUFX2_insert242 gnd vdd FILL
XFILL_4__15641_ gnd vdd FILL
XSFILL59800x35050 gnd vdd FILL
XSFILL59000x16050 gnd vdd FILL
X_16366_ _16432_/Q gnd _16368_/A vdd INVX1
XFILL_4_CLKBUF1_insert197 gnd vdd FILL
XFILL_0_BUFX2_insert253 gnd vdd FILL
XFILL_0__7970_ gnd vdd FILL
XFILL_4__12853_ gnd vdd FILL
X_13578_ _13578_/A _13578_/B gnd _13582_/C vdd NOR2X1
XFILL_3__10514_ gnd vdd FILL
XFILL_0__13122_ gnd vdd FILL
XFILL_0_BUFX2_insert264 gnd vdd FILL
XFILL_3__14282_ gnd vdd FILL
XFILL_2__8886_ gnd vdd FILL
XFILL_5__7615_ gnd vdd FILL
XFILL_6__16201_ gnd vdd FILL
XFILL_3__11494_ gnd vdd FILL
XFILL_1__15461_ gnd vdd FILL
XSFILL99400x21050 gnd vdd FILL
X_15317_ _15317_/A _15378_/B gnd _15317_/Y vdd NOR2X1
XFILL_6__13413_ gnd vdd FILL
XFILL_0_BUFX2_insert275 gnd vdd FILL
XFILL_0__6921_ gnd vdd FILL
XFILL_3__16021_ gnd vdd FILL
XFILL_0_BUFX2_insert286 gnd vdd FILL
XFILL_5__12054_ gnd vdd FILL
X_12529_ _12107_/B gnd _12529_/Y vdd INVX1
XFILL_5__8595_ gnd vdd FILL
XFILL_4__11804_ gnd vdd FILL
XFILL_3__13233_ gnd vdd FILL
XFILL_4__15572_ gnd vdd FILL
X_16297_ _15550_/A _14947_/Y _15550_/C gnd _16297_/Y vdd NOR3X1
XFILL_0_BUFX2_insert297 gnd vdd FILL
XFILL_4__12784_ gnd vdd FILL
XFILL_3__10445_ gnd vdd FILL
XFILL_2__7837_ gnd vdd FILL
XFILL_1__11624_ gnd vdd FILL
XFILL_1__14412_ gnd vdd FILL
XFILL_1__15392_ gnd vdd FILL
XFILL_2__13963_ gnd vdd FILL
XFILL_0__10265_ gnd vdd FILL
XFILL_5__7546_ gnd vdd FILL
XFILL_5__11005_ gnd vdd FILL
XFILL_0__9640_ gnd vdd FILL
X_15248_ _7682_/A gnd _15248_/Y vdd INVX1
XFILL_4__14523_ gnd vdd FILL
XFILL_2__15702_ gnd vdd FILL
XFILL_0__6852_ gnd vdd FILL
XFILL_4__11735_ gnd vdd FILL
XFILL_3__10376_ gnd vdd FILL
XFILL_3__13164_ gnd vdd FILL
XFILL_0__12004_ gnd vdd FILL
XFILL_1__14343_ gnd vdd FILL
XFILL_2__12914_ gnd vdd FILL
XFILL_1__11555_ gnd vdd FILL
XFILL_2__13894_ gnd vdd FILL
XFILL_6__13275_ gnd vdd FILL
XFILL_5__7477_ gnd vdd FILL
X_7130_ _7130_/Q _8541_/CLK _7140_/R vdd _7130_/D gnd vdd DFFSR
XFILL_2_BUFX2_insert13 gnd vdd FILL
XFILL_0__10196_ gnd vdd FILL
XFILL_5__15813_ gnd vdd FILL
XFILL_6__16063_ gnd vdd FILL
XFILL_2__9507_ gnd vdd FILL
XFILL_4__14454_ gnd vdd FILL
X_15179_ _8447_/A gnd _15179_/Y vdd INVX1
XFILL_3__12115_ gnd vdd FILL
XFILL_2_BUFX2_insert24 gnd vdd FILL
XFILL_1__10506_ gnd vdd FILL
XFILL_2__15633_ gnd vdd FILL
XSFILL43800x4050 gnd vdd FILL
XFILL_4__11666_ gnd vdd FILL
XFILL_3__9280_ gnd vdd FILL
XFILL_5__9216_ gnd vdd FILL
XFILL_2_BUFX2_insert35 gnd vdd FILL
XFILL_2__12845_ gnd vdd FILL
XFILL_3__13095_ gnd vdd FILL
XFILL_1__14274_ gnd vdd FILL
XFILL_2_BUFX2_insert46 gnd vdd FILL
XFILL_6__15014_ gnd vdd FILL
XFILL_1__11486_ gnd vdd FILL
XFILL_2__7699_ gnd vdd FILL
XFILL_2_BUFX2_insert57 gnd vdd FILL
XSFILL89320x73050 gnd vdd FILL
XFILL_4__13405_ gnd vdd FILL
XFILL_0__8522_ gnd vdd FILL
XFILL_2_BUFX2_insert68 gnd vdd FILL
XFILL_4__10617_ gnd vdd FILL
X_7061_ _7061_/A _7061_/B gnd _7061_/Y vdd NAND2X1
XFILL_5__15744_ gnd vdd FILL
XFILL_1__13225_ gnd vdd FILL
XFILL_1__16013_ gnd vdd FILL
XFILL_2_BUFX2_insert79 gnd vdd FILL
XFILL_3__8231_ gnd vdd FILL
XFILL_3__12046_ gnd vdd FILL
XFILL_4__14385_ gnd vdd FILL
XSFILL3560x14050 gnd vdd FILL
XFILL_5__12956_ gnd vdd FILL
XSFILL109480x79050 gnd vdd FILL
XFILL_1__10437_ gnd vdd FILL
XFILL_2__15564_ gnd vdd FILL
XFILL_4__11597_ gnd vdd FILL
XFILL_5__9147_ gnd vdd FILL
XFILL_2__12776_ gnd vdd FILL
XFILL_0__13955_ gnd vdd FILL
XFILL_6__12157_ gnd vdd FILL
XFILL_4__16124_ gnd vdd FILL
XFILL_4__13336_ gnd vdd FILL
XSFILL3000x57050 gnd vdd FILL
XFILL_5__11907_ gnd vdd FILL
XFILL_0__8453_ gnd vdd FILL
XSFILL28760x26050 gnd vdd FILL
.ends

