/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module mips(
    inout vdd,
    inout gnd,
    output MemRead,
    output MemWrite,
    input clk,
    output [31:0] memoryAddress,
    input [31:0] memoryOutData,
    output [31:0] memoryWriteData,
    input rst
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf2  ;
wire _1677_ ;
wire _1257_ ;
wire _5090_ ;
wire [31:0] _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire IRWrite_bF$buf0 ;
wire IRWrite_bF$buf1 ;
wire _1486_ ;
wire IRWrite_bF$buf2 ;
wire _1066_ ;
wire IRWrite_bF$buf3 ;
wire IRWrite_bF$buf4 ;
wire IRWrite_bF$buf5 ;
wire IRWrite_bF$buf6 ;
wire IRWrite_bF$buf7 ;
wire _397_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _2712_ ;
wire _5515__bF$buf0 ;
wire _5515__bF$buf1 ;
wire _5515__bF$buf2 ;
wire _5515__bF$buf3 ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf1  ;
wire \datapath_1.mux_wd3.dout_11_bF$buf4  ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _1830_ ;
wire _1410_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf0  ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf0  ;
wire _57_ ;
wire _6504_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _3884__bF$buf0 ;
wire _3884__bF$buf1 ;
wire _3884__bF$buf2 ;
wire _3884__bF$buf3 ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf4  ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf2  ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6542_ ;
wire _6122_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf3  ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _5813_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf0  ;
wire _6771_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf7  ;
wire _6351_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf3  ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf7  ;
wire _6580_ ;
wire _6160_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf5  ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _5907_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _3947__bF$buf0 ;
wire _3947__bF$buf1 ;
wire _3947__bF$buf2 ;
wire _3947__bF$buf3 ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf3  ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _2594_ ;
wire _2174_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire [31:0] \datapath_1.regfile_1.regOut[13]  ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _5503__bF$buf0 ;
wire _5503__bF$buf1 ;
wire _5503__bF$buf2 ;
wire _5503__bF$buf3 ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire \datapath_1.PCJump_27_bF$buf2  ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _2341__bF$buf0 ;
wire _2341__bF$buf1 ;
wire _2341__bF$buf2 ;
wire _2341__bF$buf3 ;
wire _4643_ ;
wire _4223_ ;
wire [31:0] \datapath_1.regfile_1.regOut[7]  ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf2  ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _5495__bF$buf0 ;
wire _5495__bF$buf1 ;
wire _5495__bF$buf2 ;
wire _5495__bF$buf3 ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf1  ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _3966__bF$buf0 ;
wire _3966__bF$buf1 ;
wire _3966__bF$buf2 ;
wire _3966__bF$buf3 ;
wire _1386_ ;
wire _297_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf5  ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _5518__bF$buf0 ;
wire _5518__bF$buf1 ;
wire _5518__bF$buf2 ;
wire _5518__bF$buf3 ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf1  ;
wire _54_ ;
wire _6501_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf4  ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _4584_ ;
wire _4164_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf1  ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf0  ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf0  ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire PCWrite ;
wire _4678_ ;
wire _4258_ ;
wire _6824_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf4  ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf2  ;
wire _3282_ ;
wire RegWrite_bF$buf0 ;
wire RegWrite_bF$buf1 ;
wire RegWrite_bF$buf2 ;
wire RegWrite_bF$buf3 ;
wire RegWrite_bF$buf4 ;
wire RegWrite_bF$buf5 ;
wire RegWrite_bF$buf6 ;
wire RegWrite_bF$buf7 ;
wire _4487_ ;
wire _4067_ ;
wire _3891__bF$buf0 ;
wire _3891__bF$buf1 ;
wire _3891__bF$buf2 ;
wire _3891__bF$buf3 ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _5904_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6442_ ;
wire _6022_ ;
wire _2782_ ;
wire _2362_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf0  ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf3  ;
wire _5713_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _2591_ ;
wire _2171_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf7  ;
wire _3796_ ;
wire _3376_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf3  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire \datapath_1.PCJump_22_bF$buf3  ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf7  ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _5807_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf3  ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _4831_ ;
wire _3954__bF$buf0 ;
wire _4411_ ;
wire _3954__bF$buf1 ;
wire _3954__bF$buf2 ;
wire _3954__bF$buf3 ;
wire _3954__bF$buf4 ;
wire \datapath_1.regfile_1.regEn_8_bF$buf7  ;
wire _5616_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6574_ ;
wire _6154_ ;
wire _2494_ ;
wire _2074_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _3088_ ;
wire _5654_ ;
wire _5234_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _4734_ ;
wire _4314_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf2  ;
wire _5939_ ;
wire _5519_ ;
wire _2344__bF$buf0 ;
wire _2344__bF$buf1 ;
wire _2344__bF$buf2 ;
wire _2344__bF$buf3 ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf2  ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf1  ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf5  ;
wire _1286_ ;
wire _197_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _2932_ ;
wire _2512_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf1  ;
wire _3717_ ;
wire _6189_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf4  ;
wire _3902__bF$buf0 ;
wire _3902__bF$buf1 ;
wire _3902__bF$buf2 ;
wire _3902__bF$buf3 ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _2741_ ;
wire _2321_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf1  ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf4  ;
wire _7_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _1821_ ;
wire _1401_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf0  ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf4  ;
wire _3793_ ;
wire _3373_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf0  ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire Branch ;
wire \datapath_1.PCJump_22_bF$buf0  ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf4  ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6533_ ;
wire _6113_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _5804_ ;
wire _1724_ ;
wire _1304_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf3  ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf0  ;
wire _6762_ ;
wire _6342_ ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf4  ;
wire _5613_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf7  ;
wire _6818_ ;
wire [31:0] _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6571_ ;
wire _6151_ ;
wire _2491_ ;
wire _2071_ ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire rst_bF$buf110 ;
wire rst_bF$buf111 ;
wire rst_bF$buf112 ;
wire rst_bF$buf113 ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _5707_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _4731_ ;
wire _4311_ ;
wire RegDst ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6474_ ;
wire _6054_ ;
wire _2394_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire clk_bF$buf80 ;
wire clk_bF$buf81 ;
wire clk_bF$buf82 ;
wire clk_bF$buf83 ;
wire clk_bF$buf84 ;
wire clk_bF$buf85 ;
wire clk_bF$buf86 ;
wire [31:0] _3620_ ;
wire clk_bF$buf87 ;
wire _3200_ ;
wire clk_bF$buf88 ;
wire clk_bF$buf89 ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _5783_ ;
wire _5363_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf2  ;
wire _2347__bF$buf0 ;
wire _2347__bF$buf1 ;
wire _2347__bF$buf2 ;
wire _2347__bF$buf3 ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf1  ;
wire _4919_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf5  ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf1  ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf5  ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire _3905__bF$buf0 ;
wire _3905__bF$buf1 ;
wire _3905__bF$buf2 ;
wire _3905__bF$buf3 ;
wire _45_ ;
wire _5532__bF$buf0 ;
wire _5532__bF$buf1 ;
wire _5532__bF$buf2 ;
wire _5532__bF$buf3 ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf1  ;
wire _3790_ ;
wire _3370_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf4  ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _2641_ ;
wire _2221_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf5  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf1  ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _1721_ ;
wire _1301_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf0  ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf1  ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf4  ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _670_ ;
wire _250_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6433_ ;
wire _6013_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _5704_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire _1853_ ;
wire [31:0] _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6471_ ;
wire _6051_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf2  ;
wire [31:0] \datapath_1.regfile_1.regOut[2]  ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire clk_bF$buf50 ;
wire clk_bF$buf51 ;
wire clk_bF$buf52 ;
wire clk_bF$buf53 ;
wire clk_bF$buf54 ;
wire clk_bF$buf55 ;
wire clk_bF$buf56 ;
wire clk_bF$buf57 ;
wire clk_bF$buf58 ;
wire clk_bF$buf59 ;
wire _4822_ ;
wire _4402_ ;
wire _5607_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6565_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf2  ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _2294_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire [31:0] \datapath_1.regfile_1.regOut[25]  ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf2  ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire [31:0] _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _5683_ ;
wire _5263_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf2  ;
wire _2388_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _4763_ ;
wire _4343_ ;
wire rst_bF$buf0 ;
wire rst_bF$buf1 ;
wire rst_bF$buf2 ;
wire rst_bF$buf3 ;
wire rst_bF$buf4 ;
wire rst_bF$buf5 ;
wire _5968_ ;
wire rst_bF$buf6 ;
wire _5548_ ;
wire rst_bF$buf7 ;
wire _5128_ ;
wire rst_bF$buf8 ;
wire rst_bF$buf9 ;
wire _42_ ;
wire [31:0] _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf1  ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf2  ;
wire _4628_ ;
wire _4208_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf5  ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _3983__bF$buf0 ;
wire _3983__bF$buf1 ;
wire _3983__bF$buf2 ;
wire _3983__bF$buf3 ;
wire _3983__bF$buf4 ;
wire _1086_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _5535__bF$buf0 ;
wire _5535__bF$buf1 ;
wire _5535__bF$buf2 ;
wire _5535__bF$buf3 ;
wire _5535__bF$buf4 ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf1  ;
wire _6812_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf4  ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf5  ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf4  ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire _1812_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6430_ ;
wire _6010_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire [31:0] _3555_ ;
wire _3135_ ;
wire rst_bF$buf90 ;
wire rst_bF$buf91 ;
wire rst_bF$buf92 ;
wire rst_bF$buf93 ;
wire rst_bF$buf94 ;
wire rst_bF$buf95 ;
wire rst_bF$buf96 ;
wire rst_bF$buf97 ;
wire rst_bF$buf98 ;
wire rst_bF$buf99 ;
wire _5701_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire IorD ;
wire clk ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6524_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _2673_ ;
wire _2253_ ;
wire clk_bF$buf20 ;
wire clk_bF$buf21 ;
wire clk_bF$buf22 ;
wire clk_bF$buf23 ;
wire clk_bF$buf24 ;
wire clk_bF$buf25 ;
wire clk_bF$buf26 ;
wire clk_bF$buf27 ;
wire clk_bF$buf28 ;
wire clk_bF$buf29 ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _5604_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6562_ ;
wire _6142_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf2  ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _4722_ ;
wire _4302_ ;
wire _3967__bF$buf0 ;
wire _3967__bF$buf1 ;
wire _3967__bF$buf2 ;
wire _3967__bF$buf3 ;
wire _5927_ ;
wire _5507_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf5  ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _2385_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _2194_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire [31:0] \datapath_1.regfile_1.regOut[15]  ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf4  ;
wire _4816_ ;
wire _5774_ ;
wire _5354_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf2  ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf6  ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _4663_ ;
wire _4243_ ;
wire [31:0] \datapath_1.regfile_1.regOut[9]  ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf1  ;
wire _1788_ ;
wire [31:0] _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf2  ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf1  ;
wire _1597_ ;
wire _1177_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf5  ;
wire _5486_ ;
wire _5066_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire rst_bF$buf60 ;
wire rst_bF$buf61 ;
wire rst_bF$buf62 ;
wire rst_bF$buf63 ;
wire rst_bF$buf64 ;
wire rst_bF$buf65 ;
wire rst_bF$buf66 ;
wire rst_bF$buf67 ;
wire rst_bF$buf68 ;
wire rst_bF$buf69 ;
wire _4757_ ;
wire _4337_ ;
wire _36_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf5  ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire RegWrite ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6521_ ;
wire _6101_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _1712_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf3  ;
wire _5601_ ;
wire [31:0] \datapath_1.mux_pcsrc.dout  ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _5459__bF$buf0 ;
wire _5459__bF$buf1 ;
wire _5459__bF$buf2 ;
wire _4910_ ;
wire _5459__bF$buf3 ;
wire [31:0] \datapath_1.regfile_1.regOut[30]  ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _5463__bF$buf0 ;
wire _5463__bF$buf1 ;
wire _5463__bF$buf2 ;
wire _5463__bF$buf3 ;
wire [5:0] \control_1.op  ;
wire _3778_ ;
wire _3358_ ;
wire _5924_ ;
wire _5504_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _3032__bF$buf0 ;
wire _3032__bF$buf1 ;
wire _3032__bF$buf2 ;
wire _3032__bF$buf3 ;
wire _3032__bF$buf4 ;
wire _755_ ;
wire _335_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf2  ;
wire _2629_ ;
wire _2209_ ;
wire _6462_ ;
wire _6042_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _2191_ ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf1  ;
wire _4813_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf5  ;
wire _4622_ ;
wire _4202_ ;
wire _5827_ ;
wire _5407_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf2  ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf3  ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _5526__bF$buf0 ;
wire _5526__bF$buf1 ;
wire _5526__bF$buf2 ;
wire _5526__bF$buf3 ;
wire _5526__bF$buf4 ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _2094_ ;
wire _3299_ ;
wire _4660_ ;
wire _4240_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf4  ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _5530__bF$buf0 ;
wire _5530__bF$buf1 ;
wire _5530__bF$buf2 ;
wire _5530__bF$buf3 ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _5674_ ;
wire _5254_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf2  ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_31_bF$buf2  ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire rst_bF$buf30 ;
wire rst_bF$buf31 ;
wire rst_bF$buf32 ;
wire rst_bF$buf33 ;
wire rst_bF$buf34 ;
wire rst_bF$buf35 ;
wire rst_bF$buf36 ;
wire rst_bF$buf37 ;
wire rst_bF$buf38 ;
wire rst_bF$buf39 ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _2462__bF$buf0 ;
wire _2462__bF$buf1 ;
wire _2462__bF$buf2 ;
wire _2462__bF$buf3 ;
wire _6497_ ;
wire _6077_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _1688_ ;
wire _1268_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf2  ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf0  ;
wire _4657_ ;
wire _4237_ ;
wire _6803_ ;
wire _5545__bF$buf0 ;
wire _5545__bF$buf1 ;
wire _5545__bF$buf2 ;
wire _5545__bF$buf3 ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire [31:0] _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6421_ ;
wire _6001_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf3  ;
wire _1612_ ;
wire _4084_ ;
wire _943_ ;
wire [31:0] _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf2  ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire [31:0] _68_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf6  ;
wire [31:0] \datapath_1.Data  ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire [31:0] \datapath_1.regfile_1.regOut[20]  ;
wire _5466__bF$buf0 ;
wire _5466__bF$buf1 ;
wire _5466__bF$buf2 ;
wire _5466__bF$buf3 ;
wire _5466__bF$buf4 ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6553_ ;
wire _6133_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf2  ;
wire _3678_ ;
wire _3258_ ;
wire _5824_ ;
wire _5404_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf0  ;
wire _5633_ ;
wire _5213_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _2091_ ;
wire _3296_ ;
wire _1609_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf1  ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _5918_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf5  ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6456_ ;
wire _6036_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf2  ;
wire _1591_ ;
wire _1171_ ;
wire _3977__bF$buf0 ;
wire _3977__bF$buf1 ;
wire _3977__bF$buf2 ;
wire _3977__bF$buf3 ;
wire _3977__bF$buf4 ;
wire _2796_ ;
wire _2376_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf5  ;
wire _5727_ ;
wire _5307_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf3  ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire [31:0] _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _2185_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire MemRead ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _3199_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire \datapath_1.PCJump_17_bF$buf4  ;
wire _4616_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _3200__bF$buf0 ;
wire _3200__bF$buf1 ;
wire \datapath_1.regfile_1.regEn_7_bF$buf6  ;
wire _3200__bF$buf2 ;
wire _3200__bF$buf3 ;
wire _3200__bF$buf4 ;
wire _2699_ ;
wire _2279_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire clk_hier0_bF$buf0 ;
wire clk_hier0_bF$buf1 ;
wire clk_hier0_bF$buf2 ;
wire clk_hier0_bF$buf3 ;
wire clk_hier0_bF$buf4 ;
wire clk_hier0_bF$buf5 ;
wire clk_hier0_bF$buf6 ;
wire clk_hier0_bF$buf7 ;
wire clk_hier0_bF$buf8 ;
wire clk_hier0_bF$buf9 ;
wire _2088_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf4  ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _1800_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _27_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf0  ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire clk_bF$buf110 ;
wire clk_bF$buf111 ;
wire clk_bF$buf112 ;
wire clk_bF$buf113 ;
wire _5548__bF$buf0 ;
wire _5548__bF$buf1 ;
wire _5548__bF$buf2 ;
wire _5548__bF$buf3 ;
wire _5548__bF$buf4 ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _6703_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _3828_ ;
wire _3408_ ;
wire _5552__bF$buf0 ;
wire _5552__bF$buf1 ;
wire _5552__bF$buf2 ;
wire _5552__bF$buf3 ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6512_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf3  ;
wire _3637_ ;
wire _3217_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf3  ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6550_ ;
wire _6130_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf2  ;
wire _5821_ ;
wire _5401_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf6  ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _4901_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _5469__bF$buf0 ;
wire _5469__bF$buf1 ;
wire _5469__bF$buf2 ;
wire _5469__bF$buf3 ;
wire _690_ ;
wire _270_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _5915_ ;
wire [31:0] \datapath_1.regfile_1.regOut[10]  ;
wire \datapath_1.regfile_1.regEn_18_bF$buf2  ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6453_ ;
wire _6033_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf2  ;
wire _5724_ ;
wire _5304_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf0  ;
wire _6509_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf7  ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _3196_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _4005__bF$buf0 ;
wire _2047_ ;
wire _4005__bF$buf1 ;
wire _4005__bF$buf2 ;
wire _4005__bF$buf3 ;
wire \datapath_1.PCJump_17_bF$buf1  ;
wire _4613_ ;
wire [31:0] \datapath_1.regfile_1.regOut[4]  ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf5  ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf3  ;
wire _2696_ ;
wire _2276_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire [31:0] _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf4  ;
wire _4707_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf1  ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire [31:0] \datapath_1.regfile_1.regOut[27]  ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf4  ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf0  ;
wire _399_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _1700_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf0  ;
wire _1297_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _6603_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf3  ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire MemToReg ;
wire _6641_ ;
wire _6221_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _1832_ ;
wire _1412_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf2  ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6450_ ;
wire _6030_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf6  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf2  ;
wire _59_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf6  ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf4  ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _3193_ ;
wire [31:0] \datapath_1.rd1  ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _5815_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf2  ;
wire _6773_ ;
wire _6353_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf0  ;
wire _2693_ ;
wire _2273_ ;
wire _5480__bF$buf0 ;
wire _5480__bF$buf1 ;
wire _5480__bF$buf2 ;
wire _5480__bF$buf3 ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _4079__bF$buf0 ;
wire _4079__bF$buf1 ;
wire _4079__bF$buf2 ;
wire _4079__bF$buf3 ;
wire _5624_ ;
wire _5204_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire [5:0] \aluControl_1.inst  ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf7  ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf1  ;
wire _4704_ ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf5  ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire PCEn_bF$buf0 ;
wire PCEn_bF$buf1 ;
wire PCEn_bF$buf2 ;
wire PCEn_bF$buf3 ;
wire PCEn_bF$buf4 ;
wire PCEn_bF$buf5 ;
wire PCEn_bF$buf6 ;
wire PCEn_bF$buf7 ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _5539__bF$buf0 ;
wire _5539__bF$buf1 ;
wire _5539__bF$buf2 ;
wire _5539__bF$buf3 ;
wire _5539__bF$buf4 ;
wire _6485_ ;
wire _6065_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf1  ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire [31:0] \datapath_1.regfile_1.regOut[17]  ;
wire \datapath_1.PCJump_27_bF$buf4  ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf4  ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_11_bF$buf3  ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _299_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf7  ;
wire _3198__bF$buf0 ;
wire _3198__bF$buf1 ;
wire _3198__bF$buf2 ;
wire _3198__bF$buf3 ;
wire _3198__bF$buf4 ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _3935__bF$buf0 ;
wire _3935__bF$buf1 ;
wire _3935__bF$buf2 ;
wire _3935__bF$buf3 ;
wire _4777_ ;
wire _3935__bF$buf4 ;
wire _4357_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf3  ;
wire _56_ ;
wire _6503_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf3  ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf1  ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6541_ ;
wire _6121_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf2  ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire [31:0] \datapath_1.alu_1.ALUInB  ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf6  ;
wire _6350_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf2  ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _5621_ ;
wire _5201_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_5_bF$buf4  ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire [3:0] \control_1.reg_state.dout  ;
wire _4701_ ;
wire _5906_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf2  ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _5483__bF$buf0 ;
wire _5483__bF$buf1 ;
wire _5483__bF$buf2 ;
wire _5483__bF$buf3 ;
wire _5483__bF$buf4 ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire \datapath_1.PCJump_27_bF$buf1  ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire [31:0] _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf1  ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf0  ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _296_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf4  ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _2399_ ;
wire _3760_ ;
wire _3340_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf4  ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _4774_ ;
wire _4354_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf0  ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6500_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf3  ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _4583_ ;
wire _4163_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf0  ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf7  ;
wire _1288_ ;
wire _199_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf3  ;
wire _3719_ ;
wire _5565__bF$buf0 ;
wire _5565__bF$buf1 ;
wire _5565__bF$buf2 ;
wire _5565__bF$buf3 ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _6823_ ;
wire _6403_ ;
wire _3942__bF$buf0 ;
wire _3942__bF$buf1 ;
wire _3942__bF$buf2 ;
wire _3942__bF$buf3 ;
wire _2743_ ;
wire _2323_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf3  ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf1  ;
wire _9_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _5903_ ;
wire _3090_ ;
wire [31:0] _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire ALUOp_0_bF$buf0 ;
wire ALUOp_0_bF$buf1 ;
wire ALUOp_0_bF$buf2 ;
wire ALUOp_0_bF$buf3 ;
wire ALUOp_0_bF$buf4 ;
wire _2608_ ;
wire ALUOp_0_bF$buf5 ;
wire _6441_ ;
wire _6021_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf2  ;
wire _5712_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _2590_ ;
wire _2170_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf6  ;
wire _3795_ ;
wire _3375_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf2  ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire \datapath_1.PCJump_22_bF$buf2  ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf6  ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _5806_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf2  ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _3201__bF$buf0 ;
wire _3201__bF$buf1 ;
wire _3201__bF$buf2 ;
wire \datapath_1.regfile_1.regEn_8_bF$buf6  ;
wire _3201__bF$buf3 ;
wire _3201__bF$buf4 ;
wire _5615_ ;
wire [31:0] \datapath_1.regfile_1.regOut[22]  ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _6573_ ;
wire _6153_ ;
wire _2493_ ;
wire _2073_ ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _2470__bF$buf0 ;
wire _2470__bF$buf1 ;
wire _2470__bF$buf2 ;
wire _2470__bF$buf3 ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _5709_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _4733_ ;
wire _4313_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf1  ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf1  ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5549__bF$buf0 ;
wire _5549__bF$buf1 ;
wire _5549__bF$buf2 ;
wire _5747_ ;
wire _5549__bF$buf3 ;
wire _5327_ ;
wire _5549__bF$buf4 ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf0  ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf4  ;
wire _1285_ ;
wire _196_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _3882__bF$buf0 ;
wire _3882__bF$buf1 ;
wire _3882__bF$buf2 ;
wire _3882__bF$buf3 ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _2299_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _2931_ ;
wire _2511_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf0  ;
wire _3716_ ;
wire _6188_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf3  ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf0  ;
wire \datapath_1.regfile_1.regEn_17_bF$buf7  ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf3  ;
wire _6_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf7  ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _1820_ ;
wire _1400_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf3  ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _2643_ ;
wire _2223_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf7  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf3  ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6532_ ;
wire _6112_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _5803_ ;
wire _1723_ ;
wire [31:0] _1303_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf2  ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _2681_ ;
wire _2261_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf3  ;
wire _5612_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf6  ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6570_ ;
wire _6150_ ;
wire _2490_ ;
wire _2070_ ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire rst_bF$buf100 ;
wire rst_bF$buf101 ;
wire rst_bF$buf102 ;
wire rst_bF$buf103 ;
wire rst_bF$buf104 ;
wire rst_bF$buf105 ;
wire rst_bF$buf106 ;
wire rst_bF$buf107 ;
wire rst_bF$buf108 ;
wire rst_bF$buf109 ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _5489__bF$buf0 ;
wire _5489__bF$buf1 ;
wire _5489__bF$buf2 ;
wire _5489__bF$buf3 ;
wire _4921_ ;
wire _4501_ ;
wire _5706_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire rst ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire [31:0] \datapath_1.regfile_1.regOut[12]  ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6473_ ;
wire _6053_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf4  ;
wire MemWrite ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire clk_bF$buf70 ;
wire clk_bF$buf71 ;
wire clk_bF$buf72 ;
wire clk_bF$buf73 ;
wire clk_bF$buf74 ;
wire clk_bF$buf75 ;
wire clk_bF$buf76 ;
wire clk_bF$buf77 ;
wire clk_bF$buf78 ;
wire clk_bF$buf79 ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _5609_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf1  ;
wire _6567_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf4  ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _4633_ ;
wire _4213_ ;
wire [31:0] \datapath_1.regfile_1.regOut[6]  ;
wire _5838_ ;
wire _5418_ ;
wire [31:0] _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf0  ;
wire _4918_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf4  ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf0  ;
wire [31:0] _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire [31:0] \datapath_1.regfile_1.regOut[29]  ;
wire _1185_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf4  ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _2199_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_24_bF$buf3  ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _3845_ ;
wire [31:0] _3425_ ;
wire _3005_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf4  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf0  ;
wire \datapath_1.regfile_1.regEn_24_bF$buf7  ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _1720_ ;
wire _1300_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf0  ;
wire _4668_ ;
wire _4248_ ;
wire [4:0] \datapath_1.a3  ;
wire \datapath_1.regfile_1.regEn_29_bF$buf3  ;
wire _6814_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf7  ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _5504__bF$buf0 ;
wire _5504__bF$buf1 ;
wire _5504__bF$buf2 ;
wire _5504__bF$buf3 ;
wire _5504__bF$buf4 ;
wire _6432_ ;
wire _6012_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _5703_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6470_ ;
wire _6050_ ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf1  ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire clk_bF$buf40 ;
wire clk_bF$buf41 ;
wire clk_bF$buf42 ;
wire clk_bF$buf43 ;
wire clk_bF$buf44 ;
wire clk_bF$buf45 ;
wire clk_bF$buf46 ;
wire clk_bF$buf47 ;
wire clk_bF$buf48 ;
wire clk_bF$buf49 ;
wire _4821_ ;
wire _4401_ ;
wire _5606_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6564_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf1  ;
wire _6144_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _2293_ ;
wire _3971__bF$buf0 ;
wire _3971__bF$buf1 ;
wire _3971__bF$buf2 ;
wire _3971__bF$buf3 ;
wire _3971__bF$buf4 ;
wire _3498_ ;
wire _3078_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf4  ;
wire _5644_ ;
wire _5224_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf1  ;
wire _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf7  ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf1  ;
wire _2387_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _1658_ ;
wire [31:0] _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire \datapath_1.mux_wd3.dout_24_bF$buf0  ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf1  ;
wire _4627_ ;
wire _4207_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf4  ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire [31:0] \datapath_1.regfile_1.regOut[19]  ;
wire _1085_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _2099_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf0  ;
wire _6811_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf3  ;
wire _2731_ ;
wire _2311_ ;
wire _3936_ ;
wire _3516_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf4  ;
wire [31:0] _913_ ;
wire _5679_ ;
wire _5259_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf7  ;
wire _6620_ ;
wire _6200_ ;
wire \datapath_1.mux_wd3.dout_31_bF$buf3  ;
wire _1599_ ;
wire _1179_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire _1811_ ;
wire _4051__bF$buf0 ;
wire _4051__bF$buf1 ;
wire _4283_ ;
wire _4051__bF$buf2 ;
wire _4051__bF$buf3 ;
wire _722_ ;
wire _302_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf7  ;
wire _5488_ ;
wire _5068_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire rst_bF$buf80 ;
wire rst_bF$buf81 ;
wire rst_bF$buf82 ;
wire rst_bF$buf83 ;
wire rst_bF$buf84 ;
wire rst_bF$buf85 ;
wire rst_bF$buf86 ;
wire rst_bF$buf87 ;
wire rst_bF$buf88 ;
wire rst_bF$buf89 ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _6714_ ;
wire _3955__bF$buf0 ;
wire _3955__bF$buf1 ;
wire _3955__bF$buf2 ;
wire _3955__bF$buf3 ;
wire _3955__bF$buf4 ;
wire _760_ ;
wire _340_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf7  ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6523_ ;
wire _6103_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _2672_ ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire clk_bF$buf11 ;
wire clk_bF$buf12 ;
wire clk_bF$buf13 ;
wire clk_bF$buf14 ;
wire clk_bF$buf15 ;
wire clk_bF$buf16 ;
wire clk_bF$buf17 ;
wire clk_bF$buf18 ;
wire clk_bF$buf19 ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _5603_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6561_ ;
wire _6141_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf1  ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _4912_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _5499__bF$buf0 ;
wire _5499__bF$buf1 ;
wire _6655_ ;
wire _5499__bF$buf2 ;
wire _6235_ ;
wire _5499__bF$buf3 ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _4721_ ;
wire _4301_ ;
wire _5926_ ;
wire _5506_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf4  ;
wire _6464_ ;
wire _6044_ ;
wire _2384_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _2193_ ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf3  ;
wire _4815_ ;
wire _5773_ ;
wire _5353_ ;
wire _6558_ ;
wire _6138_ ;
wire [31:0] _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf7  ;
wire _4624_ ;
wire _4204_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf1  ;
wire _5829_ ;
wire _5409_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf4  ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf5  ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf0  ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf1  ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf4  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf0  ;
wire _1596_ ;
wire _1176_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _4280_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf4  ;
wire _5485_ ;
wire _5065_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire rst_bF$buf50 ;
wire rst_bF$buf51 ;
wire rst_bF$buf52 ;
wire rst_bF$buf53 ;
wire rst_bF$buf54 ;
wire rst_bF$buf55 ;
wire rst_bF$buf56 ;
wire rst_bF$buf57 ;
wire rst_bF$buf58 ;
wire rst_bF$buf59 ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _3780_ ;
wire [31:0] _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf4  ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _1711_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf2  ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _660_ ;
wire _240_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6423_ ;
wire _6003_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _5923_ ;
wire _5503_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf1  ;
wire _2628_ ;
wire _2208_ ;
wire _6461_ ;
wire _6041_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf4  ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _2190_ ;
wire [31:0] \datapath_1.regfile_1.regOut[1]  ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf0  ;
wire _4812_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire [31:0] _848_ ;
wire _428_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf4  ;
wire _4621_ ;
wire _4201_ ;
wire _5826_ ;
wire _5406_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf1  ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6784_ ;
wire _6364_ ;
wire _2284_ ;
wire _3489_ ;
wire _3069_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf2  ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire [31:0] \datapath_1.regfile_1.regOut[24]  ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _2093_ ;
wire _3298_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf3  ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _4038__bF$buf0 ;
wire _4038__bF$buf1 ;
wire _4038__bF$buf2 ;
wire _4038__bF$buf3 ;
wire \datapath_1.regfile_1.regEn_18_bF$buf7  ;
wire _5673_ ;
wire _5253_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf1  ;
wire _6458_ ;
wire _6038_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf4  ;
wire _1593_ ;
wire [31:0] _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf7  ;
wire _5729_ ;
wire _5309_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf5  ;
wire _1649_ ;
wire _1229_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf1  ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire rst_bF$buf20 ;
wire rst_bF$buf21 ;
wire rst_bF$buf22 ;
wire rst_bF$buf23 ;
wire rst_bF$buf24 ;
wire rst_bF$buf25 ;
wire rst_bF$buf26 ;
wire rst_bF$buf27 ;
wire rst_bF$buf28 ;
wire rst_bF$buf29 ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _4809_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire [31:0] \datapath_1.mux_wd3.dout  ;
wire _1687_ ;
wire _1267_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf1  ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire _1802_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _29_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf2  ;
wire _1611_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf1  ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf5  ;
wire _3639_ ;
wire _3219_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _1934_ ;
wire _1514_ ;
wire _5521__bF$buf0 ;
wire _5521__bF$buf1 ;
wire _5521__bF$buf2 ;
wire _5521__bF$buf3 ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6552_ ;
wire _6132_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf1  ;
wire _3677_ ;
wire _3257_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf4  ;
wire _5823_ ;
wire _5403_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _2090_ ;
wire _3295_ ;
wire _1608_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf0  ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _5917_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf4  ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire [31:0] _328_ ;
wire _6455_ ;
wire _6035_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf1  ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf4  ;
wire _5726_ ;
wire _5306_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf2  ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _2184_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire [31:0] \datapath_1.regfile_1.regOut[14]  ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _3198_ ;
wire _5764_ ;
wire _5344_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire \datapath_1.PCJump_17_bF$buf3  ;
wire _4615_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf7  ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf5  ;
wire _2698_ ;
wire _2278_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire _4653_ ;
wire [31:0] memoryWriteData ;
wire _4233_ ;
wire [31:0] \datapath_1.regfile_1.regOut[8]  ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf3  ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire clk_bF$buf100 ;
wire clk_bF$buf101 ;
wire clk_bF$buf102 ;
wire clk_bF$buf103 ;
wire clk_bF$buf104 ;
wire clk_bF$buf105 ;
wire clk_bF$buf106 ;
wire clk_bF$buf107 ;
wire clk_bF$buf108 ;
wire clk_bF$buf109 ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6511_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf2  ;
wire _3636_ ;
wire _3216_ ;
wire _1702_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf2  ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _3674_ ;
wire _3254_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf1  ;
wire ALUSrcA ;
wire [1:0] ALUSrcB ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf5  ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _3972__bF$buf0 ;
wire _3972__bF$buf1 ;
wire _3972__bF$buf2 ;
wire _3972__bF$buf3 ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _5524__bF$buf0 ;
wire _5524__bF$buf1 ;
wire _5524__bF$buf2 ;
wire _5524__bF$buf3 ;
wire _3768_ ;
wire _3348_ ;
wire _5914_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf1  ;
wire _1834_ ;
wire _1414_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf4  ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6452_ ;
wire _6032_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf1  ;
wire _5723_ ;
wire _5303_ ;
wire \datapath_1.mux_wd3.dout_20_bF$buf4  ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf6  ;
wire PCSource_1_bF$buf0 ;
wire _1032_ ;
wire PCSource_1_bF$buf1 ;
wire PCSource_1_bF$buf2 ;
wire PCSource_1_bF$buf3 ;
wire PCSource_1_bF$buf4 ;
wire [31:0] _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _3195_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire \datapath_1.PCJump_17_bF$buf0  ;
wire _4612_ ;
wire _5817_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf4  ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf2  ;
wire _2695_ ;
wire _2275_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _3893__bF$buf0 ;
wire _3893__bF$buf1 ;
wire _3893__bF$buf2 ;
wire _3893__bF$buf3 ;
wire _5626_ ;
wire _5206_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _2084_ ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf3  ;
wire _4706_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf0  ;
wire _3098_ ;
wire _5664_ ;
wire _5244_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf7  ;
wire _4935_ ;
wire _4515_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf3  ;
wire _1678_ ;
wire _1258_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire BranchNe ;
wire _1296_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf2  ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire ALUZero ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _1831_ ;
wire _1411_ ;
wire \datapath_1.mux_wd3.dout_16_bF$buf1  ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf1  ;
wire _58_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf5  ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf3  ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _5527__bF$buf0 ;
wire _5527__bF$buf1 ;
wire _5527__bF$buf2 ;
wire _5527__bF$buf3 ;
wire _5527__bF$buf4 ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6543_ ;
wire _6123_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf4  ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _5531__bF$buf0 ;
wire _5531__bF$buf1 ;
wire _5531__bF$buf2 ;
wire _5531__bF$buf3 ;
wire _5531__bF$buf4 ;
wire _5814_ ;
wire _1734_ ;
wire _1314_ ;
wire [31:0] \datapath_1.a  ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf1  ;
wire _6772_ ;
wire _6352_ ;
wire \datapath_1.mux_wd3.dout_23_bF$buf4  ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf6  ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire [31:0] _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf0  ;
wire _4703_ ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf4  ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire \datapath_1.mux_wd3.dout_3_bF$buf0  ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire \datapath_1.PCJump_27_bF$buf3  ;
wire [31:0] _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf3  ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire \datapath_1.mux_wd3.dout_11_bF$buf2  ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _298_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf6  ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire [31:0] ALUOut ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _3036__bF$buf0 ;
wire _3036__bF$buf1 ;
wire _3036__bF$buf2 ;
wire _3036__bF$buf3 ;
wire _3036__bF$buf4 ;
wire \datapath_1.regfile_1.regEn_16_bF$buf2  ;
wire _55_ ;
wire _6502_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _5471__bF$buf0 ;
wire _5471__bF$buf1 ;
wire _5471__bF$buf2 ;
wire _5471__bF$buf3 ;
wire _5471__bF$buf4 ;
wire _5471__bF$buf5 ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf2  ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf0  ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire \datapath_1.mux_wd3.dout_19_bF$buf1  ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire [31:0] \datapath_1.alu_1.ALUInA  ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf5  ;
wire \datapath_1.mux_wd3.dout_23_bF$buf1  ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf5  ;
wire \datapath_1.regfile_1.regEn_5_bF$buf3  ;
wire ALUSrcB_1_bF$buf0 ;
wire ALUSrcB_1_bF$buf1 ;
wire ALUSrcB_1_bF$buf2 ;
wire ALUSrcB_1_bF$buf3 ;
wire ALUSrcB_1_bF$buf4 ;
wire _3283_ ;
wire _3982__bF$buf0 ;
wire _3982__bF$buf1 ;
wire _3982__bF$buf2 ;
wire _3982__bF$buf3 ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _5905_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _5534__bF$buf0 ;
wire _5534__bF$buf1 ;
wire _5534__bF$buf2 ;
wire _5534__bF$buf3 ;
wire _5534__bF$buf4 ;
wire _736_ ;
wire _316_ ;
wire _6443_ ;
wire _6023_ ;
wire _2783_ ;
wire _2363_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf1  ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf4  ;
wire _5714_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf4  ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire [31:0] \datapath_1.regfile_1.regOut[3]  ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire \datapath_1.PCJump_27_bF$buf0  ;
wire \datapath_1.mux_wd3.dout_1_bF$buf4  ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire [1:0] PCSource ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _3997__bF$buf0 ;
wire _3997__bF$buf1 ;
wire _3997__bF$buf2 ;
wire _3997__bF$buf3 ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire \datapath_1.mux_wd3.dout_6_bF$buf0  ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire [3:0] ALUControl ;
wire _5655_ ;
wire _5235_ ;
wire [31:0] \datapath_1.regfile_1.regOut[26]  ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _3930__bF$buf0 ;
wire _3930__bF$buf1 ;
wire _3930__bF$buf2 ;
wire _3930__bF$buf3 ;
wire _4735_ ;
wire _4315_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf3  ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf3  ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire \datapath_1.mux_wd3.dout_14_bF$buf2  ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf6  ;
wire _1287_ ;
wire [31:0] _198_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _2933_ ;
wire _2513_ ;
wire \datapath_1.regfile_1.regEn_19_bF$buf2  ;
wire _3718_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _2742_ ;
wire _2322_ ;
wire \datapath_1.regfile_1.regEn_23_bF$buf2  ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire \datapath_1.regfile_1.regEn_5_bF$buf0  ;
wire _8_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _1822_ ;
wire _1402_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6440_ ;
wire _6020_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire \datapath_1.mux_wd3.dout_26_bF$buf1  ;
wire _5711_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf5  ;
wire _3794_ ;
wire _3374_ ;
wire \datapath_1.mux_wd3.dout_30_bF$buf1  ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire \datapath_1.PCJump_22_bF$buf1  ;
wire MemToReg_bF$buf0 ;
wire MemToReg_bF$buf1 ;
wire MemToReg_bF$buf2 ;
wire MemToReg_bF$buf3 ;
wire MemToReg_bF$buf4 ;
wire MemToReg_bF$buf5 ;
wire MemToReg_bF$buf6 ;
wire MemToReg_bF$buf7 ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire \datapath_1.regfile_1.regEn_30_bF$buf5  ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6534_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _5805_ ;
wire _1725_ ;
wire _1305_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf4  ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire \datapath_1.mux_wd3.dout_1_bF$buf1  ;
wire _6763_ ;
wire _6343_ ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf5  ;
wire _5614_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6572_ ;
wire _6152_ ;
wire _2492_ ;
wire _2072_ ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _5708_ ;
wire [31:0] _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _4732_ ;
wire _4312_ ;
wire \datapath_1.regfile_1.regEn_11_bF$buf0  ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire \datapath_1.mux_wd3.dout_9_bF$buf0  ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _3196__bF$buf0 ;
wire _5326_ ;
wire _3196__bF$buf1 ;
wire _3196__bF$buf2 ;
wire _3196__bF$buf3 ;
wire _3196__bF$buf4 ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire [31:0] \datapath_1.regfile_1.regOut[16]  ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire clk_bF$buf90 ;
wire clk_bF$buf91 ;
wire clk_bF$buf92 ;
wire clk_bF$buf93 ;
wire clk_bF$buf94 ;
wire clk_bF$buf95 ;
wire clk_bF$buf96 ;
wire _3621_ ;
wire clk_bF$buf97 ;
wire _3201_ ;
wire clk_bF$buf98 ;
wire clk_bF$buf99 ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _5784_ ;
wire _5364_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf3  ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire \datapath_1.mux_wd3.dout_17_bF$buf2  ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf6  ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire \datapath_1.mux_wd3.dout_21_bF$buf2  ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf6  ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _46_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire \datapath_1.regfile_1.regEn_26_bF$buf2  ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _2642_ ;
wire _2222_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf6  ;
wire \datapath_1.regfile_1.regEn_30_bF$buf2  ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6531_ ;
wire _6111_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _1722_ ;
wire _1302_ ;
wire \datapath_1.mux_wd3.dout_29_bF$buf1  ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _2680_ ;
wire _2260_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire \datapath_1.regfile_1.regEn_8_bF$buf2  ;
wire _5611_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf5  ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6434_ ;
wire _6014_ ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _5544__bF$buf0 ;
wire _5544__bF$buf1 ;
wire _5544__bF$buf2 ;
wire _5544__bF$buf3 ;
wire _5705_ ;
wire [31:0] \datapath_1.regfile_1.regOut[31]  ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6472_ ;
wire _6052_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf3  ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire clk_bF$buf60 ;
wire clk_bF$buf61 ;
wire clk_bF$buf62 ;
wire clk_bF$buf63 ;
wire clk_bF$buf64 ;
wire clk_bF$buf65 ;
wire clk_bF$buf66 ;
wire clk_bF$buf67 ;
wire clk_bF$buf68 ;
wire clk_bF$buf69 ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _5608_ ;
wire _1948_ ;
wire _1528_ ;
wire [31:0] _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire \datapath_1.regfile_1.regEn_14_bF$buf0  ;
wire _859_ ;
wire _439_ ;
wire _6566_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf3  ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire IRWrite ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire _4670_ ;
wire _4250_ ;
wire _3034__bF$buf0 ;
wire _3034__bF$buf1 ;
wire _3034__bF$buf2 ;
wire _3034__bF$buf3 ;
wire _3034__bF$buf4 ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _3936__bF$buf0 ;
wire _3936__bF$buf1 ;
wire _3936__bF$buf2 ;
wire _3936__bF$buf3 ;
wire _3936__bF$buf4 ;
wire _286_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf3  ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire [31:0] _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _5684_ ;
wire _5264_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf3  ;
wire _2389_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire rst_hier0_bF$buf0 ;
wire rst_hier0_bF$buf1 ;
wire rst_hier0_bF$buf2 ;
wire rst_hier0_bF$buf3 ;
wire rst_hier0_bF$buf4 ;
wire rst_hier0_bF$buf5 ;
wire rst_hier0_bF$buf6 ;
wire rst_hier0_bF$buf7 ;
wire rst_hier0_bF$buf8 ;
wire rst_hier0_bF$buf9 ;
wire _4001__bF$buf0 ;
wire _4001__bF$buf1 ;
wire _4001__bF$buf2 ;
wire _4001__bF$buf3 ;
wire \datapath_1.mux_wd3.dout_24_bF$buf2  ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf3  ;
wire _4629_ ;
wire _4209_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf6  ;
wire ALUSrcB_0_bF$buf0 ;
wire ALUSrcB_0_bF$buf1 ;
wire ALUSrcB_0_bF$buf2 ;
wire ALUSrcB_0_bF$buf3 ;
wire ALUSrcB_0_bF$buf4 ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire \datapath_1.regfile_1.regEn_29_bF$buf2  ;
wire _6813_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf6  ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _3080_ ;
wire [3:0] \control_1.next  ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6431_ ;
wire _6011_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire _953_ ;
wire ALUSrcA_bF$buf0 ;
wire _533_ ;
wire ALUSrcA_bF$buf1 ;
wire _113_ ;
wire ALUSrcA_bF$buf2 ;
wire ALUSrcA_bF$buf3 ;
wire ALUSrcA_bF$buf4 ;
wire ALUSrcA_bF$buf5 ;
wire ALUSrcA_bF$buf6 ;
wire _2827_ ;
wire ALUSrcA_bF$buf7 ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _3594_ ;
wire _3174_ ;
wire _3995__bF$buf0 ;
wire _3995__bF$buf1 ;
wire _3995__bF$buf2 ;
wire _3995__bF$buf3 ;
wire _3995__bF$buf4 ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire \datapath_1.mux_wd3.dout_4_bF$buf0  ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire clk_bF$buf30 ;
wire clk_bF$buf31 ;
wire clk_bF$buf32 ;
wire clk_bF$buf33 ;
wire clk_bF$buf34 ;
wire clk_bF$buf35 ;
wire clk_bF$buf36 ;
wire clk_bF$buf37 ;
wire clk_bF$buf38 ;
wire clk_bF$buf39 ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _3924__bF$buf0 ;
wire _3924__bF$buf1 ;
wire _3924__bF$buf2 ;
wire _3924__bF$buf3 ;
wire _5605_ ;
wire [31:0] \datapath_1.regfile_1.regOut[21]  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6563_ ;
wire \datapath_1.mux_wd3.dout_12_bF$buf0  ;
wire _6143_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf3  ;
wire _5643_ ;
wire _5223_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire [31:0] _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire \datapath_1.regfile_1.regEn_17_bF$buf0  ;
wire _4723_ ;
wire _4303_ ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf6  ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire \datapath_1.regfile_1.regEn_21_bF$buf0  ;
wire _2386_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3037__bF$buf0 ;
wire _3037__bF$buf1 ;
wire _3037__bF$buf2 ;
wire _3037__bF$buf3 ;
wire _3037__bF$buf4 ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _5472__bF$buf0 ;
wire _5472__bF$buf1 ;
wire _5472__bF$buf2 ;
wire _5472__bF$buf3 ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire \datapath_1.regfile_1.regEn_3_bF$buf0  ;
wire _4626_ ;
wire _4206_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf3  ;
wire _5570__bF$buf0 ;
wire _5570__bF$buf1 ;
wire _5570__bF$buf2 ;
wire _5570__bF$buf3 ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _2289_ ;
wire _3650_ ;
wire _3230_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf7  ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire [3:0] _2098_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire \datapath_1.mux_wd3.dout_27_bF$buf2  ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf3  ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf6  ;
wire \datapath_1.mux_wd3.dout_31_bF$buf2  ;
wire _1598_ ;
wire _1178_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _1810_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf6  ;
wire _5487_ ;
wire _5067_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire rst_bF$buf70 ;
wire rst_bF$buf71 ;
wire rst_bF$buf72 ;
wire rst_bF$buf73 ;
wire rst_bF$buf74 ;
wire rst_bF$buf75 ;
wire rst_bF$buf76 ;
wire rst_bF$buf77 ;
wire rst_bF$buf78 ;
wire rst_bF$buf79 ;
wire [31:0] \datapath_1.regfile_1.regEn  ;
wire _4758_ ;
wire _4338_ ;
wire _37_ ;
wire _4091_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf6  ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6522_ ;
wire _6102_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6751_ ;
wire _6331_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf4  ;
wire _5602_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6560_ ;
wire _6140_ ;
wire _2480_ ;
wire _2060_ ;
wire [31:0] _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _3998__bF$buf0 ;
wire _3998__bF$buf1 ;
wire _3998__bF$buf2 ;
wire _3998__bF$buf3 ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _3494_ ;
wire _3074_ ;
wire \datapath_1.mux_wd3.dout_7_bF$buf0  ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire [31:0] _718_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _5925_ ;
wire _5505_ ;
wire [31:0] \datapath_1.regfile_1.regOut[11]  ;
wire _3931__bF$buf0 ;
wire _1845_ ;
wire _3931__bF$buf1 ;
wire _1425_ ;
wire _3931__bF$buf2 ;
wire _1005_ ;
wire _3931__bF$buf3 ;
wire _756_ ;
wire _336_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf3  ;
wire _6463_ ;
wire _6043_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _2192_ ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire [31:0] _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire \datapath_1.mux_wd3.dout_15_bF$buf2  ;
wire _4814_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf6  ;
wire _4623_ ;
wire _4203_ ;
wire \datapath_1.regfile_1.regEn_24_bF$buf0  ;
wire [31:0] \datapath_1.regfile_1.regOut[5]  ;
wire _5828_ ;
wire _5408_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf3  ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf4  ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire [31:0] \datapath_1.ALUResult  ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire \datapath_1.regfile_1.regEn_6_bF$buf0  ;
wire _5675_ ;
wire _5255_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf3  ;
wire [31:0] \datapath_1.regfile_1.regOut[28]  ;
wire _1595_ ;
wire _1175_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _3950__bF$buf0 ;
wire _3950__bF$buf1 ;
wire _3950__bF$buf2 ;
wire _3950__bF$buf3 ;
wire \datapath_1.regfile_1.regEn_4_bF$buf7  ;
wire \datapath_1.regfile_1.regEn_31_bF$buf3  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _2189_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire rst_bF$buf40 ;
wire rst_bF$buf41 ;
wire rst_bF$buf42 ;
wire rst_bF$buf43 ;
wire rst_bF$buf44 ;
wire rst_bF$buf45 ;
wire rst_bF$buf46 ;
wire rst_bF$buf47 ;
wire rst_bF$buf48 ;
wire rst_bF$buf49 ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _1689_ ;
wire _1269_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf3  ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire [31:0] _1498_ ;
wire _1078_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _1710_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire [31:0] memoryAddress ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire \datapath_1.mux_wd3.dout_2_bF$buf1  ;
wire _4658_ ;
wire _4238_ ;
wire _6804_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire PCEn ;
wire _906_ ;
wire _6613_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6422_ ;
wire _6002_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf4  ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire \datapath_1.regfile_1.regEn_12_bF$buf0  ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6460_ ;
wire _6040_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf3  ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf7  ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire [31:0] \datapath_1.PCJump  ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf3  ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _5825_ ;
wire _5405_ ;
wire \datapath_1.mux_wd3.dout_22_bF$buf0  ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire \datapath_1.regfile_1.regEn_1_bF$buf1  ;
wire _5634_ ;
wire _5214_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _2092_ ;
wire _3297_ ;
wire \datapath_1.mux_wd3.dout_18_bF$buf2  ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _5919_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf6  ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire \datapath_1.regfile_1.regEn_27_bF$buf0  ;
wire _6457_ ;
wire _6037_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf3  ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf6  ;
wire _5728_ ;
wire _5308_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf4  ;
wire _1648_ ;
wire _1228_ ;
wire \datapath_1.regfile_1.regEn_31_bF$buf0  ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire rst_bF$buf10 ;
wire rst_bF$buf11 ;
wire rst_bF$buf12 ;
wire rst_bF$buf13 ;
wire rst_bF$buf14 ;
wire rst_bF$buf15 ;
wire rst_bF$buf16 ;
wire rst_bF$buf17 ;
wire rst_bF$buf18 ;
wire rst_bF$buf19 ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _5478__bF$buf0 ;
wire _5478__bF$buf1 ;
wire _5478__bF$buf2 ;
wire _5478__bF$buf3 ;
wire _4808_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire \datapath_1.regfile_1.regEn_9_bF$buf0  ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire [31:0] \datapath_1.regfile_1.regOut[18]  ;
wire _1495_ ;
wire _1075_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf7  ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _2089_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _1589_ ;
wire _1169_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire _1801_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _28_ ;
wire \datapath_1.mux_wd3.dout_5_bF$buf1  ;
wire _1610_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire [31:0] \datapath_1.mux_iord.din0  ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _6704_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire \datapath_1.mux_wd3.dout_10_bF$buf0  ;
wire _3829_ ;
wire _3409_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6513_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf4  ;
wire _3638_ ;
wire _3218_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf4  ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _2481__bF$buf0 ;
wire _2481__bF$buf1 ;
wire _2481__bF$buf2 ;
wire _6551_ ;
wire _2481__bF$buf3 ;
wire _6131_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire \datapath_1.regfile_1.regEn_15_bF$buf0  ;
wire _3676_ ;
wire _3256_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf3  ;
wire _5822_ ;
wire _5402_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire [31:0] _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _2280_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf7  ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _3294_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _5916_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf3  ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6454_ ;
wire _6034_ ;
wire \datapath_1.mux_wd3.dout_25_bF$buf0  ;
wire _2794_ ;
wire _2374_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf3  ;
wire _5725_ ;
wire _5305_ ;
wire \datapath_1.regfile_1.regEn_4_bF$buf1  ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire _3197_ ;
wire _5763_ ;
wire _5343_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire \datapath_1.PCJump_17_bF$buf2  ;
wire _4614_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf6  ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf4  ;
wire _2697_ ;
wire _2277_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire \datapath_1.mux_wd3.dout_0_bF$buf2  ;
wire _5485__bF$buf0 ;
wire _5485__bF$buf1 ;
wire _5485__bF$buf2 ;
wire _5485__bF$buf3 ;
wire _5485__bF$buf4 ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire \datapath_1.regfile_1.regEn_10_bF$buf1  ;
wire _3635_ ;
wire _3215_ ;
wire _1701_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire \datapath_1.mux_wd3.dout_8_bF$buf1  ;
wire _1298_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _3673_ ;
wire _3253_ ;
wire \datapath_1.mux_wd3.dout_13_bF$buf0  ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _6604_ ;
wire _650_ ;
wire _230_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire \datapath_1.regfile_1.regEn_13_bF$buf4  ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _5913_ ;
wire \datapath_1.regfile_1.regEn_18_bF$buf0  ;
wire _1833_ ;
wire _1413_ ;
wire IorD_bF$buf0 ;
wire IorD_bF$buf1 ;
wire IorD_bF$buf2 ;
wire IorD_bF$buf3 ;
wire IorD_bF$buf4 ;
wire \datapath_1.mux_wd3.dout_16_bF$buf3  ;
wire IorD_bF$buf5 ;
wire IorD_bF$buf6 ;
wire IorD_bF$buf7 ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6451_ ;
wire _6031_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire \datapath_1.regfile_1.regEn_22_bF$buf0  ;
wire _5722_ ;
wire _5302_ ;
wire \datapath_1.regfile_1.regEn_16_bF$buf7  ;
wire \datapath_1.mux_wd3.dout_20_bF$buf3  ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire [31:0] _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _2180_ ;
wire [31:0] \datapath_1.regfile_1.regOut[0]  ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire \datapath_1.regfile_1.regEn_20_bF$buf7  ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire \datapath_1.regfile_1.regEn_2_bF$buf5  ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _3194_ ;
wire [31:0] \datapath_1.rd2  ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _5816_ ;
wire _1736_ ;
wire _1316_ ;
wire _3944__bF$buf0 ;
wire _3944__bF$buf1 ;
wire _3944__bF$buf2 ;
wire _3944__bF$buf3 ;
wire _3944__bF$buf4 ;
wire _647_ ;
wire _227_ ;
wire \datapath_1.regfile_1.regEn_25_bF$buf3  ;
wire _6774_ ;
wire _6354_ ;
wire \datapath_1.regfile_1.regEn_7_bF$buf1  ;
wire _2694_ ;
wire _2274_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire [31:0] \datapath_1.regfile_1.regOut[23]  ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire [31:0] memoryOutData ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire [1:0] ALUOp ;
wire _5500__bF$buf0 ;
wire _5500__bF$buf1 ;
wire _685_ ;
wire _5500__bF$buf2 ;
wire _265_ ;
wire _5500__bF$buf3 ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire \datapath_1.mux_wd3.dout_28_bF$buf2  ;
wire _4705_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire \datapath_1.regfile_1.regEn_28_bF$buf6  ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _1639_ ;
wire _1219_ ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;

BUFX2 BUFX2_insert1093 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf0)
);

BUFX2 BUFX2_insert1092 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf1)
);

BUFX2 BUFX2_insert1091 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf2)
);

BUFX2 BUFX2_insert1090 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf3)
);

BUFX2 BUFX2_insert1089 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf4)
);

BUFX2 BUFX2_insert1088 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf5)
);

BUFX2 BUFX2_insert1087 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf6)
);

BUFX2 BUFX2_insert1086 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf7)
);

BUFX2 BUFX2_insert1085 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf8)
);

BUFX2 BUFX2_insert1084 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst),
    .Y(rst_hier0_bF$buf9)
);

CLKBUF1 CLKBUF1_insert1083 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert1082 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert1081 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1080 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1079 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1078 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1077 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1076 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf7)
);

CLKBUF1 CLKBUF1_insert1075 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf8)
);

CLKBUF1 CLKBUF1_insert1074 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_hier0_bF$buf9)
);

BUFX2 BUFX2_insert1073 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf0 )
);

BUFX2 BUFX2_insert1072 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf1 )
);

BUFX2 BUFX2_insert1071 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf2 )
);

BUFX2 BUFX2_insert1070 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf3 )
);

BUFX2 BUFX2_insert1069 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf4 )
);

BUFX2 BUFX2_insert1068 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf5 )
);

BUFX2 BUFX2_insert1067 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf6 )
);

BUFX2 BUFX2_insert1066 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [16]),
    .Y(\datapath_1.regfile_1.regEn_16_bF$buf7 )
);

BUFX2 BUFX2_insert1065 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf0)
);

BUFX2 BUFX2_insert1064 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf1)
);

BUFX2 BUFX2_insert1063 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf2)
);

BUFX2 BUFX2_insert1062 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf3)
);

BUFX2 BUFX2_insert1061 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5531_),
    .Y(_5531__bF$buf0)
);

BUFX2 BUFX2_insert1060 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5531_),
    .Y(_5531__bF$buf1)
);

BUFX2 BUFX2_insert1059 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5531_),
    .Y(_5531__bF$buf2)
);

BUFX2 BUFX2_insert1058 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5531_),
    .Y(_5531__bF$buf3)
);

BUFX2 BUFX2_insert1057 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5531_),
    .Y(_5531__bF$buf4)
);

BUFX2 BUFX2_insert1056 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .Y(_4038__bF$buf0)
);

BUFX2 BUFX2_insert1055 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .Y(_4038__bF$buf1)
);

BUFX2 BUFX2_insert1054 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .Y(_4038__bF$buf2)
);

BUFX2 BUFX2_insert1053 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .Y(_4038__bF$buf3)
);

BUFX2 BUFX2_insert1052 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf0 )
);

BUFX2 BUFX2_insert1051 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf1 )
);

BUFX2 BUFX2_insert1050 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf2 )
);

BUFX2 BUFX2_insert1049 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf3 )
);

BUFX2 BUFX2_insert1048 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [17]),
    .Y(\datapath_1.PCJump_17_bF$buf4 )
);

BUFX2 BUFX2_insert1047 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf0 )
);

BUFX2 BUFX2_insert1046 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf1 )
);

BUFX2 BUFX2_insert1045 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf2 )
);

BUFX2 BUFX2_insert1044 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf3 )
);

BUFX2 BUFX2_insert1043 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf4 )
);

BUFX2 BUFX2_insert1042 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf5 )
);

BUFX2 BUFX2_insert1041 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf6 )
);

BUFX2 BUFX2_insert1040 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [7]),
    .Y(\datapath_1.regfile_1.regEn_7_bF$buf7 )
);

BUFX2 BUFX2_insert1039 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf0 )
);

BUFX2 BUFX2_insert1038 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf1 )
);

BUFX2 BUFX2_insert1037 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf2 )
);

BUFX2 BUFX2_insert1036 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf3 )
);

BUFX2 BUFX2_insert1035 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [15]),
    .Y(\datapath_1.mux_wd3.dout_15_bF$buf4 )
);

BUFX2 BUFX2_insert1034 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf0 )
);

BUFX2 BUFX2_insert1033 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf1 )
);

BUFX2 BUFX2_insert1032 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf2 )
);

BUFX2 BUFX2_insert1031 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf3 )
);

BUFX2 BUFX2_insert1030 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf4 )
);

BUFX2 BUFX2_insert1029 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf5 )
);

BUFX2 BUFX2_insert1028 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf6 )
);

BUFX2 BUFX2_insert1027 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [19]),
    .Y(\datapath_1.regfile_1.regEn_19_bF$buf7 )
);

BUFX2 BUFX2_insert1026 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf0 )
);

BUFX2 BUFX2_insert1025 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf1 )
);

BUFX2 BUFX2_insert1024 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf2 )
);

BUFX2 BUFX2_insert1023 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf3 )
);

BUFX2 BUFX2_insert1022 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf4 )
);

BUFX2 BUFX2_insert1021 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf5 )
);

BUFX2 BUFX2_insert1020 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf6 )
);

BUFX2 BUFX2_insert1019 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [22]),
    .Y(\datapath_1.regfile_1.regEn_22_bF$buf7 )
);

BUFX2 BUFX2_insert1018 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534_),
    .Y(_5534__bF$buf0)
);

BUFX2 BUFX2_insert1017 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534_),
    .Y(_5534__bF$buf1)
);

BUFX2 BUFX2_insert1016 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534_),
    .Y(_5534__bF$buf2)
);

BUFX2 BUFX2_insert1015 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534_),
    .Y(_5534__bF$buf3)
);

BUFX2 BUFX2_insert1014 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534_),
    .Y(_5534__bF$buf4)
);

BUFX2 BUFX2_insert1013 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4079_),
    .Y(_4079__bF$buf0)
);

BUFX2 BUFX2_insert1012 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4079_),
    .Y(_4079__bF$buf1)
);

BUFX2 BUFX2_insert1011 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4079_),
    .Y(_4079__bF$buf2)
);

BUFX2 BUFX2_insert1010 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4079_),
    .Y(_4079__bF$buf3)
);

BUFX2 BUFX2_insert1009 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf0)
);

BUFX2 BUFX2_insert1008 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf1)
);

BUFX2 BUFX2_insert1007 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf2)
);

BUFX2 BUFX2_insert1006 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf3)
);

BUFX2 BUFX2_insert1005 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[1]),
    .Y(ALUSrcB_1_bF$buf4)
);

BUFX2 BUFX2_insert1004 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf0 )
);

BUFX2 BUFX2_insert1003 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf1 )
);

BUFX2 BUFX2_insert1002 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf2 )
);

BUFX2 BUFX2_insert1001 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf3 )
);

BUFX2 BUFX2_insert1000 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [18]),
    .Y(\datapath_1.mux_wd3.dout_18_bF$buf4 )
);

BUFX2 BUFX2_insert999 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf0)
);

BUFX2 BUFX2_insert998 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf1)
);

BUFX2 BUFX2_insert997 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf2)
);

BUFX2 BUFX2_insert996 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf3)
);

BUFX2 BUFX2_insert995 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf0 )
);

BUFX2 BUFX2_insert994 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf1 )
);

BUFX2 BUFX2_insert993 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf2 )
);

BUFX2 BUFX2_insert992 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf3 )
);

BUFX2 BUFX2_insert991 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [21]),
    .Y(\datapath_1.mux_wd3.dout_21_bF$buf4 )
);

BUFX2 BUFX2_insert990 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf0 )
);

BUFX2 BUFX2_insert989 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf1 )
);

BUFX2 BUFX2_insert988 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf2 )
);

BUFX2 BUFX2_insert987 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf3 )
);

BUFX2 BUFX2_insert986 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf4 )
);

BUFX2 BUFX2_insert985 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf5 )
);

BUFX2 BUFX2_insert984 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf6 )
);

BUFX2 BUFX2_insert983 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [25]),
    .Y(\datapath_1.regfile_1.regEn_25_bF$buf7 )
);

BUFX2 BUFX2_insert982 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .Y(_3967__bF$buf0)
);

BUFX2 BUFX2_insert981 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .Y(_3967__bF$buf1)
);

BUFX2 BUFX2_insert980 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .Y(_3967__bF$buf2)
);

BUFX2 BUFX2_insert979 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .Y(_3967__bF$buf3)
);

BUFX2 BUFX2_insert978 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf0)
);

BUFX2 BUFX2_insert977 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf1)
);

BUFX2 BUFX2_insert976 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf2)
);

BUFX2 BUFX2_insert975 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf3)
);

BUFX2 BUFX2_insert974 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf4)
);

BUFX2 BUFX2_insert973 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf5)
);

BUFX2 BUFX2_insert972 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf6)
);

BUFX2 BUFX2_insert971 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn),
    .Y(PCEn_bF$buf7)
);

BUFX2 BUFX2_insert970 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf0 )
);

BUFX2 BUFX2_insert969 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf1 )
);

BUFX2 BUFX2_insert968 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf2 )
);

BUFX2 BUFX2_insert967 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf3 )
);

BUFX2 BUFX2_insert966 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [24]),
    .Y(\datapath_1.mux_wd3.dout_24_bF$buf4 )
);

BUFX2 BUFX2_insert965 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf0 )
);

BUFX2 BUFX2_insert964 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf1 )
);

BUFX2 BUFX2_insert963 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf2 )
);

BUFX2 BUFX2_insert962 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf3 )
);

BUFX2 BUFX2_insert961 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf4 )
);

BUFX2 BUFX2_insert960 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf5 )
);

BUFX2 BUFX2_insert959 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf6 )
);

BUFX2 BUFX2_insert958 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [28]),
    .Y(\datapath_1.regfile_1.regEn_28_bF$buf7 )
);

BUFX2 BUFX2_insert957 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf0 )
);

BUFX2 BUFX2_insert956 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf1 )
);

BUFX2 BUFX2_insert955 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf2 )
);

BUFX2 BUFX2_insert954 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf3 )
);

BUFX2 BUFX2_insert953 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf4 )
);

BUFX2 BUFX2_insert952 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf5 )
);

BUFX2 BUFX2_insert951 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf6 )
);

BUFX2 BUFX2_insert950 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [31]),
    .Y(\datapath_1.regfile_1.regEn_31_bF$buf7 )
);

BUFX2 BUFX2_insert949 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3036_),
    .Y(_3036__bF$buf0)
);

BUFX2 BUFX2_insert948 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3036_),
    .Y(_3036__bF$buf1)
);

BUFX2 BUFX2_insert947 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3036_),
    .Y(_3036__bF$buf2)
);

BUFX2 BUFX2_insert946 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3036_),
    .Y(_3036__bF$buf3)
);

BUFX2 BUFX2_insert945 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3036_),
    .Y(_3036__bF$buf4)
);

BUFX2 BUFX2_insert944 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf0 )
);

BUFX2 BUFX2_insert943 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf1 )
);

BUFX2 BUFX2_insert942 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf2 )
);

BUFX2 BUFX2_insert941 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf3 )
);

BUFX2 BUFX2_insert940 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [27]),
    .Y(\datapath_1.mux_wd3.dout_27_bF$buf4 )
);

BUFX2 BUFX2_insert939 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935_),
    .Y(_3935__bF$buf0)
);

BUFX2 BUFX2_insert938 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935_),
    .Y(_3935__bF$buf1)
);

BUFX2 BUFX2_insert937 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935_),
    .Y(_3935__bF$buf2)
);

BUFX2 BUFX2_insert936 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935_),
    .Y(_3935__bF$buf3)
);

BUFX2 BUFX2_insert935 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935_),
    .Y(_3935__bF$buf4)
);

BUFX2 BUFX2_insert934 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf0 )
);

BUFX2 BUFX2_insert933 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf1 )
);

BUFX2 BUFX2_insert932 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf2 )
);

BUFX2 BUFX2_insert931 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf3 )
);

BUFX2 BUFX2_insert930 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [30]),
    .Y(\datapath_1.mux_wd3.dout_30_bF$buf4 )
);

BUFX2 BUFX2_insert929 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf0 )
);

BUFX2 BUFX2_insert928 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf1 )
);

BUFX2 BUFX2_insert927 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf2 )
);

BUFX2 BUFX2_insert926 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf3 )
);

BUFX2 BUFX2_insert925 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [2]),
    .Y(\datapath_1.mux_wd3.dout_2_bF$buf4 )
);

BUFX2 BUFX2_insert924 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882_),
    .Y(_3882__bF$buf0)
);

BUFX2 BUFX2_insert923 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882_),
    .Y(_3882__bF$buf1)
);

BUFX2 BUFX2_insert922 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882_),
    .Y(_3882__bF$buf2)
);

BUFX2 BUFX2_insert921 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882_),
    .Y(_3882__bF$buf3)
);

BUFX2 BUFX2_insert920 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .Y(_5549__bF$buf0)
);

BUFX2 BUFX2_insert919 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .Y(_5549__bF$buf1)
);

BUFX2 BUFX2_insert918 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .Y(_5549__bF$buf2)
);

BUFX2 BUFX2_insert917 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .Y(_5549__bF$buf3)
);

BUFX2 BUFX2_insert916 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .Y(_5549__bF$buf4)
);

BUFX2 BUFX2_insert915 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf0 )
);

BUFX2 BUFX2_insert914 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf1 )
);

BUFX2 BUFX2_insert913 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf2 )
);

BUFX2 BUFX2_insert912 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf3 )
);

BUFX2 BUFX2_insert911 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [5]),
    .Y(\datapath_1.mux_wd3.dout_5_bF$buf4 )
);

BUFX2 BUFX2_insert910 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf0)
);

BUFX2 BUFX2_insert909 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf1)
);

BUFX2 BUFX2_insert908 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf2)
);

BUFX2 BUFX2_insert907 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf3)
);

BUFX2 BUFX2_insert906 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf4)
);

BUFX2 BUFX2_insert905 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf5)
);

BUFX2 BUFX2_insert904 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf6)
);

BUFX2 BUFX2_insert903 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite),
    .Y(IRWrite_bF$buf7)
);

BUFX2 BUFX2_insert902 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552_),
    .Y(_5552__bF$buf0)
);

BUFX2 BUFX2_insert901 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552_),
    .Y(_5552__bF$buf1)
);

BUFX2 BUFX2_insert900 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552_),
    .Y(_5552__bF$buf2)
);

BUFX2 BUFX2_insert899 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552_),
    .Y(_5552__bF$buf3)
);

BUFX2 BUFX2_insert898 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982_),
    .Y(_3982__bF$buf0)
);

BUFX2 BUFX2_insert897 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982_),
    .Y(_3982__bF$buf1)
);

BUFX2 BUFX2_insert896 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982_),
    .Y(_3982__bF$buf2)
);

BUFX2 BUFX2_insert895 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982_),
    .Y(_3982__bF$buf3)
);

BUFX2 BUFX2_insert894 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf0 )
);

BUFX2 BUFX2_insert893 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf1 )
);

BUFX2 BUFX2_insert892 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf2 )
);

BUFX2 BUFX2_insert891 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf3 )
);

BUFX2 BUFX2_insert890 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [8]),
    .Y(\datapath_1.mux_wd3.dout_8_bF$buf4 )
);

BUFX2 BUFX2_insert889 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .Y(_3944__bF$buf0)
);

BUFX2 BUFX2_insert888 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .Y(_3944__bF$buf1)
);

BUFX2 BUFX2_insert887 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .Y(_3944__bF$buf2)
);

BUFX2 BUFX2_insert886 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .Y(_3944__bF$buf3)
);

BUFX2 BUFX2_insert885 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .Y(_3944__bF$buf4)
);

BUFX2 BUFX2_insert884 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3201_),
    .Y(_3201__bF$buf0)
);

BUFX2 BUFX2_insert883 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3201_),
    .Y(_3201__bF$buf1)
);

BUFX2 BUFX2_insert882 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3201_),
    .Y(_3201__bF$buf2)
);

BUFX2 BUFX2_insert881 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3201_),
    .Y(_3201__bF$buf3)
);

BUFX2 BUFX2_insert880 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3201_),
    .Y(_3201__bF$buf4)
);

BUFX2 BUFX2_insert879 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499_),
    .Y(_5499__bF$buf0)
);

BUFX2 BUFX2_insert878 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499_),
    .Y(_5499__bF$buf1)
);

BUFX2 BUFX2_insert877 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499_),
    .Y(_5499__bF$buf2)
);

BUFX2 BUFX2_insert876 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499_),
    .Y(_5499__bF$buf3)
);

BUFX2 BUFX2_insert875 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947_),
    .Y(_3947__bF$buf0)
);

BUFX2 BUFX2_insert874 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947_),
    .Y(_3947__bF$buf1)
);

BUFX2 BUFX2_insert873 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947_),
    .Y(_3947__bF$buf2)
);

BUFX2 BUFX2_insert872 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947_),
    .Y(_3947__bF$buf3)
);

BUFX2 BUFX2_insert871 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891_),
    .Y(_3891__bF$buf0)
);

BUFX2 BUFX2_insert870 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891_),
    .Y(_3891__bF$buf1)
);

BUFX2 BUFX2_insert869 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891_),
    .Y(_3891__bF$buf2)
);

BUFX2 BUFX2_insert868 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891_),
    .Y(_3891__bF$buf3)
);

BUFX2 BUFX2_insert867 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .Y(_3950__bF$buf0)
);

BUFX2 BUFX2_insert866 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .Y(_3950__bF$buf1)
);

BUFX2 BUFX2_insert865 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .Y(_3950__bF$buf2)
);

BUFX2 BUFX2_insert864 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .Y(_3950__bF$buf3)
);

BUFX2 BUFX2_insert863 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf0 )
);

BUFX2 BUFX2_insert862 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf1 )
);

BUFX2 BUFX2_insert861 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf2 )
);

BUFX2 BUFX2_insert860 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf3 )
);

BUFX2 BUFX2_insert859 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf4 )
);

BUFX2 BUFX2_insert858 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf5 )
);

BUFX2 BUFX2_insert857 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf6 )
);

BUFX2 BUFX2_insert856 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [11]),
    .Y(\datapath_1.regfile_1.regEn_11_bF$buf7 )
);

BUFX2 BUFX2_insert855 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf0 )
);

BUFX2 BUFX2_insert854 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf1 )
);

BUFX2 BUFX2_insert853 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf2 )
);

BUFX2 BUFX2_insert852 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf3 )
);

BUFX2 BUFX2_insert851 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf4 )
);

BUFX2 BUFX2_insert850 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf5 )
);

BUFX2 BUFX2_insert849 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf6 )
);

BUFX2 BUFX2_insert848 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [2]),
    .Y(\datapath_1.regfile_1.regEn_2_bF$buf7 )
);

BUFX2 BUFX2_insert847 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf0 )
);

BUFX2 BUFX2_insert846 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf1 )
);

BUFX2 BUFX2_insert845 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf2 )
);

BUFX2 BUFX2_insert844 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf3 )
);

BUFX2 BUFX2_insert843 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [10]),
    .Y(\datapath_1.mux_wd3.dout_10_bF$buf4 )
);

BUFX2 BUFX2_insert842 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf0 )
);

BUFX2 BUFX2_insert841 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf1 )
);

BUFX2 BUFX2_insert840 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf2 )
);

BUFX2 BUFX2_insert839 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf3 )
);

BUFX2 BUFX2_insert838 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf4 )
);

BUFX2 BUFX2_insert837 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf5 )
);

BUFX2 BUFX2_insert836 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf6 )
);

BUFX2 BUFX2_insert835 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [14]),
    .Y(\datapath_1.regfile_1.regEn_14_bF$buf7 )
);

BUFX2 BUFX2_insert834 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526_),
    .Y(_5526__bF$buf0)
);

BUFX2 BUFX2_insert833 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526_),
    .Y(_5526__bF$buf1)
);

BUFX2 BUFX2_insert832 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526_),
    .Y(_5526__bF$buf2)
);

BUFX2 BUFX2_insert831 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526_),
    .Y(_5526__bF$buf3)
);

BUFX2 BUFX2_insert830 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526_),
    .Y(_5526__bF$buf4)
);

BUFX2 BUFX2_insert829 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf0 )
);

BUFX2 BUFX2_insert828 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf1 )
);

BUFX2 BUFX2_insert827 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf2 )
);

BUFX2 BUFX2_insert826 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf3 )
);

BUFX2 BUFX2_insert825 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf4 )
);

BUFX2 BUFX2_insert824 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf5 )
);

BUFX2 BUFX2_insert823 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf6 )
);

BUFX2 BUFX2_insert822 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [5]),
    .Y(\datapath_1.regfile_1.regEn_5_bF$buf7 )
);

BUFX2 BUFX2_insert821 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf0 )
);

BUFX2 BUFX2_insert820 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf1 )
);

BUFX2 BUFX2_insert819 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf2 )
);

BUFX2 BUFX2_insert818 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf3 )
);

BUFX2 BUFX2_insert817 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [13]),
    .Y(\datapath_1.mux_wd3.dout_13_bF$buf4 )
);

BUFX2 BUFX2_insert816 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf0 )
);

BUFX2 BUFX2_insert815 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf1 )
);

BUFX2 BUFX2_insert814 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf2 )
);

BUFX2 BUFX2_insert813 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf3 )
);

BUFX2 BUFX2_insert812 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf4 )
);

BUFX2 BUFX2_insert811 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf5 )
);

BUFX2 BUFX2_insert810 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf6 )
);

BUFX2 BUFX2_insert809 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [17]),
    .Y(\datapath_1.regfile_1.regEn_17_bF$buf7 )
);

BUFX2 BUFX2_insert808 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .Y(_4001__bF$buf0)
);

BUFX2 BUFX2_insert807 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .Y(_4001__bF$buf1)
);

BUFX2 BUFX2_insert806 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .Y(_4001__bF$buf2)
);

BUFX2 BUFX2_insert805 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .Y(_4001__bF$buf3)
);

BUFX2 BUFX2_insert804 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570_),
    .Y(_5570__bF$buf0)
);

BUFX2 BUFX2_insert803 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570_),
    .Y(_5570__bF$buf1)
);

BUFX2 BUFX2_insert802 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570_),
    .Y(_5570__bF$buf2)
);

BUFX2 BUFX2_insert801 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570_),
    .Y(_5570__bF$buf3)
);

BUFX2 BUFX2_insert800 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf0 )
);

BUFX2 BUFX2_insert799 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf1 )
);

BUFX2 BUFX2_insert798 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf2 )
);

BUFX2 BUFX2_insert797 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf3 )
);

BUFX2 BUFX2_insert796 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf4 )
);

BUFX2 BUFX2_insert795 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf5 )
);

BUFX2 BUFX2_insert794 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf6 )
);

BUFX2 BUFX2_insert793 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [20]),
    .Y(\datapath_1.regfile_1.regEn_20_bF$buf7 )
);

BUFX2 BUFX2_insert792 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5532_),
    .Y(_5532__bF$buf0)
);

BUFX2 BUFX2_insert791 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5532_),
    .Y(_5532__bF$buf1)
);

BUFX2 BUFX2_insert790 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5532_),
    .Y(_5532__bF$buf2)
);

BUFX2 BUFX2_insert789 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5532_),
    .Y(_5532__bF$buf3)
);

BUFX2 BUFX2_insert788 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3997_),
    .Y(_3997__bF$buf0)
);

BUFX2 BUFX2_insert787 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3997_),
    .Y(_3997__bF$buf1)
);

BUFX2 BUFX2_insert786 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3997_),
    .Y(_3997__bF$buf2)
);

BUFX2 BUFX2_insert785 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3997_),
    .Y(_3997__bF$buf3)
);

BUFX2 BUFX2_insert784 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf0)
);

BUFX2 BUFX2_insert783 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf1)
);

BUFX2 BUFX2_insert782 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf2)
);

BUFX2 BUFX2_insert781 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf3)
);

BUFX2 BUFX2_insert780 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf4)
);

BUFX2 BUFX2_insert779 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf5)
);

BUFX2 BUFX2_insert778 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf6)
);

BUFX2 BUFX2_insert777 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA),
    .Y(ALUSrcA_bF$buf7)
);

BUFX2 BUFX2_insert776 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf0 )
);

BUFX2 BUFX2_insert775 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf1 )
);

BUFX2 BUFX2_insert774 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf2 )
);

BUFX2 BUFX2_insert773 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf3 )
);

BUFX2 BUFX2_insert772 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf4 )
);

BUFX2 BUFX2_insert771 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf5 )
);

BUFX2 BUFX2_insert770 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf6 )
);

BUFX2 BUFX2_insert769 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [8]),
    .Y(\datapath_1.regfile_1.regEn_8_bF$buf7 )
);

BUFX2 BUFX2_insert768 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf0 )
);

BUFX2 BUFX2_insert767 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf1 )
);

BUFX2 BUFX2_insert766 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf2 )
);

BUFX2 BUFX2_insert765 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf3 )
);

BUFX2 BUFX2_insert764 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [16]),
    .Y(\datapath_1.mux_wd3.dout_16_bF$buf4 )
);

BUFX2 BUFX2_insert763 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3924_),
    .Y(_3924__bF$buf0)
);

BUFX2 BUFX2_insert762 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3924_),
    .Y(_3924__bF$buf1)
);

BUFX2 BUFX2_insert761 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3924_),
    .Y(_3924__bF$buf2)
);

BUFX2 BUFX2_insert760 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3924_),
    .Y(_3924__bF$buf3)
);

BUFX2 BUFX2_insert759 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3198_),
    .Y(_3198__bF$buf0)
);

BUFX2 BUFX2_insert758 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3198_),
    .Y(_3198__bF$buf1)
);

BUFX2 BUFX2_insert757 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3198_),
    .Y(_3198__bF$buf2)
);

BUFX2 BUFX2_insert756 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3198_),
    .Y(_3198__bF$buf3)
);

BUFX2 BUFX2_insert755 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3198_),
    .Y(_3198__bF$buf4)
);

BUFX2 BUFX2_insert754 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf0 )
);

BUFX2 BUFX2_insert753 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf1 )
);

BUFX2 BUFX2_insert752 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf2 )
);

BUFX2 BUFX2_insert751 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf3 )
);

BUFX2 BUFX2_insert750 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf4 )
);

BUFX2 BUFX2_insert749 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf5 )
);

BUFX2 BUFX2_insert748 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf6 )
);

BUFX2 BUFX2_insert747 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [23]),
    .Y(\datapath_1.regfile_1.regEn_23_bF$buf7 )
);

BUFX2 BUFX2_insert746 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5535_),
    .Y(_5535__bF$buf0)
);

BUFX2 BUFX2_insert745 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5535_),
    .Y(_5535__bF$buf1)
);

BUFX2 BUFX2_insert744 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5535_),
    .Y(_5535__bF$buf2)
);

BUFX2 BUFX2_insert743 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5535_),
    .Y(_5535__bF$buf3)
);

BUFX2 BUFX2_insert742 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5535_),
    .Y(_5535__bF$buf4)
);

BUFX2 BUFX2_insert741 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf0 )
);

BUFX2 BUFX2_insert740 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf1 )
);

BUFX2 BUFX2_insert739 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf2 )
);

BUFX2 BUFX2_insert738 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf3 )
);

BUFX2 BUFX2_insert737 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [19]),
    .Y(\datapath_1.mux_wd3.dout_19_bF$buf4 )
);

BUFX2 BUFX2_insert736 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .Y(_5500__bF$buf0)
);

BUFX2 BUFX2_insert735 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .Y(_5500__bF$buf1)
);

BUFX2 BUFX2_insert734 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .Y(_5500__bF$buf2)
);

BUFX2 BUFX2_insert733 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .Y(_5500__bF$buf3)
);

BUFX2 BUFX2_insert732 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf0 )
);

BUFX2 BUFX2_insert731 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf1 )
);

BUFX2 BUFX2_insert730 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf2 )
);

BUFX2 BUFX2_insert729 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf3 )
);

BUFX2 BUFX2_insert728 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [22]),
    .Y(\datapath_1.mux_wd3.dout_22_bF$buf4 )
);

BUFX2 BUFX2_insert727 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf0 )
);

BUFX2 BUFX2_insert726 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf1 )
);

BUFX2 BUFX2_insert725 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf2 )
);

BUFX2 BUFX2_insert724 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf3 )
);

BUFX2 BUFX2_insert723 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf4 )
);

BUFX2 BUFX2_insert722 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf5 )
);

BUFX2 BUFX2_insert721 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf6 )
);

BUFX2 BUFX2_insert720 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [26]),
    .Y(\datapath_1.regfile_1.regEn_26_bF$buf7 )
);

BUFX2 BUFX2_insert719 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .Y(_3930__bF$buf0)
);

BUFX2 BUFX2_insert718 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .Y(_3930__bF$buf1)
);

BUFX2 BUFX2_insert717 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .Y(_3930__bF$buf2)
);

BUFX2 BUFX2_insert716 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .Y(_3930__bF$buf3)
);

BUFX2 BUFX2_insert715 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .Y(_5503__bF$buf0)
);

BUFX2 BUFX2_insert714 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .Y(_5503__bF$buf1)
);

BUFX2 BUFX2_insert713 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .Y(_5503__bF$buf2)
);

BUFX2 BUFX2_insert712 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .Y(_5503__bF$buf3)
);

BUFX2 BUFX2_insert711 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf0 )
);

BUFX2 BUFX2_insert710 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf1 )
);

BUFX2 BUFX2_insert709 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf2 )
);

BUFX2 BUFX2_insert708 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf3 )
);

BUFX2 BUFX2_insert707 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [27]),
    .Y(\datapath_1.PCJump_27_bF$buf4 )
);

BUFX2 BUFX2_insert706 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .Y(_3034__bF$buf0)
);

BUFX2 BUFX2_insert705 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .Y(_3034__bF$buf1)
);

BUFX2 BUFX2_insert704 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .Y(_3034__bF$buf2)
);

BUFX2 BUFX2_insert703 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .Y(_3034__bF$buf3)
);

BUFX2 BUFX2_insert702 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .Y(_3034__bF$buf4)
);

BUFX2 BUFX2_insert701 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf0 )
);

BUFX2 BUFX2_insert700 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf1 )
);

BUFX2 BUFX2_insert699 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf2 )
);

BUFX2 BUFX2_insert698 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf3 )
);

BUFX2 BUFX2_insert697 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [25]),
    .Y(\datapath_1.mux_wd3.dout_25_bF$buf4 )
);

BUFX2 BUFX2_insert696 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf0 )
);

BUFX2 BUFX2_insert695 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf1 )
);

BUFX2 BUFX2_insert694 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf2 )
);

BUFX2 BUFX2_insert693 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf3 )
);

BUFX2 BUFX2_insert692 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf4 )
);

BUFX2 BUFX2_insert691 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf5 )
);

BUFX2 BUFX2_insert690 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf6 )
);

BUFX2 BUFX2_insert689 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [29]),
    .Y(\datapath_1.regfile_1.regEn_29_bF$buf7 )
);

BUFX2 BUFX2_insert688 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3971_),
    .Y(_3971__bF$buf0)
);

BUFX2 BUFX2_insert687 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3971_),
    .Y(_3971__bF$buf1)
);

BUFX2 BUFX2_insert686 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3971_),
    .Y(_3971__bF$buf2)
);

BUFX2 BUFX2_insert685 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3971_),
    .Y(_3971__bF$buf3)
);

BUFX2 BUFX2_insert684 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3971_),
    .Y(_3971__bF$buf4)
);

BUFX2 BUFX2_insert683 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .Y(_5485__bF$buf0)
);

BUFX2 BUFX2_insert682 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .Y(_5485__bF$buf1)
);

BUFX2 BUFX2_insert681 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .Y(_5485__bF$buf2)
);

BUFX2 BUFX2_insert680 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .Y(_5485__bF$buf3)
);

BUFX2 BUFX2_insert679 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .Y(_5485__bF$buf4)
);

BUFX2 BUFX2_insert678 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051_),
    .Y(_4051__bF$buf0)
);

BUFX2 BUFX2_insert677 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051_),
    .Y(_4051__bF$buf1)
);

BUFX2 BUFX2_insert676 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051_),
    .Y(_4051__bF$buf2)
);

BUFX2 BUFX2_insert675 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051_),
    .Y(_4051__bF$buf3)
);

BUFX2 BUFX2_insert674 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .Y(_5544__bF$buf0)
);

BUFX2 BUFX2_insert673 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .Y(_5544__bF$buf1)
);

BUFX2 BUFX2_insert672 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .Y(_5544__bF$buf2)
);

BUFX2 BUFX2_insert671 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .Y(_5544__bF$buf3)
);

BUFX2 BUFX2_insert670 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf0 )
);

BUFX2 BUFX2_insert669 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf1 )
);

BUFX2 BUFX2_insert668 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf2 )
);

BUFX2 BUFX2_insert667 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf3 )
);

BUFX2 BUFX2_insert666 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [0]),
    .Y(\datapath_1.mux_wd3.dout_0_bF$buf4 )
);

BUFX2 BUFX2_insert665 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .Y(_2481__bF$buf0)
);

BUFX2 BUFX2_insert664 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .Y(_2481__bF$buf1)
);

BUFX2 BUFX2_insert663 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .Y(_2481__bF$buf2)
);

BUFX2 BUFX2_insert662 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .Y(_2481__bF$buf3)
);

BUFX2 BUFX2_insert661 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .Y(_3037__bF$buf0)
);

BUFX2 BUFX2_insert660 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .Y(_3037__bF$buf1)
);

BUFX2 BUFX2_insert659 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .Y(_3037__bF$buf2)
);

BUFX2 BUFX2_insert658 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .Y(_3037__bF$buf3)
);

BUFX2 BUFX2_insert657 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3037_),
    .Y(_3037__bF$buf4)
);

BUFX2 BUFX2_insert656 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf0 )
);

BUFX2 BUFX2_insert655 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf1 )
);

BUFX2 BUFX2_insert654 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf2 )
);

BUFX2 BUFX2_insert653 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf3 )
);

BUFX2 BUFX2_insert652 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [28]),
    .Y(\datapath_1.mux_wd3.dout_28_bF$buf4 )
);

BUFX2 BUFX2_insert651 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf0)
);

BUFX2 BUFX2_insert650 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf1)
);

BUFX2 BUFX2_insert649 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf2)
);

BUFX2 BUFX2_insert648 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf3)
);

BUFX2 BUFX2_insert647 (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource[1]),
    .Y(PCSource_1_bF$buf4)
);

BUFX2 BUFX2_insert646 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .Y(_3936__bF$buf0)
);

BUFX2 BUFX2_insert645 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .Y(_3936__bF$buf1)
);

BUFX2 BUFX2_insert644 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .Y(_3936__bF$buf2)
);

BUFX2 BUFX2_insert643 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .Y(_3936__bF$buf3)
);

BUFX2 BUFX2_insert642 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .Y(_3936__bF$buf4)
);

BUFX2 BUFX2_insert641 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf0 )
);

BUFX2 BUFX2_insert640 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf1 )
);

BUFX2 BUFX2_insert639 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf2 )
);

BUFX2 BUFX2_insert638 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf3 )
);

BUFX2 BUFX2_insert637 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [31]),
    .Y(\datapath_1.mux_wd3.dout_31_bF$buf4 )
);

BUFX2 BUFX2_insert636 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf0 )
);

BUFX2 BUFX2_insert635 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf1 )
);

BUFX2 BUFX2_insert634 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf2 )
);

BUFX2 BUFX2_insert633 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf3 )
);

BUFX2 BUFX2_insert632 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [3]),
    .Y(\datapath_1.mux_wd3.dout_3_bF$buf4 )
);

BUFX2 BUFX2_insert631 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3977_),
    .Y(_3977__bF$buf0)
);

BUFX2 BUFX2_insert630 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3977_),
    .Y(_3977__bF$buf1)
);

BUFX2 BUFX2_insert629 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3977_),
    .Y(_3977__bF$buf2)
);

BUFX2 BUFX2_insert628 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3977_),
    .Y(_3977__bF$buf3)
);

BUFX2 BUFX2_insert627 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3977_),
    .Y(_3977__bF$buf4)
);

BUFX2 BUFX2_insert626 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf0 )
);

BUFX2 BUFX2_insert625 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf1 )
);

BUFX2 BUFX2_insert624 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf2 )
);

BUFX2 BUFX2_insert623 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf3 )
);

BUFX2 BUFX2_insert622 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [6]),
    .Y(\datapath_1.mux_wd3.dout_6_bF$buf4 )
);

BUFX2 BUFX2_insert621 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3942_),
    .Y(_3942__bF$buf0)
);

BUFX2 BUFX2_insert620 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3942_),
    .Y(_3942__bF$buf1)
);

BUFX2 BUFX2_insert619 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3942_),
    .Y(_3942__bF$buf2)
);

BUFX2 BUFX2_insert618 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3942_),
    .Y(_3942__bF$buf3)
);

BUFX2 BUFX2_insert617 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf0)
);

BUFX2 BUFX2_insert616 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf1)
);

BUFX2 BUFX2_insert615 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf2)
);

BUFX2 BUFX2_insert614 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf3)
);

BUFX2 BUFX2_insert613 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf4)
);

BUFX2 BUFX2_insert612 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[0]),
    .Y(ALUOp_0_bF$buf5)
);

BUFX2 BUFX2_insert611 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .Y(_5515__bF$buf0)
);

BUFX2 BUFX2_insert610 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .Y(_5515__bF$buf1)
);

BUFX2 BUFX2_insert609 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .Y(_5515__bF$buf2)
);

BUFX2 BUFX2_insert608 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .Y(_5515__bF$buf3)
);

BUFX2 BUFX2_insert607 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf0)
);

BUFX2 BUFX2_insert606 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf1)
);

BUFX2 BUFX2_insert605 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf2)
);

BUFX2 BUFX2_insert604 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf3)
);

BUFX2 BUFX2_insert603 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf4)
);

BUFX2 BUFX2_insert602 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf5)
);

BUFX2 BUFX2_insert601 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf6)
);

BUFX2 BUFX2_insert600 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf7)
);

BUFX2 BUFX2_insert599 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf8)
);

BUFX2 BUFX2_insert598 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf9)
);

BUFX2 BUFX2_insert597 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf10)
);

BUFX2 BUFX2_insert596 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf11)
);

BUFX2 BUFX2_insert595 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf12)
);

BUFX2 BUFX2_insert594 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf13)
);

BUFX2 BUFX2_insert593 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf14)
);

BUFX2 BUFX2_insert592 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf15)
);

BUFX2 BUFX2_insert591 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf16)
);

BUFX2 BUFX2_insert590 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf17)
);

BUFX2 BUFX2_insert589 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf18)
);

BUFX2 BUFX2_insert588 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf19)
);

BUFX2 BUFX2_insert587 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf20)
);

BUFX2 BUFX2_insert586 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf21)
);

BUFX2 BUFX2_insert585 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf22)
);

BUFX2 BUFX2_insert584 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf23)
);

BUFX2 BUFX2_insert583 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf24)
);

BUFX2 BUFX2_insert582 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf25)
);

BUFX2 BUFX2_insert581 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf26)
);

BUFX2 BUFX2_insert580 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf27)
);

BUFX2 BUFX2_insert579 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf28)
);

BUFX2 BUFX2_insert578 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf29)
);

BUFX2 BUFX2_insert577 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf30)
);

BUFX2 BUFX2_insert576 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf31)
);

BUFX2 BUFX2_insert575 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf32)
);

BUFX2 BUFX2_insert574 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf33)
);

BUFX2 BUFX2_insert573 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf34)
);

BUFX2 BUFX2_insert572 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf35)
);

BUFX2 BUFX2_insert571 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf36)
);

BUFX2 BUFX2_insert570 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf37)
);

BUFX2 BUFX2_insert569 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf38)
);

BUFX2 BUFX2_insert568 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf39)
);

BUFX2 BUFX2_insert567 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf40)
);

BUFX2 BUFX2_insert566 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf41)
);

BUFX2 BUFX2_insert565 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf42)
);

BUFX2 BUFX2_insert564 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf43)
);

BUFX2 BUFX2_insert563 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf44)
);

BUFX2 BUFX2_insert562 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf45)
);

BUFX2 BUFX2_insert561 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf46)
);

BUFX2 BUFX2_insert560 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf47)
);

BUFX2 BUFX2_insert559 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf48)
);

BUFX2 BUFX2_insert558 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf49)
);

BUFX2 BUFX2_insert557 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf50)
);

BUFX2 BUFX2_insert556 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf51)
);

BUFX2 BUFX2_insert555 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf52)
);

BUFX2 BUFX2_insert554 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf53)
);

BUFX2 BUFX2_insert553 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf54)
);

BUFX2 BUFX2_insert552 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf55)
);

BUFX2 BUFX2_insert551 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf56)
);

BUFX2 BUFX2_insert550 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf57)
);

BUFX2 BUFX2_insert549 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf58)
);

BUFX2 BUFX2_insert548 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf59)
);

BUFX2 BUFX2_insert547 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf60)
);

BUFX2 BUFX2_insert546 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf61)
);

BUFX2 BUFX2_insert545 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf62)
);

BUFX2 BUFX2_insert544 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf63)
);

BUFX2 BUFX2_insert543 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf64)
);

BUFX2 BUFX2_insert542 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf65)
);

BUFX2 BUFX2_insert541 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf66)
);

BUFX2 BUFX2_insert540 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf67)
);

BUFX2 BUFX2_insert539 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf68)
);

BUFX2 BUFX2_insert538 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf69)
);

BUFX2 BUFX2_insert537 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf70)
);

BUFX2 BUFX2_insert536 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf71)
);

BUFX2 BUFX2_insert535 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf72)
);

BUFX2 BUFX2_insert534 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf73)
);

BUFX2 BUFX2_insert533 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf74)
);

BUFX2 BUFX2_insert532 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf75)
);

BUFX2 BUFX2_insert531 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf76)
);

BUFX2 BUFX2_insert530 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf77)
);

BUFX2 BUFX2_insert529 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf78)
);

BUFX2 BUFX2_insert528 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf79)
);

BUFX2 BUFX2_insert527 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf80)
);

BUFX2 BUFX2_insert526 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf81)
);

BUFX2 BUFX2_insert525 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf82)
);

BUFX2 BUFX2_insert524 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf83)
);

BUFX2 BUFX2_insert523 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf84)
);

BUFX2 BUFX2_insert522 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf85)
);

BUFX2 BUFX2_insert521 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf86)
);

BUFX2 BUFX2_insert520 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf87)
);

BUFX2 BUFX2_insert519 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf88)
);

BUFX2 BUFX2_insert518 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf89)
);

BUFX2 BUFX2_insert517 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf90)
);

BUFX2 BUFX2_insert516 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf91)
);

BUFX2 BUFX2_insert515 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf92)
);

BUFX2 BUFX2_insert514 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf93)
);

BUFX2 BUFX2_insert513 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf94)
);

BUFX2 BUFX2_insert512 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf95)
);

BUFX2 BUFX2_insert511 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf96)
);

BUFX2 BUFX2_insert510 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf97)
);

BUFX2 BUFX2_insert509 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf98)
);

BUFX2 BUFX2_insert508 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf99)
);

BUFX2 BUFX2_insert507 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf100)
);

BUFX2 BUFX2_insert506 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf101)
);

BUFX2 BUFX2_insert505 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf102)
);

BUFX2 BUFX2_insert504 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf103)
);

BUFX2 BUFX2_insert503 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf5),
    .Y(rst_bF$buf104)
);

BUFX2 BUFX2_insert502 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf4),
    .Y(rst_bF$buf105)
);

BUFX2 BUFX2_insert501 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf3),
    .Y(rst_bF$buf106)
);

BUFX2 BUFX2_insert500 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf2),
    .Y(rst_bF$buf107)
);

BUFX2 BUFX2_insert499 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf1),
    .Y(rst_bF$buf108)
);

BUFX2 BUFX2_insert498 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf0),
    .Y(rst_bF$buf109)
);

BUFX2 BUFX2_insert497 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf9),
    .Y(rst_bF$buf110)
);

BUFX2 BUFX2_insert496 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf8),
    .Y(rst_bF$buf111)
);

BUFX2 BUFX2_insert495 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf7),
    .Y(rst_bF$buf112)
);

BUFX2 BUFX2_insert494 (
    .gnd(gnd),
    .vdd(vdd),
    .A(rst_hier0_bF$buf6),
    .Y(rst_bF$buf113)
);

BUFX2 BUFX2_insert493 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983_),
    .Y(_3983__bF$buf0)
);

BUFX2 BUFX2_insert492 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983_),
    .Y(_3983__bF$buf1)
);

BUFX2 BUFX2_insert491 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983_),
    .Y(_3983__bF$buf2)
);

BUFX2 BUFX2_insert490 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983_),
    .Y(_3983__bF$buf3)
);

BUFX2 BUFX2_insert489 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983_),
    .Y(_3983__bF$buf4)
);

BUFX2 BUFX2_insert488 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf0 )
);

BUFX2 BUFX2_insert487 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf1 )
);

BUFX2 BUFX2_insert486 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf2 )
);

BUFX2 BUFX2_insert485 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf3 )
);

BUFX2 BUFX2_insert484 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [9]),
    .Y(\datapath_1.mux_wd3.dout_9_bF$buf4 )
);

BUFX2 BUFX2_insert483 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459_),
    .Y(_5459__bF$buf0)
);

BUFX2 BUFX2_insert482 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459_),
    .Y(_5459__bF$buf1)
);

BUFX2 BUFX2_insert481 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459_),
    .Y(_5459__bF$buf2)
);

BUFX2 BUFX2_insert480 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459_),
    .Y(_5459__bF$buf3)
);

BUFX2 BUFX2_insert479 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518_),
    .Y(_5518__bF$buf0)
);

BUFX2 BUFX2_insert478 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518_),
    .Y(_5518__bF$buf1)
);

BUFX2 BUFX2_insert477 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518_),
    .Y(_5518__bF$buf2)
);

BUFX2 BUFX2_insert476 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518_),
    .Y(_5518__bF$buf3)
);

BUFX2 BUFX2_insert475 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5521_),
    .Y(_5521__bF$buf0)
);

BUFX2 BUFX2_insert474 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5521_),
    .Y(_5521__bF$buf1)
);

BUFX2 BUFX2_insert473 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5521_),
    .Y(_5521__bF$buf2)
);

BUFX2 BUFX2_insert472 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5521_),
    .Y(_5521__bF$buf3)
);

BUFX2 BUFX2_insert471 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf0 )
);

BUFX2 BUFX2_insert470 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf1 )
);

BUFX2 BUFX2_insert469 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf2 )
);

BUFX2 BUFX2_insert468 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf3 )
);

BUFX2 BUFX2_insert467 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf4 )
);

BUFX2 BUFX2_insert466 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf5 )
);

BUFX2 BUFX2_insert465 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf6 )
);

BUFX2 BUFX2_insert464 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [12]),
    .Y(\datapath_1.regfile_1.regEn_12_bF$buf7 )
);

BUFX2 BUFX2_insert463 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524_),
    .Y(_5524__bF$buf0)
);

BUFX2 BUFX2_insert462 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524_),
    .Y(_5524__bF$buf1)
);

BUFX2 BUFX2_insert461 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524_),
    .Y(_5524__bF$buf2)
);

BUFX2 BUFX2_insert460 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524_),
    .Y(_5524__bF$buf3)
);

BUFX2 BUFX2_insert459 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .Y(_3954__bF$buf0)
);

BUFX2 BUFX2_insert458 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .Y(_3954__bF$buf1)
);

BUFX2 BUFX2_insert457 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .Y(_3954__bF$buf2)
);

BUFX2 BUFX2_insert456 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .Y(_3954__bF$buf3)
);

BUFX2 BUFX2_insert455 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .Y(_3954__bF$buf4)
);

BUFX2 BUFX2_insert454 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf0 )
);

BUFX2 BUFX2_insert453 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf1 )
);

BUFX2 BUFX2_insert452 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf2 )
);

BUFX2 BUFX2_insert451 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf3 )
);

BUFX2 BUFX2_insert450 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf4 )
);

BUFX2 BUFX2_insert449 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf5 )
);

BUFX2 BUFX2_insert448 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf6 )
);

BUFX2 BUFX2_insert447 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [3]),
    .Y(\datapath_1.regfile_1.regEn_3_bF$buf7 )
);

BUFX2 BUFX2_insert446 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf0 )
);

BUFX2 BUFX2_insert445 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf1 )
);

BUFX2 BUFX2_insert444 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf2 )
);

BUFX2 BUFX2_insert443 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf3 )
);

BUFX2 BUFX2_insert442 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [11]),
    .Y(\datapath_1.mux_wd3.dout_11_bF$buf4 )
);

BUFX2 BUFX2_insert441 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565_),
    .Y(_5565__bF$buf0)
);

BUFX2 BUFX2_insert440 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565_),
    .Y(_5565__bF$buf1)
);

BUFX2 BUFX2_insert439 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565_),
    .Y(_5565__bF$buf2)
);

BUFX2 BUFX2_insert438 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565_),
    .Y(_5565__bF$buf3)
);

BUFX2 BUFX2_insert437 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf0 )
);

BUFX2 BUFX2_insert436 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf1 )
);

BUFX2 BUFX2_insert435 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf2 )
);

BUFX2 BUFX2_insert434 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf3 )
);

BUFX2 BUFX2_insert433 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf4 )
);

BUFX2 BUFX2_insert432 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf5 )
);

BUFX2 BUFX2_insert431 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf6 )
);

BUFX2 BUFX2_insert430 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [15]),
    .Y(\datapath_1.regfile_1.regEn_15_bF$buf7 )
);

BUFX2 BUFX2_insert429 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527_),
    .Y(_5527__bF$buf0)
);

BUFX2 BUFX2_insert428 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527_),
    .Y(_5527__bF$buf1)
);

BUFX2 BUFX2_insert427 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527_),
    .Y(_5527__bF$buf2)
);

BUFX2 BUFX2_insert426 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527_),
    .Y(_5527__bF$buf3)
);

BUFX2 BUFX2_insert425 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527_),
    .Y(_5527__bF$buf4)
);

BUFX2 BUFX2_insert424 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5471_),
    .Y(_5471__bF$buf0)
);

BUFX2 BUFX2_insert423 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5471_),
    .Y(_5471__bF$buf1)
);

BUFX2 BUFX2_insert422 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5471_),
    .Y(_5471__bF$buf2)
);

BUFX2 BUFX2_insert421 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5471_),
    .Y(_5471__bF$buf3)
);

BUFX2 BUFX2_insert420 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5471_),
    .Y(_5471__bF$buf4)
);

BUFX2 BUFX2_insert419 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5471_),
    .Y(_5471__bF$buf5)
);

BUFX2 BUFX2_insert418 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .Y(_5530__bF$buf0)
);

BUFX2 BUFX2_insert417 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .Y(_5530__bF$buf1)
);

BUFX2 BUFX2_insert416 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .Y(_5530__bF$buf2)
);

BUFX2 BUFX2_insert415 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .Y(_5530__bF$buf3)
);

BUFX2 BUFX2_insert414 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995_),
    .Y(_3995__bF$buf0)
);

BUFX2 BUFX2_insert413 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995_),
    .Y(_3995__bF$buf1)
);

BUFX2 BUFX2_insert412 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995_),
    .Y(_3995__bF$buf2)
);

BUFX2 BUFX2_insert411 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995_),
    .Y(_3995__bF$buf3)
);

BUFX2 BUFX2_insert410 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995_),
    .Y(_3995__bF$buf4)
);

BUFX2 BUFX2_insert409 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf0)
);

BUFX2 BUFX2_insert408 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf1)
);

BUFX2 BUFX2_insert407 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf2)
);

BUFX2 BUFX2_insert406 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf3)
);

BUFX2 BUFX2_insert405 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf4)
);

BUFX2 BUFX2_insert404 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf5)
);

BUFX2 BUFX2_insert403 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf6)
);

BUFX2 BUFX2_insert402 (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg),
    .Y(MemToReg_bF$buf7)
);

BUFX2 BUFX2_insert401 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf0 )
);

BUFX2 BUFX2_insert400 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf1 )
);

BUFX2 BUFX2_insert399 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf2 )
);

BUFX2 BUFX2_insert398 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf3 )
);

BUFX2 BUFX2_insert397 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf4 )
);

BUFX2 BUFX2_insert396 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf5 )
);

BUFX2 BUFX2_insert395 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf6 )
);

BUFX2 BUFX2_insert394 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [6]),
    .Y(\datapath_1.regfile_1.regEn_6_bF$buf7 )
);

BUFX2 BUFX2_insert393 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf0 )
);

BUFX2 BUFX2_insert392 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf1 )
);

BUFX2 BUFX2_insert391 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf2 )
);

BUFX2 BUFX2_insert390 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf3 )
);

BUFX2 BUFX2_insert389 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [14]),
    .Y(\datapath_1.mux_wd3.dout_14_bF$buf4 )
);

BUFX2 BUFX2_insert388 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf0 )
);

BUFX2 BUFX2_insert387 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf1 )
);

BUFX2 BUFX2_insert386 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf2 )
);

BUFX2 BUFX2_insert385 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf3 )
);

BUFX2 BUFX2_insert384 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf4 )
);

BUFX2 BUFX2_insert383 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf5 )
);

BUFX2 BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf6 )
);

BUFX2 BUFX2_insert381 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [18]),
    .Y(\datapath_1.regfile_1.regEn_18_bF$buf7 )
);

BUFX2 BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3196_),
    .Y(_3196__bF$buf0)
);

BUFX2 BUFX2_insert379 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3196_),
    .Y(_3196__bF$buf1)
);

BUFX2 BUFX2_insert378 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3196_),
    .Y(_3196__bF$buf2)
);

BUFX2 BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3196_),
    .Y(_3196__bF$buf3)
);

BUFX2 BUFX2_insert376 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3196_),
    .Y(_3196__bF$buf4)
);

BUFX2 BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf0 )
);

BUFX2 BUFX2_insert374 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf1 )
);

BUFX2 BUFX2_insert373 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf2 )
);

BUFX2 BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf3 )
);

BUFX2 BUFX2_insert371 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf4 )
);

BUFX2 BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf5 )
);

BUFX2 BUFX2_insert369 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf6 )
);

BUFX2 BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [21]),
    .Y(\datapath_1.regfile_1.regEn_21_bF$buf7 )
);

BUFX2 BUFX2_insert367 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3998_),
    .Y(_3998__bF$buf0)
);

BUFX2 BUFX2_insert366 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3998_),
    .Y(_3998__bF$buf1)
);

BUFX2 BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3998_),
    .Y(_3998__bF$buf2)
);

BUFX2 BUFX2_insert364 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3998_),
    .Y(_3998__bF$buf3)
);

BUFX2 BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .Y(_2470__bF$buf0)
);

BUFX2 BUFX2_insert362 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .Y(_2470__bF$buf1)
);

BUFX2 BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .Y(_2470__bF$buf2)
);

BUFX2 BUFX2_insert360 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .Y(_2470__bF$buf3)
);

BUFX2 BUFX2_insert359 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf0 )
);

BUFX2 BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf1 )
);

BUFX2 BUFX2_insert357 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf2 )
);

BUFX2 BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf3 )
);

BUFX2 BUFX2_insert355 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf4 )
);

BUFX2 BUFX2_insert354 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf5 )
);

BUFX2 BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf6 )
);

BUFX2 BUFX2_insert352 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [9]),
    .Y(\datapath_1.regfile_1.regEn_9_bF$buf7 )
);

BUFX2 BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf0)
);

BUFX2 BUFX2_insert350 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf1)
);

BUFX2 BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf2)
);

BUFX2 BUFX2_insert348 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf3)
);

BUFX2 BUFX2_insert347 (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB[0]),
    .Y(ALUSrcB_0_bF$buf4)
);

BUFX2 BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf0 )
);

BUFX2 BUFX2_insert345 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf1 )
);

BUFX2 BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf2 )
);

BUFX2 BUFX2_insert343 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf3 )
);

BUFX2 BUFX2_insert342 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [17]),
    .Y(\datapath_1.mux_wd3.dout_17_bF$buf4 )
);

BUFX2 BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf0 )
);

BUFX2 BUFX2_insert340 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf1 )
);

BUFX2 BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf2 )
);

BUFX2 BUFX2_insert338 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [22]),
    .Y(\datapath_1.PCJump_22_bF$buf3 )
);

BUFX2 BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4005_),
    .Y(_4005__bF$buf0)
);

BUFX2 BUFX2_insert336 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4005_),
    .Y(_4005__bF$buf1)
);

BUFX2 BUFX2_insert335 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4005_),
    .Y(_4005__bF$buf2)
);

BUFX2 BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4005_),
    .Y(_4005__bF$buf3)
);

BUFX2 BUFX2_insert333 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf0 )
);

BUFX2 BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf1 )
);

BUFX2 BUFX2_insert331 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf2 )
);

BUFX2 BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf3 )
);

BUFX2 BUFX2_insert329 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [20]),
    .Y(\datapath_1.mux_wd3.dout_20_bF$buf4 )
);

BUFX2 BUFX2_insert328 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf0 )
);

BUFX2 BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf1 )
);

BUFX2 BUFX2_insert326 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf2 )
);

BUFX2 BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf3 )
);

BUFX2 BUFX2_insert324 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf4 )
);

BUFX2 BUFX2_insert323 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf5 )
);

BUFX2 BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf6 )
);

BUFX2 BUFX2_insert321 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [24]),
    .Y(\datapath_1.regfile_1.regEn_24_bF$buf7 )
);

BUFX2 BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf0)
);

BUFX2 BUFX2_insert319 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf1)
);

BUFX2 BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf2)
);

BUFX2 BUFX2_insert317 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf3)
);

BUFX2 BUFX2_insert316 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3966_),
    .Y(_3966__bF$buf0)
);

BUFX2 BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3966_),
    .Y(_3966__bF$buf1)
);

BUFX2 BUFX2_insert314 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3966_),
    .Y(_3966__bF$buf2)
);

BUFX2 BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3966_),
    .Y(_3966__bF$buf3)
);

BUFX2 BUFX2_insert312 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .Y(_2341__bF$buf0)
);

BUFX2 BUFX2_insert311 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .Y(_2341__bF$buf1)
);

BUFX2 BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .Y(_2341__bF$buf2)
);

BUFX2 BUFX2_insert309 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .Y(_2341__bF$buf3)
);

BUFX2 BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .Y(_3032__bF$buf0)
);

BUFX2 BUFX2_insert307 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .Y(_3032__bF$buf1)
);

BUFX2 BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .Y(_3032__bF$buf2)
);

BUFX2 BUFX2_insert305 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .Y(_3032__bF$buf3)
);

BUFX2 BUFX2_insert304 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .Y(_3032__bF$buf4)
);

BUFX2 BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf0 )
);

BUFX2 BUFX2_insert302 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf1 )
);

BUFX2 BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf2 )
);

BUFX2 BUFX2_insert300 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf3 )
);

BUFX2 BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [23]),
    .Y(\datapath_1.mux_wd3.dout_23_bF$buf4 )
);

BUFX2 BUFX2_insert298 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf0 )
);

BUFX2 BUFX2_insert297 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf1 )
);

BUFX2 BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf2 )
);

BUFX2 BUFX2_insert295 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf3 )
);

BUFX2 BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf4 )
);

BUFX2 BUFX2_insert293 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf5 )
);

BUFX2 BUFX2_insert292 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf6 )
);

BUFX2 BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [27]),
    .Y(\datapath_1.regfile_1.regEn_27_bF$buf7 )
);

BUFX2 BUFX2_insert290 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .Y(_5539__bF$buf0)
);

BUFX2 BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .Y(_5539__bF$buf1)
);

BUFX2 BUFX2_insert288 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .Y(_5539__bF$buf2)
);

BUFX2 BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .Y(_5539__bF$buf3)
);

BUFX2 BUFX2_insert286 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .Y(_5539__bF$buf4)
);

BUFX2 BUFX2_insert285 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .Y(_5483__bF$buf0)
);

BUFX2 BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .Y(_5483__bF$buf1)
);

BUFX2 BUFX2_insert283 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .Y(_5483__bF$buf2)
);

BUFX2 BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .Y(_5483__bF$buf3)
);

BUFX2 BUFX2_insert281 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .Y(_5483__bF$buf4)
);

BUFX2 BUFX2_insert280 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .Y(_3931__bF$buf0)
);

BUFX2 BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .Y(_3931__bF$buf1)
);

BUFX2 BUFX2_insert278 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .Y(_3931__bF$buf2)
);

BUFX2 BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .Y(_3931__bF$buf3)
);

BUFX2 BUFX2_insert276 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf0 )
);

BUFX2 BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf1 )
);

BUFX2 BUFX2_insert274 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf2 )
);

BUFX2 BUFX2_insert273 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf3 )
);

BUFX2 BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf4 )
);

BUFX2 BUFX2_insert271 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf5 )
);

BUFX2 BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf6 )
);

BUFX2 BUFX2_insert269 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [30]),
    .Y(\datapath_1.regfile_1.regEn_30_bF$buf7 )
);

BUFX2 BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .Y(_5504__bF$buf0)
);

BUFX2 BUFX2_insert267 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .Y(_5504__bF$buf1)
);

BUFX2 BUFX2_insert266 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .Y(_5504__bF$buf2)
);

BUFX2 BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .Y(_5504__bF$buf3)
);

BUFX2 BUFX2_insert264 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .Y(_5504__bF$buf4)
);

BUFX2 BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344_),
    .Y(_2344__bF$buf0)
);

BUFX2 BUFX2_insert262 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344_),
    .Y(_2344__bF$buf1)
);

BUFX2 BUFX2_insert261 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344_),
    .Y(_2344__bF$buf2)
);

BUFX2 BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344_),
    .Y(_2344__bF$buf3)
);

BUFX2 BUFX2_insert259 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf0 )
);

BUFX2 BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf1 )
);

BUFX2 BUFX2_insert257 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf2 )
);

BUFX2 BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf3 )
);

BUFX2 BUFX2_insert255 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [26]),
    .Y(\datapath_1.mux_wd3.dout_26_bF$buf4 )
);

BUFX2 BUFX2_insert254 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf0)
);

BUFX2 BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf1)
);

BUFX2 BUFX2_insert252 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf2)
);

BUFX2 BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf3)
);

BUFX2 BUFX2_insert250 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf4)
);

BUFX2 BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf5)
);

BUFX2 BUFX2_insert248 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf6)
);

BUFX2 BUFX2_insert247 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite),
    .Y(RegWrite_bF$buf7)
);

BUFX2 BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972_),
    .Y(_3972__bF$buf0)
);

BUFX2 BUFX2_insert245 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972_),
    .Y(_3972__bF$buf1)
);

BUFX2 BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972_),
    .Y(_3972__bF$buf2)
);

BUFX2 BUFX2_insert243 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972_),
    .Y(_3972__bF$buf3)
);

BUFX2 BUFX2_insert242 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf0)
);

BUFX2 BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf1)
);

BUFX2 BUFX2_insert240 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf2)
);

BUFX2 BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf3)
);

BUFX2 BUFX2_insert238 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf0 )
);

BUFX2 BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf1 )
);

BUFX2 BUFX2_insert236 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf2 )
);

BUFX2 BUFX2_insert235 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf3 )
);

BUFX2 BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [1]),
    .Y(\datapath_1.mux_wd3.dout_1_bF$buf4 )
);

BUFX2 BUFX2_insert233 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347_),
    .Y(_2347__bF$buf0)
);

BUFX2 BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347_),
    .Y(_2347__bF$buf1)
);

BUFX2 BUFX2_insert231 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347_),
    .Y(_2347__bF$buf2)
);

BUFX2 BUFX2_insert230 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347_),
    .Y(_2347__bF$buf3)
);

BUFX2 BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf0 )
);

BUFX2 BUFX2_insert228 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf1 )
);

BUFX2 BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf2 )
);

BUFX2 BUFX2_insert226 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf3 )
);

BUFX2 BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [29]),
    .Y(\datapath_1.mux_wd3.dout_29_bF$buf4 )
);

CLKBUF1 CLKBUF1_insert224 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert223 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert222 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert221 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert220 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert219 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert218 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert217 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert216 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert215 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert214 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert213 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert212 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf12)
);

CLKBUF1 CLKBUF1_insert211 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf13)
);

CLKBUF1 CLKBUF1_insert210 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf14)
);

CLKBUF1 CLKBUF1_insert209 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf15)
);

CLKBUF1 CLKBUF1_insert208 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf16)
);

CLKBUF1 CLKBUF1_insert207 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf17)
);

CLKBUF1 CLKBUF1_insert206 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf18)
);

CLKBUF1 CLKBUF1_insert205 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf19)
);

CLKBUF1 CLKBUF1_insert204 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf20)
);

CLKBUF1 CLKBUF1_insert203 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf21)
);

CLKBUF1 CLKBUF1_insert202 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf22)
);

CLKBUF1 CLKBUF1_insert201 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf23)
);

CLKBUF1 CLKBUF1_insert200 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf24)
);

CLKBUF1 CLKBUF1_insert199 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf25)
);

CLKBUF1 CLKBUF1_insert198 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf26)
);

CLKBUF1 CLKBUF1_insert197 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf27)
);

CLKBUF1 CLKBUF1_insert196 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf28)
);

CLKBUF1 CLKBUF1_insert195 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf29)
);

CLKBUF1 CLKBUF1_insert194 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf30)
);

CLKBUF1 CLKBUF1_insert193 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf31)
);

CLKBUF1 CLKBUF1_insert192 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf32)
);

CLKBUF1 CLKBUF1_insert191 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf33)
);

CLKBUF1 CLKBUF1_insert190 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf34)
);

CLKBUF1 CLKBUF1_insert189 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf35)
);

CLKBUF1 CLKBUF1_insert188 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf36)
);

CLKBUF1 CLKBUF1_insert187 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf37)
);

CLKBUF1 CLKBUF1_insert186 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf38)
);

CLKBUF1 CLKBUF1_insert185 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf39)
);

CLKBUF1 CLKBUF1_insert184 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf40)
);

CLKBUF1 CLKBUF1_insert183 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf41)
);

CLKBUF1 CLKBUF1_insert182 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf42)
);

CLKBUF1 CLKBUF1_insert181 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf43)
);

CLKBUF1 CLKBUF1_insert180 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf44)
);

CLKBUF1 CLKBUF1_insert179 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf45)
);

CLKBUF1 CLKBUF1_insert178 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf46)
);

CLKBUF1 CLKBUF1_insert177 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf47)
);

CLKBUF1 CLKBUF1_insert176 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf48)
);

CLKBUF1 CLKBUF1_insert175 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf49)
);

CLKBUF1 CLKBUF1_insert174 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf50)
);

CLKBUF1 CLKBUF1_insert173 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf51)
);

CLKBUF1 CLKBUF1_insert172 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf52)
);

CLKBUF1 CLKBUF1_insert171 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf53)
);

CLKBUF1 CLKBUF1_insert170 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf54)
);

CLKBUF1 CLKBUF1_insert169 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf55)
);

CLKBUF1 CLKBUF1_insert168 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf56)
);

CLKBUF1 CLKBUF1_insert167 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf57)
);

CLKBUF1 CLKBUF1_insert166 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf58)
);

CLKBUF1 CLKBUF1_insert165 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf59)
);

CLKBUF1 CLKBUF1_insert164 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf60)
);

CLKBUF1 CLKBUF1_insert163 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf61)
);

CLKBUF1 CLKBUF1_insert162 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf62)
);

CLKBUF1 CLKBUF1_insert161 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf63)
);

CLKBUF1 CLKBUF1_insert160 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf64)
);

CLKBUF1 CLKBUF1_insert159 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf65)
);

CLKBUF1 CLKBUF1_insert158 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf66)
);

CLKBUF1 CLKBUF1_insert157 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf67)
);

CLKBUF1 CLKBUF1_insert156 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf68)
);

CLKBUF1 CLKBUF1_insert155 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf69)
);

CLKBUF1 CLKBUF1_insert154 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf70)
);

CLKBUF1 CLKBUF1_insert153 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf71)
);

CLKBUF1 CLKBUF1_insert152 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf72)
);

CLKBUF1 CLKBUF1_insert151 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf73)
);

CLKBUF1 CLKBUF1_insert150 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf74)
);

CLKBUF1 CLKBUF1_insert149 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf75)
);

CLKBUF1 CLKBUF1_insert148 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf76)
);

CLKBUF1 CLKBUF1_insert147 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf77)
);

CLKBUF1 CLKBUF1_insert146 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf78)
);

CLKBUF1 CLKBUF1_insert145 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf79)
);

CLKBUF1 CLKBUF1_insert144 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf80)
);

CLKBUF1 CLKBUF1_insert143 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf81)
);

CLKBUF1 CLKBUF1_insert142 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf82)
);

CLKBUF1 CLKBUF1_insert141 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf83)
);

CLKBUF1 CLKBUF1_insert140 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf84)
);

CLKBUF1 CLKBUF1_insert139 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf85)
);

CLKBUF1 CLKBUF1_insert138 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf86)
);

CLKBUF1 CLKBUF1_insert137 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf87)
);

CLKBUF1 CLKBUF1_insert136 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf88)
);

CLKBUF1 CLKBUF1_insert135 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf89)
);

CLKBUF1 CLKBUF1_insert134 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf90)
);

CLKBUF1 CLKBUF1_insert133 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf91)
);

CLKBUF1 CLKBUF1_insert132 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf92)
);

CLKBUF1 CLKBUF1_insert131 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf93)
);

CLKBUF1 CLKBUF1_insert130 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf94)
);

CLKBUF1 CLKBUF1_insert129 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf95)
);

CLKBUF1 CLKBUF1_insert128 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf96)
);

CLKBUF1 CLKBUF1_insert127 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf97)
);

CLKBUF1 CLKBUF1_insert126 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf98)
);

CLKBUF1 CLKBUF1_insert125 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf99)
);

CLKBUF1 CLKBUF1_insert124 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf100)
);

CLKBUF1 CLKBUF1_insert123 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf101)
);

CLKBUF1 CLKBUF1_insert122 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf102)
);

CLKBUF1 CLKBUF1_insert121 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf103)
);

CLKBUF1 CLKBUF1_insert120 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf5),
    .Y(clk_bF$buf104)
);

CLKBUF1 CLKBUF1_insert119 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf4),
    .Y(clk_bF$buf105)
);

CLKBUF1 CLKBUF1_insert118 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf3),
    .Y(clk_bF$buf106)
);

CLKBUF1 CLKBUF1_insert117 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf2),
    .Y(clk_bF$buf107)
);

CLKBUF1 CLKBUF1_insert116 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf1),
    .Y(clk_bF$buf108)
);

CLKBUF1 CLKBUF1_insert115 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf0),
    .Y(clk_bF$buf109)
);

CLKBUF1 CLKBUF1_insert114 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf9),
    .Y(clk_bF$buf110)
);

CLKBUF1 CLKBUF1_insert113 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf8),
    .Y(clk_bF$buf111)
);

CLKBUF1 CLKBUF1_insert112 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf7),
    .Y(clk_bF$buf112)
);

CLKBUF1 CLKBUF1_insert111 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk_hier0_bF$buf6),
    .Y(clk_bF$buf113)
);

BUFX2 BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf0)
);

BUFX2 BUFX2_insert109 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf1)
);

BUFX2 BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf2)
);

BUFX2 BUFX2_insert107 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf3)
);

BUFX2 BUFX2_insert106 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf4)
);

BUFX2 BUFX2_insert105 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf5)
);

BUFX2 BUFX2_insert104 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf6)
);

BUFX2 BUFX2_insert103 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD),
    .Y(IorD_bF$buf7)
);

BUFX2 BUFX2_insert102 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489_),
    .Y(_5489__bF$buf0)
);

BUFX2 BUFX2_insert101 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489_),
    .Y(_5489__bF$buf1)
);

BUFX2 BUFX2_insert100 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489_),
    .Y(_5489__bF$buf2)
);

BUFX2 BUFX2_insert99 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489_),
    .Y(_5489__bF$buf3)
);

BUFX2 BUFX2_insert98 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5548_),
    .Y(_5548__bF$buf0)
);

BUFX2 BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5548_),
    .Y(_5548__bF$buf1)
);

BUFX2 BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5548_),
    .Y(_5548__bF$buf2)
);

BUFX2 BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5548_),
    .Y(_5548__bF$buf3)
);

BUFX2 BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5548_),
    .Y(_5548__bF$buf4)
);

BUFX2 BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf0 )
);

BUFX2 BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf1 )
);

BUFX2 BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf2 )
);

BUFX2 BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf3 )
);

BUFX2 BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [4]),
    .Y(\datapath_1.mux_wd3.dout_4_bF$buf4 )
);

BUFX2 BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .Y(_3902__bF$buf0)
);

BUFX2 BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .Y(_3902__bF$buf1)
);

BUFX2 BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .Y(_3902__bF$buf2)
);

BUFX2 BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .Y(_3902__bF$buf3)
);

BUFX2 BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884_),
    .Y(_3884__bF$buf0)
);

BUFX2 BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884_),
    .Y(_3884__bF$buf1)
);

BUFX2 BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884_),
    .Y(_3884__bF$buf2)
);

BUFX2 BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884_),
    .Y(_3884__bF$buf3)
);

BUFX2 BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495_),
    .Y(_5495__bF$buf0)
);

BUFX2 BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495_),
    .Y(_5495__bF$buf1)
);

BUFX2 BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495_),
    .Y(_5495__bF$buf2)
);

BUFX2 BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495_),
    .Y(_5495__bF$buf3)
);

BUFX2 BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf0 )
);

BUFX2 BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf1 )
);

BUFX2 BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf2 )
);

BUFX2 BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf3 )
);

BUFX2 BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [7]),
    .Y(\datapath_1.mux_wd3.dout_7_bF$buf4 )
);

BUFX2 BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905_),
    .Y(_3905__bF$buf0)
);

BUFX2 BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905_),
    .Y(_3905__bF$buf1)
);

BUFX2 BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905_),
    .Y(_3905__bF$buf2)
);

BUFX2 BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905_),
    .Y(_3905__bF$buf3)
);

BUFX2 BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .Y(_3200__bF$buf0)
);

BUFX2 BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .Y(_3200__bF$buf1)
);

BUFX2 BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .Y(_3200__bF$buf2)
);

BUFX2 BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .Y(_3200__bF$buf3)
);

BUFX2 BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .Y(_3200__bF$buf4)
);

BUFX2 BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463_),
    .Y(_5463__bF$buf0)
);

BUFX2 BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463_),
    .Y(_5463__bF$buf1)
);

BUFX2 BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463_),
    .Y(_5463__bF$buf2)
);

BUFX2 BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463_),
    .Y(_5463__bF$buf3)
);

BUFX2 BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf0 )
);

BUFX2 BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf1 )
);

BUFX2 BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf2 )
);

BUFX2 BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf3 )
);

BUFX2 BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf4 )
);

BUFX2 BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf5 )
);

BUFX2 BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf6 )
);

BUFX2 BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [10]),
    .Y(\datapath_1.regfile_1.regEn_10_bF$buf7 )
);

BUFX2 BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893_),
    .Y(_3893__bF$buf0)
);

BUFX2 BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893_),
    .Y(_3893__bF$buf1)
);

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893_),
    .Y(_3893__bF$buf2)
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893_),
    .Y(_3893__bF$buf3)
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf0)
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf4)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf0 )
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf1 )
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf2 )
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf3 )
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf4 )
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf5 )
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf6 )
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [1]),
    .Y(\datapath_1.regfile_1.regEn_1_bF$buf7 )
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf0 )
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf1 )
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf2 )
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf3 )
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf4 )
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf5 )
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf6 )
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [13]),
    .Y(\datapath_1.regfile_1.regEn_13_bF$buf7 )
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .Y(_2462__bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .Y(_2462__bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .Y(_2462__bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .Y(_2462__bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3955_),
    .Y(_3955__bF$buf0)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3955_),
    .Y(_3955__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3955_),
    .Y(_3955__bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3955_),
    .Y(_3955__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3955_),
    .Y(_3955__bF$buf4)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5469_),
    .Y(_5469__bF$buf0)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5469_),
    .Y(_5469__bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5469_),
    .Y(_5469__bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5469_),
    .Y(_5469__bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf0 )
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf1 )
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf2 )
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf3 )
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf4 )
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf5 )
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf6 )
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn [4]),
    .Y(\datapath_1.regfile_1.regEn_4_bF$buf7 )
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf0 )
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf1 )
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf2 )
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf3 )
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout [12]),
    .Y(\datapath_1.mux_wd3.dout_12_bF$buf4 )
);

OAI21X1 _10000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1578_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1579_),
    .Y(_1563_[8])
);

INVX1 _10001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_1580_)
);

NAND2X1 _10002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1581_)
);

OAI21X1 _10003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1580_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1581_),
    .Y(_1563_[9])
);

INVX1 _10004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_1582_)
);

NAND2X1 _10005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1583_)
);

OAI21X1 _10006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1583_),
    .Y(_1563_[10])
);

INVX1 _10007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_1584_)
);

NAND2X1 _10008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1585_)
);

OAI21X1 _10009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1584_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1585_),
    .Y(_1563_[11])
);

INVX1 _10010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_1586_)
);

NAND2X1 _10011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1587_)
);

OAI21X1 _10012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1586_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1587_),
    .Y(_1563_[12])
);

INVX1 _10013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_1588_)
);

NAND2X1 _10014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1589_)
);

OAI21X1 _10015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1589_),
    .Y(_1563_[13])
);

INVX1 _10016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_1590_)
);

NAND2X1 _10017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1591_)
);

OAI21X1 _10018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1591_),
    .Y(_1563_[14])
);

INVX1 _10019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_1592_)
);

NAND2X1 _10020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1593_)
);

OAI21X1 _10021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1593_),
    .Y(_1563_[15])
);

INVX1 _10022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_1594_)
);

NAND2X1 _10023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1595_)
);

OAI21X1 _10024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1594_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1595_),
    .Y(_1563_[16])
);

INVX1 _10025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_1596_)
);

NAND2X1 _10026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1597_)
);

OAI21X1 _10027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1597_),
    .Y(_1563_[17])
);

INVX1 _10028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_1598_)
);

NAND2X1 _10029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1599_)
);

OAI21X1 _10030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1599_),
    .Y(_1563_[18])
);

INVX1 _10031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_1600_)
);

NAND2X1 _10032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1601_)
);

OAI21X1 _10033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1600_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1601_),
    .Y(_1563_[19])
);

INVX1 _10034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_1602_)
);

NAND2X1 _10035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1603_)
);

OAI21X1 _10036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1602_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1603_),
    .Y(_1563_[20])
);

INVX1 _10037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_1604_)
);

NAND2X1 _10038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1605_)
);

OAI21X1 _10039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1604_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1605_),
    .Y(_1563_[21])
);

INVX1 _10040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_1606_)
);

NAND2X1 _10041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1607_)
);

OAI21X1 _10042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1607_),
    .Y(_1563_[22])
);

INVX1 _10043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_1608_)
);

NAND2X1 _10044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1609_)
);

OAI21X1 _10045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1608_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1609_),
    .Y(_1563_[23])
);

INVX1 _10046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_1610_)
);

NAND2X1 _10047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1611_)
);

OAI21X1 _10048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1610_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1611_),
    .Y(_1563_[24])
);

INVX1 _10049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_1612_)
);

NAND2X1 _10050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1613_)
);

OAI21X1 _10051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1613_),
    .Y(_1563_[25])
);

INVX1 _10052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_1614_)
);

NAND2X1 _10053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1615_)
);

OAI21X1 _10054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1614_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1615_),
    .Y(_1563_[26])
);

INVX1 _10055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_1616_)
);

NAND2X1 _10056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1617_)
);

OAI21X1 _10057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1617_),
    .Y(_1563_[27])
);

INVX1 _10058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_1618_)
);

NAND2X1 _10059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1619_)
);

OAI21X1 _10060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1619_),
    .Y(_1563_[28])
);

INVX1 _10061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_1620_)
);

NAND2X1 _10062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1621_)
);

OAI21X1 _10063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1621_),
    .Y(_1563_[29])
);

INVX1 _10064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_1622_)
);

NAND2X1 _10065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1623_)
);

OAI21X1 _10066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1622_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1623_),
    .Y(_1563_[30])
);

INVX1 _10067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_1624_)
);

NAND2X1 _10068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1625_)
);

OAI21X1 _10069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1624_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1625_),
    .Y(_1563_[31])
);

DFFSR _10070_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_1563_[0]),
    .Q(\datapath_1.regfile_1.regOut[25] [0]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _10071_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_1563_[1]),
    .Q(\datapath_1.regfile_1.regOut[25] [1]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _10072_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_1563_[2]),
    .Q(\datapath_1.regfile_1.regOut[25] [2]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _10073_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_1563_[3]),
    .Q(\datapath_1.regfile_1.regOut[25] [3]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _10074_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_1563_[4]),
    .Q(\datapath_1.regfile_1.regOut[25] [4]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _10075_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_1563_[5]),
    .Q(\datapath_1.regfile_1.regOut[25] [5]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _10076_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_1563_[6]),
    .Q(\datapath_1.regfile_1.regOut[25] [6]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _10077_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_1563_[7]),
    .Q(\datapath_1.regfile_1.regOut[25] [7]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _10078_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_1563_[8]),
    .Q(\datapath_1.regfile_1.regOut[25] [8]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _10079_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_1563_[9]),
    .Q(\datapath_1.regfile_1.regOut[25] [9]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _10080_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_1563_[10]),
    .Q(\datapath_1.regfile_1.regOut[25] [10]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _10081_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_1563_[11]),
    .Q(\datapath_1.regfile_1.regOut[25] [11]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _10082_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_1563_[12]),
    .Q(\datapath_1.regfile_1.regOut[25] [12]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _10083_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_1563_[13]),
    .Q(\datapath_1.regfile_1.regOut[25] [13]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _10084_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_1563_[14]),
    .Q(\datapath_1.regfile_1.regOut[25] [14]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _10085_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_1563_[15]),
    .Q(\datapath_1.regfile_1.regOut[25] [15]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _10086_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_1563_[16]),
    .Q(\datapath_1.regfile_1.regOut[25] [16]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _10087_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_1563_[17]),
    .Q(\datapath_1.regfile_1.regOut[25] [17]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _10088_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_1563_[18]),
    .Q(\datapath_1.regfile_1.regOut[25] [18]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _10089_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_1563_[19]),
    .Q(\datapath_1.regfile_1.regOut[25] [19]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _10090_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_1563_[20]),
    .Q(\datapath_1.regfile_1.regOut[25] [20]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _10091_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_1563_[21]),
    .Q(\datapath_1.regfile_1.regOut[25] [21]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _10092_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_1563_[22]),
    .Q(\datapath_1.regfile_1.regOut[25] [22]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _10093_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_1563_[23]),
    .Q(\datapath_1.regfile_1.regOut[25] [23]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _10094_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_1563_[24]),
    .Q(\datapath_1.regfile_1.regOut[25] [24]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _10095_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_1563_[25]),
    .Q(\datapath_1.regfile_1.regOut[25] [25]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _10096_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_1563_[26]),
    .Q(\datapath_1.regfile_1.regOut[25] [26]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _10097_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_1563_[27]),
    .Q(\datapath_1.regfile_1.regOut[25] [27]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _10098_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_1563_[28]),
    .Q(\datapath_1.regfile_1.regOut[25] [28]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _10099_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_1563_[29]),
    .Q(\datapath_1.regfile_1.regOut[25] [29]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _10100_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_1563_[30]),
    .Q(\datapath_1.regfile_1.regOut[25] [30]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _10101_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_1563_[31]),
    .Q(\datapath_1.regfile_1.regOut[25] [31]),
    .R(rst_bF$buf82),
    .S(vdd)
);

INVX1 _10102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_1691_)
);

NAND2X1 _10103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .Y(_1692_)
);

OAI21X1 _10104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1691_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1692_),
    .Y(_1628_[0])
);

INVX1 _10105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_1629_)
);

NAND2X1 _10106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1630_)
);

OAI21X1 _10107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1629_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1630_),
    .Y(_1628_[1])
);

INVX1 _10108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_1631_)
);

NAND2X1 _10109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1632_)
);

OAI21X1 _10110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1631_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1632_),
    .Y(_1628_[2])
);

INVX1 _10111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_1633_)
);

NAND2X1 _10112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1634_)
);

OAI21X1 _10113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1633_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1634_),
    .Y(_1628_[3])
);

INVX1 _10114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_1635_)
);

NAND2X1 _10115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1636_)
);

OAI21X1 _10116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1635_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1636_),
    .Y(_1628_[4])
);

INVX1 _10117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_1637_)
);

NAND2X1 _10118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1638_)
);

OAI21X1 _10119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1637_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1638_),
    .Y(_1628_[5])
);

INVX1 _10120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_1639_)
);

NAND2X1 _10121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1640_)
);

OAI21X1 _10122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1639_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1640_),
    .Y(_1628_[6])
);

INVX1 _10123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_1641_)
);

NAND2X1 _10124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1642_)
);

OAI21X1 _10125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1641_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1642_),
    .Y(_1628_[7])
);

INVX1 _10126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_1643_)
);

NAND2X1 _10127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1644_)
);

OAI21X1 _10128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1644_),
    .Y(_1628_[8])
);

INVX1 _10129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_1645_)
);

NAND2X1 _10130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1646_)
);

OAI21X1 _10131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1645_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1646_),
    .Y(_1628_[9])
);

INVX1 _10132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_1647_)
);

NAND2X1 _10133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1648_)
);

OAI21X1 _10134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1648_),
    .Y(_1628_[10])
);

INVX1 _10135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_1649_)
);

NAND2X1 _10136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1650_)
);

OAI21X1 _10137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1650_),
    .Y(_1628_[11])
);

INVX1 _10138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_1651_)
);

NAND2X1 _10139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1652_)
);

OAI21X1 _10140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1652_),
    .Y(_1628_[12])
);

INVX1 _10141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_1653_)
);

NAND2X1 _10142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1654_)
);

OAI21X1 _10143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1654_),
    .Y(_1628_[13])
);

INVX1 _10144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_1655_)
);

NAND2X1 _10145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1656_)
);

OAI21X1 _10146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1655_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1656_),
    .Y(_1628_[14])
);

INVX1 _10147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_1657_)
);

NAND2X1 _10148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1658_)
);

OAI21X1 _10149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1658_),
    .Y(_1628_[15])
);

INVX1 _10150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_1659_)
);

NAND2X1 _10151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1660_)
);

OAI21X1 _10152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1660_),
    .Y(_1628_[16])
);

INVX1 _10153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_1661_)
);

NAND2X1 _10154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1662_)
);

OAI21X1 _10155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1662_),
    .Y(_1628_[17])
);

INVX1 _10156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_1663_)
);

NAND2X1 _10157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1664_)
);

OAI21X1 _10158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1663_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1664_),
    .Y(_1628_[18])
);

INVX1 _10159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_1665_)
);

NAND2X1 _10160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1666_)
);

OAI21X1 _10161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1665_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1666_),
    .Y(_1628_[19])
);

INVX1 _10162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_1667_)
);

NAND2X1 _10163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1668_)
);

OAI21X1 _10164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1667_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1668_),
    .Y(_1628_[20])
);

INVX1 _10165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_1669_)
);

NAND2X1 _10166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1670_)
);

OAI21X1 _10167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1669_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1670_),
    .Y(_1628_[21])
);

INVX1 _10168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_1671_)
);

NAND2X1 _10169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1672_)
);

OAI21X1 _10170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1671_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1672_),
    .Y(_1628_[22])
);

INVX1 _10171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_1673_)
);

NAND2X1 _10172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1674_)
);

OAI21X1 _10173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1674_),
    .Y(_1628_[23])
);

INVX1 _10174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_1675_)
);

NAND2X1 _10175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1676_)
);

OAI21X1 _10176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1676_),
    .Y(_1628_[24])
);

INVX1 _10177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_1677_)
);

NAND2X1 _10178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_1678_)
);

OAI21X1 _10179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1678_),
    .Y(_1628_[25])
);

INVX1 _10180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_1679_)
);

NAND2X1 _10181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1680_)
);

OAI21X1 _10182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1679_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1680_),
    .Y(_1628_[26])
);

INVX1 _10183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_1681_)
);

NAND2X1 _10184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1682_)
);

OAI21X1 _10185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1681_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1682_),
    .Y(_1628_[27])
);

INVX1 _10186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_1683_)
);

NAND2X1 _10187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1684_)
);

OAI21X1 _10188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1683_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf6 ),
    .C(_1684_),
    .Y(_1628_[28])
);

INVX1 _10189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_1685_)
);

NAND2X1 _10190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_1686_)
);

OAI21X1 _10191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf4 ),
    .C(_1686_),
    .Y(_1628_[29])
);

INVX1 _10192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_1687_)
);

NAND2X1 _10193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1688_)
);

OAI21X1 _10194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1687_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf2 ),
    .C(_1688_),
    .Y(_1628_[30])
);

INVX1 _10195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_1689_)
);

NAND2X1 _10196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_26_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_1690_)
);

OAI21X1 _10197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1689_),
    .B(\datapath_1.regfile_1.regEn_26_bF$buf0 ),
    .C(_1690_),
    .Y(_1628_[31])
);

DFFSR _10198_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_1628_[0]),
    .Q(\datapath_1.regfile_1.regOut[26] [0]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _10199_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_1628_[1]),
    .Q(\datapath_1.regfile_1.regOut[26] [1]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _10200_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_1628_[2]),
    .Q(\datapath_1.regfile_1.regOut[26] [2]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _10201_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_1628_[3]),
    .Q(\datapath_1.regfile_1.regOut[26] [3]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _10202_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_1628_[4]),
    .Q(\datapath_1.regfile_1.regOut[26] [4]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _10203_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_1628_[5]),
    .Q(\datapath_1.regfile_1.regOut[26] [5]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _10204_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_1628_[6]),
    .Q(\datapath_1.regfile_1.regOut[26] [6]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _10205_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_1628_[7]),
    .Q(\datapath_1.regfile_1.regOut[26] [7]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _10206_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_1628_[8]),
    .Q(\datapath_1.regfile_1.regOut[26] [8]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _10207_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_1628_[9]),
    .Q(\datapath_1.regfile_1.regOut[26] [9]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _10208_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_1628_[10]),
    .Q(\datapath_1.regfile_1.regOut[26] [10]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _10209_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_1628_[11]),
    .Q(\datapath_1.regfile_1.regOut[26] [11]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _10210_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_1628_[12]),
    .Q(\datapath_1.regfile_1.regOut[26] [12]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _10211_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_1628_[13]),
    .Q(\datapath_1.regfile_1.regOut[26] [13]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _10212_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_1628_[14]),
    .Q(\datapath_1.regfile_1.regOut[26] [14]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _10213_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_1628_[15]),
    .Q(\datapath_1.regfile_1.regOut[26] [15]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _10214_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_1628_[16]),
    .Q(\datapath_1.regfile_1.regOut[26] [16]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _10215_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_1628_[17]),
    .Q(\datapath_1.regfile_1.regOut[26] [17]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _10216_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_1628_[18]),
    .Q(\datapath_1.regfile_1.regOut[26] [18]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _10217_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_1628_[19]),
    .Q(\datapath_1.regfile_1.regOut[26] [19]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _10218_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_1628_[20]),
    .Q(\datapath_1.regfile_1.regOut[26] [20]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _10219_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_1628_[21]),
    .Q(\datapath_1.regfile_1.regOut[26] [21]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _10220_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_1628_[22]),
    .Q(\datapath_1.regfile_1.regOut[26] [22]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _10221_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_1628_[23]),
    .Q(\datapath_1.regfile_1.regOut[26] [23]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _10222_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_1628_[24]),
    .Q(\datapath_1.regfile_1.regOut[26] [24]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _10223_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_1628_[25]),
    .Q(\datapath_1.regfile_1.regOut[26] [25]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _10224_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_1628_[26]),
    .Q(\datapath_1.regfile_1.regOut[26] [26]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _10225_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_1628_[27]),
    .Q(\datapath_1.regfile_1.regOut[26] [27]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _10226_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_1628_[28]),
    .Q(\datapath_1.regfile_1.regOut[26] [28]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _10227_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_1628_[29]),
    .Q(\datapath_1.regfile_1.regOut[26] [29]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _10228_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_1628_[30]),
    .Q(\datapath_1.regfile_1.regOut[26] [30]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _10229_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_1628_[31]),
    .Q(\datapath_1.regfile_1.regOut[26] [31]),
    .R(rst_bF$buf50),
    .S(vdd)
);

INVX1 _10230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_1756_)
);

NAND2X1 _10231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .Y(_1757_)
);

OAI21X1 _10232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1756_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1757_),
    .Y(_1693_[0])
);

INVX1 _10233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_1694_)
);

NAND2X1 _10234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1695_)
);

OAI21X1 _10235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1695_),
    .Y(_1693_[1])
);

INVX1 _10236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_1696_)
);

NAND2X1 _10237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1697_)
);

OAI21X1 _10238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1696_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1697_),
    .Y(_1693_[2])
);

INVX1 _10239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_1698_)
);

NAND2X1 _10240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_1699_)
);

OAI21X1 _10241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1698_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1699_),
    .Y(_1693_[3])
);

INVX1 _10242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_1700_)
);

NAND2X1 _10243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1701_)
);

OAI21X1 _10244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1700_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1701_),
    .Y(_1693_[4])
);

INVX1 _10245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_1702_)
);

NAND2X1 _10246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1703_)
);

OAI21X1 _10247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1702_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1703_),
    .Y(_1693_[5])
);

INVX1 _10248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_1704_)
);

NAND2X1 _10249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1705_)
);

OAI21X1 _10250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1704_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1705_),
    .Y(_1693_[6])
);

INVX1 _10251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_1706_)
);

NAND2X1 _10252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1707_)
);

OAI21X1 _10253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1706_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1707_),
    .Y(_1693_[7])
);

INVX1 _10254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_1708_)
);

NAND2X1 _10255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1709_)
);

OAI21X1 _10256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1708_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1709_),
    .Y(_1693_[8])
);

INVX1 _10257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_1710_)
);

NAND2X1 _10258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1711_)
);

OAI21X1 _10259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1710_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1711_),
    .Y(_1693_[9])
);

INVX1 _10260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_1712_)
);

NAND2X1 _10261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1713_)
);

OAI21X1 _10262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1713_),
    .Y(_1693_[10])
);

INVX1 _10263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_1714_)
);

NAND2X1 _10264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1715_)
);

OAI21X1 _10265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1714_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1715_),
    .Y(_1693_[11])
);

INVX1 _10266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [12]),
    .Y(_1716_)
);

NAND2X1 _10267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1717_)
);

OAI21X1 _10268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1716_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1717_),
    .Y(_1693_[12])
);

INVX1 _10269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_1718_)
);

NAND2X1 _10270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1719_)
);

OAI21X1 _10271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1718_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1719_),
    .Y(_1693_[13])
);

INVX1 _10272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_1720_)
);

NAND2X1 _10273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1721_)
);

OAI21X1 _10274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1720_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1721_),
    .Y(_1693_[14])
);

INVX1 _10275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [15]),
    .Y(_1722_)
);

NAND2X1 _10276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1723_)
);

OAI21X1 _10277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1722_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1723_),
    .Y(_1693_[15])
);

INVX1 _10278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_1724_)
);

NAND2X1 _10279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1725_)
);

OAI21X1 _10280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1725_),
    .Y(_1693_[16])
);

INVX1 _10281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_1726_)
);

NAND2X1 _10282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1727_)
);

OAI21X1 _10283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1726_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1727_),
    .Y(_1693_[17])
);

INVX1 _10284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_1728_)
);

NAND2X1 _10285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1729_)
);

OAI21X1 _10286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1728_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1729_),
    .Y(_1693_[18])
);

INVX1 _10287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_1730_)
);

NAND2X1 _10288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1731_)
);

OAI21X1 _10289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1730_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1731_),
    .Y(_1693_[19])
);

INVX1 _10290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [20]),
    .Y(_1732_)
);

NAND2X1 _10291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1733_)
);

OAI21X1 _10292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1732_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1733_),
    .Y(_1693_[20])
);

INVX1 _10293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_1734_)
);

NAND2X1 _10294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1735_)
);

OAI21X1 _10295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1734_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1735_),
    .Y(_1693_[21])
);

INVX1 _10296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_1736_)
);

NAND2X1 _10297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1737_)
);

OAI21X1 _10298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1736_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1737_),
    .Y(_1693_[22])
);

INVX1 _10299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_1738_)
);

NAND2X1 _10300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1739_)
);

OAI21X1 _10301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1739_),
    .Y(_1693_[23])
);

INVX1 _10302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_1740_)
);

NAND2X1 _10303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1741_)
);

OAI21X1 _10304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1740_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1741_),
    .Y(_1693_[24])
);

INVX1 _10305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .Y(_1742_)
);

NAND2X1 _10306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1743_)
);

OAI21X1 _10307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1742_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1743_),
    .Y(_1693_[25])
);

INVX1 _10308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_1744_)
);

NAND2X1 _10309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1745_)
);

OAI21X1 _10310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1744_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1745_),
    .Y(_1693_[26])
);

INVX1 _10311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_1746_)
);

NAND2X1 _10312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1747_)
);

OAI21X1 _10313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1746_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1747_),
    .Y(_1693_[27])
);

INVX1 _10314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [28]),
    .Y(_1748_)
);

NAND2X1 _10315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1749_)
);

OAI21X1 _10316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1748_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf6 ),
    .C(_1749_),
    .Y(_1693_[28])
);

INVX1 _10317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_1750_)
);

NAND2X1 _10318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1751_)
);

OAI21X1 _10319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1750_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf4 ),
    .C(_1751_),
    .Y(_1693_[29])
);

INVX1 _10320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_1752_)
);

NAND2X1 _10321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1753_)
);

OAI21X1 _10322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1752_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf2 ),
    .C(_1753_),
    .Y(_1693_[30])
);

INVX1 _10323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_1754_)
);

NAND2X1 _10324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_27_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1755_)
);

OAI21X1 _10325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1754_),
    .B(\datapath_1.regfile_1.regEn_27_bF$buf0 ),
    .C(_1755_),
    .Y(_1693_[31])
);

DFFSR _10326_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_1693_[0]),
    .Q(\datapath_1.regfile_1.regOut[27] [0]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _10327_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_1693_[1]),
    .Q(\datapath_1.regfile_1.regOut[27] [1]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _10328_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_1693_[2]),
    .Q(\datapath_1.regfile_1.regOut[27] [2]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _10329_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_1693_[3]),
    .Q(\datapath_1.regfile_1.regOut[27] [3]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _10330_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_1693_[4]),
    .Q(\datapath_1.regfile_1.regOut[27] [4]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _10331_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_1693_[5]),
    .Q(\datapath_1.regfile_1.regOut[27] [5]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _10332_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_1693_[6]),
    .Q(\datapath_1.regfile_1.regOut[27] [6]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _10333_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_1693_[7]),
    .Q(\datapath_1.regfile_1.regOut[27] [7]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _10334_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_1693_[8]),
    .Q(\datapath_1.regfile_1.regOut[27] [8]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _10335_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_1693_[9]),
    .Q(\datapath_1.regfile_1.regOut[27] [9]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _10336_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_1693_[10]),
    .Q(\datapath_1.regfile_1.regOut[27] [10]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _10337_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_1693_[11]),
    .Q(\datapath_1.regfile_1.regOut[27] [11]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _10338_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_1693_[12]),
    .Q(\datapath_1.regfile_1.regOut[27] [12]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _10339_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_1693_[13]),
    .Q(\datapath_1.regfile_1.regOut[27] [13]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _10340_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_1693_[14]),
    .Q(\datapath_1.regfile_1.regOut[27] [14]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _10341_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_1693_[15]),
    .Q(\datapath_1.regfile_1.regOut[27] [15]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _10342_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_1693_[16]),
    .Q(\datapath_1.regfile_1.regOut[27] [16]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _10343_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_1693_[17]),
    .Q(\datapath_1.regfile_1.regOut[27] [17]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _10344_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_1693_[18]),
    .Q(\datapath_1.regfile_1.regOut[27] [18]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _10345_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_1693_[19]),
    .Q(\datapath_1.regfile_1.regOut[27] [19]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _10346_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_1693_[20]),
    .Q(\datapath_1.regfile_1.regOut[27] [20]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _10347_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_1693_[21]),
    .Q(\datapath_1.regfile_1.regOut[27] [21]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _10348_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_1693_[22]),
    .Q(\datapath_1.regfile_1.regOut[27] [22]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _10349_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_1693_[23]),
    .Q(\datapath_1.regfile_1.regOut[27] [23]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _10350_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_1693_[24]),
    .Q(\datapath_1.regfile_1.regOut[27] [24]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _10351_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_1693_[25]),
    .Q(\datapath_1.regfile_1.regOut[27] [25]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _10352_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_1693_[26]),
    .Q(\datapath_1.regfile_1.regOut[27] [26]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _10353_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_1693_[27]),
    .Q(\datapath_1.regfile_1.regOut[27] [27]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _10354_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_1693_[28]),
    .Q(\datapath_1.regfile_1.regOut[27] [28]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _10355_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_1693_[29]),
    .Q(\datapath_1.regfile_1.regOut[27] [29]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _10356_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_1693_[30]),
    .Q(\datapath_1.regfile_1.regOut[27] [30]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _10357_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_1693_[31]),
    .Q(\datapath_1.regfile_1.regOut[27] [31]),
    .R(rst_bF$buf18),
    .S(vdd)
);

INVX1 _10358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_1821_)
);

NAND2X1 _10359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .Y(_1822_)
);

OAI21X1 _10360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1821_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1822_),
    .Y(_1758_[0])
);

INVX1 _10361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .Y(_1759_)
);

NAND2X1 _10362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1760_)
);

OAI21X1 _10363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1759_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1760_),
    .Y(_1758_[1])
);

INVX1 _10364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_1761_)
);

NAND2X1 _10365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1762_)
);

OAI21X1 _10366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1762_),
    .Y(_1758_[2])
);

INVX1 _10367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .Y(_1763_)
);

NAND2X1 _10368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1764_)
);

OAI21X1 _10369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1763_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1764_),
    .Y(_1758_[3])
);

INVX1 _10370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_1765_)
);

NAND2X1 _10371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1766_)
);

OAI21X1 _10372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1765_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1766_),
    .Y(_1758_[4])
);

INVX1 _10373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_1767_)
);

NAND2X1 _10374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1768_)
);

OAI21X1 _10375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1767_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1768_),
    .Y(_1758_[5])
);

INVX1 _10376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_1769_)
);

NAND2X1 _10377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1770_)
);

OAI21X1 _10378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1769_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1770_),
    .Y(_1758_[6])
);

INVX1 _10379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .Y(_1771_)
);

NAND2X1 _10380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1772_)
);

OAI21X1 _10381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1771_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1772_),
    .Y(_1758_[7])
);

INVX1 _10382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_1773_)
);

NAND2X1 _10383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1774_)
);

OAI21X1 _10384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1773_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1774_),
    .Y(_1758_[8])
);

INVX1 _10385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_1775_)
);

NAND2X1 _10386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1776_)
);

OAI21X1 _10387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1775_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1776_),
    .Y(_1758_[9])
);

INVX1 _10388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .Y(_1777_)
);

NAND2X1 _10389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1778_)
);

OAI21X1 _10390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1777_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1778_),
    .Y(_1758_[10])
);

INVX1 _10391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_1779_)
);

NAND2X1 _10392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1780_)
);

OAI21X1 _10393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1779_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1780_),
    .Y(_1758_[11])
);

INVX1 _10394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_1781_)
);

NAND2X1 _10395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1782_)
);

OAI21X1 _10396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1781_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1782_),
    .Y(_1758_[12])
);

INVX1 _10397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_1783_)
);

NAND2X1 _10398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1784_)
);

OAI21X1 _10399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1783_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1784_),
    .Y(_1758_[13])
);

INVX1 _10400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_1785_)
);

NAND2X1 _10401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1786_)
);

OAI21X1 _10402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1785_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1786_),
    .Y(_1758_[14])
);

INVX1 _10403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_1787_)
);

NAND2X1 _10404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1788_)
);

OAI21X1 _10405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1787_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1788_),
    .Y(_1758_[15])
);

INVX1 _10406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_1789_)
);

NAND2X1 _10407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1790_)
);

OAI21X1 _10408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1789_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1790_),
    .Y(_1758_[16])
);

INVX1 _10409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_1791_)
);

NAND2X1 _10410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1792_)
);

OAI21X1 _10411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1791_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1792_),
    .Y(_1758_[17])
);

INVX1 _10412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_1793_)
);

NAND2X1 _10413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1794_)
);

OAI21X1 _10414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1793_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1794_),
    .Y(_1758_[18])
);

INVX1 _10415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [19]),
    .Y(_1795_)
);

NAND2X1 _10416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1796_)
);

OAI21X1 _10417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1795_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1796_),
    .Y(_1758_[19])
);

INVX1 _10418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_1797_)
);

NAND2X1 _10419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1798_)
);

OAI21X1 _10420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1797_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1798_),
    .Y(_1758_[20])
);

INVX1 _10421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .Y(_1799_)
);

NAND2X1 _10422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1800_)
);

OAI21X1 _10423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1800_),
    .Y(_1758_[21])
);

INVX1 _10424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_1801_)
);

NAND2X1 _10425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_1802_)
);

OAI21X1 _10426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1801_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1802_),
    .Y(_1758_[22])
);

INVX1 _10427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_1803_)
);

NAND2X1 _10428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1804_)
);

OAI21X1 _10429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1803_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1804_),
    .Y(_1758_[23])
);

INVX1 _10430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_1805_)
);

NAND2X1 _10431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1806_)
);

OAI21X1 _10432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1805_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1806_),
    .Y(_1758_[24])
);

INVX1 _10433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_1807_)
);

NAND2X1 _10434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1808_)
);

OAI21X1 _10435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1807_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1808_),
    .Y(_1758_[25])
);

INVX1 _10436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_1809_)
);

NAND2X1 _10437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1810_)
);

OAI21X1 _10438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1810_),
    .Y(_1758_[26])
);

INVX1 _10439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_1811_)
);

NAND2X1 _10440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1812_)
);

OAI21X1 _10441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1812_),
    .Y(_1758_[27])
);

INVX1 _10442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [28]),
    .Y(_1813_)
);

NAND2X1 _10443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1814_)
);

OAI21X1 _10444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf6 ),
    .C(_1814_),
    .Y(_1758_[28])
);

INVX1 _10445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_1815_)
);

NAND2X1 _10446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1816_)
);

OAI21X1 _10447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf4 ),
    .C(_1816_),
    .Y(_1758_[29])
);

INVX1 _10448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_1817_)
);

NAND2X1 _10449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1818_)
);

OAI21X1 _10450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1817_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf2 ),
    .C(_1818_),
    .Y(_1758_[30])
);

INVX1 _10451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_1819_)
);

NAND2X1 _10452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_28_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1820_)
);

OAI21X1 _10453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1819_),
    .B(\datapath_1.regfile_1.regEn_28_bF$buf0 ),
    .C(_1820_),
    .Y(_1758_[31])
);

DFFSR _10454_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_1758_[0]),
    .Q(\datapath_1.regfile_1.regOut[28] [0]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _10455_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_1758_[1]),
    .Q(\datapath_1.regfile_1.regOut[28] [1]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _10456_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_1758_[2]),
    .Q(\datapath_1.regfile_1.regOut[28] [2]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _10457_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_1758_[3]),
    .Q(\datapath_1.regfile_1.regOut[28] [3]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _10458_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_1758_[4]),
    .Q(\datapath_1.regfile_1.regOut[28] [4]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _10459_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_1758_[5]),
    .Q(\datapath_1.regfile_1.regOut[28] [5]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _10460_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_1758_[6]),
    .Q(\datapath_1.regfile_1.regOut[28] [6]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _10461_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_1758_[7]),
    .Q(\datapath_1.regfile_1.regOut[28] [7]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _10462_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_1758_[8]),
    .Q(\datapath_1.regfile_1.regOut[28] [8]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _10463_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_1758_[9]),
    .Q(\datapath_1.regfile_1.regOut[28] [9]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _10464_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1758_[10]),
    .Q(\datapath_1.regfile_1.regOut[28] [10]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _10465_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1758_[11]),
    .Q(\datapath_1.regfile_1.regOut[28] [11]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _10466_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1758_[12]),
    .Q(\datapath_1.regfile_1.regOut[28] [12]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _10467_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1758_[13]),
    .Q(\datapath_1.regfile_1.regOut[28] [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _10468_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1758_[14]),
    .Q(\datapath_1.regfile_1.regOut[28] [14]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _10469_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1758_[15]),
    .Q(\datapath_1.regfile_1.regOut[28] [15]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _10470_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1758_[16]),
    .Q(\datapath_1.regfile_1.regOut[28] [16]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _10471_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1758_[17]),
    .Q(\datapath_1.regfile_1.regOut[28] [17]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _10472_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_1758_[18]),
    .Q(\datapath_1.regfile_1.regOut[28] [18]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _10473_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_1758_[19]),
    .Q(\datapath_1.regfile_1.regOut[28] [19]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _10474_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_1758_[20]),
    .Q(\datapath_1.regfile_1.regOut[28] [20]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _10475_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_1758_[21]),
    .Q(\datapath_1.regfile_1.regOut[28] [21]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _10476_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_1758_[22]),
    .Q(\datapath_1.regfile_1.regOut[28] [22]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _10477_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_1758_[23]),
    .Q(\datapath_1.regfile_1.regOut[28] [23]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _10478_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_1758_[24]),
    .Q(\datapath_1.regfile_1.regOut[28] [24]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _10479_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_1758_[25]),
    .Q(\datapath_1.regfile_1.regOut[28] [25]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _10480_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_1758_[26]),
    .Q(\datapath_1.regfile_1.regOut[28] [26]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _10481_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_1758_[27]),
    .Q(\datapath_1.regfile_1.regOut[28] [27]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _10482_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_1758_[28]),
    .Q(\datapath_1.regfile_1.regOut[28] [28]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _10483_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_1758_[29]),
    .Q(\datapath_1.regfile_1.regOut[28] [29]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _10484_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_1758_[30]),
    .Q(\datapath_1.regfile_1.regOut[28] [30]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _10485_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_1758_[31]),
    .Q(\datapath_1.regfile_1.regOut[28] [31]),
    .R(rst_bF$buf100),
    .S(vdd)
);

INVX1 _10486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_1886_)
);

NAND2X1 _10487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .Y(_1887_)
);

OAI21X1 _10488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1886_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1887_),
    .Y(_1823_[0])
);

INVX1 _10489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_1824_)
);

NAND2X1 _10490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1825_)
);

OAI21X1 _10491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1825_),
    .Y(_1823_[1])
);

INVX1 _10492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_1826_)
);

NAND2X1 _10493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1827_)
);

OAI21X1 _10494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1827_),
    .Y(_1823_[2])
);

INVX1 _10495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_1828_)
);

NAND2X1 _10496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1829_)
);

OAI21X1 _10497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1828_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1829_),
    .Y(_1823_[3])
);

INVX1 _10498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_1830_)
);

NAND2X1 _10499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1831_)
);

OAI21X1 _10500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1830_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1831_),
    .Y(_1823_[4])
);

INVX1 _10501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_1832_)
);

NAND2X1 _10502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1833_)
);

OAI21X1 _10503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1832_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1833_),
    .Y(_1823_[5])
);

INVX1 _10504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_1834_)
);

NAND2X1 _10505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1835_)
);

OAI21X1 _10506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1835_),
    .Y(_1823_[6])
);

INVX1 _10507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_1836_)
);

NAND2X1 _10508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1837_)
);

OAI21X1 _10509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1836_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1837_),
    .Y(_1823_[7])
);

INVX1 _10510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_1838_)
);

NAND2X1 _10511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1839_)
);

OAI21X1 _10512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1838_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1839_),
    .Y(_1823_[8])
);

INVX1 _10513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_1840_)
);

NAND2X1 _10514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1841_)
);

OAI21X1 _10515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1840_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1841_),
    .Y(_1823_[9])
);

INVX1 _10516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_1842_)
);

NAND2X1 _10517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1843_)
);

OAI21X1 _10518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1842_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1843_),
    .Y(_1823_[10])
);

INVX1 _10519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_1844_)
);

NAND2X1 _10520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1845_)
);

OAI21X1 _10521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1844_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1845_),
    .Y(_1823_[11])
);

INVX1 _10522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_1846_)
);

NAND2X1 _10523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1847_)
);

OAI21X1 _10524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1846_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1847_),
    .Y(_1823_[12])
);

INVX1 _10525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_1848_)
);

NAND2X1 _10526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1849_)
);

OAI21X1 _10527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1849_),
    .Y(_1823_[13])
);

INVX1 _10528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_1850_)
);

NAND2X1 _10529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1851_)
);

OAI21X1 _10530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1850_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1851_),
    .Y(_1823_[14])
);

INVX1 _10531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_1852_)
);

NAND2X1 _10532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1853_)
);

OAI21X1 _10533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1853_),
    .Y(_1823_[15])
);

INVX1 _10534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_1854_)
);

NAND2X1 _10535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1855_)
);

OAI21X1 _10536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1854_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1855_),
    .Y(_1823_[16])
);

INVX1 _10537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_1856_)
);

NAND2X1 _10538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1857_)
);

OAI21X1 _10539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1856_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1857_),
    .Y(_1823_[17])
);

INVX1 _10540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_1858_)
);

NAND2X1 _10541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1859_)
);

OAI21X1 _10542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1858_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1859_),
    .Y(_1823_[18])
);

INVX1 _10543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_1860_)
);

NAND2X1 _10544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1861_)
);

OAI21X1 _10545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1860_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1861_),
    .Y(_1823_[19])
);

INVX1 _10546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_1862_)
);

NAND2X1 _10547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1863_)
);

OAI21X1 _10548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1862_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1863_),
    .Y(_1823_[20])
);

INVX1 _10549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_1864_)
);

NAND2X1 _10550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1865_)
);

OAI21X1 _10551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1864_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1865_),
    .Y(_1823_[21])
);

INVX1 _10552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_1866_)
);

NAND2X1 _10553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1867_)
);

OAI21X1 _10554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1867_),
    .Y(_1823_[22])
);

INVX1 _10555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_1868_)
);

NAND2X1 _10556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1869_)
);

OAI21X1 _10557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1868_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1869_),
    .Y(_1823_[23])
);

INVX1 _10558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_1870_)
);

NAND2X1 _10559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1871_)
);

OAI21X1 _10560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1870_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1871_),
    .Y(_1823_[24])
);

INVX1 _10561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_1872_)
);

NAND2X1 _10562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1873_)
);

OAI21X1 _10563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1873_),
    .Y(_1823_[25])
);

INVX1 _10564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_1874_)
);

NAND2X1 _10565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1875_)
);

OAI21X1 _10566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1874_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1875_),
    .Y(_1823_[26])
);

INVX1 _10567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_1876_)
);

NAND2X1 _10568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1877_)
);

OAI21X1 _10569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1876_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1877_),
    .Y(_1823_[27])
);

INVX1 _10570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_1878_)
);

NAND2X1 _10571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1879_)
);

OAI21X1 _10572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf6 ),
    .C(_1879_),
    .Y(_1823_[28])
);

INVX1 _10573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_1880_)
);

NAND2X1 _10574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1881_)
);

OAI21X1 _10575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1880_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf4 ),
    .C(_1881_),
    .Y(_1823_[29])
);

INVX1 _10576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_1882_)
);

NAND2X1 _10577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1883_)
);

OAI21X1 _10578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1882_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf2 ),
    .C(_1883_),
    .Y(_1823_[30])
);

INVX1 _10579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_1884_)
);

NAND2X1 _10580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_29_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1885_)
);

OAI21X1 _10581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(\datapath_1.regfile_1.regEn_29_bF$buf0 ),
    .C(_1885_),
    .Y(_1823_[31])
);

DFFSR _10582_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_1823_[0]),
    .Q(\datapath_1.regfile_1.regOut[29] [0]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _10583_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_1823_[1]),
    .Q(\datapath_1.regfile_1.regOut[29] [1]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _10584_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_1823_[2]),
    .Q(\datapath_1.regfile_1.regOut[29] [2]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _10585_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_1823_[3]),
    .Q(\datapath_1.regfile_1.regOut[29] [3]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _10586_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_1823_[4]),
    .Q(\datapath_1.regfile_1.regOut[29] [4]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _10587_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_1823_[5]),
    .Q(\datapath_1.regfile_1.regOut[29] [5]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _10588_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_1823_[6]),
    .Q(\datapath_1.regfile_1.regOut[29] [6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _10589_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_1823_[7]),
    .Q(\datapath_1.regfile_1.regOut[29] [7]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _10590_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_1823_[8]),
    .Q(\datapath_1.regfile_1.regOut[29] [8]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _10591_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_1823_[9]),
    .Q(\datapath_1.regfile_1.regOut[29] [9]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _10592_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_1823_[10]),
    .Q(\datapath_1.regfile_1.regOut[29] [10]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _10593_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_1823_[11]),
    .Q(\datapath_1.regfile_1.regOut[29] [11]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _10594_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_1823_[12]),
    .Q(\datapath_1.regfile_1.regOut[29] [12]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _10595_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_1823_[13]),
    .Q(\datapath_1.regfile_1.regOut[29] [13]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _10596_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_1823_[14]),
    .Q(\datapath_1.regfile_1.regOut[29] [14]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _10597_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_1823_[15]),
    .Q(\datapath_1.regfile_1.regOut[29] [15]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _10598_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_1823_[16]),
    .Q(\datapath_1.regfile_1.regOut[29] [16]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _10599_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_1823_[17]),
    .Q(\datapath_1.regfile_1.regOut[29] [17]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _10600_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_1823_[18]),
    .Q(\datapath_1.regfile_1.regOut[29] [18]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _10601_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_1823_[19]),
    .Q(\datapath_1.regfile_1.regOut[29] [19]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _10602_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_1823_[20]),
    .Q(\datapath_1.regfile_1.regOut[29] [20]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _10603_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_1823_[21]),
    .Q(\datapath_1.regfile_1.regOut[29] [21]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _10604_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_1823_[22]),
    .Q(\datapath_1.regfile_1.regOut[29] [22]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _10605_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_1823_[23]),
    .Q(\datapath_1.regfile_1.regOut[29] [23]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _10606_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_1823_[24]),
    .Q(\datapath_1.regfile_1.regOut[29] [24]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _10607_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_1823_[25]),
    .Q(\datapath_1.regfile_1.regOut[29] [25]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _10608_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_1823_[26]),
    .Q(\datapath_1.regfile_1.regOut[29] [26]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _10609_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_1823_[27]),
    .Q(\datapath_1.regfile_1.regOut[29] [27]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _10610_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_1823_[28]),
    .Q(\datapath_1.regfile_1.regOut[29] [28]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _10611_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_1823_[29]),
    .Q(\datapath_1.regfile_1.regOut[29] [29]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _10612_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_1823_[30]),
    .Q(\datapath_1.regfile_1.regOut[29] [30]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _10613_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_1823_[31]),
    .Q(\datapath_1.regfile_1.regOut[29] [31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

INVX1 _10614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .Y(_1951_)
);

NAND2X1 _10615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .Y(_1952_)
);

OAI21X1 _10616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1951_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1952_),
    .Y(_1888_[0])
);

INVX1 _10617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_1889_)
);

NAND2X1 _10618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1890_)
);

OAI21X1 _10619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1889_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1890_),
    .Y(_1888_[1])
);

INVX1 _10620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [2]),
    .Y(_1891_)
);

NAND2X1 _10621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1892_)
);

OAI21X1 _10622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1891_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1892_),
    .Y(_1888_[2])
);

INVX1 _10623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_1893_)
);

NAND2X1 _10624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1894_)
);

OAI21X1 _10625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1894_),
    .Y(_1888_[3])
);

INVX1 _10626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_1895_)
);

NAND2X1 _10627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1896_)
);

OAI21X1 _10628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1895_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1896_),
    .Y(_1888_[4])
);

INVX1 _10629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_1897_)
);

NAND2X1 _10630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1898_)
);

OAI21X1 _10631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1897_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1898_),
    .Y(_1888_[5])
);

INVX1 _10632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_1899_)
);

NAND2X1 _10633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1900_)
);

OAI21X1 _10634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1899_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1900_),
    .Y(_1888_[6])
);

INVX1 _10635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_1901_)
);

NAND2X1 _10636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1902_)
);

OAI21X1 _10637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1902_),
    .Y(_1888_[7])
);

INVX1 _10638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_1903_)
);

NAND2X1 _10639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1904_)
);

OAI21X1 _10640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1903_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1904_),
    .Y(_1888_[8])
);

INVX1 _10641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_1905_)
);

NAND2X1 _10642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1906_)
);

OAI21X1 _10643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1905_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1906_),
    .Y(_1888_[9])
);

INVX1 _10644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_1907_)
);

NAND2X1 _10645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1908_)
);

OAI21X1 _10646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1908_),
    .Y(_1888_[10])
);

INVX1 _10647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_1909_)
);

NAND2X1 _10648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1910_)
);

OAI21X1 _10649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1909_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1910_),
    .Y(_1888_[11])
);

INVX1 _10650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_1911_)
);

NAND2X1 _10651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1912_)
);

OAI21X1 _10652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1911_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1912_),
    .Y(_1888_[12])
);

INVX1 _10653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_1913_)
);

NAND2X1 _10654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1914_)
);

OAI21X1 _10655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1913_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1914_),
    .Y(_1888_[13])
);

INVX1 _10656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_1915_)
);

NAND2X1 _10657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1916_)
);

OAI21X1 _10658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1915_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1916_),
    .Y(_1888_[14])
);

INVX1 _10659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_1917_)
);

NAND2X1 _10660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1918_)
);

OAI21X1 _10661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1918_),
    .Y(_1888_[15])
);

INVX1 _10662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_1919_)
);

NAND2X1 _10663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1920_)
);

OAI21X1 _10664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1920_),
    .Y(_1888_[16])
);

INVX1 _10665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_1921_)
);

NAND2X1 _10666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1922_)
);

OAI21X1 _10667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1921_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1922_),
    .Y(_1888_[17])
);

INVX1 _10668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_1923_)
);

NAND2X1 _10669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1924_)
);

OAI21X1 _10670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1924_),
    .Y(_1888_[18])
);

INVX1 _10671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_1925_)
);

NAND2X1 _10672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1926_)
);

OAI21X1 _10673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1926_),
    .Y(_1888_[19])
);

INVX1 _10674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_1927_)
);

NAND2X1 _10675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1928_)
);

OAI21X1 _10676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1927_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1928_),
    .Y(_1888_[20])
);

INVX1 _10677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [21]),
    .Y(_1929_)
);

NAND2X1 _10678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1930_)
);

OAI21X1 _10679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1929_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1930_),
    .Y(_1888_[21])
);

INVX1 _10680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_1931_)
);

NAND2X1 _10681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1932_)
);

OAI21X1 _10682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1931_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1932_),
    .Y(_1888_[22])
);

INVX1 _10683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_1933_)
);

NAND2X1 _10684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1934_)
);

OAI21X1 _10685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1933_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1934_),
    .Y(_1888_[23])
);

INVX1 _10686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_1935_)
);

NAND2X1 _10687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1936_)
);

OAI21X1 _10688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1935_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1936_),
    .Y(_1888_[24])
);

INVX1 _10689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [25]),
    .Y(_1937_)
);

NAND2X1 _10690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1938_)
);

OAI21X1 _10691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1937_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1938_),
    .Y(_1888_[25])
);

INVX1 _10692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_1939_)
);

NAND2X1 _10693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1940_)
);

OAI21X1 _10694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1940_),
    .Y(_1888_[26])
);

INVX1 _10695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_1941_)
);

NAND2X1 _10696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1942_)
);

OAI21X1 _10697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1941_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1942_),
    .Y(_1888_[27])
);

INVX1 _10698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_1943_)
);

NAND2X1 _10699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1944_)
);

OAI21X1 _10700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1943_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf6 ),
    .C(_1944_),
    .Y(_1888_[28])
);

INVX1 _10701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_1945_)
);

NAND2X1 _10702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1946_)
);

OAI21X1 _10703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1945_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf4 ),
    .C(_1946_),
    .Y(_1888_[29])
);

INVX1 _10704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_1947_)
);

NAND2X1 _10705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1948_)
);

OAI21X1 _10706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1947_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf2 ),
    .C(_1948_),
    .Y(_1888_[30])
);

INVX1 _10707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_1949_)
);

NAND2X1 _10708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_30_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1950_)
);

OAI21X1 _10709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1949_),
    .B(\datapath_1.regfile_1.regEn_30_bF$buf0 ),
    .C(_1950_),
    .Y(_1888_[31])
);

DFFSR _10710_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_1888_[0]),
    .Q(\datapath_1.regfile_1.regOut[30] [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _10711_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_1888_[1]),
    .Q(\datapath_1.regfile_1.regOut[30] [1]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _10712_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_1888_[2]),
    .Q(\datapath_1.regfile_1.regOut[30] [2]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _10713_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_1888_[3]),
    .Q(\datapath_1.regfile_1.regOut[30] [3]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _10714_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_1888_[4]),
    .Q(\datapath_1.regfile_1.regOut[30] [4]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _10715_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_1888_[5]),
    .Q(\datapath_1.regfile_1.regOut[30] [5]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _10716_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_1888_[6]),
    .Q(\datapath_1.regfile_1.regOut[30] [6]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _10717_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_1888_[7]),
    .Q(\datapath_1.regfile_1.regOut[30] [7]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _10718_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_1888_[8]),
    .Q(\datapath_1.regfile_1.regOut[30] [8]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _10719_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_1888_[9]),
    .Q(\datapath_1.regfile_1.regOut[30] [9]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _10720_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_1888_[10]),
    .Q(\datapath_1.regfile_1.regOut[30] [10]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _10721_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_1888_[11]),
    .Q(\datapath_1.regfile_1.regOut[30] [11]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _10722_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_1888_[12]),
    .Q(\datapath_1.regfile_1.regOut[30] [12]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _10723_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_1888_[13]),
    .Q(\datapath_1.regfile_1.regOut[30] [13]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _10724_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_1888_[14]),
    .Q(\datapath_1.regfile_1.regOut[30] [14]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _10725_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_1888_[15]),
    .Q(\datapath_1.regfile_1.regOut[30] [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _10726_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_1888_[16]),
    .Q(\datapath_1.regfile_1.regOut[30] [16]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _10727_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_1888_[17]),
    .Q(\datapath_1.regfile_1.regOut[30] [17]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _10728_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_1888_[18]),
    .Q(\datapath_1.regfile_1.regOut[30] [18]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _10729_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_1888_[19]),
    .Q(\datapath_1.regfile_1.regOut[30] [19]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _10730_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_1888_[20]),
    .Q(\datapath_1.regfile_1.regOut[30] [20]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _10731_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_1888_[21]),
    .Q(\datapath_1.regfile_1.regOut[30] [21]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _10732_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_1888_[22]),
    .Q(\datapath_1.regfile_1.regOut[30] [22]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _10733_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_1888_[23]),
    .Q(\datapath_1.regfile_1.regOut[30] [23]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _10734_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_1888_[24]),
    .Q(\datapath_1.regfile_1.regOut[30] [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _10735_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_1888_[25]),
    .Q(\datapath_1.regfile_1.regOut[30] [25]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _10736_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_1888_[26]),
    .Q(\datapath_1.regfile_1.regOut[30] [26]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _10737_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_1888_[27]),
    .Q(\datapath_1.regfile_1.regOut[30] [27]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _10738_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_1888_[28]),
    .Q(\datapath_1.regfile_1.regOut[30] [28]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _10739_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_1888_[29]),
    .Q(\datapath_1.regfile_1.regOut[30] [29]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _10740_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_1888_[30]),
    .Q(\datapath_1.regfile_1.regOut[30] [30]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _10741_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_1888_[31]),
    .Q(\datapath_1.regfile_1.regOut[30] [31]),
    .R(rst_bF$buf36),
    .S(vdd)
);

INVX1 _10742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_2016_)
);

NAND2X1 _10743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .Y(_2017_)
);

OAI21X1 _10744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_2017_),
    .Y(_1953_[0])
);

INVX1 _10745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .Y(_1954_)
);

NAND2X1 _10746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1955_)
);

OAI21X1 _10747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1955_),
    .Y(_1953_[1])
);

INVX1 _10748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_1956_)
);

NAND2X1 _10749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1957_)
);

OAI21X1 _10750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1956_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1957_),
    .Y(_1953_[2])
);

INVX1 _10751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_1958_)
);

NAND2X1 _10752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1959_)
);

OAI21X1 _10753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1958_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1959_),
    .Y(_1953_[3])
);

INVX1 _10754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_1960_)
);

NAND2X1 _10755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1961_)
);

OAI21X1 _10756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1960_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1961_),
    .Y(_1953_[4])
);

INVX1 _10757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_1962_)
);

NAND2X1 _10758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1963_)
);

OAI21X1 _10759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1962_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1963_),
    .Y(_1953_[5])
);

INVX1 _10760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [6]),
    .Y(_1964_)
);

NAND2X1 _10761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1965_)
);

OAI21X1 _10762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1964_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1965_),
    .Y(_1953_[6])
);

INVX1 _10763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [7]),
    .Y(_1966_)
);

NAND2X1 _10764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1967_)
);

OAI21X1 _10765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1966_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1967_),
    .Y(_1953_[7])
);

INVX1 _10766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_1968_)
);

NAND2X1 _10767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1969_)
);

OAI21X1 _10768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1968_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1969_),
    .Y(_1953_[8])
);

INVX1 _10769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_1970_)
);

NAND2X1 _10770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1971_)
);

OAI21X1 _10771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1970_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1971_),
    .Y(_1953_[9])
);

INVX1 _10772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_1972_)
);

NAND2X1 _10773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1973_)
);

OAI21X1 _10774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1972_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1973_),
    .Y(_1953_[10])
);

INVX1 _10775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [11]),
    .Y(_1974_)
);

NAND2X1 _10776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1975_)
);

OAI21X1 _10777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1974_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1975_),
    .Y(_1953_[11])
);

INVX1 _10778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_1976_)
);

NAND2X1 _10779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1977_)
);

OAI21X1 _10780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1976_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1977_),
    .Y(_1953_[12])
);

INVX1 _10781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_1978_)
);

NAND2X1 _10782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1979_)
);

OAI21X1 _10783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1978_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1979_),
    .Y(_1953_[13])
);

INVX1 _10784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_1980_)
);

NAND2X1 _10785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1981_)
);

OAI21X1 _10786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1980_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1981_),
    .Y(_1953_[14])
);

INVX1 _10787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_1982_)
);

NAND2X1 _10788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1983_)
);

OAI21X1 _10789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1982_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1983_),
    .Y(_1953_[15])
);

INVX1 _10790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_1984_)
);

NAND2X1 _10791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1985_)
);

OAI21X1 _10792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1984_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1985_),
    .Y(_1953_[16])
);

INVX1 _10793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_1986_)
);

NAND2X1 _10794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1987_)
);

OAI21X1 _10795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1986_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1987_),
    .Y(_1953_[17])
);

INVX1 _10796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_1988_)
);

NAND2X1 _10797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1989_)
);

OAI21X1 _10798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1989_),
    .Y(_1953_[18])
);

INVX1 _10799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [19]),
    .Y(_1990_)
);

NAND2X1 _10800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1991_)
);

OAI21X1 _10801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1991_),
    .Y(_1953_[19])
);

INVX1 _10802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_1992_)
);

NAND2X1 _10803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1993_)
);

OAI21X1 _10804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1992_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_1993_),
    .Y(_1953_[20])
);

INVX1 _10805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_1994_)
);

NAND2X1 _10806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1995_)
);

OAI21X1 _10807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1994_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_1995_),
    .Y(_1953_[21])
);

INVX1 _10808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .Y(_1996_)
);

NAND2X1 _10809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1997_)
);

OAI21X1 _10810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_1997_),
    .Y(_1953_[22])
);

INVX1 _10811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_1998_)
);

NAND2X1 _10812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1999_)
);

OAI21X1 _10813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1998_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_1999_),
    .Y(_1953_[23])
);

INVX1 _10814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_2000_)
);

NAND2X1 _10815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_2001_)
);

OAI21X1 _10816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2000_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_2001_),
    .Y(_1953_[24])
);

INVX1 _10817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_2002_)
);

NAND2X1 _10818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_2003_)
);

OAI21X1 _10819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2002_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_2003_),
    .Y(_1953_[25])
);

INVX1 _10820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_2004_)
);

NAND2X1 _10821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_2005_)
);

OAI21X1 _10822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_2005_),
    .Y(_1953_[26])
);

INVX1 _10823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_2006_)
);

NAND2X1 _10824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_2007_)
);

OAI21X1 _10825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2006_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_2007_),
    .Y(_1953_[27])
);

INVX1 _10826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [28]),
    .Y(_2008_)
);

NAND2X1 _10827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_2009_)
);

OAI21X1 _10828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf6 ),
    .C(_2009_),
    .Y(_1953_[28])
);

INVX1 _10829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_2010_)
);

NAND2X1 _10830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_2011_)
);

OAI21X1 _10831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2010_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf4 ),
    .C(_2011_),
    .Y(_1953_[29])
);

INVX1 _10832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_2012_)
);

NAND2X1 _10833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_2013_)
);

OAI21X1 _10834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2012_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf2 ),
    .C(_2013_),
    .Y(_1953_[30])
);

INVX1 _10835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [31]),
    .Y(_2014_)
);

NAND2X1 _10836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_31_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_2015_)
);

OAI21X1 _10837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2014_),
    .B(\datapath_1.regfile_1.regEn_31_bF$buf0 ),
    .C(_2015_),
    .Y(_1953_[31])
);

DFFSR _10838_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_1953_[0]),
    .Q(\datapath_1.regfile_1.regOut[31] [0]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _10839_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_1953_[1]),
    .Q(\datapath_1.regfile_1.regOut[31] [1]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _10840_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_1953_[2]),
    .Q(\datapath_1.regfile_1.regOut[31] [2]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _10841_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_1953_[3]),
    .Q(\datapath_1.regfile_1.regOut[31] [3]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _10842_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_1953_[4]),
    .Q(\datapath_1.regfile_1.regOut[31] [4]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _10843_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_1953_[5]),
    .Q(\datapath_1.regfile_1.regOut[31] [5]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _10844_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_1953_[6]),
    .Q(\datapath_1.regfile_1.regOut[31] [6]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _10845_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_1953_[7]),
    .Q(\datapath_1.regfile_1.regOut[31] [7]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _10846_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_1953_[8]),
    .Q(\datapath_1.regfile_1.regOut[31] [8]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _10847_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_1953_[9]),
    .Q(\datapath_1.regfile_1.regOut[31] [9]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _10848_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_1953_[10]),
    .Q(\datapath_1.regfile_1.regOut[31] [10]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _10849_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_1953_[11]),
    .Q(\datapath_1.regfile_1.regOut[31] [11]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _10850_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_1953_[12]),
    .Q(\datapath_1.regfile_1.regOut[31] [12]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _10851_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_1953_[13]),
    .Q(\datapath_1.regfile_1.regOut[31] [13]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _10852_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_1953_[14]),
    .Q(\datapath_1.regfile_1.regOut[31] [14]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _10853_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_1953_[15]),
    .Q(\datapath_1.regfile_1.regOut[31] [15]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _10854_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_1953_[16]),
    .Q(\datapath_1.regfile_1.regOut[31] [16]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _10855_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_1953_[17]),
    .Q(\datapath_1.regfile_1.regOut[31] [17]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _10856_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_1953_[18]),
    .Q(\datapath_1.regfile_1.regOut[31] [18]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _10857_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_1953_[19]),
    .Q(\datapath_1.regfile_1.regOut[31] [19]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _10858_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_1953_[20]),
    .Q(\datapath_1.regfile_1.regOut[31] [20]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _10859_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_1953_[21]),
    .Q(\datapath_1.regfile_1.regOut[31] [21]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _10860_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_1953_[22]),
    .Q(\datapath_1.regfile_1.regOut[31] [22]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _10861_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_1953_[23]),
    .Q(\datapath_1.regfile_1.regOut[31] [23]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _10862_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_1953_[24]),
    .Q(\datapath_1.regfile_1.regOut[31] [24]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _10863_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_1953_[25]),
    .Q(\datapath_1.regfile_1.regOut[31] [25]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _10864_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_1953_[26]),
    .Q(\datapath_1.regfile_1.regOut[31] [26]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _10865_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_1953_[27]),
    .Q(\datapath_1.regfile_1.regOut[31] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _10866_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1953_[28]),
    .Q(\datapath_1.regfile_1.regOut[31] [28]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _10867_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1953_[29]),
    .Q(\datapath_1.regfile_1.regOut[31] [29]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _10868_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1953_[30]),
    .Q(\datapath_1.regfile_1.regOut[31] [30]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _10869_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1953_[31]),
    .Q(\datapath_1.regfile_1.regOut[31] [31]),
    .R(rst_bF$buf4),
    .S(vdd)
);

INVX1 _10870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [4]),
    .Y(_2018_)
);

NAND2X1 _10871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [5]),
    .B(_2018_),
    .Y(_2019_)
);

INVX1 _10872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [3]),
    .Y(_2020_)
);

NAND2X1 _10873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [2]),
    .B(_2020_),
    .Y(_2021_)
);

NOR2X1 _10874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2019_),
    .B(_2021_),
    .Y(_2022_)
);

INVX1 _10875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2022_),
    .Y(_2023_)
);

NAND2X1 _10876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2024_)
);

INVX1 _10877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf5),
    .Y(_2025_)
);

NAND2X1 _10878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[1]),
    .B(_2025_),
    .Y(_2026_)
);

NOR2X1 _10879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [0]),
    .B(\aluControl_1.inst [1]),
    .Y(_2027_)
);

NOR2X1 _10880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2027_),
    .B(_2026_),
    .Y(_2028_)
);

NAND2X1 _10881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2024_),
    .B(_2028_),
    .Y(_2029_)
);

NOR2X1 _10882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2023_),
    .B(_2029_),
    .Y(ALUControl[0])
);

INVX1 _10883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [1]),
    .Y(_2030_)
);

NOR2X1 _10884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [0]),
    .B(_2030_),
    .Y(_2031_)
);

OR2X2 _10885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [3]),
    .B(\aluControl_1.inst [2]),
    .Y(_2032_)
);

NOR2X1 _10886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2032_),
    .B(_2019_),
    .Y(_2033_)
);

OAI21X1 _10887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2022_),
    .B(_2033_),
    .C(_2031_),
    .Y(_2034_)
);

AOI21X1 _10888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2027_),
    .B(_2033_),
    .C(_2026_),
    .Y(_2035_)
);

NAND2X1 _10889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2035_),
    .B(_2034_),
    .Y(ALUControl[1])
);

INVX1 _10890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[1]),
    .Y(_2036_)
);

INVX1 _10891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2019_),
    .Y(_2037_)
);

NOR3X1 _10892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [0]),
    .B(_2030_),
    .C(_2032_),
    .Y(_2038_)
);

INVX1 _10893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [2]),
    .Y(_2039_)
);

NOR3X1 _10894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [3]),
    .B(_2039_),
    .C(_2024_),
    .Y(_2040_)
);

OAI21X1 _10895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2038_),
    .B(_2040_),
    .C(_2037_),
    .Y(_2041_)
);

OAI21X1 _10896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2041_),
    .B(_2036_),
    .C(_2025_),
    .Y(ALUControl[2])
);

INVX2 _10897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [2]),
    .Y(_2046_)
);

NAND2X1 _10898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [3]),
    .B(_2046_),
    .Y(_2047_)
);

INVX1 _10899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .Y(_2048_)
);

NAND2X1 _10900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [0]),
    .B(_2048_),
    .Y(_2049_)
);

NOR2X1 _10901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_2049_),
    .Y(BranchNe)
);

INVX1 _10902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [0]),
    .Y(_2050_)
);

NAND2X1 _10903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2048_),
    .B(_2050_),
    .Y(_2051_)
);

NOR2X1 _10904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_2051_),
    .Y(Branch)
);

INVX2 _10905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [3]),
    .Y(_2052_)
);

NAND2X1 _10906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [2]),
    .B(_2052_),
    .Y(_2053_)
);

NAND2X1 _10907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .B(_2050_),
    .Y(_2054_)
);

NOR2X1 _10908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .B(_2054_),
    .Y(ALUOp[1])
);

INVX2 _10909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2054_),
    .Y(_2055_)
);

OAI21X1 _10910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_2052_),
    .C(_2055_),
    .Y(_2056_)
);

OAI21X1 _10911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .B(_2047_),
    .C(_2056_),
    .Y(ALUSrcA)
);

NAND2X1 _10912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_2052_),
    .Y(_2057_)
);

NOR2X1 _10913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2051_),
    .B(_2057_),
    .Y(IRWrite)
);

NAND2X1 _10914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [2]),
    .B(\control_1.reg_state.dout [3]),
    .Y(_2058_)
);

NOR2X1 _10915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2058_),
    .B(_2051_),
    .Y(PCSource[1])
);

NAND2X1 _10916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_2053_),
    .Y(_2059_)
);

NOR2X1 _10917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2051_),
    .B(_2059_),
    .Y(PCWrite)
);

NAND2X1 _10918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .B(\control_1.reg_state.dout [0]),
    .Y(_2060_)
);

NOR2X1 _10919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2060_),
    .B(_2053_),
    .Y(RegDst)
);

NOR2X1 _10920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .B(_2051_),
    .Y(MemToReg)
);

OAI21X1 _10921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2051_),
    .B(_2053_),
    .C(_2060_),
    .Y(_2061_)
);

AND2X2 _10922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2061_),
    .B(_2059_),
    .Y(RegWrite)
);

NOR2X1 _10923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .B(_2053_),
    .Y(_0_)
);

NOR2X1 _10924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2060_),
    .B(_2057_),
    .Y(_2062_)
);

OR2X2 _10925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2062_),
    .B(_0_),
    .Y(IorD)
);

NOR2X1 _10926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .B(_2047_),
    .Y(ALUOp[0])
);

NOR2X1 _10927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .B(_2057_),
    .Y(ALUSrcB[0])
);

OAI22X1 _10928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2054_),
    .B(\control_1.reg_state.dout [2]),
    .C(_2057_),
    .D(_2049_),
    .Y(ALUSrcB[1])
);

NOR2X1 _10929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .B(_2057_),
    .Y(_2063_)
);

NOR2X1 _10930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [4]),
    .B(\control_1.op [5]),
    .Y(_2064_)
);

INVX1 _10931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .Y(_2065_)
);

INVX1 _10932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [1]),
    .Y(_2066_)
);

INVX1 _10933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [3]),
    .Y(_2067_)
);

NAND3X1 _10934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [2]),
    .B(_2066_),
    .C(_2067_),
    .Y(_2068_)
);

NOR2X1 _10935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2068_),
    .Y(_2069_)
);

NAND3X1 _10936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [0]),
    .B(_2063_),
    .C(_2069_),
    .Y(_2070_)
);

INVX2 _10937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [2]),
    .Y(_2071_)
);

NOR2X1 _10938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2054_),
    .B(_2057_),
    .Y(_2072_)
);

INVX1 _10939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [4]),
    .Y(_2073_)
);

NAND2X1 _10940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [5]),
    .B(_2073_),
    .Y(_2074_)
);

NAND2X1 _10941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [0]),
    .B(\control_1.op [1]),
    .Y(_2075_)
);

NOR2X1 _10942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2074_),
    .Y(_2076_)
);

NAND3X1 _10943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2071_),
    .B(_2076_),
    .C(_2072_),
    .Y(_2077_)
);

AOI21X1 _10944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2055_),
    .B(_2059_),
    .C(IRWrite_bF$buf7),
    .Y(_2078_)
);

NAND3X1 _10945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2078_),
    .B(_2077_),
    .C(_2070_),
    .Y(\control_1.next [0])
);

NAND2X1 _10946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2055_),
    .B(_2059_),
    .Y(_2079_)
);

NOR2X1 _10947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [0]),
    .B(\control_1.op [1]),
    .Y(_2080_)
);

NAND2X1 _10948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2080_),
    .Y(_2081_)
);

OAI21X1 _10949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2074_),
    .B(_2075_),
    .C(_2081_),
    .Y(_2082_)
);

NAND3X1 _10950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2071_),
    .B(_2063_),
    .C(_2082_),
    .Y(_2083_)
);

INVX1 _10951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2074_),
    .Y(_2084_)
);

NOR2X1 _10952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [2]),
    .B(\control_1.op [3]),
    .Y(_2085_)
);

INVX1 _10953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .Y(_2086_)
);

NOR2X1 _10954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2086_),
    .Y(_2087_)
);

NAND3X1 _10955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2084_),
    .B(_2072_),
    .C(_2087_),
    .Y(_2088_)
);

NAND3X1 _10956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2079_),
    .B(_2088_),
    .C(_2083_),
    .Y(\control_1.next [1])
);

NAND2X1 _10957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [3]),
    .B(_2071_),
    .Y(_2089_)
);

NOR2X1 _10958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2089_),
    .Y(_2090_)
);

NAND3X1 _10959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2084_),
    .B(_2090_),
    .C(_2072_),
    .Y(_2091_)
);

NAND2X1 _10960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2085_),
    .Y(_2092_)
);

NOR2X1 _10961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [0]),
    .B(_2092_),
    .Y(_2093_)
);

NAND2X1 _10962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2063_),
    .B(_2093_),
    .Y(_2094_)
);

NOR2X1 _10963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp[1]),
    .B(_2062_),
    .Y(_2095_)
);

NAND3X1 _10964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2095_),
    .C(_2094_),
    .Y(\control_1.next [2])
);

OR2X2 _10965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_2054_),
    .Y(_2096_)
);

NOR2X1 _10966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2081_),
    .Y(_2097_)
);

INVX1 _10967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [0]),
    .Y(_2042_)
);

NAND2X1 _10968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [1]),
    .B(_2042_),
    .Y(_2043_)
);

OAI22X1 _10969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2068_),
    .C(_2092_),
    .D(_2043_),
    .Y(_2044_)
);

OAI21X1 _10970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2044_),
    .B(_2097_),
    .C(_2063_),
    .Y(_2045_)
);

NAND2X1 _10971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2096_),
    .B(_2045_),
    .Y(\control_1.next [3])
);

INVX1 _10972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [0]),
    .Y(_2099_)
);

NAND2X1 _10973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.next [0]),
    .B(vdd),
    .Y(_2100_)
);

OAI21X1 _10974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(vdd),
    .C(_2100_),
    .Y(_2098_[0])
);

INVX1 _10975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [1]),
    .Y(_2101_)
);

NAND2X1 _10976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\control_1.next [1]),
    .Y(_2102_)
);

OAI21X1 _10977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2101_),
    .B(vdd),
    .C(_2102_),
    .Y(_2098_[1])
);

INVX1 _10978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [2]),
    .Y(_2103_)
);

NAND2X1 _10979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\control_1.next [2]),
    .Y(_2104_)
);

OAI21X1 _10980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2103_),
    .B(vdd),
    .C(_2104_),
    .Y(_2098_[2])
);

INVX1 _10981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.reg_state.dout [3]),
    .Y(_2105_)
);

NAND2X1 _10982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\control_1.next [3]),
    .Y(_2106_)
);

OAI21X1 _10983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2105_),
    .B(vdd),
    .C(_2106_),
    .Y(_2098_[3])
);

DFFSR _10984_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_2098_[0]),
    .Q(\control_1.reg_state.dout [0]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _10985_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_2098_[1]),
    .Q(\control_1.reg_state.dout [1]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _10986_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_2098_[2]),
    .Q(\control_1.reg_state.dout [2]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _10987_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_2098_[3]),
    .Q(\control_1.reg_state.dout [3]),
    .R(rst_bF$buf0),
    .S(vdd)
);

NOR2X1 _10988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2107_)
);

NAND2X1 _10989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [31]),
    .B(\datapath_1.alu_1.ALUInB [31]),
    .Y(_2108_)
);

INVX1 _10990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2108_),
    .Y(_2109_)
);

NOR2X1 _10991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2109_),
    .Y(_2110_)
);

INVX2 _10992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .Y(_2111_)
);

INVX1 _10993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [30]),
    .Y(_2112_)
);

INVX1 _10994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2113_)
);

NOR2X1 _10995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2112_),
    .B(_2113_),
    .Y(_2114_)
);

NOR2X1 _10996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [30]),
    .B(\datapath_1.alu_1.ALUInB [30]),
    .Y(_2115_)
);

NOR2X1 _10997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2114_),
    .Y(_2116_)
);

INVX2 _10998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .Y(_2117_)
);

INVX1 _10999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2118_)
);

NOR2X1 _11000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2118_),
    .Y(_2119_)
);

INVX1 _11001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2120_)
);

NOR2X1 _11002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(_2120_),
    .Y(_2121_)
);

NAND2X1 _11003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2122_)
);

OR2X2 _11004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2123_)
);

NAND2X1 _11005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .B(_2123_),
    .Y(_2124_)
);

AOI21X1 _11006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2121_),
    .B(_2124_),
    .C(_2119_),
    .Y(_2125_)
);

INVX1 _11007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2126_)
);

NOR2X1 _11008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(_2126_),
    .Y(_2127_)
);

INVX1 _11009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2128_)
);

NAND2X1 _11010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2129_)
);

OR2X2 _11011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2130_)
);

AOI22X1 _11012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(_2128_),
    .C(_2130_),
    .D(_2129_),
    .Y(_2131_)
);

NAND2X1 _11013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2132_)
);

OR2X2 _11014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2133_)
);

AOI22X1 _11015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2133_),
    .B(_2132_),
    .C(_2122_),
    .D(_2123_),
    .Y(_2134_)
);

OAI21X1 _11016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2131_),
    .B(_2127_),
    .C(_2134_),
    .Y(_2135_)
);

AND2X2 _11017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2136_)
);

NOR2X1 _11018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2137_)
);

AND2X2 _11019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2138_)
);

NOR2X1 _11020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2139_)
);

OAI22X1 _11021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2137_),
    .C(_2138_),
    .D(_2139_),
    .Y(_2140_)
);

AND2X2 _11022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2141_)
);

NOR2X1 _11023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2142_)
);

AND2X2 _11024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2143_)
);

NOR2X1 _11025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2144_)
);

OAI22X1 _11026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2142_),
    .C(_2143_),
    .D(_2144_),
    .Y(_2145_)
);

OR2X2 _11027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2140_),
    .B(_2145_),
    .Y(_2146_)
);

AOI21X1 _11028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .B(_2135_),
    .C(_2146_),
    .Y(_2147_)
);

XNOR2X1 _11029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2148_)
);

INVX1 _11030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2149_)
);

NOR2X1 _11031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(_2149_),
    .Y(_2150_)
);

INVX1 _11032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2151_)
);

NOR2X1 _11033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(_2151_),
    .Y(_2152_)
);

AOI21X1 _11034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2152_),
    .B(_2148_),
    .C(_2150_),
    .Y(_2153_)
);

XNOR2X1 _11035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2154_)
);

INVX1 _11036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2155_)
);

NOR2X1 _11037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(_2155_),
    .Y(_2156_)
);

INVX1 _11038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2157_)
);

NOR2X1 _11039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2157_),
    .Y(_2158_)
);

AOI21X1 _11040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .B(_2154_),
    .C(_2158_),
    .Y(_2159_)
);

OAI21X1 _11041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2153_),
    .B(_2140_),
    .C(_2159_),
    .Y(_2160_)
);

XOR2X1 _11042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2161_)
);

XOR2X1 _11043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2162_)
);

NOR2X1 _11044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2162_),
    .Y(_2163_)
);

XOR2X1 _11045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2164_)
);

XOR2X1 _11046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2165_)
);

NOR2X1 _11047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .B(_2165_),
    .Y(_2166_)
);

NAND2X1 _11048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .B(_2166_),
    .Y(_2167_)
);

XOR2X1 _11049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2168_)
);

XOR2X1 _11050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2169_)
);

NOR2X1 _11051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2169_),
    .Y(_2170_)
);

XOR2X1 _11052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2171_)
);

XOR2X1 _11053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2172_)
);

NOR2X1 _11054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2172_),
    .Y(_2173_)
);

NAND2X1 _11055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2170_),
    .B(_2173_),
    .Y(_2174_)
);

NOR2X1 _11056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2167_),
    .B(_2174_),
    .Y(_2175_)
);

OAI21X1 _11057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2147_),
    .B(_2160_),
    .C(_2175_),
    .Y(_2176_)
);

XNOR2X1 _11058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2177_)
);

AND2X2 _11059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2178_)
);

NOR2X1 _11060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2179_)
);

OAI21X1 _11061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .B(_2179_),
    .C(_2177_),
    .Y(_2180_)
);

XNOR2X1 _11062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2181_)
);

INVX1 _11063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [12]),
    .Y(_2182_)
);

INVX2 _11064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2183_)
);

NOR2X1 _11065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2183_),
    .Y(_2184_)
);

NOR2X1 _11066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(\datapath_1.alu_1.ALUInA [12]),
    .Y(_2185_)
);

OAI21X1 _11067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2184_),
    .B(_2185_),
    .C(_2181_),
    .Y(_2186_)
);

NOR2X1 _11068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2180_),
    .B(_2186_),
    .Y(_2187_)
);

XNOR2X1 _11069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2188_)
);

INVX1 _11070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [10]),
    .Y(_2189_)
);

INVX2 _11071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2190_)
);

NOR2X1 _11072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2189_),
    .B(_2190_),
    .Y(_2191_)
);

NOR2X1 _11073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(\datapath_1.alu_1.ALUInA [10]),
    .Y(_2192_)
);

OAI21X1 _11074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2191_),
    .B(_2192_),
    .C(_2188_),
    .Y(_2193_)
);

XNOR2X1 _11075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2194_)
);

INVX1 _11076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2195_)
);

NOR2X1 _11077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(_2195_),
    .Y(_2196_)
);

INVX2 _11078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [8]),
    .Y(_2197_)
);

NAND2X1 _11079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [8]),
    .B(_2197_),
    .Y(_2198_)
);

INVX1 _11080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .Y(_2199_)
);

AOI21X1 _11081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2194_),
    .B(_2199_),
    .C(_2196_),
    .Y(_2200_)
);

NOR2X1 _11082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2190_),
    .Y(_2201_)
);

INVX2 _11083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [11]),
    .Y(_2202_)
);

NOR2X1 _11084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(_2202_),
    .Y(_2203_)
);

AOI21X1 _11085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2201_),
    .B(_2188_),
    .C(_2203_),
    .Y(_2204_)
);

OAI21X1 _11086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2200_),
    .B(_2193_),
    .C(_2204_),
    .Y(_2205_)
);

INVX2 _11087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2206_)
);

NOR2X1 _11088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(_2206_),
    .Y(_2207_)
);

NOR2X1 _11089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(_2183_),
    .Y(_2208_)
);

AOI21X1 _11090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2208_),
    .B(_2181_),
    .C(_2207_),
    .Y(_2209_)
);

INVX1 _11091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [14]),
    .Y(_2210_)
);

NOR2X1 _11092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [14]),
    .B(_2210_),
    .Y(_2211_)
);

INVX1 _11093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2212_)
);

NOR2X1 _11094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(_2212_),
    .Y(_2213_)
);

AOI21X1 _11095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .B(_2177_),
    .C(_2213_),
    .Y(_2214_)
);

OAI21X1 _11096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2209_),
    .B(_2180_),
    .C(_2214_),
    .Y(_2215_)
);

AOI21X1 _11097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2187_),
    .B(_2205_),
    .C(_2215_),
    .Y(_2216_)
);

NOR2X1 _11098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2217_)
);

NAND2X1 _11099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [22]),
    .B(\datapath_1.alu_1.ALUInB [22]),
    .Y(_2218_)
);

INVX2 _11100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2218_),
    .Y(_2219_)
);

NOR2X1 _11101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .B(_2219_),
    .Y(_2220_)
);

INVX1 _11102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [23]),
    .Y(_2221_)
);

INVX1 _11103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2222_)
);

NOR2X1 _11104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(_2222_),
    .Y(_2223_)
);

NOR2X1 _11105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [23]),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .Y(_2224_)
);

NOR2X1 _11106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .B(_2223_),
    .Y(_2225_)
);

NOR2X1 _11107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2220_),
    .B(_2225_),
    .Y(_2226_)
);

INVX1 _11108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [21]),
    .Y(_2227_)
);

INVX1 _11109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2228_)
);

NOR2X1 _11110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(_2228_),
    .Y(_2229_)
);

NOR2X1 _11111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [21]),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .Y(_2230_)
);

NOR2X1 _11112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2230_),
    .B(_2229_),
    .Y(_2231_)
);

INVX1 _11113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [20]),
    .Y(_2232_)
);

INVX1 _11114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2233_)
);

NOR2X1 _11115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2232_),
    .B(_2233_),
    .Y(_2234_)
);

NOR2X1 _11116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [20]),
    .B(\datapath_1.alu_1.ALUInB [20]),
    .Y(_2235_)
);

NOR2X1 _11117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2234_),
    .Y(_2236_)
);

NOR2X1 _11118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2236_),
    .Y(_2237_)
);

AND2X2 _11119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2237_),
    .B(_2226_),
    .Y(_2238_)
);

NOR2X1 _11120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2239_)
);

NAND2X1 _11121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [18]),
    .B(\datapath_1.alu_1.ALUInB [18]),
    .Y(_2240_)
);

INVX2 _11122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .Y(_2241_)
);

INVX1 _11123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [19]),
    .Y(_2242_)
);

INVX1 _11124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2243_)
);

NOR2X1 _11125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2242_),
    .B(_2243_),
    .Y(_2244_)
);

INVX2 _11126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2244_),
    .Y(_2245_)
);

NOR2X1 _11127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [19]),
    .B(\datapath_1.alu_1.ALUInB [19]),
    .Y(_2246_)
);

INVX1 _11128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .Y(_2247_)
);

NAND2X1 _11129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2247_),
    .B(_2245_),
    .Y(_2248_)
);

OAI21X1 _11130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_2241_),
    .C(_2248_),
    .Y(_2249_)
);

NAND2X1 _11131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2250_)
);

INVX1 _11132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2250_),
    .Y(_2251_)
);

NOR2X1 _11133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [17]),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .Y(_2252_)
);

NAND2X1 _11134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2253_)
);

INVX2 _11135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [16]),
    .Y(_2254_)
);

INVX1 _11136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [16]),
    .Y(_2255_)
);

NAND2X1 _11137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(_2255_),
    .Y(_2256_)
);

NAND2X1 _11138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2253_),
    .B(_2256_),
    .Y(_2257_)
);

OAI21X1 _11139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2251_),
    .B(_2252_),
    .C(_2257_),
    .Y(_2258_)
);

NOR2X1 _11140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2249_),
    .Y(_2259_)
);

NAND2X1 _11141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2238_),
    .B(_2259_),
    .Y(_2260_)
);

AOI21X1 _11142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2216_),
    .B(_2176_),
    .C(_2260_),
    .Y(_2261_)
);

NAND2X1 _11143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2237_),
    .Y(_2262_)
);

NOR2X1 _11144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_2241_),
    .Y(_2263_)
);

NOR2X1 _11145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .B(_2244_),
    .Y(_2264_)
);

NOR2X1 _11146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2264_),
    .Y(_2265_)
);

INVX1 _11147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [17]),
    .Y(_2266_)
);

NOR2X1 _11148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [16]),
    .B(_2254_),
    .Y(_2267_)
);

OAI21X1 _11149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2251_),
    .B(_2252_),
    .C(_2267_),
    .Y(_2268_)
);

OAI21X1 _11150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2266_),
    .B(\datapath_1.alu_1.ALUInB [17]),
    .C(_2268_),
    .Y(_2269_)
);

NAND2X1 _11151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .B(_2265_),
    .Y(_2270_)
);

INVX1 _11152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [18]),
    .Y(_2271_)
);

NOR2X1 _11153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [18]),
    .B(_2271_),
    .Y(_2272_)
);

NOR2X1 _11154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [19]),
    .B(_2242_),
    .Y(_2273_)
);

AOI21X1 _11155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2272_),
    .B(_2248_),
    .C(_2273_),
    .Y(_2274_)
);

AND2X2 _11156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2270_),
    .B(_2274_),
    .Y(_2275_)
);

NOR2X1 _11157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [20]),
    .B(_2232_),
    .Y(_2276_)
);

OAI21X1 _11158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .B(_2230_),
    .C(_2276_),
    .Y(_2277_)
);

OAI21X1 _11159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(\datapath_1.alu_1.ALUInB [21]),
    .C(_2277_),
    .Y(_2278_)
);

INVX1 _11160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [22]),
    .Y(_2279_)
);

NOR2X1 _11161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [22]),
    .B(_2279_),
    .Y(_2280_)
);

OAI21X1 _11162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2223_),
    .B(_2224_),
    .C(_2280_),
    .Y(_2281_)
);

OAI21X1 _11163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(\datapath_1.alu_1.ALUInB [23]),
    .C(_2281_),
    .Y(_2282_)
);

AOI21X1 _11164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2278_),
    .C(_2282_),
    .Y(_2283_)
);

OAI21X1 _11165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2275_),
    .B(_2262_),
    .C(_2283_),
    .Y(_2284_)
);

NOR2X1 _11166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2285_)
);

NAND2X1 _11167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [26]),
    .B(\datapath_1.alu_1.ALUInB [26]),
    .Y(_2286_)
);

INVX1 _11168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2286_),
    .Y(_2287_)
);

NOR2X1 _11169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2285_),
    .B(_2287_),
    .Y(_2288_)
);

INVX4 _11170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .Y(_2289_)
);

NAND2X1 _11171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2290_)
);

INVX2 _11172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2290_),
    .Y(_2291_)
);

NOR2X1 _11173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [27]),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .Y(_2292_)
);

OAI21X1 _11174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2291_),
    .B(_2292_),
    .C(_2289_),
    .Y(_2293_)
);

AND2X2 _11175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2294_)
);

NOR2X1 _11176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2295_)
);

NOR2X1 _11177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2295_),
    .B(_2294_),
    .Y(_2296_)
);

INVX2 _11178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .Y(_2297_)
);

INVX1 _11179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [24]),
    .Y(_2298_)
);

INVX1 _11180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2299_)
);

NOR2X1 _11181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2298_),
    .B(_2299_),
    .Y(_2300_)
);

NOR2X1 _11182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [24]),
    .B(\datapath_1.alu_1.ALUInB [24]),
    .Y(_2301_)
);

OAI21X1 _11183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2301_),
    .C(_2297_),
    .Y(_2302_)
);

NOR2X1 _11184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .B(_2293_),
    .Y(_2303_)
);

OAI21X1 _11185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2261_),
    .B(_2284_),
    .C(_2303_),
    .Y(_2304_)
);

NAND2X1 _11186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [24]),
    .B(_2299_),
    .Y(_2305_)
);

INVX1 _11187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [25]),
    .Y(_2306_)
);

NAND2X1 _11188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [25]),
    .B(_2306_),
    .Y(_2307_)
);

OAI21X1 _11189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2305_),
    .C(_2307_),
    .Y(_2308_)
);

INVX2 _11190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2308_),
    .Y(_2309_)
);

NOR2X1 _11191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2309_),
    .B(_2293_),
    .Y(_2310_)
);

INVX1 _11192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [27]),
    .Y(_2311_)
);

INVX1 _11193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [26]),
    .Y(_2312_)
);

NOR2X1 _11194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [26]),
    .B(_2312_),
    .Y(_2313_)
);

OAI21X1 _11195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2291_),
    .B(_2292_),
    .C(_2313_),
    .Y(_2314_)
);

OAI21X1 _11196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(\datapath_1.alu_1.ALUInB [27]),
    .C(_2314_),
    .Y(_2315_)
);

NOR2X1 _11197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2315_),
    .B(_2310_),
    .Y(_2316_)
);

INVX2 _11198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [29]),
    .Y(_2317_)
);

INVX1 _11199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [29]),
    .Y(_2318_)
);

NOR2X1 _11200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2317_),
    .B(_2318_),
    .Y(_2319_)
);

NOR2X1 _11201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .Y(_2320_)
);

AND2X2 _11202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2321_)
);

NOR2X1 _11203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [28]),
    .B(\datapath_1.alu_1.ALUInB [28]),
    .Y(_2322_)
);

NOR2X1 _11204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .B(_2321_),
    .Y(_2323_)
);

INVX2 _11205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2323_),
    .Y(_2324_)
);

OAI21X1 _11206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2319_),
    .B(_2320_),
    .C(_2324_),
    .Y(_2325_)
);

AOI21X1 _11207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .B(_2304_),
    .C(_2325_),
    .Y(_2326_)
);

INVX1 _11208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [28]),
    .Y(_2327_)
);

NOR2X1 _11209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [28]),
    .B(_2327_),
    .Y(_2328_)
);

OAI21X1 _11210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2319_),
    .B(_2320_),
    .C(_2328_),
    .Y(_2329_)
);

OAI21X1 _11211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2317_),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .C(_2329_),
    .Y(_2330_)
);

OAI21X1 _11212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2326_),
    .B(_2330_),
    .C(_2117_),
    .Y(_2331_)
);

OAI21X1 _11213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2112_),
    .B(\datapath_1.alu_1.ALUInB [30]),
    .C(_2331_),
    .Y(_2332_)
);

INVX2 _11214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUControl[1]),
    .Y(_2333_)
);

NOR2X1 _11215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUControl[0]),
    .B(_2333_),
    .Y(_2334_)
);

INVX1 _11216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUControl[2]),
    .Y(_2335_)
);

NOR2X1 _11217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_2335_),
    .Y(_2336_)
);

NAND2X1 _11218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2334_),
    .B(_2336_),
    .Y(_2337_)
);

AOI21X1 _11219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_2332_),
    .C(_2337_),
    .Y(_2338_)
);

OAI21X1 _11220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_2332_),
    .C(_2338_),
    .Y(_2339_)
);

NOR2X1 _11221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUControl[1]),
    .B(ALUControl[0]),
    .Y(_2340_)
);

AND2X2 _11222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .B(_2340_),
    .Y(_2341_)
);

NAND2X1 _11223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2341__bF$buf3),
    .Y(_2342_)
);

NOR2X1 _11224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(ALUControl[2]),
    .Y(_2343_)
);

NAND3X1 _11225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUControl[1]),
    .B(ALUControl[0]),
    .C(_2343_),
    .Y(_2344_)
);

OAI21X1 _11226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_2344__bF$buf3),
    .C(_2342_),
    .Y(_2345_)
);

NAND2X1 _11227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .B(_2343_),
    .Y(_2346_)
);

NAND3X1 _11228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2333_),
    .B(ALUControl[0]),
    .C(_2343_),
    .Y(_2347_)
);

OAI22X1 _11229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2108_),
    .B(_2346_),
    .C(_2347__bF$buf3),
    .D(_2107_),
    .Y(_2348_)
);

NOR2X1 _11230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2348_),
    .B(_2345_),
    .Y(_2349_)
);

INVX1 _11231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2114_),
    .Y(_2350_)
);

AND2X2 _11232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2351_)
);

NOR2X1 _11233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(\datapath_1.alu_1.ALUInA [2]),
    .Y(_2352_)
);

NOR2X1 _11234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .B(_2351_),
    .Y(_2353_)
);

AND2X2 _11235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2354_)
);

NOR2X1 _11236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(\datapath_1.alu_1.ALUInA [3]),
    .Y(_2355_)
);

NOR2X1 _11237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2355_),
    .B(_2354_),
    .Y(_2356_)
);

NOR2X1 _11238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2357_)
);

NAND2X1 _11239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2358_)
);

OAI21X1 _11240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2358_),
    .C(_2129_),
    .Y(_2359_)
);

NAND3X1 _11241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .B(_2353_),
    .C(_2356_),
    .Y(_2360_)
);

OAI21X1 _11242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2355_),
    .B(_2132_),
    .C(_2122_),
    .Y(_2361_)
);

INVX1 _11243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2361_),
    .Y(_2362_)
);

NAND2X1 _11244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .B(_2360_),
    .Y(_2363_)
);

XOR2X1 _11245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(\datapath_1.alu_1.ALUInA [7]),
    .Y(_2364_)
);

XOR2X1 _11246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2365_)
);

NAND2X1 _11247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2365_),
    .Y(_2366_)
);

XOR2X1 _11248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(\datapath_1.alu_1.ALUInA [5]),
    .Y(_2367_)
);

XOR2X1 _11249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2368_)
);

NAND2X1 _11250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2367_),
    .B(_2368_),
    .Y(_2369_)
);

NOR2X1 _11251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2366_),
    .B(_2369_),
    .Y(_2370_)
);

INVX1 _11252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .Y(_2371_)
);

AOI21X1 _11253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2143_),
    .B(_2371_),
    .C(_2141_),
    .Y(_2372_)
);

INVX1 _11254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2137_),
    .Y(_2373_)
);

AOI21X1 _11255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_2373_),
    .C(_2136_),
    .Y(_2374_)
);

OAI21X1 _11256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2366_),
    .B(_2372_),
    .C(_2374_),
    .Y(_2375_)
);

AOI21X1 _11257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2370_),
    .B(_2363_),
    .C(_2375_),
    .Y(_2376_)
);

NAND2X1 _11258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2162_),
    .Y(_2377_)
);

NAND2X1 _11259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .B(_2165_),
    .Y(_2378_)
);

NOR2X1 _11260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2377_),
    .B(_2378_),
    .Y(_2379_)
);

NAND2X1 _11261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2169_),
    .Y(_2380_)
);

NAND2X1 _11262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2172_),
    .Y(_2381_)
);

NOR2X1 _11263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .B(_2381_),
    .Y(_2382_)
);

NAND2X1 _11264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2382_),
    .Y(_2383_)
);

INVX1 _11265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [9]),
    .Y(_2384_)
);

NOR2X1 _11266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2384_),
    .B(_2195_),
    .Y(_2385_)
);

NOR2X1 _11267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [9]),
    .B(\datapath_1.alu_1.ALUInA [9]),
    .Y(_2386_)
);

INVX1 _11268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .Y(_2387_)
);

INVX2 _11269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2388_)
);

NOR2X1 _11270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2197_),
    .B(_2388_),
    .Y(_2389_)
);

AOI21X1 _11271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .B(_2389_),
    .C(_2385_),
    .Y(_2390_)
);

INVX1 _11272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [11]),
    .Y(_2391_)
);

NOR2X1 _11273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2202_),
    .Y(_2392_)
);

NAND2X1 _11274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2202_),
    .Y(_2393_)
);

AOI21X1 _11275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2393_),
    .B(_2191_),
    .C(_2392_),
    .Y(_2394_)
);

OAI21X1 _11276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .B(_2390_),
    .C(_2394_),
    .Y(_2395_)
);

INVX1 _11277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [13]),
    .Y(_2396_)
);

NOR2X1 _11278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2396_),
    .B(_2206_),
    .Y(_2397_)
);

NOR2X1 _11279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(\datapath_1.alu_1.ALUInA [13]),
    .Y(_2398_)
);

INVX1 _11280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .Y(_2399_)
);

AOI21X1 _11281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2399_),
    .B(_2184_),
    .C(_2397_),
    .Y(_2400_)
);

INVX1 _11282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [15]),
    .Y(_2401_)
);

NOR2X1 _11283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2401_),
    .B(_2212_),
    .Y(_2402_)
);

NOR2X1 _11284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [15]),
    .B(\datapath_1.alu_1.ALUInA [15]),
    .Y(_2403_)
);

INVX2 _11285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2403_),
    .Y(_2404_)
);

AOI21X1 _11286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .B(_2404_),
    .C(_2402_),
    .Y(_2405_)
);

OAI21X1 _11287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2377_),
    .B(_2400_),
    .C(_2405_),
    .Y(_2406_)
);

AOI21X1 _11288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2395_),
    .C(_2406_),
    .Y(_2407_)
);

OAI21X1 _11289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2383_),
    .C(_2407_),
    .Y(_2408_)
);

INVX1 _11290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .Y(_2409_)
);

NAND2X1 _11291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2218_),
    .B(_2409_),
    .Y(_2410_)
);

OR2X2 _11292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2223_),
    .B(_2224_),
    .Y(_2411_)
);

NOR2X1 _11293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2411_),
    .Y(_2412_)
);

NAND2X1 _11294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2236_),
    .Y(_2413_)
);

INVX1 _11295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2413_),
    .Y(_2414_)
);

NAND2X1 _11296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2412_),
    .B(_2414_),
    .Y(_2415_)
);

NAND2X1 _11297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2264_),
    .Y(_2416_)
);

INVX1 _11298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2416_),
    .Y(_2417_)
);

INVX1 _11299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2252_),
    .Y(_2418_)
);

NAND2X1 _11300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2250_),
    .B(_2418_),
    .Y(_2419_)
);

NOR2X1 _11301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .B(_2419_),
    .Y(_2420_)
);

NAND2X1 _11302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2420_),
    .B(_2417_),
    .Y(_2421_)
);

NOR2X1 _11303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2421_),
    .B(_2415_),
    .Y(_2422_)
);

OAI21X1 _11304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2252_),
    .B(_2253_),
    .C(_2250_),
    .Y(_2423_)
);

INVX2 _11305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2423_),
    .Y(_2424_)
);

OAI21X1 _11306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .B(_2240_),
    .C(_2245_),
    .Y(_2425_)
);

INVX1 _11307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2425_),
    .Y(_2426_)
);

OAI21X1 _11308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2416_),
    .B(_2424_),
    .C(_2426_),
    .Y(_2427_)
);

INVX1 _11309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2427_),
    .Y(_2428_)
);

INVX1 _11310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .Y(_2429_)
);

INVX2 _11311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .Y(_2430_)
);

OAI21X1 _11312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .B(_2230_),
    .C(_2429_),
    .Y(_2431_)
);

NAND2X1 _11313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2412_),
    .Y(_2432_)
);

INVX1 _11314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .Y(_2433_)
);

AOI21X1 _11315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2219_),
    .B(_2433_),
    .C(_2223_),
    .Y(_2434_)
);

AND2X2 _11316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .B(_2434_),
    .Y(_2435_)
);

OAI21X1 _11317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2428_),
    .C(_2435_),
    .Y(_2436_)
);

AOI21X1 _11318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2408_),
    .B(_2422_),
    .C(_2436_),
    .Y(_2437_)
);

NOR2X1 _11319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2292_),
    .B(_2291_),
    .Y(_2438_)
);

INVX2 _11320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2438_),
    .Y(_2439_)
);

NOR2X1 _11321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2289_),
    .B(_2439_),
    .Y(_2440_)
);

INVX1 _11322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2440_),
    .Y(_2441_)
);

NOR2X1 _11323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2301_),
    .B(_2300_),
    .Y(_2442_)
);

NAND2X1 _11324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2442_),
    .Y(_2443_)
);

NOR2X1 _11325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2443_),
    .B(_2441_),
    .Y(_2444_)
);

INVX1 _11326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .Y(_2445_)
);

AOI21X1 _11327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2296_),
    .C(_2294_),
    .Y(_2446_)
);

INVX1 _11328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2446_),
    .Y(_2447_)
);

OAI21X1 _11329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2292_),
    .B(_2286_),
    .C(_2290_),
    .Y(_2448_)
);

AOI21X1 _11330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2440_),
    .C(_2448_),
    .Y(_2449_)
);

OAI21X1 _11331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2445_),
    .C(_2449_),
    .Y(_2450_)
);

NOR2X1 _11332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .B(_2319_),
    .Y(_2451_)
);

INVX2 _11333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .Y(_2452_)
);

NOR2X1 _11334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2324_),
    .B(_2452_),
    .Y(_2453_)
);

OAI21X1 _11335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [29]),
    .B(\datapath_1.alu_1.ALUInB [29]),
    .C(_2321_),
    .Y(_2454_)
);

OAI21X1 _11336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2317_),
    .B(_2318_),
    .C(_2454_),
    .Y(_2455_)
);

AOI21X1 _11337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2453_),
    .B(_2450_),
    .C(_2455_),
    .Y(_2456_)
);

OAI21X1 _11338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2115_),
    .C(_2350_),
    .Y(_2457_)
);

NAND2X1 _11339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2343_),
    .B(_2334_),
    .Y(_2458_)
);

AOI21X1 _11340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .B(_2457_),
    .C(_2458_),
    .Y(_2459_)
);

OAI21X1 _11341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .B(_2457_),
    .C(_2459_),
    .Y(_2460_)
);

NAND3X1 _11342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2460_),
    .C(_2339_),
    .Y(\datapath_1.ALUResult [31])
);

NOR2X1 _11343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2330_),
    .B(_2326_),
    .Y(_2461_)
);

INVX8 _11344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .Y(_2462_)
);

OAI21X1 _11345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(_2116_),
    .C(_2462__bF$buf3),
    .Y(_2463_)
);

AOI21X1 _11346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_2461_),
    .C(_2463_),
    .Y(_2464_)
);

NAND2X1 _11347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2341__bF$buf2),
    .Y(_2465_)
);

OAI21X1 _11348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2117_),
    .B(_2344__bF$buf2),
    .C(_2465_),
    .Y(_2466_)
);

OAI22X1 _11349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2347__bF$buf2),
    .C(_2350_),
    .D(_2346_),
    .Y(_2467_)
);

NOR2X1 _11350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2466_),
    .Y(_2468_)
);

AND2X2 _11351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2117_),
    .Y(_2469_)
);

INVX8 _11352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2458_),
    .Y(_2470_)
);

OAI21X1 _11353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2117_),
    .C(_2470__bF$buf3),
    .Y(_2471_)
);

OAI21X1 _11354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2471_),
    .C(_2468_),
    .Y(_2472_)
);

NOR2X1 _11355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2472_),
    .B(_2464_),
    .Y(_2473_)
);

INVX1 _11356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2473_),
    .Y(\datapath_1.ALUResult [30])
);

INVX1 _11357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .Y(_2474_)
);

AOI21X1 _11358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2450_),
    .C(_2321_),
    .Y(_2475_)
);

AND2X2 _11359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(_2452_),
    .Y(_2476_)
);

OAI21X1 _11360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(_2452_),
    .C(_2470__bF$buf2),
    .Y(_2477_)
);

INVX4 _11361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344__bF$buf1),
    .Y(_2478_)
);

INVX1 _11362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .Y(_2479_)
);

NAND2X1 _11363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .B(_2336_),
    .Y(_2480_)
);

INVX8 _11364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2346_),
    .Y(_2481_)
);

NAND2X1 _11365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2319_),
    .B(_2481__bF$buf3),
    .Y(_2482_)
);

OAI21X1 _11366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2480_),
    .C(_2482_),
    .Y(_2483_)
);

AOI21X1 _11367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2478_),
    .C(_2483_),
    .Y(_2484_)
);

OAI21X1 _11368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .B(_2347__bF$buf1),
    .C(_2484_),
    .Y(_2485_)
);

INVX1 _11369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2328_),
    .Y(_2486_)
);

OAI21X1 _11370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2354_),
    .B(_2355_),
    .C(_2121_),
    .Y(_2487_)
);

OAI21X1 _11371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [3]),
    .B(_2118_),
    .C(_2487_),
    .Y(_2488_)
);

INVX1 _11372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2127_),
    .Y(_2489_)
);

INVX1 _11373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .Y(_2490_)
);

AND2X2 _11374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(\datapath_1.alu_1.ALUInA [1]),
    .Y(_2491_)
);

OAI22X1 _11375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2490_),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .C(_2491_),
    .D(_2357_),
    .Y(_2492_)
);

OAI22X1 _11376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2351_),
    .B(_2352_),
    .C(_2354_),
    .D(_2355_),
    .Y(_2493_)
);

AOI21X1 _11377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2489_),
    .C(_2493_),
    .Y(_2494_)
);

NOR2X1 _11378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2140_),
    .B(_2145_),
    .Y(_2495_)
);

OAI21X1 _11379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2494_),
    .B(_2488_),
    .C(_2495_),
    .Y(_2496_)
);

INVX1 _11380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2140_),
    .Y(_2497_)
);

OAI21X1 _11381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2142_),
    .C(_2152_),
    .Y(_2498_)
);

OAI21X1 _11382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [5]),
    .B(_2149_),
    .C(_2498_),
    .Y(_2499_)
);

OAI21X1 _11383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2137_),
    .C(_2156_),
    .Y(_2500_)
);

OAI21X1 _11384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [7]),
    .B(_2157_),
    .C(_2500_),
    .Y(_2501_)
);

AOI21X1 _11385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .B(_2499_),
    .C(_2501_),
    .Y(_2502_)
);

XNOR2X1 _11386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [8]),
    .B(\datapath_1.alu_1.ALUInA [8]),
    .Y(_2503_)
);

OAI21X1 _11387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2386_),
    .C(_2503_),
    .Y(_2504_)
);

NOR2X1 _11388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(_2193_),
    .Y(_2505_)
);

NAND2X1 _11389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2187_),
    .B(_2505_),
    .Y(_2506_)
);

AOI21X1 _11390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2496_),
    .B(_2502_),
    .C(_2506_),
    .Y(_2507_)
);

INVX1 _11391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2196_),
    .Y(_2508_)
);

OAI21X1 _11392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2198_),
    .C(_2508_),
    .Y(_2509_)
);

INVX1 _11393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2201_),
    .Y(_2510_)
);

INVX1 _11394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2203_),
    .Y(_2511_)
);

OAI21X1 _11395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .B(_2171_),
    .C(_2511_),
    .Y(_2512_)
);

AOI21X1 _11396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2509_),
    .C(_2512_),
    .Y(_2513_)
);

OAI21X1 _11397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2397_),
    .B(_2398_),
    .C(_2208_),
    .Y(_2514_)
);

OAI21X1 _11398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [13]),
    .B(_2206_),
    .C(_2514_),
    .Y(_2515_)
);

INVX1 _11399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2214_),
    .Y(_2516_)
);

AOI21X1 _11400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .B(_2515_),
    .C(_2516_),
    .Y(_2517_)
);

OAI21X1 _11401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2167_),
    .B(_2513_),
    .C(_2517_),
    .Y(_2518_)
);

INVX1 _11402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .Y(_2519_)
);

NAND2X1 _11403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2265_),
    .B(_2519_),
    .Y(_2520_)
);

NOR2X1 _11404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2520_),
    .Y(_2521_)
);

OAI21X1 _11405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2507_),
    .B(_2518_),
    .C(_2521_),
    .Y(_2522_)
);

INVX2 _11406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .Y(_2523_)
);

OAI21X1 _11407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2249_),
    .C(_2274_),
    .Y(_2524_)
);

INVX1 _11408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2283_),
    .Y(_2525_)
);

AOI21X1 _11409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2238_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_)
);

INVX1 _11410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2303_),
    .Y(_2527_)
);

AOI21X1 _11411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2526_),
    .B(_2522_),
    .C(_2527_),
    .Y(_2528_)
);

INVX1 _11412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .Y(_2529_)
);

OAI21X1 _11413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2528_),
    .B(_2529_),
    .C(_2324_),
    .Y(_2530_)
);

NAND3X1 _11414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2486_),
    .C(_2530_),
    .Y(_2531_)
);

OAI21X1 _11415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2486_),
    .C(_2462__bF$buf2),
    .Y(_2532_)
);

NOR2X1 _11416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_2326_),
    .Y(_2533_)
);

AOI21X1 _11417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2531_),
    .B(_2533_),
    .C(_2485_),
    .Y(_2534_)
);

OAI21X1 _11418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2476_),
    .B(_2477_),
    .C(_2534_),
    .Y(\datapath_1.ALUResult [29])
);

NAND3X1 _11419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .B(_2323_),
    .C(_2304_),
    .Y(_2535_)
);

NAND3X1 _11420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf1),
    .B(_2535_),
    .C(_2530_),
    .Y(_2536_)
);

OAI22X1 _11421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2480_),
    .C(_2324_),
    .D(_2344__bF$buf0),
    .Y(_2537_)
);

NAND2X1 _11422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2321_),
    .B(_2481__bF$buf2),
    .Y(_2538_)
);

OAI21X1 _11423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .B(_2347__bF$buf0),
    .C(_2538_),
    .Y(_2539_)
);

NOR2X1 _11424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2537_),
    .B(_2539_),
    .Y(_2540_)
);

NAND2X1 _11425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2132_),
    .B(_2133_),
    .Y(_2541_)
);

AND2X2 _11426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2542_)
);

AOI21X1 _11427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2542_),
    .B(_2130_),
    .C(_2491_),
    .Y(_2543_)
);

NOR3X1 _11428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2541_),
    .B(_2124_),
    .C(_2543_),
    .Y(_2544_)
);

OAI21X1 _11429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2544_),
    .B(_2361_),
    .C(_2370_),
    .Y(_2545_)
);

INVX1 _11430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2375_),
    .Y(_2546_)
);

AOI21X1 _11431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .B(_2545_),
    .C(_2383_),
    .Y(_2547_)
);

INVX2 _11432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2407_),
    .Y(_2548_)
);

OAI21X1 _11433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2548_),
    .C(_2422_),
    .Y(_2549_)
);

NAND2X1 _11434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2220_),
    .B(_2225_),
    .Y(_2550_)
);

NOR2X1 _11435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2550_),
    .B(_2413_),
    .Y(_2551_)
);

INVX2 _11436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .Y(_2552_)
);

OAI21X1 _11437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2552_),
    .B(_2550_),
    .C(_2434_),
    .Y(_2553_)
);

AOI21X1 _11438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(_2427_),
    .C(_2553_),
    .Y(_2554_)
);

AOI21X1 _11439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2549_),
    .C(_2445_),
    .Y(_2555_)
);

INVX1 _11440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .Y(_2556_)
);

OAI21X1 _11441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2555_),
    .B(_2556_),
    .C(_2323_),
    .Y(_2557_)
);

XNOR2X1 _11442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [6]),
    .B(\datapath_1.alu_1.ALUInA [6]),
    .Y(_2558_)
);

NOR2X1 _11443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2154_),
    .B(_2558_),
    .Y(_2559_)
);

XNOR2X1 _11444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(\datapath_1.alu_1.ALUInA [4]),
    .Y(_2560_)
);

NOR2X1 _11445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2148_),
    .B(_2560_),
    .Y(_2561_)
);

NAND2X1 _11446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2559_),
    .B(_2561_),
    .Y(_2562_)
);

AOI21X1 _11447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2362_),
    .C(_2562_),
    .Y(_2563_)
);

AND2X2 _11448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2382_),
    .Y(_2564_)
);

OAI21X1 _11449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2563_),
    .B(_2375_),
    .C(_2564_),
    .Y(_2565_)
);

INVX1 _11450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2420_),
    .Y(_2566_)
);

NOR2X1 _11451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2416_),
    .B(_2566_),
    .Y(_2567_)
);

NAND2X1 _11452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(_2567_),
    .Y(_2568_)
);

AOI21X1 _11453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2407_),
    .B(_2565_),
    .C(_2568_),
    .Y(_2569_)
);

OAI21X1 _11454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2569_),
    .B(_2436_),
    .C(_2444_),
    .Y(_2570_)
);

NAND3X1 _11455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2324_),
    .B(_2449_),
    .C(_2570_),
    .Y(_2571_)
);

NAND3X1 _11456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf1),
    .B(_2557_),
    .C(_2571_),
    .Y(_2572_)
);

NAND3X1 _11457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_2536_),
    .C(_2572_),
    .Y(\datapath_1.ALUResult [28])
);

INVX1 _11458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2313_),
    .Y(_2573_)
);

AOI21X1 _11459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2526_),
    .B(_2522_),
    .C(_2302_),
    .Y(_2574_)
);

OAI21X1 _11460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2574_),
    .B(_2308_),
    .C(_2289_),
    .Y(_2575_)
);

NAND3X1 _11461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2438_),
    .B(_2573_),
    .C(_2575_),
    .Y(_2576_)
);

INVX1 _11462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .Y(_2577_)
);

OAI21X1 _11463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2261_),
    .B(_2284_),
    .C(_2577_),
    .Y(_2578_)
);

AOI21X1 _11464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2309_),
    .B(_2578_),
    .C(_2288_),
    .Y(_2579_)
);

OAI21X1 _11465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2579_),
    .B(_2313_),
    .C(_2439_),
    .Y(_2580_)
);

NAND3X1 _11466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf0),
    .B(_2576_),
    .C(_2580_),
    .Y(_2581_)
);

INVX1 _11467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2292_),
    .Y(_2582_)
);

OAI22X1 _11468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2290_),
    .B(_2346_),
    .C(_2480_),
    .D(_2582_),
    .Y(_2583_)
);

OAI21X1 _11469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344__bF$buf3),
    .B(_2291_),
    .C(_2347__bF$buf3),
    .Y(_2584_)
);

AOI21X1 _11470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2582_),
    .B(_2584_),
    .C(_2583_),
    .Y(_2585_)
);

AOI21X1 _11471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2549_),
    .C(_2443_),
    .Y(_2586_)
);

OAI21X1 _11472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .B(_2447_),
    .C(_2288_),
    .Y(_2587_)
);

NAND3X1 _11473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2286_),
    .B(_2439_),
    .C(_2587_),
    .Y(_2588_)
);

INVX1 _11474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2443_),
    .Y(_2589_)
);

OAI21X1 _11475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2569_),
    .B(_2436_),
    .C(_2589_),
    .Y(_2590_)
);

AOI21X1 _11476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2446_),
    .B(_2590_),
    .C(_2289_),
    .Y(_2591_)
);

OAI21X1 _11477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2591_),
    .B(_2287_),
    .C(_2438_),
    .Y(_2592_)
);

NAND3X1 _11478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf0),
    .B(_2588_),
    .C(_2592_),
    .Y(_2593_)
);

NAND3X1 _11479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2581_),
    .B(_2585_),
    .C(_2593_),
    .Y(\datapath_1.ALUResult [27])
);

NAND3X1 _11480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .B(_2309_),
    .C(_2578_),
    .Y(_2594_)
);

NAND3X1 _11481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf3),
    .B(_2594_),
    .C(_2575_),
    .Y(_2595_)
);

NAND2X1 _11482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2285_),
    .B(_2341__bF$buf1),
    .Y(_2596_)
);

OAI21X1 _11483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2289_),
    .B(_2344__bF$buf2),
    .C(_2596_),
    .Y(_2597_)
);

OAI22X1 _11484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2286_),
    .B(_2346_),
    .C(_2347__bF$buf2),
    .D(_2285_),
    .Y(_2598_)
);

NOR2X1 _11485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2598_),
    .B(_2597_),
    .Y(_2599_)
);

NAND3X1 _11486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2289_),
    .B(_2446_),
    .C(_2590_),
    .Y(_2600_)
);

NAND3X1 _11487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf3),
    .B(_2587_),
    .C(_2600_),
    .Y(_2601_)
);

NAND3X1 _11488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_2595_),
    .C(_2601_),
    .Y(\datapath_1.ALUResult [26])
);

INVX1 _11489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2301_),
    .Y(_2602_)
);

NAND2X1 _11490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2549_),
    .Y(_2603_)
);

AOI21X1 _11491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2603_),
    .C(_2300_),
    .Y(_2604_)
);

AND2X2 _11492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .B(_2297_),
    .Y(_2605_)
);

OAI21X1 _11493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .B(_2297_),
    .C(_2470__bF$buf2),
    .Y(_2606_)
);

NAND2X1 _11494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2478_),
    .Y(_2607_)
);

AOI22X1 _11495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2294_),
    .B(_2481__bF$buf1),
    .C(_2341__bF$buf0),
    .D(_2295_),
    .Y(_2608_)
);

AND2X2 _11496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2608_),
    .B(_2607_),
    .Y(_2609_)
);

OAI21X1 _11497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2295_),
    .B(_2347__bF$buf1),
    .C(_2609_),
    .Y(_2610_)
);

INVX2 _11498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .Y(_2611_)
);

OAI21X1 _11499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2261_),
    .B(_2284_),
    .C(_2611_),
    .Y(_2612_)
);

NAND3X1 _11500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2305_),
    .C(_2612_),
    .Y(_2613_)
);

OAI21X1 _11501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2305_),
    .C(_2462__bF$buf2),
    .Y(_2614_)
);

NOR2X1 _11502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2614_),
    .B(_2574_),
    .Y(_2615_)
);

AOI21X1 _11503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2615_),
    .B(_2613_),
    .C(_2610_),
    .Y(_2616_)
);

OAI21X1 _11504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2605_),
    .B(_2606_),
    .C(_2616_),
    .Y(\datapath_1.ALUResult [25])
);

NOR2X1 _11505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2284_),
    .B(_2261_),
    .Y(_2617_)
);

NAND2X1 _11506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf1),
    .B(_2612_),
    .Y(_2618_)
);

AOI21X1 _11507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2617_),
    .B(_2442_),
    .C(_2618_),
    .Y(_2619_)
);

INVX8 _11508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347__bF$buf0),
    .Y(_2620_)
);

AOI22X1 _11509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2481__bF$buf0),
    .C(_2341__bF$buf3),
    .D(_2301_),
    .Y(_2621_)
);

OAI21X1 _11510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2611_),
    .B(_2344__bF$buf1),
    .C(_2621_),
    .Y(_2622_)
);

AOI21X1 _11511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2620_),
    .C(_2622_),
    .Y(_2623_)
);

NOR2X1 _11512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .B(_2603_),
    .Y(_2624_)
);

OAI21X1 _11513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2611_),
    .C(_2470__bF$buf1),
    .Y(_2625_)
);

OAI21X1 _11514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2625_),
    .B(_2624_),
    .C(_2623_),
    .Y(_2626_)
);

NOR2X1 _11515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2619_),
    .B(_2626_),
    .Y(_2627_)
);

INVX1 _11516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2627_),
    .Y(\datapath_1.ALUResult [24])
);

INVX1 _11517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2280_),
    .Y(_2628_)
);

INVX1 _11518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2237_),
    .Y(_2629_)
);

OAI21X1 _11519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2507_),
    .B(_2518_),
    .C(_2259_),
    .Y(_2630_)
);

AOI21X1 _11520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2275_),
    .B(_2630_),
    .C(_2629_),
    .Y(_2631_)
);

OAI21X1 _11521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_2278_),
    .C(_2410_),
    .Y(_2632_)
);

NAND3X1 _11522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2225_),
    .B(_2628_),
    .C(_2632_),
    .Y(_2633_)
);

INVX1 _11523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2278_),
    .Y(_2634_)
);

AOI21X1 _11524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2216_),
    .B(_2176_),
    .C(_2520_),
    .Y(_2635_)
);

OAI21X1 _11525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2635_),
    .B(_2524_),
    .C(_2237_),
    .Y(_2636_)
);

AOI21X1 _11526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2634_),
    .B(_2636_),
    .C(_2220_),
    .Y(_2637_)
);

OAI21X1 _11527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2637_),
    .B(_2280_),
    .C(_2411_),
    .Y(_2638_)
);

NAND3X1 _11528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf0),
    .B(_2633_),
    .C(_2638_),
    .Y(_2639_)
);

AOI22X1 _11529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2223_),
    .B(_2481__bF$buf3),
    .C(_2341__bF$buf2),
    .D(_2224_),
    .Y(_2640_)
);

OAI21X1 _11530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2411_),
    .B(_2344__bF$buf0),
    .C(_2640_),
    .Y(_2641_)
);

AOI21X1 _11531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(_2620_),
    .C(_2641_),
    .Y(_2642_)
);

OAI21X1 _11532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2548_),
    .C(_2567_),
    .Y(_2643_)
);

AOI21X1 _11533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2428_),
    .B(_2643_),
    .C(_2413_),
    .Y(_2644_)
);

OAI21X1 _11534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2644_),
    .B(_2431_),
    .C(_2220_),
    .Y(_2645_)
);

NAND3X1 _11535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2218_),
    .B(_2411_),
    .C(_2645_),
    .Y(_2646_)
);

AOI21X1 _11536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2407_),
    .B(_2565_),
    .C(_2421_),
    .Y(_2647_)
);

OAI21X1 _11537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2647_),
    .B(_2427_),
    .C(_2414_),
    .Y(_2648_)
);

AOI21X1 _11538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2552_),
    .B(_2648_),
    .C(_2410_),
    .Y(_2649_)
);

OAI21X1 _11539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .B(_2219_),
    .C(_2225_),
    .Y(_2650_)
);

NAND3X1 _11540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf0),
    .B(_2646_),
    .C(_2650_),
    .Y(_2651_)
);

NAND3X1 _11541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2639_),
    .B(_2642_),
    .C(_2651_),
    .Y(\datapath_1.ALUResult [23])
);

NAND3X1 _11542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2220_),
    .B(_2634_),
    .C(_2636_),
    .Y(_2652_)
);

NAND3X1 _11543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf3),
    .B(_2652_),
    .C(_2632_),
    .Y(_2653_)
);

AOI22X1 _11544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2219_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf1),
    .D(_2217_),
    .Y(_2654_)
);

OAI21X1 _11545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2344__bF$buf3),
    .C(_2654_),
    .Y(_2655_)
);

AOI21X1 _11546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2409_),
    .B(_2620_),
    .C(_2655_),
    .Y(_2656_)
);

NAND3X1 _11547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2552_),
    .C(_2648_),
    .Y(_2657_)
);

NAND3X1 _11548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf3),
    .B(_2645_),
    .C(_2657_),
    .Y(_2658_)
);

NAND3X1 _11549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2653_),
    .B(_2656_),
    .C(_2658_),
    .Y(\datapath_1.ALUResult [22])
);

AOI21X1 _11550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2567_),
    .B(_2408_),
    .C(_2427_),
    .Y(_2659_)
);

OAI21X1 _11551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .B(_2235_),
    .C(_2430_),
    .Y(_2660_)
);

AND2X2 _11552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2660_),
    .B(_2231_),
    .Y(_2661_)
);

OAI21X1 _11553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2660_),
    .B(_2231_),
    .C(_2470__bF$buf2),
    .Y(_2662_)
);

AOI22X1 _11554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2231_),
    .C(_2230_),
    .D(_2341__bF$buf0),
    .Y(_2663_)
);

NOR2X1 _11555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2230_),
    .B(_2347__bF$buf3),
    .Y(_2664_)
);

AOI21X1 _11556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .B(_2481__bF$buf1),
    .C(_2664_),
    .Y(_2665_)
);

AND2X2 _11557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2663_),
    .B(_2665_),
    .Y(_2666_)
);

INVX1 _11558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .Y(_2667_)
);

INVX1 _11559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2276_),
    .Y(_2668_)
);

INVX1 _11560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .Y(_2669_)
);

NAND2X1 _11561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .B(_2430_),
    .Y(_2670_)
);

OAI21X1 _11562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2635_),
    .B(_2524_),
    .C(_2670_),
    .Y(_2671_)
);

NAND3X1 _11563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2668_),
    .C(_2671_),
    .Y(_2672_)
);

OAI21X1 _11564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2668_),
    .C(_2462__bF$buf2),
    .Y(_2673_)
);

NOR2X1 _11565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2673_),
    .B(_2631_),
    .Y(_2674_)
);

AOI21X1 _11566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2674_),
    .B(_2672_),
    .C(_2667_),
    .Y(_2675_)
);

OAI21X1 _11567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2662_),
    .C(_2675_),
    .Y(\datapath_1.ALUResult [21])
);

NOR2X1 _11568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2518_),
    .B(_2507_),
    .Y(_2676_)
);

OAI21X1 _11569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2676_),
    .B(_2520_),
    .C(_2275_),
    .Y(_2677_)
);

INVX1 _11570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .Y(_2678_)
);

NAND2X1 _11571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf1),
    .B(_2671_),
    .Y(_2679_)
);

AOI21X1 _11572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2236_),
    .B(_2678_),
    .C(_2679_),
    .Y(_2680_)
);

AOI22X1 _11573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .B(_2481__bF$buf0),
    .C(_2341__bF$buf3),
    .D(_2235_),
    .Y(_2681_)
);

OAI21X1 _11574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2670_),
    .B(_2344__bF$buf2),
    .C(_2681_),
    .Y(_2682_)
);

AOI21X1 _11575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .B(_2620_),
    .C(_2682_),
    .Y(_2683_)
);

AND2X2 _11576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .B(_2670_),
    .Y(_2684_)
);

OAI21X1 _11577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .B(_2670_),
    .C(_2470__bF$buf1),
    .Y(_2685_)
);

OAI21X1 _11578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2684_),
    .B(_2685_),
    .C(_2683_),
    .Y(_2686_)
);

NOR2X1 _11579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .B(_2680_),
    .Y(_2687_)
);

INVX1 _11580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2687_),
    .Y(\datapath_1.ALUResult [20])
);

OAI21X1 _11581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2507_),
    .B(_2518_),
    .C(_2519_),
    .Y(_2688_)
);

AOI21X1 _11582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2688_),
    .C(_2263_),
    .Y(_2689_)
);

OAI21X1 _11583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_2272_),
    .C(_2248_),
    .Y(_2690_)
);

INVX1 _11584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2272_),
    .Y(_2691_)
);

INVX2 _11585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .Y(_2692_)
);

AOI21X1 _11586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2216_),
    .B(_2176_),
    .C(_2258_),
    .Y(_2693_)
);

OAI21X1 _11587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2693_),
    .B(_2269_),
    .C(_2692_),
    .Y(_2694_)
);

NAND3X1 _11588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2264_),
    .B(_2691_),
    .C(_2694_),
    .Y(_2695_)
);

NAND3X1 _11589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf0),
    .B(_2695_),
    .C(_2690_),
    .Y(_2696_)
);

OAI22X1 _11590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2247_),
    .B(_2480_),
    .C(_2248_),
    .D(_2344__bF$buf1),
    .Y(_2697_)
);

OAI22X1 _11591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .B(_2347__bF$buf2),
    .C(_2245_),
    .D(_2346_),
    .Y(_2698_)
);

NOR2X1 _11592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2698_),
    .B(_2697_),
    .Y(_2699_)
);

AOI21X1 _11593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2407_),
    .B(_2565_),
    .C(_2566_),
    .Y(_2700_)
);

OAI21X1 _11594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2423_),
    .C(_2263_),
    .Y(_2701_)
);

NAND3X1 _11595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .B(_2248_),
    .C(_2701_),
    .Y(_2702_)
);

OAI21X1 _11596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2548_),
    .C(_2420_),
    .Y(_2703_)
);

AOI21X1 _11597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2703_),
    .C(_2692_),
    .Y(_2704_)
);

OAI21X1 _11598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2704_),
    .B(_2241_),
    .C(_2264_),
    .Y(_2705_)
);

NAND3X1 _11599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf0),
    .B(_2705_),
    .C(_2702_),
    .Y(_2706_)
);

NAND3X1 _11600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2696_),
    .B(_2699_),
    .C(_2706_),
    .Y(\datapath_1.ALUResult [19])
);

OAI21X1 _11601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2676_),
    .B(_2258_),
    .C(_2523_),
    .Y(_2707_)
);

INVX1 _11602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .Y(_2708_)
);

NAND2X1 _11603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf3),
    .B(_2694_),
    .Y(_2709_)
);

AOI21X1 _11604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2708_),
    .C(_2709_),
    .Y(_2710_)
);

NAND2X1 _11605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_2341__bF$buf2),
    .Y(_2711_)
);

OAI21X1 _11606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2344__bF$buf0),
    .C(_2711_),
    .Y(_2712_)
);

OAI22X1 _11607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .B(_2346_),
    .C(_2347__bF$buf1),
    .D(_2239_),
    .Y(_2713_)
);

NOR2X1 _11608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2713_),
    .B(_2712_),
    .Y(_2714_)
);

NAND3X1 _11609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2424_),
    .C(_2703_),
    .Y(_2715_)
);

NAND2X1 _11610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2715_),
    .B(_2701_),
    .Y(_2716_)
);

OAI21X1 _11611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2716_),
    .B(_2458_),
    .C(_2714_),
    .Y(_2717_)
);

NOR2X1 _11612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2710_),
    .B(_2717_),
    .Y(_2718_)
);

INVX1 _11613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2718_),
    .Y(\datapath_1.ALUResult [18])
);

INVX1 _11614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2419_),
    .Y(_2719_)
);

INVX2 _11615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .Y(_2720_)
);

OAI21X1 _11616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2548_),
    .C(_2720_),
    .Y(_2721_)
);

OAI21X1 _11617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(_2255_),
    .C(_2721_),
    .Y(_2722_)
);

OR2X2 _11618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2722_),
    .B(_2719_),
    .Y(_2723_)
);

AOI21X1 _11619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2719_),
    .B(_2722_),
    .C(_2458_),
    .Y(_2724_)
);

OAI22X1 _11620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .B(_2418_),
    .C(_2419_),
    .D(_2344__bF$buf3),
    .Y(_2725_)
);

OAI22X1 _11621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2250_),
    .B(_2346_),
    .C(_2347__bF$buf0),
    .D(_2252_),
    .Y(_2726_)
);

NOR2X1 _11622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2726_),
    .B(_2725_),
    .Y(_2727_)
);

OAI21X1 _11623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2507_),
    .B(_2518_),
    .C(_2257_),
    .Y(_2728_)
);

OAI21X1 _11624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .C(_2728_),
    .Y(_2729_)
);

NOR2X1 _11625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2419_),
    .B(_2729_),
    .Y(_2730_)
);

NAND3X1 _11626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2268_),
    .B(_2462__bF$buf2),
    .C(_2688_),
    .Y(_2731_)
);

OAI21X1 _11627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2730_),
    .B(_2731_),
    .C(_2727_),
    .Y(_2732_)
);

AOI21X1 _11628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2723_),
    .B(_2724_),
    .C(_2732_),
    .Y(_2733_)
);

INVX1 _11629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .Y(\datapath_1.ALUResult [17])
);

NAND2X1 _11630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2720_),
    .B(_2676_),
    .Y(_2734_)
);

NAND3X1 _11631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf1),
    .B(_2728_),
    .C(_2734_),
    .Y(_2735_)
);

OAI22X1 _11632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .B(_2344__bF$buf2),
    .C(_2480_),
    .D(_2256_),
    .Y(_2736_)
);

OAI21X1 _11633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [16]),
    .B(\datapath_1.alu_1.ALUInB [16]),
    .C(_2620_),
    .Y(_2737_)
);

OAI21X1 _11634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2253_),
    .B(_2346_),
    .C(_2737_),
    .Y(_2738_)
);

NOR2X1 _11635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .B(_2738_),
    .Y(_2739_)
);

AOI21X1 _11636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2720_),
    .B(_2408_),
    .C(_2458_),
    .Y(_2740_)
);

OAI21X1 _11637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2720_),
    .B(_2408_),
    .C(_2740_),
    .Y(_2741_)
);

NAND3X1 _11638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2739_),
    .B(_2741_),
    .C(_2735_),
    .Y(\datapath_1.ALUResult [16])
);

AOI21X1 _11639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2496_),
    .C(_2174_),
    .Y(_2742_)
);

OAI21X1 _11640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2742_),
    .B(_2205_),
    .C(_2166_),
    .Y(_2743_)
);

AOI21X1 _11641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2209_),
    .B(_2743_),
    .C(_2162_),
    .Y(_2744_)
);

NOR2X1 _11642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .B(_2744_),
    .Y(_2745_)
);

AOI21X1 _11643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2745_),
    .C(_2337_),
    .Y(_2746_)
);

OAI21X1 _11644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2745_),
    .C(_2746_),
    .Y(_2747_)
);

NAND2X1 _11645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2402_),
    .B(_2481__bF$buf3),
    .Y(_2748_)
);

OAI21X1 _11646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .B(_2480_),
    .C(_2748_),
    .Y(_2749_)
);

OAI21X1 _11647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344__bF$buf1),
    .B(_2402_),
    .C(_2347__bF$buf3),
    .Y(_2750_)
);

AOI21X1 _11648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .B(_2750_),
    .C(_2749_),
    .Y(_2751_)
);

INVX2 _11649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2162_),
    .Y(_2752_)
);

INVX1 _11650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .Y(_2753_)
);

INVX1 _11651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2400_),
    .Y(_2754_)
);

INVX1 _11652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2382_),
    .Y(_2755_)
);

INVX1 _11653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2395_),
    .Y(_2756_)
);

OAI21X1 _11654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2755_),
    .C(_2756_),
    .Y(_2757_)
);

AOI21X1 _11655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2753_),
    .B(_2757_),
    .C(_2754_),
    .Y(_2758_)
);

NOR2X1 _11656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2758_),
    .Y(_2759_)
);

NOR2X1 _11657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .B(_2759_),
    .Y(_2760_)
);

OAI21X1 _11658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2402_),
    .B(_2403_),
    .C(_2760_),
    .Y(_2761_)
);

OAI21X1 _11659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2759_),
    .B(_2178_),
    .C(_2161_),
    .Y(_2762_)
);

NAND3X1 _11660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470__bF$buf3),
    .B(_2762_),
    .C(_2761_),
    .Y(_2763_)
);

NAND3X1 _11661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2747_),
    .B(_2751_),
    .C(_2763_),
    .Y(\datapath_1.ALUResult [15])
);

NOR2X1 _11662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2205_),
    .B(_2742_),
    .Y(_2764_)
);

OAI21X1 _11663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2764_),
    .B(_2186_),
    .C(_2209_),
    .Y(_2765_)
);

NOR2X1 _11664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2765_),
    .Y(_2766_)
);

NOR3X1 _11665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2744_),
    .C(_2766_),
    .Y(_2767_)
);

NAND2X1 _11666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2179_),
    .B(_2341__bF$buf1),
    .Y(_2768_)
);

OAI21X1 _11667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2344__bF$buf0),
    .C(_2768_),
    .Y(_2769_)
);

NAND2X1 _11668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .B(_2481__bF$buf2),
    .Y(_2770_)
);

OAI21X1 _11669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2179_),
    .B(_2347__bF$buf2),
    .C(_2770_),
    .Y(_2771_)
);

NOR2X1 _11670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2771_),
    .B(_2769_),
    .Y(_2772_)
);

AND2X2 _11671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(_2752_),
    .Y(_2773_)
);

OAI21X1 _11672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(_2752_),
    .C(_2470__bF$buf2),
    .Y(_2774_)
);

OAI21X1 _11673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2773_),
    .B(_2774_),
    .C(_2772_),
    .Y(_2775_)
);

NOR2X1 _11674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2775_),
    .B(_2767_),
    .Y(_2776_)
);

INVX1 _11675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2776_),
    .Y(\datapath_1.ALUResult [14])
);

NAND2X1 _11676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2757_),
    .Y(_2777_)
);

OAI21X1 _11677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2183_),
    .C(_2777_),
    .Y(_2778_)
);

OR2X2 _11678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2778_),
    .B(_2164_),
    .Y(_2779_)
);

AOI21X1 _11679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .B(_2778_),
    .C(_2458_),
    .Y(_2780_)
);

OAI22X1 _11680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2181_),
    .B(_2344__bF$buf3),
    .C(_2480_),
    .D(_2399_),
    .Y(_2781_)
);

NAND2X1 _11681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2397_),
    .B(_2481__bF$buf1),
    .Y(_2782_)
);

OAI21X1 _11682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .B(_2347__bF$buf1),
    .C(_2782_),
    .Y(_2783_)
);

NOR2X1 _11683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2781_),
    .B(_2783_),
    .Y(_2784_)
);

NOR2X1 _11684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2764_),
    .Y(_2785_)
);

OAI21X1 _11685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [12]),
    .B(_2183_),
    .C(_2164_),
    .Y(_2786_)
);

NOR2X1 _11686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2786_),
    .B(_2785_),
    .Y(_2787_)
);

NAND3X1 _11687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2514_),
    .B(_2462__bF$buf0),
    .C(_2743_),
    .Y(_2788_)
);

OAI21X1 _11688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2787_),
    .B(_2788_),
    .C(_2784_),
    .Y(_2789_)
);

AOI21X1 _11689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2779_),
    .B(_2780_),
    .C(_2789_),
    .Y(_2790_)
);

INVX1 _11690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2790_),
    .Y(\datapath_1.ALUResult [13])
);

OAI21X1 _11691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2764_),
    .B(_2165_),
    .C(_2462__bF$buf3),
    .Y(_2791_)
);

AOI21X1 _11692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2764_),
    .C(_2791_),
    .Y(_2792_)
);

NAND2X1 _11693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2480_),
    .Y(_2793_)
);

OAI21X1 _11694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2620_),
    .C(_2793_),
    .Y(_2794_)
);

AOI22X1 _11695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2184_),
    .B(_2481__bF$buf0),
    .C(_2478_),
    .D(_2165_),
    .Y(_2795_)
);

AOI21X1 _11696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2757_),
    .C(_2458_),
    .Y(_2796_)
);

OAI21X1 _11697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2165_),
    .B(_2757_),
    .C(_2796_),
    .Y(_2797_)
);

NAND3X1 _11698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2794_),
    .B(_2795_),
    .C(_2797_),
    .Y(_2798_)
);

NOR2X1 _11699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_2798_),
    .Y(_2799_)
);

INVX1 _11700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .Y(\datapath_1.ALUResult [12])
);

INVX1 _11701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .Y(_2800_)
);

AOI21X1 _11702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2496_),
    .C(_2504_),
    .Y(_2801_)
);

OAI21X1 _11703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2509_),
    .C(_2800_),
    .Y(_2802_)
);

OAI21X1 _11704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [10]),
    .B(_2190_),
    .C(_2802_),
    .Y(_2803_)
);

OAI21X1 _11705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2803_),
    .B(_2188_),
    .C(_2462__bF$buf2),
    .Y(_2804_)
);

AOI21X1 _11706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2188_),
    .B(_2803_),
    .C(_2804_),
    .Y(_2805_)
);

OAI21X1 _11707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [11]),
    .B(\datapath_1.alu_1.ALUInA [11]),
    .C(_2347__bF$buf0),
    .Y(_2806_)
);

OAI21X1 _11708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341__bF$buf0),
    .B(_2393_),
    .C(_2806_),
    .Y(_2807_)
);

AOI22X1 _11709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2481__bF$buf3),
    .C(_2478_),
    .D(_2171_),
    .Y(_2808_)
);

AND2X2 _11710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2807_),
    .B(_2808_),
    .Y(_2809_)
);

INVX1 _11711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2192_),
    .Y(_2810_)
);

OAI21X1 _11712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2380_),
    .C(_2390_),
    .Y(_2811_)
);

AOI21X1 _11713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(_2811_),
    .C(_2191_),
    .Y(_2812_)
);

AND2X2 _11714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2812_),
    .B(_2188_),
    .Y(_2813_)
);

OAI21X1 _11715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2812_),
    .B(_2188_),
    .C(_2470__bF$buf1),
    .Y(_2814_)
);

OAI21X1 _11716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2813_),
    .B(_2814_),
    .C(_2809_),
    .Y(_2815_)
);

NOR2X1 _11717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2815_),
    .B(_2805_),
    .Y(_2816_)
);

INVX1 _11718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_),
    .Y(\datapath_1.ALUResult [11])
);

NOR2X1 _11719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2509_),
    .B(_2801_),
    .Y(_2817_)
);

NAND2X1 _11720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2817_),
    .Y(_2818_)
);

NAND3X1 _11721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf1),
    .B(_2802_),
    .C(_2818_),
    .Y(_2819_)
);

AOI22X1 _11722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2191_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf3),
    .D(_2192_),
    .Y(_2820_)
);

OAI21X1 _11723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2800_),
    .B(_2344__bF$buf2),
    .C(_2820_),
    .Y(_2821_)
);

AOI21X1 _11724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(_2620_),
    .C(_2821_),
    .Y(_2822_)
);

AOI21X1 _11725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2811_),
    .C(_2458_),
    .Y(_2823_)
);

OAI21X1 _11726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2811_),
    .C(_2823_),
    .Y(_2824_)
);

NAND3X1 _11727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2822_),
    .B(_2824_),
    .C(_2819_),
    .Y(\datapath_1.ALUResult [10])
);

OAI21X1 _11728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2563_),
    .B(_2375_),
    .C(_2169_),
    .Y(_2825_)
);

OAI21X1 _11729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2197_),
    .B(_2388_),
    .C(_2825_),
    .Y(_2826_)
);

AND2X2 _11730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2168_),
    .Y(_2827_)
);

OAI21X1 _11731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2168_),
    .C(_2470__bF$buf0),
    .Y(_2828_)
);

NAND2X1 _11732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2481__bF$buf1),
    .Y(_2829_)
);

OAI21X1 _11733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .B(_2480_),
    .C(_2829_),
    .Y(_2830_)
);

AOI21X1 _11734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2478_),
    .C(_2830_),
    .Y(_2831_)
);

OAI21X1 _11735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .B(_2347__bF$buf3),
    .C(_2831_),
    .Y(_2832_)
);

OAI21X1 _11736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2147_),
    .B(_2160_),
    .C(_2503_),
    .Y(_2833_)
);

NAND3X1 _11737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2198_),
    .C(_2833_),
    .Y(_2834_)
);

OAI21X1 _11738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2198_),
    .C(_2462__bF$buf0),
    .Y(_2835_)
);

NOR2X1 _11739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2835_),
    .B(_2801_),
    .Y(_2836_)
);

AOI21X1 _11740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2836_),
    .B(_2834_),
    .C(_2832_),
    .Y(_2837_)
);

OAI21X1 _11741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2827_),
    .B(_2828_),
    .C(_2837_),
    .Y(\datapath_1.ALUResult [9])
);

NOR2X1 _11742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2160_),
    .B(_2147_),
    .Y(_2838_)
);

NAND2X1 _11743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf3),
    .B(_2833_),
    .Y(_2839_)
);

AOI21X1 _11744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2838_),
    .B(_2169_),
    .C(_2839_),
    .Y(_2840_)
);

NAND2X1 _11745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2197_),
    .B(_2388_),
    .Y(_2841_)
);

NAND2X1 _11746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2389_),
    .B(_2481__bF$buf0),
    .Y(_2842_)
);

OAI21X1 _11747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2480_),
    .C(_2842_),
    .Y(_2843_)
);

OAI21X1 _11748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344__bF$buf1),
    .B(_2389_),
    .C(_2347__bF$buf2),
    .Y(_2844_)
);

AOI21X1 _11749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2844_),
    .C(_2843_),
    .Y(_2845_)
);

AND2X2 _11750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2503_),
    .Y(_2846_)
);

OAI21X1 _11751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2503_),
    .C(_2470__bF$buf3),
    .Y(_2847_)
);

OAI21X1 _11752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2846_),
    .B(_2847_),
    .C(_2845_),
    .Y(_2848_)
);

NOR2X1 _11753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2848_),
    .B(_2840_),
    .Y(_2849_)
);

INVX1 _11754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2849_),
    .Y(\datapath_1.ALUResult [8])
);

NOR2X1 _11755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2488_),
    .B(_2494_),
    .Y(_2850_)
);

OAI21X1 _11756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2850_),
    .B(_2145_),
    .C(_2153_),
    .Y(_2851_)
);

AND2X2 _11757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2851_),
    .B(_2558_),
    .Y(_2852_)
);

NOR2X1 _11758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .B(_2852_),
    .Y(_2853_)
);

INVX1 _11759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .Y(_2854_)
);

OAI21X1 _11760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_2139_),
    .C(_2851_),
    .Y(_2855_)
);

AOI21X1 _11761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2854_),
    .B(_2855_),
    .C(_2364_),
    .Y(_2856_)
);

OR2X2 _11762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2856_),
    .B(_2337_),
    .Y(_2857_)
);

AOI21X1 _11763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2853_),
    .C(_2857_),
    .Y(_2858_)
);

AOI22X1 _11764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2364_),
    .C(_2137_),
    .D(_2341__bF$buf2),
    .Y(_2859_)
);

AOI22X1 _11765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2481__bF$buf3),
    .C(_2620_),
    .D(_2373_),
    .Y(_2860_)
);

INVX1 _11766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .Y(_2861_)
);

INVX1 _11767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2372_),
    .Y(_2862_)
);

AOI21X1 _11768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2561_),
    .B(_2363_),
    .C(_2862_),
    .Y(_2863_)
);

OAI21X1 _11769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2863_),
    .B(_2139_),
    .C(_2861_),
    .Y(_2864_)
);

AOI21X1 _11770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2864_),
    .C(_2458_),
    .Y(_2865_)
);

OAI21X1 _11771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2864_),
    .C(_2865_),
    .Y(_2866_)
);

NAND3X1 _11772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2859_),
    .B(_2860_),
    .C(_2866_),
    .Y(_2867_)
);

NOR2X1 _11773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2867_),
    .B(_2858_),
    .Y(_2868_)
);

INVX1 _11774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2868_),
    .Y(\datapath_1.ALUResult [7])
);

NOR2X1 _11775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2852_),
    .Y(_2869_)
);

OAI21X1 _11776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2851_),
    .C(_2869_),
    .Y(_2870_)
);

NAND2X1 _11777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2139_),
    .B(_2341__bF$buf1),
    .Y(_2871_)
);

OAI21X1 _11778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2344__bF$buf0),
    .C(_2871_),
    .Y(_2872_)
);

OAI22X1 _11779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2861_),
    .B(_2346_),
    .C(_2347__bF$buf1),
    .D(_2139_),
    .Y(_2873_)
);

NOR2X1 _11780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2873_),
    .B(_2872_),
    .Y(_2874_)
);

AND2X2 _11781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2863_),
    .B(_2558_),
    .Y(_2875_)
);

OAI21X1 _11782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2863_),
    .B(_2558_),
    .C(_2470__bF$buf2),
    .Y(_2876_)
);

OR2X2 _11783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2875_),
    .B(_2876_),
    .Y(_2877_)
);

NAND3X1 _11784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2874_),
    .B(_2877_),
    .C(_2870_),
    .Y(\datapath_1.ALUResult [6])
);

INVX1 _11785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2152_),
    .Y(_2878_)
);

OAI21X1 _11786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2494_),
    .B(_2488_),
    .C(_2560_),
    .Y(_2879_)
);

AOI21X1 _11787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2878_),
    .B(_2879_),
    .C(_2367_),
    .Y(_2880_)
);

OAI21X1 _11788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [4]),
    .B(_2151_),
    .C(_2879_),
    .Y(_2881_)
);

NOR2X1 _11789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2148_),
    .B(_2881_),
    .Y(_2882_)
);

NOR3X1 _11790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2880_),
    .C(_2882_),
    .Y(_2883_)
);

AOI22X1 _11791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2481__bF$buf2),
    .C(_2341__bF$buf0),
    .D(_2142_),
    .Y(_2884_)
);

OAI21X1 _11792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2148_),
    .B(_2344__bF$buf3),
    .C(_2884_),
    .Y(_2885_)
);

AOI21X1 _11793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2371_),
    .B(_2620_),
    .C(_2885_),
    .Y(_2886_)
);

INVX1 _11794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2144_),
    .Y(_2887_)
);

AOI21X1 _11795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2887_),
    .B(_2363_),
    .C(_2143_),
    .Y(_2888_)
);

AND2X2 _11796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2888_),
    .B(_2148_),
    .Y(_2889_)
);

OAI21X1 _11797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2888_),
    .B(_2148_),
    .C(_2470__bF$buf1),
    .Y(_2890_)
);

OAI21X1 _11798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2889_),
    .B(_2890_),
    .C(_2886_),
    .Y(_2891_)
);

NOR2X1 _11799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2891_),
    .B(_2883_),
    .Y(_2892_)
);

INVX1 _11800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2892_),
    .Y(\datapath_1.ALUResult [5])
);

NAND2X1 _11801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2368_),
    .B(_2850_),
    .Y(_2893_)
);

NAND3X1 _11802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462__bF$buf2),
    .B(_2879_),
    .C(_2893_),
    .Y(_2894_)
);

AOI22X1 _11803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2143_),
    .B(_2481__bF$buf1),
    .C(_2341__bF$buf3),
    .D(_2144_),
    .Y(_2895_)
);

OAI21X1 _11804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .B(_2344__bF$buf2),
    .C(_2895_),
    .Y(_2896_)
);

AOI21X1 _11805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2887_),
    .B(_2620_),
    .C(_2896_),
    .Y(_2897_)
);

AOI21X1 _11806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2368_),
    .B(_2363_),
    .C(_2458_),
    .Y(_2898_)
);

OAI21X1 _11807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2368_),
    .B(_2363_),
    .C(_2898_),
    .Y(_2899_)
);

NAND3X1 _11808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2897_),
    .B(_2899_),
    .C(_2894_),
    .Y(\datapath_1.ALUResult [4])
);

OAI21X1 _11809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2131_),
    .B(_2127_),
    .C(_2541_),
    .Y(_2900_)
);

OAI21X1 _11810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [2]),
    .B(_2120_),
    .C(_2900_),
    .Y(_2901_)
);

AND2X2 _11811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2901_),
    .B(_2124_),
    .Y(_2902_)
);

OAI21X1 _11812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2901_),
    .B(_2124_),
    .C(_2462__bF$buf1),
    .Y(_2903_)
);

OAI22X1 _11813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2124_),
    .B(_2344__bF$buf1),
    .C(_2480_),
    .D(_2123_),
    .Y(_2904_)
);

OAI22X1 _11814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .B(_2346_),
    .C(_2347__bF$buf0),
    .D(_2355_),
    .Y(_2905_)
);

NOR2X1 _11815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2905_),
    .B(_2904_),
    .Y(_2906_)
);

AOI21X1 _11816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2133_),
    .B(_2359_),
    .C(_2351_),
    .Y(_2907_)
);

AOI21X1 _11817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2124_),
    .B(_2907_),
    .C(_2458_),
    .Y(_2908_)
);

OAI21X1 _11818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2124_),
    .B(_2907_),
    .C(_2908_),
    .Y(_2909_)
);

AND2X2 _11819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2909_),
    .B(_2906_),
    .Y(_2910_)
);

OAI21X1 _11820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2903_),
    .B(_2902_),
    .C(_2910_),
    .Y(\datapath_1.ALUResult [3])
);

OAI21X1 _11821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [1]),
    .B(_2126_),
    .C(_2492_),
    .Y(_2911_)
);

OAI21X1 _11822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2911_),
    .B(_2541_),
    .C(_2462__bF$buf0),
    .Y(_2912_)
);

AOI21X1 _11823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2911_),
    .B(_2541_),
    .C(_2912_),
    .Y(_2913_)
);

AOI22X1 _11824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2353_),
    .C(_2352_),
    .D(_2341__bF$buf2),
    .Y(_2914_)
);

AOI22X1 _11825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2351_),
    .B(_2481__bF$buf0),
    .C(_2620_),
    .D(_2133_),
    .Y(_2915_)
);

AOI21X1 _11826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2353_),
    .B(_2359_),
    .C(_2458_),
    .Y(_2916_)
);

OAI21X1 _11827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2353_),
    .B(_2359_),
    .C(_2916_),
    .Y(_2917_)
);

NAND3X1 _11828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2914_),
    .B(_2915_),
    .C(_2917_),
    .Y(_2918_)
);

NOR2X1 _11829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2913_),
    .B(_2918_),
    .Y(_2919_)
);

INVX1 _11830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2919_),
    .Y(\datapath_1.ALUResult [2])
);

NOR2X1 _11831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2491_),
    .Y(_2920_)
);

AOI22X1 _11832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2920_),
    .C(_2357_),
    .D(_2341__bF$buf1),
    .Y(_2921_)
);

AOI22X1 _11833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2491_),
    .B(_2481__bF$buf3),
    .C(_2620_),
    .D(_2130_),
    .Y(_2922_)
);

NAND2X1 _11834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2922_),
    .B(_2921_),
    .Y(_2923_)
);

AOI21X1 _11835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2920_),
    .B(_2542_),
    .C(_2458_),
    .Y(_2924_)
);

OAI21X1 _11836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2920_),
    .B(_2542_),
    .C(_2924_),
    .Y(_2925_)
);

NOR2X1 _11837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInA [0]),
    .B(_2490_),
    .Y(_2926_)
);

NAND2X1 _11838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2926_),
    .B(_2920_),
    .Y(_2927_)
);

NAND2X1 _11839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2927_),
    .Y(_2928_)
);

OAI21X1 _11840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2928_),
    .B(_2337_),
    .C(_2925_),
    .Y(_2929_)
);

OR2X2 _11841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2929_),
    .B(_2923_),
    .Y(\datapath_1.ALUResult [1])
);

NOR2X1 _11842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(_2128_),
    .Y(_2930_)
);

OR2X2 _11843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2333_),
    .B(ALUControl[0]),
    .Y(_2931_)
);

OAI21X1 _11844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .B(gnd),
    .C(_2344__bF$buf0),
    .Y(_2932_)
);

OAI21X1 _11845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2926_),
    .B(_2930_),
    .C(_2932_),
    .Y(_2933_)
);

OAI21X1 _11846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .C(_2620_),
    .Y(_2934_)
);

NOR2X1 _11847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.alu_1.ALUInB [0]),
    .B(\datapath_1.alu_1.ALUInA [0]),
    .Y(_2935_)
);

AOI22X1 _11848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481__bF$buf2),
    .B(_2542_),
    .C(_2341__bF$buf0),
    .D(_2935_),
    .Y(_2936_)
);

NAND3X1 _11849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2934_),
    .B(_2933_),
    .C(_2936_),
    .Y(\datapath_1.ALUResult [0])
);

NOR3X1 _11850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2923_),
    .B(\datapath_1.ALUResult [0]),
    .C(_2929_),
    .Y(_2937_)
);

NAND2X1 _11851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2919_),
    .B(_2937_),
    .Y(_2938_)
);

NOR3X1 _11852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [4]),
    .B(\datapath_1.ALUResult [3]),
    .C(_2938_),
    .Y(_2939_)
);

NAND3X1 _11853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2849_),
    .B(_2892_),
    .C(_2939_),
    .Y(_2940_)
);

NOR2X1 _11854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [9]),
    .B(_2940_),
    .Y(_2941_)
);

NAND3X1 _11855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .B(_2941_),
    .C(_2733_),
    .Y(_2942_)
);

OR2X2 _11856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2662_),
    .Y(_2943_)
);

NAND3X1 _11857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(_2675_),
    .C(_2776_),
    .Y(_2944_)
);

NOR3X1 _11858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2942_),
    .B(\datapath_1.ALUResult [25]),
    .C(_2944_),
    .Y(_2945_)
);

NAND3X1 _11859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2868_),
    .B(_2790_),
    .C(_2816_),
    .Y(_2946_)
);

NAND2X1 _11860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2687_),
    .B(_2718_),
    .Y(_2947_)
);

NOR3X1 _11861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [10]),
    .B(\datapath_1.ALUResult [6]),
    .C(\datapath_1.ALUResult [16]),
    .Y(_2948_)
);

NAND2X1 _11862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2627_),
    .B(_2948_),
    .Y(_2949_)
);

NOR3X1 _11863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2946_),
    .B(_2949_),
    .C(_2947_),
    .Y(_2950_)
);

NOR2X1 _11864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [29]),
    .B(\datapath_1.ALUResult [15]),
    .Y(_2951_)
);

NAND3X1 _11865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2950_),
    .B(_2951_),
    .C(_2945_),
    .Y(_2952_)
);

NOR2X1 _11866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [28]),
    .B(\datapath_1.ALUResult [26]),
    .Y(_2953_)
);

NOR2X1 _11867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [22]),
    .B(\datapath_1.ALUResult [19]),
    .Y(_2954_)
);

AND2X2 _11868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2953_),
    .B(_2954_),
    .Y(_2955_)
);

NOR2X1 _11869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [27]),
    .B(\datapath_1.ALUResult [23]),
    .Y(_2956_)
);

NAND3X1 _11870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2473_),
    .B(_2955_),
    .C(_2956_),
    .Y(_2957_)
);

NOR3X1 _11871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [31]),
    .B(_2952_),
    .C(_2957_),
    .Y(ALUZero)
);

INVX1 _11872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [18]),
    .Y(_2958_)
);

NAND2X1 _11873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [13]),
    .B(RegDst),
    .Y(_2959_)
);

OAI21X1 _11874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2958_),
    .B(RegDst),
    .C(_2959_),
    .Y(\datapath_1.a3 [0])
);

INVX1 _11875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [19]),
    .Y(_2960_)
);

NAND2X1 _11876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegDst),
    .B(\datapath_1.PCJump [14]),
    .Y(_2961_)
);

OAI21X1 _11877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2960_),
    .B(RegDst),
    .C(_2961_),
    .Y(\datapath_1.a3 [1])
);

INVX1 _11878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [20]),
    .Y(_2962_)
);

NAND2X1 _11879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegDst),
    .B(\datapath_1.PCJump [15]),
    .Y(_2963_)
);

OAI21X1 _11880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2962_),
    .B(RegDst),
    .C(_2963_),
    .Y(\datapath_1.a3 [2])
);

INVX1 _11881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .Y(_2964_)
);

NAND2X1 _11882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegDst),
    .B(\datapath_1.PCJump [16]),
    .Y(_2965_)
);

OAI21X1 _11883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2964_),
    .B(RegDst),
    .C(_2965_),
    .Y(\datapath_1.a3 [3])
);

INVX1 _11884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .Y(_2966_)
);

NAND2X1 _11885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegDst),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_2967_)
);

OAI21X1 _11886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2966_),
    .B(RegDst),
    .C(_2967_),
    .Y(\datapath_1.a3 [4])
);

INVX1 _11887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3030_)
);

NAND2X1 _11888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[0]),
    .B(IorD_bF$buf7),
    .Y(_3031_)
);

OAI21X1 _11889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3030_),
    .B(IorD_bF$buf6),
    .C(_3031_),
    .Y(_1_[0])
);

INVX1 _11890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_2968_)
);

NAND2X1 _11891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[1]),
    .Y(_2969_)
);

OAI21X1 _11892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2968_),
    .B(IorD_bF$buf4),
    .C(_2969_),
    .Y(_1_[1])
);

INVX1 _11893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_2970_)
);

NAND2X1 _11894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[2]),
    .Y(_2971_)
);

OAI21X1 _11895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2970_),
    .B(IorD_bF$buf2),
    .C(_2971_),
    .Y(_1_[2])
);

INVX1 _11896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_2972_)
);

NAND2X1 _11897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[3]),
    .Y(_2973_)
);

OAI21X1 _11898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2972_),
    .B(IorD_bF$buf0),
    .C(_2973_),
    .Y(_1_[3])
);

INVX1 _11899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_2974_)
);

NAND2X1 _11900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[4]),
    .Y(_2975_)
);

OAI21X1 _11901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2974_),
    .B(IorD_bF$buf6),
    .C(_2975_),
    .Y(_1_[4])
);

INVX1 _11902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_2976_)
);

NAND2X1 _11903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[5]),
    .Y(_2977_)
);

OAI21X1 _11904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2976_),
    .B(IorD_bF$buf4),
    .C(_2977_),
    .Y(_1_[5])
);

INVX1 _11905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_2978_)
);

NAND2X1 _11906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[6]),
    .Y(_2979_)
);

OAI21X1 _11907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2978_),
    .B(IorD_bF$buf2),
    .C(_2979_),
    .Y(_1_[6])
);

INVX1 _11908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_2980_)
);

NAND2X1 _11909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[7]),
    .Y(_2981_)
);

OAI21X1 _11910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2980_),
    .B(IorD_bF$buf0),
    .C(_2981_),
    .Y(_1_[7])
);

INVX1 _11911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_2982_)
);

NAND2X1 _11912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[8]),
    .Y(_2983_)
);

OAI21X1 _11913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2982_),
    .B(IorD_bF$buf6),
    .C(_2983_),
    .Y(_1_[8])
);

INVX1 _11914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_2984_)
);

NAND2X1 _11915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[9]),
    .Y(_2985_)
);

OAI21X1 _11916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2984_),
    .B(IorD_bF$buf4),
    .C(_2985_),
    .Y(_1_[9])
);

INVX1 _11917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_2986_)
);

NAND2X1 _11918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[10]),
    .Y(_2987_)
);

OAI21X1 _11919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2986_),
    .B(IorD_bF$buf2),
    .C(_2987_),
    .Y(_1_[10])
);

INVX1 _11920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_2988_)
);

NAND2X1 _11921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[11]),
    .Y(_2989_)
);

OAI21X1 _11922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2988_),
    .B(IorD_bF$buf0),
    .C(_2989_),
    .Y(_1_[11])
);

INVX1 _11923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_2990_)
);

NAND2X1 _11924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[12]),
    .Y(_2991_)
);

OAI21X1 _11925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2990_),
    .B(IorD_bF$buf6),
    .C(_2991_),
    .Y(_1_[12])
);

INVX1 _11926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_2992_)
);

NAND2X1 _11927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[13]),
    .Y(_2993_)
);

OAI21X1 _11928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2992_),
    .B(IorD_bF$buf4),
    .C(_2993_),
    .Y(_1_[13])
);

INVX1 _11929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_2994_)
);

NAND2X1 _11930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[14]),
    .Y(_2995_)
);

OAI21X1 _11931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2994_),
    .B(IorD_bF$buf2),
    .C(_2995_),
    .Y(_1_[14])
);

INVX1 _11932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_2996_)
);

NAND2X1 _11933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[15]),
    .Y(_2997_)
);

OAI21X1 _11934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2996_),
    .B(IorD_bF$buf0),
    .C(_2997_),
    .Y(_1_[15])
);

INVX1 _11935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_2998_)
);

NAND2X1 _11936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[16]),
    .Y(_2999_)
);

OAI21X1 _11937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2998_),
    .B(IorD_bF$buf6),
    .C(_2999_),
    .Y(_1_[16])
);

INVX1 _11938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3000_)
);

NAND2X1 _11939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[17]),
    .Y(_3001_)
);

OAI21X1 _11940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3000_),
    .B(IorD_bF$buf4),
    .C(_3001_),
    .Y(_1_[17])
);

INVX1 _11941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3002_)
);

NAND2X1 _11942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[18]),
    .Y(_3003_)
);

OAI21X1 _11943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3002_),
    .B(IorD_bF$buf2),
    .C(_3003_),
    .Y(_1_[18])
);

INVX1 _11944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3004_)
);

NAND2X1 _11945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[19]),
    .Y(_3005_)
);

OAI21X1 _11946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3004_),
    .B(IorD_bF$buf0),
    .C(_3005_),
    .Y(_1_[19])
);

INVX1 _11947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3006_)
);

NAND2X1 _11948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[20]),
    .Y(_3007_)
);

OAI21X1 _11949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3006_),
    .B(IorD_bF$buf6),
    .C(_3007_),
    .Y(_1_[20])
);

INVX1 _11950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3008_)
);

NAND2X1 _11951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[21]),
    .Y(_3009_)
);

OAI21X1 _11952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3008_),
    .B(IorD_bF$buf4),
    .C(_3009_),
    .Y(_1_[21])
);

INVX1 _11953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3010_)
);

NAND2X1 _11954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[22]),
    .Y(_3011_)
);

OAI21X1 _11955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3010_),
    .B(IorD_bF$buf2),
    .C(_3011_),
    .Y(_1_[22])
);

INVX1 _11956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3012_)
);

NAND2X1 _11957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[23]),
    .Y(_3013_)
);

OAI21X1 _11958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3012_),
    .B(IorD_bF$buf0),
    .C(_3013_),
    .Y(_1_[23])
);

INVX1 _11959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3014_)
);

NAND2X1 _11960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[24]),
    .Y(_3015_)
);

OAI21X1 _11961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3014_),
    .B(IorD_bF$buf6),
    .C(_3015_),
    .Y(_1_[24])
);

INVX1 _11962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3016_)
);

NAND2X1 _11963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[25]),
    .Y(_3017_)
);

OAI21X1 _11964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3016_),
    .B(IorD_bF$buf4),
    .C(_3017_),
    .Y(_1_[25])
);

INVX1 _11965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3018_)
);

NAND2X1 _11966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[26]),
    .Y(_3019_)
);

OAI21X1 _11967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3018_),
    .B(IorD_bF$buf2),
    .C(_3019_),
    .Y(_1_[26])
);

INVX1 _11968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3020_)
);

NAND2X1 _11969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[27]),
    .Y(_3021_)
);

OAI21X1 _11970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3020_),
    .B(IorD_bF$buf0),
    .C(_3021_),
    .Y(_1_[27])
);

INVX1 _11971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [28]),
    .Y(_3022_)
);

NAND2X1 _11972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf7),
    .B(ALUOut[28]),
    .Y(_3023_)
);

OAI21X1 _11973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3022_),
    .B(IorD_bF$buf6),
    .C(_3023_),
    .Y(_1_[28])
);

INVX1 _11974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [29]),
    .Y(_3024_)
);

NAND2X1 _11975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf5),
    .B(ALUOut[29]),
    .Y(_3025_)
);

OAI21X1 _11976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3024_),
    .B(IorD_bF$buf4),
    .C(_3025_),
    .Y(_1_[29])
);

INVX1 _11977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [30]),
    .Y(_3026_)
);

NAND2X1 _11978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf3),
    .B(ALUOut[30]),
    .Y(_3027_)
);

OAI21X1 _11979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3026_),
    .B(IorD_bF$buf2),
    .C(_3027_),
    .Y(_1_[30])
);

INVX1 _11980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [31]),
    .Y(_3028_)
);

NAND2X1 _11981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IorD_bF$buf1),
    .B(ALUOut[31]),
    .Y(_3029_)
);

OAI21X1 _11982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3028_),
    .B(IorD_bF$buf0),
    .C(_3029_),
    .Y(_1_[31])
);

INVX8 _11983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .Y(_3032_)
);

NAND3X1 _11984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[0]),
    .C(_3032__bF$buf4),
    .Y(_3033_)
);

INVX8 _11985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf3),
    .Y(_3034_)
);

NAND3X1 _11986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(gnd),
    .C(_3034__bF$buf4),
    .Y(_3035_)
);

NOR2X1 _11987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf2),
    .B(PCSource_1_bF$buf2),
    .Y(_3036_)
);

AND2X2 _11988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf1),
    .B(PCSource_1_bF$buf1),
    .Y(_3037_)
);

AOI22X1 _11989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [0]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3038_)
);

NAND3X1 _11990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3033_),
    .B(_3035_),
    .C(_3038_),
    .Y(\datapath_1.mux_pcsrc.dout [0])
);

NAND3X1 _11991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[1]),
    .C(_3032__bF$buf3),
    .Y(_3039_)
);

NAND3X1 _11992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(gnd),
    .C(_3034__bF$buf3),
    .Y(_3040_)
);

AOI22X1 _11993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [1]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3041_)
);

NAND3X1 _11994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3039_),
    .B(_3040_),
    .C(_3041_),
    .Y(\datapath_1.mux_pcsrc.dout [1])
);

NAND3X1 _11995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[2]),
    .C(_3032__bF$buf2),
    .Y(_3042_)
);

NAND3X1 _11996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .B(\aluControl_1.inst [0]),
    .C(_3034__bF$buf2),
    .Y(_3043_)
);

AOI22X1 _11997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [2]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3044_)
);

NAND3X1 _11998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3042_),
    .B(_3043_),
    .C(_3044_),
    .Y(\datapath_1.mux_pcsrc.dout [2])
);

NAND3X1 _11999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[3]),
    .C(_3032__bF$buf1),
    .Y(_3045_)
);

NAND3X1 _12000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(\aluControl_1.inst [1]),
    .C(_3034__bF$buf1),
    .Y(_3046_)
);

AOI22X1 _12001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [3]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3047_)
);

NAND3X1 _12002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3045_),
    .B(_3046_),
    .C(_3047_),
    .Y(\datapath_1.mux_pcsrc.dout [3])
);

NAND3X1 _12003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[4]),
    .C(_3032__bF$buf0),
    .Y(_3048_)
);

NAND3X1 _12004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf2),
    .B(\aluControl_1.inst [2]),
    .C(_3034__bF$buf0),
    .Y(_3049_)
);

AOI22X1 _12005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [4]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3050_)
);

NAND3X1 _12006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3048_),
    .B(_3049_),
    .C(_3050_),
    .Y(\datapath_1.mux_pcsrc.dout [4])
);

NAND3X1 _12007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[5]),
    .C(_3032__bF$buf4),
    .Y(_3051_)
);

NAND3X1 _12008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf1),
    .B(\aluControl_1.inst [3]),
    .C(_3034__bF$buf4),
    .Y(_3052_)
);

AOI22X1 _12009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [5]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3053_)
);

NAND3X1 _12010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3051_),
    .B(_3052_),
    .C(_3053_),
    .Y(\datapath_1.mux_pcsrc.dout [5])
);

NAND3X1 _12011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[6]),
    .C(_3032__bF$buf3),
    .Y(_3054_)
);

NAND3X1 _12012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(\aluControl_1.inst [4]),
    .C(_3034__bF$buf3),
    .Y(_3055_)
);

AOI22X1 _12013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [6]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3056_)
);

NAND3X1 _12014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3054_),
    .B(_3055_),
    .C(_3056_),
    .Y(\datapath_1.mux_pcsrc.dout [6])
);

NAND3X1 _12015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[7]),
    .C(_3032__bF$buf2),
    .Y(_3057_)
);

NAND3X1 _12016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .B(\aluControl_1.inst [5]),
    .C(_3034__bF$buf2),
    .Y(_3058_)
);

AOI22X1 _12017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [7]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3059_)
);

NAND3X1 _12018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3057_),
    .B(_3058_),
    .C(_3059_),
    .Y(\datapath_1.mux_pcsrc.dout [7])
);

NAND3X1 _12019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[8]),
    .C(_3032__bF$buf1),
    .Y(_3060_)
);

NAND3X1 _12020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [8]),
    .C(_3034__bF$buf1),
    .Y(_3061_)
);

AOI22X1 _12021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [8]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3062_)
);

NAND3X1 _12022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3060_),
    .B(_3061_),
    .C(_3062_),
    .Y(\datapath_1.mux_pcsrc.dout [8])
);

NAND3X1 _12023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[9]),
    .C(_3032__bF$buf0),
    .Y(_3063_)
);

NAND3X1 _12024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [9]),
    .C(_3034__bF$buf0),
    .Y(_3064_)
);

AOI22X1 _12025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [9]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3065_)
);

NAND3X1 _12026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3063_),
    .B(_3064_),
    .C(_3065_),
    .Y(\datapath_1.mux_pcsrc.dout [9])
);

NAND3X1 _12027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[10]),
    .C(_3032__bF$buf4),
    .Y(_3066_)
);

NAND3X1 _12028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [10]),
    .C(_3034__bF$buf4),
    .Y(_3067_)
);

AOI22X1 _12029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [10]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3068_)
);

NAND3X1 _12030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3066_),
    .B(_3067_),
    .C(_3068_),
    .Y(\datapath_1.mux_pcsrc.dout [10])
);

NAND3X1 _12031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[11]),
    .C(_3032__bF$buf3),
    .Y(_3069_)
);

NAND3X1 _12032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [11]),
    .C(_3034__bF$buf3),
    .Y(_3070_)
);

AOI22X1 _12033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [11]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3071_)
);

NAND3X1 _12034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3069_),
    .B(_3070_),
    .C(_3071_),
    .Y(\datapath_1.mux_pcsrc.dout [11])
);

NAND3X1 _12035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[12]),
    .C(_3032__bF$buf2),
    .Y(_3072_)
);

NAND3X1 _12036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump [12]),
    .C(_3034__bF$buf2),
    .Y(_3073_)
);

AOI22X1 _12037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [12]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3074_)
);

NAND3X1 _12038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3072_),
    .B(_3073_),
    .C(_3074_),
    .Y(\datapath_1.mux_pcsrc.dout [12])
);

NAND3X1 _12039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[13]),
    .C(_3032__bF$buf1),
    .Y(_3075_)
);

NAND3X1 _12040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [13]),
    .C(_3034__bF$buf1),
    .Y(_3076_)
);

AOI22X1 _12041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [13]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3077_)
);

NAND3X1 _12042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3075_),
    .B(_3076_),
    .C(_3077_),
    .Y(\datapath_1.mux_pcsrc.dout [13])
);

NAND3X1 _12043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[14]),
    .C(_3032__bF$buf0),
    .Y(_3078_)
);

NAND3X1 _12044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [14]),
    .C(_3034__bF$buf0),
    .Y(_3079_)
);

AOI22X1 _12045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [14]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3080_)
);

NAND3X1 _12046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3078_),
    .B(_3079_),
    .C(_3080_),
    .Y(\datapath_1.mux_pcsrc.dout [14])
);

NAND3X1 _12047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[15]),
    .C(_3032__bF$buf4),
    .Y(_3081_)
);

NAND3X1 _12048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [15]),
    .C(_3034__bF$buf4),
    .Y(_3082_)
);

AOI22X1 _12049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [15]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3083_)
);

NAND3X1 _12050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3081_),
    .B(_3082_),
    .C(_3083_),
    .Y(\datapath_1.mux_pcsrc.dout [15])
);

NAND3X1 _12051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[16]),
    .C(_3032__bF$buf3),
    .Y(_3084_)
);

NAND3X1 _12052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [16]),
    .C(_3034__bF$buf3),
    .Y(_3085_)
);

AOI22X1 _12053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [16]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3086_)
);

NAND3X1 _12054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3084_),
    .B(_3085_),
    .C(_3086_),
    .Y(\datapath_1.mux_pcsrc.dout [16])
);

NAND3X1 _12055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[17]),
    .C(_3032__bF$buf2),
    .Y(_3087_)
);

NAND3X1 _12056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3034__bF$buf2),
    .Y(_3088_)
);

AOI22X1 _12057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [17]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3089_)
);

NAND3X1 _12058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3087_),
    .B(_3088_),
    .C(_3089_),
    .Y(\datapath_1.mux_pcsrc.dout [17])
);

NAND3X1 _12059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[18]),
    .C(_3032__bF$buf1),
    .Y(_3090_)
);

NAND3X1 _12060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [18]),
    .C(_3034__bF$buf1),
    .Y(_3091_)
);

AOI22X1 _12061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [18]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3092_)
);

NAND3X1 _12062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3090_),
    .B(_3091_),
    .C(_3092_),
    .Y(\datapath_1.mux_pcsrc.dout [18])
);

NAND3X1 _12063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[19]),
    .C(_3032__bF$buf0),
    .Y(_3093_)
);

NAND3X1 _12064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [19]),
    .C(_3034__bF$buf0),
    .Y(_3094_)
);

AOI22X1 _12065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [19]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3095_)
);

NAND3X1 _12066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3093_),
    .B(_3094_),
    .C(_3095_),
    .Y(\datapath_1.mux_pcsrc.dout [19])
);

NAND3X1 _12067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[20]),
    .C(_3032__bF$buf4),
    .Y(_3096_)
);

NAND3X1 _12068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [20]),
    .C(_3034__bF$buf4),
    .Y(_3097_)
);

AOI22X1 _12069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [20]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3098_)
);

NAND3X1 _12070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3096_),
    .B(_3097_),
    .C(_3098_),
    .Y(\datapath_1.mux_pcsrc.dout [20])
);

NAND3X1 _12071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[21]),
    .C(_3032__bF$buf3),
    .Y(_3099_)
);

NAND3X1 _12072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [21]),
    .C(_3034__bF$buf3),
    .Y(_3100_)
);

AOI22X1 _12073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [21]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3101_)
);

NAND3X1 _12074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3099_),
    .B(_3100_),
    .C(_3101_),
    .Y(\datapath_1.mux_pcsrc.dout [21])
);

NAND3X1 _12075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[22]),
    .C(_3032__bF$buf2),
    .Y(_3102_)
);

NAND3X1 _12076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_22_bF$buf2 ),
    .C(_3034__bF$buf2),
    .Y(_3103_)
);

AOI22X1 _12077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [22]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3104_)
);

NAND3X1 _12078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3102_),
    .B(_3103_),
    .C(_3104_),
    .Y(\datapath_1.mux_pcsrc.dout [22])
);

NAND3X1 _12079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[23]),
    .C(_3032__bF$buf1),
    .Y(_3105_)
);

NAND3X1 _12080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [23]),
    .C(_3034__bF$buf1),
    .Y(_3106_)
);

AOI22X1 _12081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [23]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3107_)
);

NAND3X1 _12082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3105_),
    .B(_3106_),
    .C(_3107_),
    .Y(\datapath_1.mux_pcsrc.dout [23])
);

NAND3X1 _12083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[24]),
    .C(_3032__bF$buf0),
    .Y(_3108_)
);

NAND3X1 _12084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [24]),
    .C(_3034__bF$buf0),
    .Y(_3109_)
);

AOI22X1 _12085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [24]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3110_)
);

NAND3X1 _12086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3108_),
    .B(_3109_),
    .C(_3110_),
    .Y(\datapath_1.mux_pcsrc.dout [24])
);

NAND3X1 _12087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[25]),
    .C(_3032__bF$buf4),
    .Y(_3111_)
);

NAND3X1 _12088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [25]),
    .C(_3034__bF$buf4),
    .Y(_3112_)
);

AOI22X1 _12089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [25]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3113_)
);

NAND3X1 _12090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3111_),
    .B(_3112_),
    .C(_3113_),
    .Y(\datapath_1.mux_pcsrc.dout [25])
);

NAND3X1 _12091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf5),
    .B(ALUOut[26]),
    .C(_3032__bF$buf3),
    .Y(_3114_)
);

NAND3X1 _12092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [26]),
    .C(_3034__bF$buf3),
    .Y(_3115_)
);

AOI22X1 _12093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [26]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3116_)
);

NAND3X1 _12094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3114_),
    .B(_3115_),
    .C(_3116_),
    .Y(\datapath_1.mux_pcsrc.dout [26])
);

NAND3X1 _12095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf4),
    .B(ALUOut[27]),
    .C(_3032__bF$buf2),
    .Y(_3117_)
);

NAND3X1 _12096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf4),
    .B(\datapath_1.PCJump_27_bF$buf4 ),
    .C(_3034__bF$buf2),
    .Y(_3118_)
);

AOI22X1 _12097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [27]),
    .B(_3036__bF$buf2),
    .C(_3037__bF$buf2),
    .D(gnd),
    .Y(_3119_)
);

NAND3X1 _12098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3117_),
    .B(_3118_),
    .C(_3119_),
    .Y(\datapath_1.mux_pcsrc.dout [27])
);

NAND3X1 _12099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf3),
    .B(ALUOut[28]),
    .C(_3032__bF$buf1),
    .Y(_3120_)
);

NAND3X1 _12100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf3),
    .B(\datapath_1.PCJump [28]),
    .C(_3034__bF$buf1),
    .Y(_3121_)
);

AOI22X1 _12101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [28]),
    .B(_3036__bF$buf1),
    .C(_3037__bF$buf1),
    .D(gnd),
    .Y(_3122_)
);

NAND3X1 _12102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3120_),
    .B(_3121_),
    .C(_3122_),
    .Y(\datapath_1.mux_pcsrc.dout [28])
);

NAND3X1 _12103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf2),
    .B(ALUOut[29]),
    .C(_3032__bF$buf0),
    .Y(_3123_)
);

NAND3X1 _12104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf2),
    .B(\datapath_1.PCJump [29]),
    .C(_3034__bF$buf0),
    .Y(_3124_)
);

AOI22X1 _12105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [29]),
    .B(_3036__bF$buf0),
    .C(_3037__bF$buf0),
    .D(gnd),
    .Y(_3125_)
);

NAND3X1 _12106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3123_),
    .B(_3124_),
    .C(_3125_),
    .Y(\datapath_1.mux_pcsrc.dout [29])
);

NAND3X1 _12107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf1),
    .B(ALUOut[30]),
    .C(_3032__bF$buf4),
    .Y(_3126_)
);

NAND3X1 _12108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf1),
    .B(\datapath_1.PCJump [30]),
    .C(_3034__bF$buf4),
    .Y(_3127_)
);

AOI22X1 _12109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [30]),
    .B(_3036__bF$buf4),
    .C(_3037__bF$buf4),
    .D(gnd),
    .Y(_3128_)
);

NAND3X1 _12110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3126_),
    .B(_3127_),
    .C(_3128_),
    .Y(\datapath_1.mux_pcsrc.dout [30])
);

NAND3X1 _12111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOp_0_bF$buf0),
    .B(ALUOut[31]),
    .C(_3032__bF$buf3),
    .Y(_3129_)
);

NAND3X1 _12112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCSource_1_bF$buf0),
    .B(\datapath_1.PCJump [31]),
    .C(_3034__bF$buf3),
    .Y(_3130_)
);

AOI22X1 _12113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [31]),
    .B(_3036__bF$buf3),
    .C(_3037__bF$buf3),
    .D(gnd),
    .Y(_3131_)
);

NAND3X1 _12114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3129_),
    .B(_3130_),
    .C(_3131_),
    .Y(\datapath_1.mux_pcsrc.dout [31])
);

INVX1 _12115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3194_)
);

NAND2X1 _12116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [0]),
    .B(ALUSrcA_bF$buf7),
    .Y(_3195_)
);

OAI21X1 _12117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3194_),
    .B(ALUSrcA_bF$buf6),
    .C(_3195_),
    .Y(\datapath_1.alu_1.ALUInA [0])
);

INVX1 _12118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_3132_)
);

NAND2X1 _12119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [1]),
    .Y(_3133_)
);

OAI21X1 _12120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3132_),
    .B(ALUSrcA_bF$buf4),
    .C(_3133_),
    .Y(\datapath_1.alu_1.ALUInA [1])
);

INVX1 _12121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_3134_)
);

NAND2X1 _12122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [2]),
    .Y(_3135_)
);

OAI21X1 _12123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3134_),
    .B(ALUSrcA_bF$buf2),
    .C(_3135_),
    .Y(\datapath_1.alu_1.ALUInA [2])
);

INVX1 _12124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_3136_)
);

NAND2X1 _12125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [3]),
    .Y(_3137_)
);

OAI21X1 _12126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3136_),
    .B(ALUSrcA_bF$buf0),
    .C(_3137_),
    .Y(\datapath_1.alu_1.ALUInA [3])
);

INVX1 _12127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_3138_)
);

NAND2X1 _12128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [4]),
    .Y(_3139_)
);

OAI21X1 _12129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3138_),
    .B(ALUSrcA_bF$buf6),
    .C(_3139_),
    .Y(\datapath_1.alu_1.ALUInA [4])
);

INVX1 _12130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_3140_)
);

NAND2X1 _12131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [5]),
    .Y(_3141_)
);

OAI21X1 _12132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3140_),
    .B(ALUSrcA_bF$buf4),
    .C(_3141_),
    .Y(\datapath_1.alu_1.ALUInA [5])
);

INVX1 _12133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_3142_)
);

NAND2X1 _12134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [6]),
    .Y(_3143_)
);

OAI21X1 _12135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3142_),
    .B(ALUSrcA_bF$buf2),
    .C(_3143_),
    .Y(\datapath_1.alu_1.ALUInA [6])
);

INVX1 _12136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_3144_)
);

NAND2X1 _12137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [7]),
    .Y(_3145_)
);

OAI21X1 _12138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3144_),
    .B(ALUSrcA_bF$buf0),
    .C(_3145_),
    .Y(\datapath_1.alu_1.ALUInA [7])
);

INVX1 _12139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_3146_)
);

NAND2X1 _12140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [8]),
    .Y(_3147_)
);

OAI21X1 _12141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146_),
    .B(ALUSrcA_bF$buf6),
    .C(_3147_),
    .Y(\datapath_1.alu_1.ALUInA [8])
);

INVX1 _12142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_3148_)
);

NAND2X1 _12143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [9]),
    .Y(_3149_)
);

OAI21X1 _12144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3148_),
    .B(ALUSrcA_bF$buf4),
    .C(_3149_),
    .Y(\datapath_1.alu_1.ALUInA [9])
);

INVX1 _12145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_3150_)
);

NAND2X1 _12146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [10]),
    .Y(_3151_)
);

OAI21X1 _12147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3150_),
    .B(ALUSrcA_bF$buf2),
    .C(_3151_),
    .Y(\datapath_1.alu_1.ALUInA [10])
);

INVX1 _12148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_3152_)
);

NAND2X1 _12149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [11]),
    .Y(_3153_)
);

OAI21X1 _12150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3152_),
    .B(ALUSrcA_bF$buf0),
    .C(_3153_),
    .Y(\datapath_1.alu_1.ALUInA [11])
);

INVX1 _12151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_3154_)
);

NAND2X1 _12152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [12]),
    .Y(_3155_)
);

OAI21X1 _12153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3154_),
    .B(ALUSrcA_bF$buf6),
    .C(_3155_),
    .Y(\datapath_1.alu_1.ALUInA [12])
);

INVX1 _12154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_3156_)
);

NAND2X1 _12155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [13]),
    .Y(_3157_)
);

OAI21X1 _12156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3156_),
    .B(ALUSrcA_bF$buf4),
    .C(_3157_),
    .Y(\datapath_1.alu_1.ALUInA [13])
);

INVX1 _12157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_3158_)
);

NAND2X1 _12158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [14]),
    .Y(_3159_)
);

OAI21X1 _12159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3158_),
    .B(ALUSrcA_bF$buf2),
    .C(_3159_),
    .Y(\datapath_1.alu_1.ALUInA [14])
);

INVX1 _12160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_3160_)
);

NAND2X1 _12161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [15]),
    .Y(_3161_)
);

OAI21X1 _12162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3160_),
    .B(ALUSrcA_bF$buf0),
    .C(_3161_),
    .Y(\datapath_1.alu_1.ALUInA [15])
);

INVX1 _12163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_3162_)
);

NAND2X1 _12164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [16]),
    .Y(_3163_)
);

OAI21X1 _12165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3162_),
    .B(ALUSrcA_bF$buf6),
    .C(_3163_),
    .Y(\datapath_1.alu_1.ALUInA [16])
);

INVX1 _12166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3164_)
);

NAND2X1 _12167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [17]),
    .Y(_3165_)
);

OAI21X1 _12168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3164_),
    .B(ALUSrcA_bF$buf4),
    .C(_3165_),
    .Y(\datapath_1.alu_1.ALUInA [17])
);

INVX1 _12169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3166_)
);

NAND2X1 _12170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [18]),
    .Y(_3167_)
);

OAI21X1 _12171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3166_),
    .B(ALUSrcA_bF$buf2),
    .C(_3167_),
    .Y(\datapath_1.alu_1.ALUInA [18])
);

INVX1 _12172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3168_)
);

NAND2X1 _12173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [19]),
    .Y(_3169_)
);

OAI21X1 _12174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3168_),
    .B(ALUSrcA_bF$buf0),
    .C(_3169_),
    .Y(\datapath_1.alu_1.ALUInA [19])
);

INVX1 _12175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3170_)
);

NAND2X1 _12176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [20]),
    .Y(_3171_)
);

OAI21X1 _12177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3170_),
    .B(ALUSrcA_bF$buf6),
    .C(_3171_),
    .Y(\datapath_1.alu_1.ALUInA [20])
);

INVX1 _12178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3172_)
);

NAND2X1 _12179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [21]),
    .Y(_3173_)
);

OAI21X1 _12180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3172_),
    .B(ALUSrcA_bF$buf4),
    .C(_3173_),
    .Y(\datapath_1.alu_1.ALUInA [21])
);

INVX1 _12181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3174_)
);

NAND2X1 _12182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [22]),
    .Y(_3175_)
);

OAI21X1 _12183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3174_),
    .B(ALUSrcA_bF$buf2),
    .C(_3175_),
    .Y(\datapath_1.alu_1.ALUInA [22])
);

INVX1 _12184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3176_)
);

NAND2X1 _12185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [23]),
    .Y(_3177_)
);

OAI21X1 _12186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3176_),
    .B(ALUSrcA_bF$buf0),
    .C(_3177_),
    .Y(\datapath_1.alu_1.ALUInA [23])
);

INVX1 _12187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3178_)
);

NAND2X1 _12188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [24]),
    .Y(_3179_)
);

OAI21X1 _12189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3178_),
    .B(ALUSrcA_bF$buf6),
    .C(_3179_),
    .Y(\datapath_1.alu_1.ALUInA [24])
);

INVX1 _12190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3180_)
);

NAND2X1 _12191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [25]),
    .Y(_3181_)
);

OAI21X1 _12192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3180_),
    .B(ALUSrcA_bF$buf4),
    .C(_3181_),
    .Y(\datapath_1.alu_1.ALUInA [25])
);

INVX1 _12193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3182_)
);

NAND2X1 _12194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [26]),
    .Y(_3183_)
);

OAI21X1 _12195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3182_),
    .B(ALUSrcA_bF$buf2),
    .C(_3183_),
    .Y(\datapath_1.alu_1.ALUInA [26])
);

INVX1 _12196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3184_)
);

NAND2X1 _12197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [27]),
    .Y(_3185_)
);

OAI21X1 _12198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3184_),
    .B(ALUSrcA_bF$buf0),
    .C(_3185_),
    .Y(\datapath_1.alu_1.ALUInA [27])
);

INVX1 _12199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [28]),
    .Y(_3186_)
);

NAND2X1 _12200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf7),
    .B(\datapath_1.a [28]),
    .Y(_3187_)
);

OAI21X1 _12201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3186_),
    .B(ALUSrcA_bF$buf6),
    .C(_3187_),
    .Y(\datapath_1.alu_1.ALUInA [28])
);

INVX1 _12202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [29]),
    .Y(_3188_)
);

NAND2X1 _12203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf5),
    .B(\datapath_1.a [29]),
    .Y(_3189_)
);

OAI21X1 _12204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3188_),
    .B(ALUSrcA_bF$buf4),
    .C(_3189_),
    .Y(\datapath_1.alu_1.ALUInA [29])
);

INVX1 _12205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [30]),
    .Y(_3190_)
);

NAND2X1 _12206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf3),
    .B(\datapath_1.a [30]),
    .Y(_3191_)
);

OAI21X1 _12207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3190_),
    .B(ALUSrcA_bF$buf2),
    .C(_3191_),
    .Y(\datapath_1.alu_1.ALUInA [30])
);

INVX1 _12208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [31]),
    .Y(_3192_)
);

NAND2X1 _12209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcA_bF$buf1),
    .B(\datapath_1.a [31]),
    .Y(_3193_)
);

OAI21X1 _12210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3192_),
    .B(ALUSrcA_bF$buf0),
    .C(_3193_),
    .Y(\datapath_1.alu_1.ALUInA [31])
);

INVX8 _12211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .Y(_3196_)
);

NAND3X1 _12212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3197_)
);

INVX8 _12213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .Y(_3198_)
);

NAND3X1 _12214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [0]),
    .C(_3198__bF$buf4),
    .Y(_3199_)
);

NOR2X1 _12215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(ALUSrcB_1_bF$buf2),
    .Y(_3200_)
);

AND2X2 _12216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(ALUSrcB_1_bF$buf1),
    .Y(_3201_)
);

AOI22X1 _12217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[0]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(gnd),
    .Y(_3202_)
);

NAND3X1 _12218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3197_),
    .B(_3199_),
    .C(_3202_),
    .Y(\datapath_1.alu_1.ALUInB [0])
);

NAND3X1 _12219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3203_)
);

NAND3X1 _12220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\aluControl_1.inst [1]),
    .C(_3198__bF$buf3),
    .Y(_3204_)
);

AOI22X1 _12221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[1]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(gnd),
    .Y(_3205_)
);

NAND3X1 _12222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3203_),
    .B(_3204_),
    .C(_3205_),
    .Y(\datapath_1.alu_1.ALUInB [1])
);

NAND3X1 _12223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(vdd),
    .C(_3196__bF$buf2),
    .Y(_3206_)
);

NAND3X1 _12224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .B(\aluControl_1.inst [2]),
    .C(_3198__bF$buf2),
    .Y(_3207_)
);

AOI22X1 _12225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[2]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf2),
    .D(\aluControl_1.inst [0]),
    .Y(_3208_)
);

NAND3X1 _12226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3206_),
    .B(_3207_),
    .C(_3208_),
    .Y(\datapath_1.alu_1.ALUInB [2])
);

NAND3X1 _12227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3209_)
);

NAND3X1 _12228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\aluControl_1.inst [3]),
    .C(_3198__bF$buf1),
    .Y(_3210_)
);

AOI22X1 _12229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[3]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf1),
    .D(\aluControl_1.inst [1]),
    .Y(_3211_)
);

NAND3X1 _12230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3209_),
    .B(_3210_),
    .C(_3211_),
    .Y(\datapath_1.alu_1.ALUInB [3])
);

NAND3X1 _12231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3212_)
);

NAND3X1 _12232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf2),
    .B(\aluControl_1.inst [4]),
    .C(_3198__bF$buf0),
    .Y(_3213_)
);

AOI22X1 _12233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[4]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf0),
    .D(\aluControl_1.inst [2]),
    .Y(_3214_)
);

NAND3X1 _12234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3212_),
    .B(_3213_),
    .C(_3214_),
    .Y(\datapath_1.alu_1.ALUInB [4])
);

NAND3X1 _12235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3215_)
);

NAND3X1 _12236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf1),
    .B(\aluControl_1.inst [5]),
    .C(_3198__bF$buf4),
    .Y(_3216_)
);

AOI22X1 _12237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[5]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(\aluControl_1.inst [3]),
    .Y(_3217_)
);

NAND3X1 _12238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3215_),
    .B(_3216_),
    .C(_3217_),
    .Y(\datapath_1.alu_1.ALUInB [5])
);

NAND3X1 _12239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3218_)
);

NAND3X1 _12240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [8]),
    .C(_3198__bF$buf3),
    .Y(_3219_)
);

AOI22X1 _12241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[6]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(\aluControl_1.inst [4]),
    .Y(_3220_)
);

NAND3X1 _12242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3218_),
    .B(_3219_),
    .C(_3220_),
    .Y(\datapath_1.alu_1.ALUInB [6])
);

NAND3X1 _12243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3221_)
);

NAND3X1 _12244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [9]),
    .C(_3198__bF$buf2),
    .Y(_3222_)
);

AOI22X1 _12245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[7]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf2),
    .D(\aluControl_1.inst [5]),
    .Y(_3223_)
);

NAND3X1 _12246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3221_),
    .B(_3222_),
    .C(_3223_),
    .Y(\datapath_1.alu_1.ALUInB [7])
);

NAND3X1 _12247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3224_)
);

NAND3X1 _12248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump [10]),
    .C(_3198__bF$buf1),
    .Y(_3225_)
);

AOI22X1 _12249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[8]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [8]),
    .Y(_3226_)
);

NAND3X1 _12250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3224_),
    .B(_3225_),
    .C(_3226_),
    .Y(\datapath_1.alu_1.ALUInB [8])
);

NAND3X1 _12251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3227_)
);

NAND3X1 _12252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump [11]),
    .C(_3198__bF$buf0),
    .Y(_3228_)
);

AOI22X1 _12253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[9]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump [9]),
    .Y(_3229_)
);

NAND3X1 _12254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3227_),
    .B(_3228_),
    .C(_3229_),
    .Y(\datapath_1.alu_1.ALUInB [9])
);

NAND3X1 _12255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3230_)
);

NAND3X1 _12256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump [12]),
    .C(_3198__bF$buf4),
    .Y(_3231_)
);

AOI22X1 _12257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[10]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump [10]),
    .Y(_3232_)
);

NAND3X1 _12258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3231_),
    .C(_3232_),
    .Y(\datapath_1.alu_1.ALUInB [10])
);

NAND3X1 _12259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3233_)
);

NAND3X1 _12260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump [13]),
    .C(_3198__bF$buf3),
    .Y(_3234_)
);

AOI22X1 _12261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[11]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump [11]),
    .Y(_3235_)
);

NAND3X1 _12262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3233_),
    .B(_3234_),
    .C(_3235_),
    .Y(\datapath_1.alu_1.ALUInB [11])
);

NAND3X1 _12263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3236_)
);

NAND3X1 _12264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump [14]),
    .C(_3198__bF$buf2),
    .Y(_3237_)
);

AOI22X1 _12265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[12]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump [12]),
    .Y(_3238_)
);

NAND3X1 _12266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3236_),
    .B(_3237_),
    .C(_3238_),
    .Y(\datapath_1.alu_1.ALUInB [12])
);

NAND3X1 _12267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3239_)
);

NAND3X1 _12268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump [15]),
    .C(_3198__bF$buf1),
    .Y(_3240_)
);

AOI22X1 _12269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[13]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump [13]),
    .Y(_3241_)
);

NAND3X1 _12270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3239_),
    .B(_3240_),
    .C(_3241_),
    .Y(\datapath_1.alu_1.ALUInB [13])
);

NAND3X1 _12271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3242_)
);

NAND3X1 _12272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump [16]),
    .C(_3198__bF$buf0),
    .Y(_3243_)
);

AOI22X1 _12273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[14]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump [14]),
    .Y(_3244_)
);

NAND3X1 _12274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3242_),
    .B(_3243_),
    .C(_3244_),
    .Y(\datapath_1.alu_1.ALUInB [14])
);

NAND3X1 _12275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3245_)
);

NAND3X1 _12276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf4),
    .Y(_3246_)
);

AOI22X1 _12277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[15]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump [15]),
    .Y(_3247_)
);

NAND3X1 _12278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3245_),
    .B(_3246_),
    .C(_3247_),
    .Y(\datapath_1.alu_1.ALUInB [15])
);

NAND3X1 _12279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3248_)
);

NAND3X1 _12280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3198__bF$buf3),
    .Y(_3249_)
);

AOI22X1 _12281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[16]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump [16]),
    .Y(_3250_)
);

NAND3X1 _12282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3248_),
    .B(_3249_),
    .C(_3250_),
    .Y(\datapath_1.alu_1.ALUInB [16])
);

NAND3X1 _12283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3251_)
);

NAND3X1 _12284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3198__bF$buf2),
    .Y(_3252_)
);

AOI22X1 _12285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[17]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3253_)
);

NAND3X1 _12286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3251_),
    .B(_3252_),
    .C(_3253_),
    .Y(\datapath_1.alu_1.ALUInB [17])
);

NAND3X1 _12287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3254_)
);

NAND3X1 _12288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf1),
    .Y(_3255_)
);

AOI22X1 _12289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[18]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3256_)
);

NAND3X1 _12290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3254_),
    .B(_3255_),
    .C(_3256_),
    .Y(\datapath_1.alu_1.ALUInB [18])
);

NAND3X1 _12291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3257_)
);

NAND3X1 _12292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3198__bF$buf0),
    .Y(_3258_)
);

AOI22X1 _12293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[19]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3259_)
);

NAND3X1 _12294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3257_),
    .B(_3258_),
    .C(_3259_),
    .Y(\datapath_1.alu_1.ALUInB [19])
);

NAND3X1 _12295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3260_)
);

NAND3X1 _12296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3198__bF$buf4),
    .Y(_3261_)
);

AOI22X1 _12297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[20]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3262_)
);

NAND3X1 _12298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3260_),
    .B(_3261_),
    .C(_3262_),
    .Y(\datapath_1.alu_1.ALUInB [20])
);

NAND3X1 _12299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3263_)
);

NAND3X1 _12300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf3),
    .Y(_3264_)
);

AOI22X1 _12301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[21]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3265_)
);

NAND3X1 _12302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3263_),
    .B(_3264_),
    .C(_3265_),
    .Y(\datapath_1.alu_1.ALUInB [21])
);

NAND3X1 _12303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3266_)
);

NAND3X1 _12304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3198__bF$buf2),
    .Y(_3267_)
);

AOI22X1 _12305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[22]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3268_)
);

NAND3X1 _12306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3266_),
    .B(_3267_),
    .C(_3268_),
    .Y(\datapath_1.alu_1.ALUInB [22])
);

NAND3X1 _12307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3269_)
);

NAND3X1 _12308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf1),
    .Y(_3270_)
);

AOI22X1 _12309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[23]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3271_)
);

NAND3X1 _12310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3269_),
    .B(_3270_),
    .C(_3271_),
    .Y(\datapath_1.alu_1.ALUInB [23])
);

NAND3X1 _12311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3272_)
);

NAND3X1 _12312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3198__bF$buf0),
    .Y(_3273_)
);

AOI22X1 _12313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[24]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3274_)
);

NAND3X1 _12314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3272_),
    .B(_3273_),
    .C(_3274_),
    .Y(\datapath_1.alu_1.ALUInB [24])
);

NAND3X1 _12315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3275_)
);

NAND3X1 _12316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3198__bF$buf4),
    .Y(_3276_)
);

AOI22X1 _12317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[25]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3277_)
);

NAND3X1 _12318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3275_),
    .B(_3276_),
    .C(_3277_),
    .Y(\datapath_1.alu_1.ALUInB [25])
);

NAND3X1 _12319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3278_)
);

NAND3X1 _12320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf3),
    .Y(_3279_)
);

AOI22X1 _12321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[26]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3280_)
);

NAND3X1 _12322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3278_),
    .B(_3279_),
    .C(_3280_),
    .Y(\datapath_1.alu_1.ALUInB [26])
);

NAND3X1 _12323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf4),
    .B(gnd),
    .C(_3196__bF$buf2),
    .Y(_3281_)
);

NAND3X1 _12324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf4),
    .B(\datapath_1.PCJump_17_bF$buf0 ),
    .C(_3198__bF$buf2),
    .Y(_3282_)
);

AOI22X1 _12325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[27]),
    .B(_3200__bF$buf2),
    .C(_3201__bF$buf2),
    .D(\datapath_1.PCJump_17_bF$buf4 ),
    .Y(_3283_)
);

NAND3X1 _12326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3281_),
    .B(_3282_),
    .C(_3283_),
    .Y(\datapath_1.alu_1.ALUInB [27])
);

NAND3X1 _12327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf3),
    .B(gnd),
    .C(_3196__bF$buf1),
    .Y(_3284_)
);

NAND3X1 _12328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf3),
    .B(\datapath_1.PCJump_17_bF$buf3 ),
    .C(_3198__bF$buf1),
    .Y(_3285_)
);

AOI22X1 _12329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[28]),
    .B(_3200__bF$buf1),
    .C(_3201__bF$buf1),
    .D(\datapath_1.PCJump_17_bF$buf2 ),
    .Y(_3286_)
);

NAND3X1 _12330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3284_),
    .B(_3285_),
    .C(_3286_),
    .Y(\datapath_1.alu_1.ALUInB [28])
);

NAND3X1 _12331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf2),
    .B(gnd),
    .C(_3196__bF$buf0),
    .Y(_3287_)
);

NAND3X1 _12332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf2),
    .B(\datapath_1.PCJump_17_bF$buf1 ),
    .C(_3198__bF$buf0),
    .Y(_3288_)
);

AOI22X1 _12333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[29]),
    .B(_3200__bF$buf0),
    .C(_3201__bF$buf0),
    .D(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3289_)
);

NAND3X1 _12334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3287_),
    .B(_3288_),
    .C(_3289_),
    .Y(\datapath_1.alu_1.ALUInB [29])
);

NAND3X1 _12335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf1),
    .B(gnd),
    .C(_3196__bF$buf4),
    .Y(_3290_)
);

NAND3X1 _12336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf1),
    .B(\datapath_1.PCJump_17_bF$buf4 ),
    .C(_3198__bF$buf4),
    .Y(_3291_)
);

AOI22X1 _12337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[30]),
    .B(_3200__bF$buf4),
    .C(_3201__bF$buf4),
    .D(\datapath_1.PCJump_17_bF$buf3 ),
    .Y(_3292_)
);

NAND3X1 _12338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3290_),
    .B(_3291_),
    .C(_3292_),
    .Y(\datapath_1.alu_1.ALUInB [30])
);

NAND3X1 _12339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_0_bF$buf0),
    .B(gnd),
    .C(_3196__bF$buf3),
    .Y(_3293_)
);

NAND3X1 _12340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUSrcB_1_bF$buf0),
    .B(\datapath_1.PCJump_17_bF$buf2 ),
    .C(_3198__bF$buf3),
    .Y(_3294_)
);

AOI22X1 _12341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[31]),
    .B(_3200__bF$buf3),
    .C(_3201__bF$buf3),
    .D(\datapath_1.PCJump_17_bF$buf1 ),
    .Y(_3295_)
);

NAND3X1 _12342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3293_),
    .B(_3294_),
    .C(_3295_),
    .Y(\datapath_1.alu_1.ALUInB [31])
);

INVX1 _12343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[0]),
    .Y(_3358_)
);

NAND2X1 _12344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [0]),
    .B(MemToReg_bF$buf7),
    .Y(_3359_)
);

OAI21X1 _12345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3358_),
    .B(MemToReg_bF$buf6),
    .C(_3359_),
    .Y(\datapath_1.mux_wd3.dout [0])
);

INVX1 _12346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[1]),
    .Y(_3296_)
);

NAND2X1 _12347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [1]),
    .Y(_3297_)
);

OAI21X1 _12348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3296_),
    .B(MemToReg_bF$buf4),
    .C(_3297_),
    .Y(\datapath_1.mux_wd3.dout [1])
);

INVX1 _12349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[2]),
    .Y(_3298_)
);

NAND2X1 _12350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [2]),
    .Y(_3299_)
);

OAI21X1 _12351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3298_),
    .B(MemToReg_bF$buf2),
    .C(_3299_),
    .Y(\datapath_1.mux_wd3.dout [2])
);

INVX1 _12352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[3]),
    .Y(_3300_)
);

NAND2X1 _12353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [3]),
    .Y(_3301_)
);

OAI21X1 _12354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3300_),
    .B(MemToReg_bF$buf0),
    .C(_3301_),
    .Y(\datapath_1.mux_wd3.dout [3])
);

INVX1 _12355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[4]),
    .Y(_3302_)
);

NAND2X1 _12356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [4]),
    .Y(_3303_)
);

OAI21X1 _12357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3302_),
    .B(MemToReg_bF$buf6),
    .C(_3303_),
    .Y(\datapath_1.mux_wd3.dout [4])
);

INVX1 _12358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[5]),
    .Y(_3304_)
);

NAND2X1 _12359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [5]),
    .Y(_3305_)
);

OAI21X1 _12360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3304_),
    .B(MemToReg_bF$buf4),
    .C(_3305_),
    .Y(\datapath_1.mux_wd3.dout [5])
);

INVX1 _12361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[6]),
    .Y(_3306_)
);

NAND2X1 _12362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [6]),
    .Y(_3307_)
);

OAI21X1 _12363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3306_),
    .B(MemToReg_bF$buf2),
    .C(_3307_),
    .Y(\datapath_1.mux_wd3.dout [6])
);

INVX1 _12364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[7]),
    .Y(_3308_)
);

NAND2X1 _12365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [7]),
    .Y(_3309_)
);

OAI21X1 _12366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3308_),
    .B(MemToReg_bF$buf0),
    .C(_3309_),
    .Y(\datapath_1.mux_wd3.dout [7])
);

INVX1 _12367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[8]),
    .Y(_3310_)
);

NAND2X1 _12368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [8]),
    .Y(_3311_)
);

OAI21X1 _12369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3310_),
    .B(MemToReg_bF$buf6),
    .C(_3311_),
    .Y(\datapath_1.mux_wd3.dout [8])
);

INVX1 _12370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[9]),
    .Y(_3312_)
);

NAND2X1 _12371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [9]),
    .Y(_3313_)
);

OAI21X1 _12372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3312_),
    .B(MemToReg_bF$buf4),
    .C(_3313_),
    .Y(\datapath_1.mux_wd3.dout [9])
);

INVX1 _12373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[10]),
    .Y(_3314_)
);

NAND2X1 _12374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [10]),
    .Y(_3315_)
);

OAI21X1 _12375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3314_),
    .B(MemToReg_bF$buf2),
    .C(_3315_),
    .Y(\datapath_1.mux_wd3.dout [10])
);

INVX1 _12376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[11]),
    .Y(_3316_)
);

NAND2X1 _12377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [11]),
    .Y(_3317_)
);

OAI21X1 _12378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3316_),
    .B(MemToReg_bF$buf0),
    .C(_3317_),
    .Y(\datapath_1.mux_wd3.dout [11])
);

INVX1 _12379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[12]),
    .Y(_3318_)
);

NAND2X1 _12380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [12]),
    .Y(_3319_)
);

OAI21X1 _12381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3318_),
    .B(MemToReg_bF$buf6),
    .C(_3319_),
    .Y(\datapath_1.mux_wd3.dout [12])
);

INVX1 _12382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[13]),
    .Y(_3320_)
);

NAND2X1 _12383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [13]),
    .Y(_3321_)
);

OAI21X1 _12384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3320_),
    .B(MemToReg_bF$buf4),
    .C(_3321_),
    .Y(\datapath_1.mux_wd3.dout [13])
);

INVX1 _12385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[14]),
    .Y(_3322_)
);

NAND2X1 _12386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [14]),
    .Y(_3323_)
);

OAI21X1 _12387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3322_),
    .B(MemToReg_bF$buf2),
    .C(_3323_),
    .Y(\datapath_1.mux_wd3.dout [14])
);

INVX1 _12388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[15]),
    .Y(_3324_)
);

NAND2X1 _12389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [15]),
    .Y(_3325_)
);

OAI21X1 _12390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3324_),
    .B(MemToReg_bF$buf0),
    .C(_3325_),
    .Y(\datapath_1.mux_wd3.dout [15])
);

INVX1 _12391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[16]),
    .Y(_3326_)
);

NAND2X1 _12392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [16]),
    .Y(_3327_)
);

OAI21X1 _12393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3326_),
    .B(MemToReg_bF$buf6),
    .C(_3327_),
    .Y(\datapath_1.mux_wd3.dout [16])
);

INVX1 _12394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[17]),
    .Y(_3328_)
);

NAND2X1 _12395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [17]),
    .Y(_3329_)
);

OAI21X1 _12396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3328_),
    .B(MemToReg_bF$buf4),
    .C(_3329_),
    .Y(\datapath_1.mux_wd3.dout [17])
);

INVX1 _12397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[18]),
    .Y(_3330_)
);

NAND2X1 _12398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [18]),
    .Y(_3331_)
);

OAI21X1 _12399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3330_),
    .B(MemToReg_bF$buf2),
    .C(_3331_),
    .Y(\datapath_1.mux_wd3.dout [18])
);

INVX1 _12400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[19]),
    .Y(_3332_)
);

NAND2X1 _12401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [19]),
    .Y(_3333_)
);

OAI21X1 _12402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3332_),
    .B(MemToReg_bF$buf0),
    .C(_3333_),
    .Y(\datapath_1.mux_wd3.dout [19])
);

INVX1 _12403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[20]),
    .Y(_3334_)
);

NAND2X1 _12404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [20]),
    .Y(_3335_)
);

OAI21X1 _12405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3334_),
    .B(MemToReg_bF$buf6),
    .C(_3335_),
    .Y(\datapath_1.mux_wd3.dout [20])
);

INVX1 _12406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[21]),
    .Y(_3336_)
);

NAND2X1 _12407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [21]),
    .Y(_3337_)
);

OAI21X1 _12408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3336_),
    .B(MemToReg_bF$buf4),
    .C(_3337_),
    .Y(\datapath_1.mux_wd3.dout [21])
);

INVX1 _12409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[22]),
    .Y(_3338_)
);

NAND2X1 _12410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [22]),
    .Y(_3339_)
);

OAI21X1 _12411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3338_),
    .B(MemToReg_bF$buf2),
    .C(_3339_),
    .Y(\datapath_1.mux_wd3.dout [22])
);

INVX1 _12412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[23]),
    .Y(_3340_)
);

NAND2X1 _12413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [23]),
    .Y(_3341_)
);

OAI21X1 _12414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3340_),
    .B(MemToReg_bF$buf0),
    .C(_3341_),
    .Y(\datapath_1.mux_wd3.dout [23])
);

INVX1 _12415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[24]),
    .Y(_3342_)
);

NAND2X1 _12416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [24]),
    .Y(_3343_)
);

OAI21X1 _12417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3342_),
    .B(MemToReg_bF$buf6),
    .C(_3343_),
    .Y(\datapath_1.mux_wd3.dout [24])
);

INVX1 _12418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[25]),
    .Y(_3344_)
);

NAND2X1 _12419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [25]),
    .Y(_3345_)
);

OAI21X1 _12420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3344_),
    .B(MemToReg_bF$buf4),
    .C(_3345_),
    .Y(\datapath_1.mux_wd3.dout [25])
);

INVX1 _12421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[26]),
    .Y(_3346_)
);

NAND2X1 _12422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [26]),
    .Y(_3347_)
);

OAI21X1 _12423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3346_),
    .B(MemToReg_bF$buf2),
    .C(_3347_),
    .Y(\datapath_1.mux_wd3.dout [26])
);

INVX1 _12424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[27]),
    .Y(_3348_)
);

NAND2X1 _12425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [27]),
    .Y(_3349_)
);

OAI21X1 _12426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3348_),
    .B(MemToReg_bF$buf0),
    .C(_3349_),
    .Y(\datapath_1.mux_wd3.dout [27])
);

INVX1 _12427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[28]),
    .Y(_3350_)
);

NAND2X1 _12428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf7),
    .B(\datapath_1.Data [28]),
    .Y(_3351_)
);

OAI21X1 _12429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3350_),
    .B(MemToReg_bF$buf6),
    .C(_3351_),
    .Y(\datapath_1.mux_wd3.dout [28])
);

INVX1 _12430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[29]),
    .Y(_3352_)
);

NAND2X1 _12431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf5),
    .B(\datapath_1.Data [29]),
    .Y(_3353_)
);

OAI21X1 _12432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3352_),
    .B(MemToReg_bF$buf4),
    .C(_3353_),
    .Y(\datapath_1.mux_wd3.dout [29])
);

INVX1 _12433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[30]),
    .Y(_3354_)
);

NAND2X1 _12434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf3),
    .B(\datapath_1.Data [30]),
    .Y(_3355_)
);

OAI21X1 _12435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3354_),
    .B(MemToReg_bF$buf2),
    .C(_3355_),
    .Y(\datapath_1.mux_wd3.dout [30])
);

INVX1 _12436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[31]),
    .Y(_3356_)
);

NAND2X1 _12437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(MemToReg_bF$buf1),
    .B(\datapath_1.Data [31]),
    .Y(_3357_)
);

OAI21X1 _12438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3356_),
    .B(MemToReg_bF$buf0),
    .C(_3357_),
    .Y(\datapath_1.mux_wd3.dout [31])
);

INVX1 _12439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[0]),
    .Y(_3423_)
);

NAND2X1 _12440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.ALUResult [0]),
    .B(vdd),
    .Y(_3424_)
);

OAI21X1 _12441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3423_),
    .B(vdd),
    .C(_3424_),
    .Y(_3360_[0])
);

INVX1 _12442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[1]),
    .Y(_3361_)
);

NAND2X1 _12443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [1]),
    .Y(_3362_)
);

OAI21X1 _12444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3361_),
    .B(vdd),
    .C(_3362_),
    .Y(_3360_[1])
);

INVX1 _12445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[2]),
    .Y(_3363_)
);

NAND2X1 _12446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [2]),
    .Y(_3364_)
);

OAI21X1 _12447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3363_),
    .B(vdd),
    .C(_3364_),
    .Y(_3360_[2])
);

INVX1 _12448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[3]),
    .Y(_3365_)
);

NAND2X1 _12449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [3]),
    .Y(_3366_)
);

OAI21X1 _12450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3365_),
    .B(vdd),
    .C(_3366_),
    .Y(_3360_[3])
);

INVX1 _12451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[4]),
    .Y(_3367_)
);

NAND2X1 _12452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [4]),
    .Y(_3368_)
);

OAI21X1 _12453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3367_),
    .B(vdd),
    .C(_3368_),
    .Y(_3360_[4])
);

INVX1 _12454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[5]),
    .Y(_3369_)
);

NAND2X1 _12455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [5]),
    .Y(_3370_)
);

OAI21X1 _12456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3369_),
    .B(vdd),
    .C(_3370_),
    .Y(_3360_[5])
);

INVX1 _12457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[6]),
    .Y(_3371_)
);

NAND2X1 _12458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [6]),
    .Y(_3372_)
);

OAI21X1 _12459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3371_),
    .B(vdd),
    .C(_3372_),
    .Y(_3360_[6])
);

INVX1 _12460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[7]),
    .Y(_3373_)
);

NAND2X1 _12461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [7]),
    .Y(_3374_)
);

OAI21X1 _12462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3373_),
    .B(vdd),
    .C(_3374_),
    .Y(_3360_[7])
);

INVX1 _12463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[8]),
    .Y(_3375_)
);

NAND2X1 _12464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [8]),
    .Y(_3376_)
);

OAI21X1 _12465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3375_),
    .B(vdd),
    .C(_3376_),
    .Y(_3360_[8])
);

INVX1 _12466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[9]),
    .Y(_3377_)
);

NAND2X1 _12467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [9]),
    .Y(_3378_)
);

OAI21X1 _12468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3377_),
    .B(vdd),
    .C(_3378_),
    .Y(_3360_[9])
);

INVX1 _12469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[10]),
    .Y(_3379_)
);

NAND2X1 _12470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [10]),
    .Y(_3380_)
);

OAI21X1 _12471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3379_),
    .B(vdd),
    .C(_3380_),
    .Y(_3360_[10])
);

INVX1 _12472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[11]),
    .Y(_3381_)
);

NAND2X1 _12473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [11]),
    .Y(_3382_)
);

OAI21X1 _12474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3381_),
    .B(vdd),
    .C(_3382_),
    .Y(_3360_[11])
);

INVX1 _12475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[12]),
    .Y(_3383_)
);

NAND2X1 _12476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [12]),
    .Y(_3384_)
);

OAI21X1 _12477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3383_),
    .B(vdd),
    .C(_3384_),
    .Y(_3360_[12])
);

INVX1 _12478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[13]),
    .Y(_3385_)
);

NAND2X1 _12479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [13]),
    .Y(_3386_)
);

OAI21X1 _12480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3385_),
    .B(vdd),
    .C(_3386_),
    .Y(_3360_[13])
);

INVX1 _12481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[14]),
    .Y(_3387_)
);

NAND2X1 _12482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [14]),
    .Y(_3388_)
);

OAI21X1 _12483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3387_),
    .B(vdd),
    .C(_3388_),
    .Y(_3360_[14])
);

INVX1 _12484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[15]),
    .Y(_3389_)
);

NAND2X1 _12485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [15]),
    .Y(_3390_)
);

OAI21X1 _12486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3389_),
    .B(vdd),
    .C(_3390_),
    .Y(_3360_[15])
);

INVX1 _12487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[16]),
    .Y(_3391_)
);

NAND2X1 _12488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [16]),
    .Y(_3392_)
);

OAI21X1 _12489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3391_),
    .B(vdd),
    .C(_3392_),
    .Y(_3360_[16])
);

INVX1 _12490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[17]),
    .Y(_3393_)
);

NAND2X1 _12491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [17]),
    .Y(_3394_)
);

OAI21X1 _12492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3393_),
    .B(vdd),
    .C(_3394_),
    .Y(_3360_[17])
);

INVX1 _12493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[18]),
    .Y(_3395_)
);

NAND2X1 _12494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [18]),
    .Y(_3396_)
);

OAI21X1 _12495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3395_),
    .B(vdd),
    .C(_3396_),
    .Y(_3360_[18])
);

INVX1 _12496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[19]),
    .Y(_3397_)
);

NAND2X1 _12497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [19]),
    .Y(_3398_)
);

OAI21X1 _12498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3397_),
    .B(vdd),
    .C(_3398_),
    .Y(_3360_[19])
);

INVX1 _12499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[20]),
    .Y(_3399_)
);

NAND2X1 _12500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [20]),
    .Y(_3400_)
);

OAI21X1 _12501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3399_),
    .B(vdd),
    .C(_3400_),
    .Y(_3360_[20])
);

INVX1 _12502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[21]),
    .Y(_3401_)
);

NAND2X1 _12503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [21]),
    .Y(_3402_)
);

OAI21X1 _12504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3401_),
    .B(vdd),
    .C(_3402_),
    .Y(_3360_[21])
);

INVX1 _12505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[22]),
    .Y(_3403_)
);

NAND2X1 _12506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [22]),
    .Y(_3404_)
);

OAI21X1 _12507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3403_),
    .B(vdd),
    .C(_3404_),
    .Y(_3360_[22])
);

INVX1 _12508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[23]),
    .Y(_3405_)
);

NAND2X1 _12509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [23]),
    .Y(_3406_)
);

OAI21X1 _12510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3405_),
    .B(vdd),
    .C(_3406_),
    .Y(_3360_[23])
);

INVX1 _12511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[24]),
    .Y(_3407_)
);

NAND2X1 _12512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [24]),
    .Y(_3408_)
);

OAI21X1 _12513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3407_),
    .B(vdd),
    .C(_3408_),
    .Y(_3360_[24])
);

INVX1 _12514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[25]),
    .Y(_3409_)
);

NAND2X1 _12515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [25]),
    .Y(_3410_)
);

OAI21X1 _12516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3409_),
    .B(vdd),
    .C(_3410_),
    .Y(_3360_[25])
);

INVX1 _12517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[26]),
    .Y(_3411_)
);

NAND2X1 _12518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [26]),
    .Y(_3412_)
);

OAI21X1 _12519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3411_),
    .B(vdd),
    .C(_3412_),
    .Y(_3360_[26])
);

INVX1 _12520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[27]),
    .Y(_3413_)
);

NAND2X1 _12521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [27]),
    .Y(_3414_)
);

OAI21X1 _12522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3413_),
    .B(vdd),
    .C(_3414_),
    .Y(_3360_[27])
);

INVX1 _12523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[28]),
    .Y(_3415_)
);

NAND2X1 _12524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [28]),
    .Y(_3416_)
);

OAI21X1 _12525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3415_),
    .B(vdd),
    .C(_3416_),
    .Y(_3360_[28])
);

INVX1 _12526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[29]),
    .Y(_3417_)
);

NAND2X1 _12527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [29]),
    .Y(_3418_)
);

OAI21X1 _12528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3417_),
    .B(vdd),
    .C(_3418_),
    .Y(_3360_[29])
);

INVX1 _12529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[30]),
    .Y(_3419_)
);

NAND2X1 _12530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [30]),
    .Y(_3420_)
);

OAI21X1 _12531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3419_),
    .B(vdd),
    .C(_3420_),
    .Y(_3360_[30])
);

INVX1 _12532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ALUOut[31]),
    .Y(_3421_)
);

NAND2X1 _12533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.ALUResult [31]),
    .Y(_3422_)
);

OAI21X1 _12534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3421_),
    .B(vdd),
    .C(_3422_),
    .Y(_3360_[31])
);

DFFSR _12535_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_3360_[0]),
    .Q(ALUOut[0]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _12536_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_3360_[1]),
    .Q(ALUOut[1]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _12537_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_3360_[2]),
    .Q(ALUOut[2]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _12538_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_3360_[3]),
    .Q(ALUOut[3]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _12539_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_3360_[4]),
    .Q(ALUOut[4]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _12540_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_3360_[5]),
    .Q(ALUOut[5]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _12541_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_3360_[6]),
    .Q(ALUOut[6]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _12542_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_3360_[7]),
    .Q(ALUOut[7]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _12543_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_3360_[8]),
    .Q(ALUOut[8]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _12544_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_3360_[9]),
    .Q(ALUOut[9]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _12545_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_3360_[10]),
    .Q(ALUOut[10]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _12546_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_3360_[11]),
    .Q(ALUOut[11]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _12547_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_3360_[12]),
    .Q(ALUOut[12]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _12548_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_3360_[13]),
    .Q(ALUOut[13]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _12549_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_3360_[14]),
    .Q(ALUOut[14]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _12550_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_3360_[15]),
    .Q(ALUOut[15]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _12551_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_3360_[16]),
    .Q(ALUOut[16]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _12552_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_3360_[17]),
    .Q(ALUOut[17]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _12553_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_3360_[18]),
    .Q(ALUOut[18]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _12554_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_3360_[19]),
    .Q(ALUOut[19]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _12555_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_3360_[20]),
    .Q(ALUOut[20]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _12556_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_3360_[21]),
    .Q(ALUOut[21]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _12557_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_3360_[22]),
    .Q(ALUOut[22]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _12558_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_3360_[23]),
    .Q(ALUOut[23]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _12559_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_3360_[24]),
    .Q(ALUOut[24]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _12560_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_3360_[25]),
    .Q(ALUOut[25]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _12561_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_3360_[26]),
    .Q(ALUOut[26]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _12562_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_3360_[27]),
    .Q(ALUOut[27]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _12563_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_3360_[28]),
    .Q(ALUOut[28]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _12564_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_3360_[29]),
    .Q(ALUOut[29]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _12565_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_3360_[30]),
    .Q(ALUOut[30]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _12566_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_3360_[31]),
    .Q(ALUOut[31]),
    .R(rst_bF$buf82),
    .S(vdd)
);

INVX1 _12567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [0]),
    .Y(_3488_)
);

NAND2X1 _12568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(memoryOutData[0]),
    .B(vdd),
    .Y(_3489_)
);

OAI21X1 _12569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3488_),
    .B(vdd),
    .C(_3489_),
    .Y(_3425_[0])
);

INVX1 _12570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [1]),
    .Y(_3426_)
);

NAND2X1 _12571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[1]),
    .Y(_3427_)
);

OAI21X1 _12572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3426_),
    .B(vdd),
    .C(_3427_),
    .Y(_3425_[1])
);

INVX1 _12573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [2]),
    .Y(_3428_)
);

NAND2X1 _12574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[2]),
    .Y(_3429_)
);

OAI21X1 _12575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3428_),
    .B(vdd),
    .C(_3429_),
    .Y(_3425_[2])
);

INVX1 _12576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [3]),
    .Y(_3430_)
);

NAND2X1 _12577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[3]),
    .Y(_3431_)
);

OAI21X1 _12578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3430_),
    .B(vdd),
    .C(_3431_),
    .Y(_3425_[3])
);

INVX1 _12579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [4]),
    .Y(_3432_)
);

NAND2X1 _12580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[4]),
    .Y(_3433_)
);

OAI21X1 _12581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3432_),
    .B(vdd),
    .C(_3433_),
    .Y(_3425_[4])
);

INVX1 _12582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [5]),
    .Y(_3434_)
);

NAND2X1 _12583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[5]),
    .Y(_3435_)
);

OAI21X1 _12584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3434_),
    .B(vdd),
    .C(_3435_),
    .Y(_3425_[5])
);

INVX1 _12585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [6]),
    .Y(_3436_)
);

NAND2X1 _12586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[6]),
    .Y(_3437_)
);

OAI21X1 _12587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3436_),
    .B(vdd),
    .C(_3437_),
    .Y(_3425_[6])
);

INVX1 _12588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [7]),
    .Y(_3438_)
);

NAND2X1 _12589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[7]),
    .Y(_3439_)
);

OAI21X1 _12590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3438_),
    .B(vdd),
    .C(_3439_),
    .Y(_3425_[7])
);

INVX1 _12591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [8]),
    .Y(_3440_)
);

NAND2X1 _12592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[8]),
    .Y(_3441_)
);

OAI21X1 _12593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(vdd),
    .C(_3441_),
    .Y(_3425_[8])
);

INVX1 _12594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [9]),
    .Y(_3442_)
);

NAND2X1 _12595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[9]),
    .Y(_3443_)
);

OAI21X1 _12596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3442_),
    .B(vdd),
    .C(_3443_),
    .Y(_3425_[9])
);

INVX1 _12597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [10]),
    .Y(_3444_)
);

NAND2X1 _12598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[10]),
    .Y(_3445_)
);

OAI21X1 _12599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3444_),
    .B(vdd),
    .C(_3445_),
    .Y(_3425_[10])
);

INVX1 _12600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [11]),
    .Y(_3446_)
);

NAND2X1 _12601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[11]),
    .Y(_3447_)
);

OAI21X1 _12602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3446_),
    .B(vdd),
    .C(_3447_),
    .Y(_3425_[11])
);

INVX1 _12603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [12]),
    .Y(_3448_)
);

NAND2X1 _12604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[12]),
    .Y(_3449_)
);

OAI21X1 _12605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .B(vdd),
    .C(_3449_),
    .Y(_3425_[12])
);

INVX1 _12606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [13]),
    .Y(_3450_)
);

NAND2X1 _12607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[13]),
    .Y(_3451_)
);

OAI21X1 _12608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3450_),
    .B(vdd),
    .C(_3451_),
    .Y(_3425_[13])
);

INVX1 _12609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [14]),
    .Y(_3452_)
);

NAND2X1 _12610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[14]),
    .Y(_3453_)
);

OAI21X1 _12611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3452_),
    .B(vdd),
    .C(_3453_),
    .Y(_3425_[14])
);

INVX1 _12612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [15]),
    .Y(_3454_)
);

NAND2X1 _12613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[15]),
    .Y(_3455_)
);

OAI21X1 _12614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3454_),
    .B(vdd),
    .C(_3455_),
    .Y(_3425_[15])
);

INVX1 _12615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [16]),
    .Y(_3456_)
);

NAND2X1 _12616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[16]),
    .Y(_3457_)
);

OAI21X1 _12617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3456_),
    .B(vdd),
    .C(_3457_),
    .Y(_3425_[16])
);

INVX1 _12618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [17]),
    .Y(_3458_)
);

NAND2X1 _12619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[17]),
    .Y(_3459_)
);

OAI21X1 _12620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3458_),
    .B(vdd),
    .C(_3459_),
    .Y(_3425_[17])
);

INVX1 _12621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [18]),
    .Y(_3460_)
);

NAND2X1 _12622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[18]),
    .Y(_3461_)
);

OAI21X1 _12623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3460_),
    .B(vdd),
    .C(_3461_),
    .Y(_3425_[18])
);

INVX1 _12624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [19]),
    .Y(_3462_)
);

NAND2X1 _12625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[19]),
    .Y(_3463_)
);

OAI21X1 _12626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3462_),
    .B(vdd),
    .C(_3463_),
    .Y(_3425_[19])
);

INVX1 _12627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [20]),
    .Y(_3464_)
);

NAND2X1 _12628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[20]),
    .Y(_3465_)
);

OAI21X1 _12629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3464_),
    .B(vdd),
    .C(_3465_),
    .Y(_3425_[20])
);

INVX1 _12630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [21]),
    .Y(_3466_)
);

NAND2X1 _12631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[21]),
    .Y(_3467_)
);

OAI21X1 _12632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3466_),
    .B(vdd),
    .C(_3467_),
    .Y(_3425_[21])
);

INVX1 _12633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [22]),
    .Y(_3468_)
);

NAND2X1 _12634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[22]),
    .Y(_3469_)
);

OAI21X1 _12635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3468_),
    .B(vdd),
    .C(_3469_),
    .Y(_3425_[22])
);

INVX1 _12636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [23]),
    .Y(_3470_)
);

NAND2X1 _12637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[23]),
    .Y(_3471_)
);

OAI21X1 _12638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3470_),
    .B(vdd),
    .C(_3471_),
    .Y(_3425_[23])
);

INVX1 _12639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [24]),
    .Y(_3472_)
);

NAND2X1 _12640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[24]),
    .Y(_3473_)
);

OAI21X1 _12641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3472_),
    .B(vdd),
    .C(_3473_),
    .Y(_3425_[24])
);

INVX1 _12642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [25]),
    .Y(_3474_)
);

NAND2X1 _12643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[25]),
    .Y(_3475_)
);

OAI21X1 _12644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3474_),
    .B(vdd),
    .C(_3475_),
    .Y(_3425_[25])
);

INVX1 _12645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [26]),
    .Y(_3476_)
);

NAND2X1 _12646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[26]),
    .Y(_3477_)
);

OAI21X1 _12647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3476_),
    .B(vdd),
    .C(_3477_),
    .Y(_3425_[26])
);

INVX1 _12648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [27]),
    .Y(_3478_)
);

NAND2X1 _12649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[27]),
    .Y(_3479_)
);

OAI21X1 _12650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3478_),
    .B(vdd),
    .C(_3479_),
    .Y(_3425_[27])
);

INVX1 _12651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [28]),
    .Y(_3480_)
);

NAND2X1 _12652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[28]),
    .Y(_3481_)
);

OAI21X1 _12653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3480_),
    .B(vdd),
    .C(_3481_),
    .Y(_3425_[28])
);

INVX1 _12654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [29]),
    .Y(_3482_)
);

NAND2X1 _12655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[29]),
    .Y(_3483_)
);

OAI21X1 _12656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3482_),
    .B(vdd),
    .C(_3483_),
    .Y(_3425_[29])
);

INVX1 _12657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [30]),
    .Y(_3484_)
);

NAND2X1 _12658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[30]),
    .Y(_3485_)
);

OAI21X1 _12659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3484_),
    .B(vdd),
    .C(_3485_),
    .Y(_3425_[30])
);

INVX1 _12660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.Data [31]),
    .Y(_3486_)
);

NAND2X1 _12661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(memoryOutData[31]),
    .Y(_3487_)
);

OAI21X1 _12662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3486_),
    .B(vdd),
    .C(_3487_),
    .Y(_3425_[31])
);

DFFSR _12663_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_3425_[0]),
    .Q(\datapath_1.Data [0]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _12664_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_3425_[1]),
    .Q(\datapath_1.Data [1]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _12665_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_3425_[2]),
    .Q(\datapath_1.Data [2]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _12666_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_3425_[3]),
    .Q(\datapath_1.Data [3]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _12667_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_3425_[4]),
    .Q(\datapath_1.Data [4]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _12668_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_3425_[5]),
    .Q(\datapath_1.Data [5]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _12669_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_3425_[6]),
    .Q(\datapath_1.Data [6]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _12670_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_3425_[7]),
    .Q(\datapath_1.Data [7]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _12671_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_3425_[8]),
    .Q(\datapath_1.Data [8]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _12672_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_3425_[9]),
    .Q(\datapath_1.Data [9]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _12673_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_3425_[10]),
    .Q(\datapath_1.Data [10]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _12674_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_3425_[11]),
    .Q(\datapath_1.Data [11]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _12675_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_3425_[12]),
    .Q(\datapath_1.Data [12]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _12676_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_3425_[13]),
    .Q(\datapath_1.Data [13]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _12677_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_3425_[14]),
    .Q(\datapath_1.Data [14]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _12678_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_3425_[15]),
    .Q(\datapath_1.Data [15]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _12679_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_3425_[16]),
    .Q(\datapath_1.Data [16]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _12680_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_3425_[17]),
    .Q(\datapath_1.Data [17]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _12681_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_3425_[18]),
    .Q(\datapath_1.Data [18]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _12682_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_3425_[19]),
    .Q(\datapath_1.Data [19]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _12683_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_3425_[20]),
    .Q(\datapath_1.Data [20]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _12684_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_3425_[21]),
    .Q(\datapath_1.Data [21]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _12685_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_3425_[22]),
    .Q(\datapath_1.Data [22]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _12686_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_3425_[23]),
    .Q(\datapath_1.Data [23]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _12687_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_3425_[24]),
    .Q(\datapath_1.Data [24]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _12688_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_3425_[25]),
    .Q(\datapath_1.Data [25]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _12689_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_3425_[26]),
    .Q(\datapath_1.Data [26]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _12690_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_3425_[27]),
    .Q(\datapath_1.Data [27]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _12691_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_3425_[28]),
    .Q(\datapath_1.Data [28]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _12692_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_3425_[29]),
    .Q(\datapath_1.Data [29]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _12693_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_3425_[30]),
    .Q(\datapath_1.Data [30]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _12694_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_3425_[31]),
    .Q(\datapath_1.Data [31]),
    .R(rst_bF$buf50),
    .S(vdd)
);

INVX1 _12695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [0]),
    .Y(_3553_)
);

NAND2X1 _12696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(memoryOutData[0]),
    .B(IRWrite_bF$buf6),
    .Y(_3554_)
);

OAI21X1 _12697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3553_),
    .B(IRWrite_bF$buf5),
    .C(_3554_),
    .Y(_3490_[0])
);

INVX1 _12698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [1]),
    .Y(_3491_)
);

NAND2X1 _12699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[1]),
    .Y(_3492_)
);

OAI21X1 _12700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(IRWrite_bF$buf3),
    .C(_3492_),
    .Y(_3490_[1])
);

INVX1 _12701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [2]),
    .Y(_3493_)
);

NAND2X1 _12702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[2]),
    .Y(_3494_)
);

OAI21X1 _12703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3493_),
    .B(IRWrite_bF$buf1),
    .C(_3494_),
    .Y(_3490_[2])
);

INVX1 _12704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [3]),
    .Y(_3495_)
);

NAND2X1 _12705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[3]),
    .Y(_3496_)
);

OAI21X1 _12706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3495_),
    .B(IRWrite_bF$buf7),
    .C(_3496_),
    .Y(_3490_[3])
);

INVX1 _12707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [4]),
    .Y(_3497_)
);

NAND2X1 _12708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[4]),
    .Y(_3498_)
);

OAI21X1 _12709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3497_),
    .B(IRWrite_bF$buf5),
    .C(_3498_),
    .Y(_3490_[4])
);

INVX1 _12710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\aluControl_1.inst [5]),
    .Y(_3499_)
);

NAND2X1 _12711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[5]),
    .Y(_3500_)
);

OAI21X1 _12712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3499_),
    .B(IRWrite_bF$buf3),
    .C(_3500_),
    .Y(_3490_[5])
);

INVX1 _12713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [8]),
    .Y(_3501_)
);

NAND2X1 _12714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[6]),
    .Y(_3502_)
);

OAI21X1 _12715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3501_),
    .B(IRWrite_bF$buf1),
    .C(_3502_),
    .Y(_3490_[6])
);

INVX1 _12716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [9]),
    .Y(_3503_)
);

NAND2X1 _12717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[7]),
    .Y(_3504_)
);

OAI21X1 _12718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3503_),
    .B(IRWrite_bF$buf7),
    .C(_3504_),
    .Y(_3490_[7])
);

INVX1 _12719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [10]),
    .Y(_3505_)
);

NAND2X1 _12720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[8]),
    .Y(_3506_)
);

OAI21X1 _12721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3505_),
    .B(IRWrite_bF$buf5),
    .C(_3506_),
    .Y(_3490_[8])
);

INVX1 _12722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [11]),
    .Y(_3507_)
);

NAND2X1 _12723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[9]),
    .Y(_3508_)
);

OAI21X1 _12724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3507_),
    .B(IRWrite_bF$buf3),
    .C(_3508_),
    .Y(_3490_[9])
);

INVX1 _12725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [12]),
    .Y(_3509_)
);

NAND2X1 _12726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[10]),
    .Y(_3510_)
);

OAI21X1 _12727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3509_),
    .B(IRWrite_bF$buf1),
    .C(_3510_),
    .Y(_3490_[10])
);

INVX1 _12728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [13]),
    .Y(_3511_)
);

NAND2X1 _12729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[11]),
    .Y(_3512_)
);

OAI21X1 _12730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3511_),
    .B(IRWrite_bF$buf7),
    .C(_3512_),
    .Y(_3490_[11])
);

INVX1 _12731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [14]),
    .Y(_3513_)
);

NAND2X1 _12732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[12]),
    .Y(_3514_)
);

OAI21X1 _12733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3513_),
    .B(IRWrite_bF$buf5),
    .C(_3514_),
    .Y(_3490_[12])
);

INVX1 _12734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [15]),
    .Y(_3515_)
);

NAND2X1 _12735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[13]),
    .Y(_3516_)
);

OAI21X1 _12736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3515_),
    .B(IRWrite_bF$buf3),
    .C(_3516_),
    .Y(_3490_[13])
);

INVX1 _12737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [16]),
    .Y(_3517_)
);

NAND2X1 _12738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[14]),
    .Y(_3518_)
);

OAI21X1 _12739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3517_),
    .B(IRWrite_bF$buf1),
    .C(_3518_),
    .Y(_3490_[14])
);

INVX1 _12740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_17_bF$buf0 ),
    .Y(_3519_)
);

NAND2X1 _12741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[15]),
    .Y(_3520_)
);

OAI21X1 _12742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3519_),
    .B(IRWrite_bF$buf7),
    .C(_3520_),
    .Y(_3490_[15])
);

INVX1 _12743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [18]),
    .Y(_3521_)
);

NAND2X1 _12744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[16]),
    .Y(_3522_)
);

OAI21X1 _12745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3521_),
    .B(IRWrite_bF$buf5),
    .C(_3522_),
    .Y(_3490_[16])
);

INVX1 _12746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [19]),
    .Y(_3523_)
);

NAND2X1 _12747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[17]),
    .Y(_3524_)
);

OAI21X1 _12748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3523_),
    .B(IRWrite_bF$buf3),
    .C(_3524_),
    .Y(_3490_[17])
);

INVX1 _12749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [20]),
    .Y(_3525_)
);

NAND2X1 _12750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[18]),
    .Y(_3526_)
);

OAI21X1 _12751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3525_),
    .B(IRWrite_bF$buf1),
    .C(_3526_),
    .Y(_3490_[18])
);

INVX1 _12752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .Y(_3527_)
);

NAND2X1 _12753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[19]),
    .Y(_3528_)
);

OAI21X1 _12754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3527_),
    .B(IRWrite_bF$buf7),
    .C(_3528_),
    .Y(_3490_[19])
);

INVX1 _12755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_3529_)
);

NAND2X1 _12756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[20]),
    .Y(_3530_)
);

OAI21X1 _12757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .B(IRWrite_bF$buf5),
    .C(_3530_),
    .Y(_3490_[20])
);

INVX1 _12758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [23]),
    .Y(_3531_)
);

NAND2X1 _12759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[21]),
    .Y(_3532_)
);

OAI21X1 _12760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3531_),
    .B(IRWrite_bF$buf3),
    .C(_3532_),
    .Y(_3490_[21])
);

INVX1 _12761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .Y(_3533_)
);

NAND2X1 _12762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[22]),
    .Y(_3534_)
);

OAI21X1 _12763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3533_),
    .B(IRWrite_bF$buf1),
    .C(_3534_),
    .Y(_3490_[22])
);

INVX1 _12764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [25]),
    .Y(_3535_)
);

NAND2X1 _12765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[23]),
    .Y(_3536_)
);

OAI21X1 _12766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3535_),
    .B(IRWrite_bF$buf7),
    .C(_3536_),
    .Y(_3490_[23])
);

INVX1 _12767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .Y(_3537_)
);

NAND2X1 _12768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[24]),
    .Y(_3538_)
);

OAI21X1 _12769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3537_),
    .B(IRWrite_bF$buf5),
    .C(_3538_),
    .Y(_3490_[24])
);

INVX1 _12770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .Y(_3539_)
);

NAND2X1 _12771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[25]),
    .Y(_3540_)
);

OAI21X1 _12772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3539_),
    .B(IRWrite_bF$buf3),
    .C(_3540_),
    .Y(_3490_[25])
);

INVX1 _12773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [0]),
    .Y(_3541_)
);

NAND2X1 _12774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[26]),
    .Y(_3542_)
);

OAI21X1 _12775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3541_),
    .B(IRWrite_bF$buf1),
    .C(_3542_),
    .Y(_3490_[26])
);

INVX1 _12776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [1]),
    .Y(_3543_)
);

NAND2X1 _12777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[27]),
    .Y(_3544_)
);

OAI21X1 _12778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3543_),
    .B(IRWrite_bF$buf7),
    .C(_3544_),
    .Y(_3490_[27])
);

INVX1 _12779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [2]),
    .Y(_3545_)
);

NAND2X1 _12780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf6),
    .B(memoryOutData[28]),
    .Y(_3546_)
);

OAI21X1 _12781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3545_),
    .B(IRWrite_bF$buf5),
    .C(_3546_),
    .Y(_3490_[28])
);

INVX1 _12782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [3]),
    .Y(_3547_)
);

NAND2X1 _12783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf4),
    .B(memoryOutData[29]),
    .Y(_3548_)
);

OAI21X1 _12784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3547_),
    .B(IRWrite_bF$buf3),
    .C(_3548_),
    .Y(_3490_[29])
);

INVX1 _12785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [4]),
    .Y(_3549_)
);

NAND2X1 _12786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf2),
    .B(memoryOutData[30]),
    .Y(_3550_)
);

OAI21X1 _12787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3549_),
    .B(IRWrite_bF$buf1),
    .C(_3550_),
    .Y(_3490_[30])
);

INVX1 _12788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\control_1.op [5]),
    .Y(_3551_)
);

NAND2X1 _12789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRWrite_bF$buf0),
    .B(memoryOutData[31]),
    .Y(_3552_)
);

OAI21X1 _12790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3551_),
    .B(IRWrite_bF$buf7),
    .C(_3552_),
    .Y(_3490_[31])
);

DFFSR _12791_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_3490_[0]),
    .Q(\aluControl_1.inst [0]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _12792_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_3490_[1]),
    .Q(\aluControl_1.inst [1]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _12793_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_3490_[2]),
    .Q(\aluControl_1.inst [2]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _12794_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_3490_[3]),
    .Q(\aluControl_1.inst [3]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _12795_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_3490_[4]),
    .Q(\aluControl_1.inst [4]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _12796_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_3490_[5]),
    .Q(\aluControl_1.inst [5]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _12797_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_3490_[6]),
    .Q(\datapath_1.PCJump [8]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _12798_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_3490_[7]),
    .Q(\datapath_1.PCJump [9]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _12799_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_3490_[8]),
    .Q(\datapath_1.PCJump [10]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _12800_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_3490_[9]),
    .Q(\datapath_1.PCJump [11]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _12801_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_3490_[10]),
    .Q(\datapath_1.PCJump [12]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _12802_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_3490_[11]),
    .Q(\datapath_1.PCJump [13]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _12803_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_3490_[12]),
    .Q(\datapath_1.PCJump [14]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _12804_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_3490_[13]),
    .Q(\datapath_1.PCJump [15]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _12805_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_3490_[14]),
    .Q(\datapath_1.PCJump [16]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _12806_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_3490_[15]),
    .Q(\datapath_1.PCJump [17]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _12807_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_3490_[16]),
    .Q(\datapath_1.PCJump [18]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _12808_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_3490_[17]),
    .Q(\datapath_1.PCJump [19]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _12809_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_3490_[18]),
    .Q(\datapath_1.PCJump [20]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _12810_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_3490_[19]),
    .Q(\datapath_1.PCJump [21]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _12811_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_3490_[20]),
    .Q(\datapath_1.PCJump [22]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _12812_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_3490_[21]),
    .Q(\datapath_1.PCJump [23]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _12813_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_3490_[22]),
    .Q(\datapath_1.PCJump [24]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _12814_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_3490_[23]),
    .Q(\datapath_1.PCJump [25]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _12815_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_3490_[24]),
    .Q(\datapath_1.PCJump [26]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _12816_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_3490_[25]),
    .Q(\datapath_1.PCJump [27]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _12817_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_3490_[26]),
    .Q(\control_1.op [0]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _12818_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_3490_[27]),
    .Q(\control_1.op [1]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _12819_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_3490_[28]),
    .Q(\control_1.op [2]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _12820_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_3490_[29]),
    .Q(\control_1.op [3]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _12821_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_3490_[30]),
    .Q(\control_1.op [4]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _12822_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_3490_[31]),
    .Q(\control_1.op [5]),
    .R(rst_bF$buf18),
    .S(vdd)
);

INVX1 _12823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [0]),
    .Y(_3618_)
);

NAND2X1 _12824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.rd1 [0]),
    .B(vdd),
    .Y(_3619_)
);

OAI21X1 _12825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3618_),
    .B(vdd),
    .C(_3619_),
    .Y(_3555_[0])
);

INVX1 _12826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [1]),
    .Y(_3556_)
);

NAND2X1 _12827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [1]),
    .Y(_3557_)
);

OAI21X1 _12828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3556_),
    .B(vdd),
    .C(_3557_),
    .Y(_3555_[1])
);

INVX1 _12829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [2]),
    .Y(_3558_)
);

NAND2X1 _12830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [2]),
    .Y(_3559_)
);

OAI21X1 _12831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3558_),
    .B(vdd),
    .C(_3559_),
    .Y(_3555_[2])
);

INVX1 _12832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [3]),
    .Y(_3560_)
);

NAND2X1 _12833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [3]),
    .Y(_3561_)
);

OAI21X1 _12834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3560_),
    .B(vdd),
    .C(_3561_),
    .Y(_3555_[3])
);

INVX1 _12835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [4]),
    .Y(_3562_)
);

NAND2X1 _12836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [4]),
    .Y(_3563_)
);

OAI21X1 _12837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3562_),
    .B(vdd),
    .C(_3563_),
    .Y(_3555_[4])
);

INVX1 _12838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [5]),
    .Y(_3564_)
);

NAND2X1 _12839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [5]),
    .Y(_3565_)
);

OAI21X1 _12840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3564_),
    .B(vdd),
    .C(_3565_),
    .Y(_3555_[5])
);

INVX1 _12841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [6]),
    .Y(_3566_)
);

NAND2X1 _12842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [6]),
    .Y(_3567_)
);

OAI21X1 _12843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3566_),
    .B(vdd),
    .C(_3567_),
    .Y(_3555_[6])
);

INVX1 _12844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [7]),
    .Y(_3568_)
);

NAND2X1 _12845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [7]),
    .Y(_3569_)
);

OAI21X1 _12846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(vdd),
    .C(_3569_),
    .Y(_3555_[7])
);

INVX1 _12847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [8]),
    .Y(_3570_)
);

NAND2X1 _12848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [8]),
    .Y(_3571_)
);

OAI21X1 _12849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3570_),
    .B(vdd),
    .C(_3571_),
    .Y(_3555_[8])
);

INVX1 _12850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [9]),
    .Y(_3572_)
);

NAND2X1 _12851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [9]),
    .Y(_3573_)
);

OAI21X1 _12852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3572_),
    .B(vdd),
    .C(_3573_),
    .Y(_3555_[9])
);

INVX1 _12853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [10]),
    .Y(_3574_)
);

NAND2X1 _12854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [10]),
    .Y(_3575_)
);

OAI21X1 _12855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3574_),
    .B(vdd),
    .C(_3575_),
    .Y(_3555_[10])
);

INVX1 _12856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [11]),
    .Y(_3576_)
);

NAND2X1 _12857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [11]),
    .Y(_3577_)
);

OAI21X1 _12858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3576_),
    .B(vdd),
    .C(_3577_),
    .Y(_3555_[11])
);

INVX1 _12859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [12]),
    .Y(_3578_)
);

NAND2X1 _12860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [12]),
    .Y(_3579_)
);

OAI21X1 _12861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3578_),
    .B(vdd),
    .C(_3579_),
    .Y(_3555_[12])
);

INVX1 _12862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [13]),
    .Y(_3580_)
);

NAND2X1 _12863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [13]),
    .Y(_3581_)
);

OAI21X1 _12864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3580_),
    .B(vdd),
    .C(_3581_),
    .Y(_3555_[13])
);

INVX1 _12865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [14]),
    .Y(_3582_)
);

NAND2X1 _12866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [14]),
    .Y(_3583_)
);

OAI21X1 _12867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3582_),
    .B(vdd),
    .C(_3583_),
    .Y(_3555_[14])
);

INVX1 _12868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [15]),
    .Y(_3584_)
);

NAND2X1 _12869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [15]),
    .Y(_3585_)
);

OAI21X1 _12870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3584_),
    .B(vdd),
    .C(_3585_),
    .Y(_3555_[15])
);

INVX1 _12871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [16]),
    .Y(_3586_)
);

NAND2X1 _12872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [16]),
    .Y(_3587_)
);

OAI21X1 _12873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3586_),
    .B(vdd),
    .C(_3587_),
    .Y(_3555_[16])
);

INVX1 _12874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [17]),
    .Y(_3588_)
);

NAND2X1 _12875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [17]),
    .Y(_3589_)
);

OAI21X1 _12876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3588_),
    .B(vdd),
    .C(_3589_),
    .Y(_3555_[17])
);

INVX1 _12877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [18]),
    .Y(_3590_)
);

NAND2X1 _12878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [18]),
    .Y(_3591_)
);

OAI21X1 _12879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3590_),
    .B(vdd),
    .C(_3591_),
    .Y(_3555_[18])
);

INVX1 _12880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [19]),
    .Y(_3592_)
);

NAND2X1 _12881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [19]),
    .Y(_3593_)
);

OAI21X1 _12882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3592_),
    .B(vdd),
    .C(_3593_),
    .Y(_3555_[19])
);

INVX1 _12883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [20]),
    .Y(_3594_)
);

NAND2X1 _12884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [20]),
    .Y(_3595_)
);

OAI21X1 _12885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3594_),
    .B(vdd),
    .C(_3595_),
    .Y(_3555_[20])
);

INVX1 _12886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [21]),
    .Y(_3596_)
);

NAND2X1 _12887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [21]),
    .Y(_3597_)
);

OAI21X1 _12888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3596_),
    .B(vdd),
    .C(_3597_),
    .Y(_3555_[21])
);

INVX1 _12889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [22]),
    .Y(_3598_)
);

NAND2X1 _12890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [22]),
    .Y(_3599_)
);

OAI21X1 _12891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3598_),
    .B(vdd),
    .C(_3599_),
    .Y(_3555_[22])
);

INVX1 _12892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [23]),
    .Y(_3600_)
);

NAND2X1 _12893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [23]),
    .Y(_3601_)
);

OAI21X1 _12894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3600_),
    .B(vdd),
    .C(_3601_),
    .Y(_3555_[23])
);

INVX1 _12895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [24]),
    .Y(_3602_)
);

NAND2X1 _12896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [24]),
    .Y(_3603_)
);

OAI21X1 _12897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3602_),
    .B(vdd),
    .C(_3603_),
    .Y(_3555_[24])
);

INVX1 _12898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [25]),
    .Y(_3604_)
);

NAND2X1 _12899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [25]),
    .Y(_3605_)
);

OAI21X1 _12900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3604_),
    .B(vdd),
    .C(_3605_),
    .Y(_3555_[25])
);

INVX1 _12901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [26]),
    .Y(_3606_)
);

NAND2X1 _12902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [26]),
    .Y(_3607_)
);

OAI21X1 _12903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3606_),
    .B(vdd),
    .C(_3607_),
    .Y(_3555_[26])
);

INVX1 _12904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [27]),
    .Y(_3608_)
);

NAND2X1 _12905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [27]),
    .Y(_3609_)
);

OAI21X1 _12906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3608_),
    .B(vdd),
    .C(_3609_),
    .Y(_3555_[27])
);

INVX1 _12907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [28]),
    .Y(_3610_)
);

NAND2X1 _12908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [28]),
    .Y(_3611_)
);

OAI21X1 _12909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3610_),
    .B(vdd),
    .C(_3611_),
    .Y(_3555_[28])
);

INVX1 _12910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [29]),
    .Y(_3612_)
);

NAND2X1 _12911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [29]),
    .Y(_3613_)
);

OAI21X1 _12912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3612_),
    .B(vdd),
    .C(_3613_),
    .Y(_3555_[29])
);

INVX1 _12913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [30]),
    .Y(_3614_)
);

NAND2X1 _12914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [30]),
    .Y(_3615_)
);

OAI21X1 _12915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3614_),
    .B(vdd),
    .C(_3615_),
    .Y(_3555_[30])
);

INVX1 _12916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a [31]),
    .Y(_3616_)
);

NAND2X1 _12917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd1 [31]),
    .Y(_3617_)
);

OAI21X1 _12918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3616_),
    .B(vdd),
    .C(_3617_),
    .Y(_3555_[31])
);

DFFSR _12919_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_3555_[0]),
    .Q(\datapath_1.a [0]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _12920_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_3555_[1]),
    .Q(\datapath_1.a [1]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _12921_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_3555_[2]),
    .Q(\datapath_1.a [2]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _12922_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_3555_[3]),
    .Q(\datapath_1.a [3]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _12923_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_3555_[4]),
    .Q(\datapath_1.a [4]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _12924_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_3555_[5]),
    .Q(\datapath_1.a [5]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _12925_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_3555_[6]),
    .Q(\datapath_1.a [6]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _12926_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_3555_[7]),
    .Q(\datapath_1.a [7]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _12927_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_3555_[8]),
    .Q(\datapath_1.a [8]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _12928_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_3555_[9]),
    .Q(\datapath_1.a [9]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _12929_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_3555_[10]),
    .Q(\datapath_1.a [10]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _12930_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_3555_[11]),
    .Q(\datapath_1.a [11]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _12931_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_3555_[12]),
    .Q(\datapath_1.a [12]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _12932_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_3555_[13]),
    .Q(\datapath_1.a [13]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _12933_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_3555_[14]),
    .Q(\datapath_1.a [14]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _12934_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_3555_[15]),
    .Q(\datapath_1.a [15]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _12935_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_3555_[16]),
    .Q(\datapath_1.a [16]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _12936_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_3555_[17]),
    .Q(\datapath_1.a [17]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _12937_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_3555_[18]),
    .Q(\datapath_1.a [18]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _12938_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_3555_[19]),
    .Q(\datapath_1.a [19]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _12939_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_3555_[20]),
    .Q(\datapath_1.a [20]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _12940_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_3555_[21]),
    .Q(\datapath_1.a [21]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _12941_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_3555_[22]),
    .Q(\datapath_1.a [22]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _12942_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_3555_[23]),
    .Q(\datapath_1.a [23]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _12943_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_3555_[24]),
    .Q(\datapath_1.a [24]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _12944_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_3555_[25]),
    .Q(\datapath_1.a [25]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _12945_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_3555_[26]),
    .Q(\datapath_1.a [26]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _12946_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_3555_[27]),
    .Q(\datapath_1.a [27]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _12947_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_3555_[28]),
    .Q(\datapath_1.a [28]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _12948_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_3555_[29]),
    .Q(\datapath_1.a [29]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _12949_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_3555_[30]),
    .Q(\datapath_1.a [30]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _12950_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_3555_[31]),
    .Q(\datapath_1.a [31]),
    .R(rst_bF$buf100),
    .S(vdd)
);

INVX1 _12951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[0]),
    .Y(_3683_)
);

NAND2X1 _12952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.rd2 [0]),
    .B(vdd),
    .Y(_3684_)
);

OAI21X1 _12953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3683_),
    .B(vdd),
    .C(_3684_),
    .Y(_3620_[0])
);

INVX1 _12954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[1]),
    .Y(_3621_)
);

NAND2X1 _12955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [1]),
    .Y(_3622_)
);

OAI21X1 _12956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3621_),
    .B(vdd),
    .C(_3622_),
    .Y(_3620_[1])
);

INVX1 _12957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[2]),
    .Y(_3623_)
);

NAND2X1 _12958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [2]),
    .Y(_3624_)
);

OAI21X1 _12959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3623_),
    .B(vdd),
    .C(_3624_),
    .Y(_3620_[2])
);

INVX1 _12960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[3]),
    .Y(_3625_)
);

NAND2X1 _12961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [3]),
    .Y(_3626_)
);

OAI21X1 _12962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3625_),
    .B(vdd),
    .C(_3626_),
    .Y(_3620_[3])
);

INVX1 _12963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[4]),
    .Y(_3627_)
);

NAND2X1 _12964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [4]),
    .Y(_3628_)
);

OAI21X1 _12965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3627_),
    .B(vdd),
    .C(_3628_),
    .Y(_3620_[4])
);

INVX1 _12966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[5]),
    .Y(_3629_)
);

NAND2X1 _12967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [5]),
    .Y(_3630_)
);

OAI21X1 _12968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3629_),
    .B(vdd),
    .C(_3630_),
    .Y(_3620_[5])
);

INVX1 _12969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[6]),
    .Y(_3631_)
);

NAND2X1 _12970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [6]),
    .Y(_3632_)
);

OAI21X1 _12971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3631_),
    .B(vdd),
    .C(_3632_),
    .Y(_3620_[6])
);

INVX1 _12972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[7]),
    .Y(_3633_)
);

NAND2X1 _12973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [7]),
    .Y(_3634_)
);

OAI21X1 _12974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3633_),
    .B(vdd),
    .C(_3634_),
    .Y(_3620_[7])
);

INVX1 _12975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[8]),
    .Y(_3635_)
);

NAND2X1 _12976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [8]),
    .Y(_3636_)
);

OAI21X1 _12977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3635_),
    .B(vdd),
    .C(_3636_),
    .Y(_3620_[8])
);

INVX1 _12978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[9]),
    .Y(_3637_)
);

NAND2X1 _12979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [9]),
    .Y(_3638_)
);

OAI21X1 _12980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3637_),
    .B(vdd),
    .C(_3638_),
    .Y(_3620_[9])
);

INVX1 _12981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[10]),
    .Y(_3639_)
);

NAND2X1 _12982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [10]),
    .Y(_3640_)
);

OAI21X1 _12983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3639_),
    .B(vdd),
    .C(_3640_),
    .Y(_3620_[10])
);

INVX1 _12984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[11]),
    .Y(_3641_)
);

NAND2X1 _12985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [11]),
    .Y(_3642_)
);

OAI21X1 _12986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3641_),
    .B(vdd),
    .C(_3642_),
    .Y(_3620_[11])
);

INVX1 _12987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[12]),
    .Y(_3643_)
);

NAND2X1 _12988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [12]),
    .Y(_3644_)
);

OAI21X1 _12989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3643_),
    .B(vdd),
    .C(_3644_),
    .Y(_3620_[12])
);

INVX1 _12990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[13]),
    .Y(_3645_)
);

NAND2X1 _12991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [13]),
    .Y(_3646_)
);

OAI21X1 _12992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3645_),
    .B(vdd),
    .C(_3646_),
    .Y(_3620_[13])
);

INVX1 _12993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[14]),
    .Y(_3647_)
);

NAND2X1 _12994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [14]),
    .Y(_3648_)
);

OAI21X1 _12995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3647_),
    .B(vdd),
    .C(_3648_),
    .Y(_3620_[14])
);

INVX1 _12996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[15]),
    .Y(_3649_)
);

NAND2X1 _12997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [15]),
    .Y(_3650_)
);

OAI21X1 _12998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3649_),
    .B(vdd),
    .C(_3650_),
    .Y(_3620_[15])
);

INVX1 _12999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[16]),
    .Y(_3651_)
);

NAND2X1 _13000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [16]),
    .Y(_3652_)
);

OAI21X1 _13001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3651_),
    .B(vdd),
    .C(_3652_),
    .Y(_3620_[16])
);

INVX1 _13002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[17]),
    .Y(_3653_)
);

NAND2X1 _13003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [17]),
    .Y(_3654_)
);

OAI21X1 _13004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3653_),
    .B(vdd),
    .C(_3654_),
    .Y(_3620_[17])
);

INVX1 _13005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[18]),
    .Y(_3655_)
);

NAND2X1 _13006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [18]),
    .Y(_3656_)
);

OAI21X1 _13007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3655_),
    .B(vdd),
    .C(_3656_),
    .Y(_3620_[18])
);

INVX1 _13008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[19]),
    .Y(_3657_)
);

NAND2X1 _13009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [19]),
    .Y(_3658_)
);

OAI21X1 _13010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3657_),
    .B(vdd),
    .C(_3658_),
    .Y(_3620_[19])
);

INVX1 _13011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[20]),
    .Y(_3659_)
);

NAND2X1 _13012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [20]),
    .Y(_3660_)
);

OAI21X1 _13013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3659_),
    .B(vdd),
    .C(_3660_),
    .Y(_3620_[20])
);

INVX1 _13014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[21]),
    .Y(_3661_)
);

NAND2X1 _13015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [21]),
    .Y(_3662_)
);

OAI21X1 _13016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3661_),
    .B(vdd),
    .C(_3662_),
    .Y(_3620_[21])
);

INVX1 _13017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[22]),
    .Y(_3663_)
);

NAND2X1 _13018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [22]),
    .Y(_3664_)
);

OAI21X1 _13019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3663_),
    .B(vdd),
    .C(_3664_),
    .Y(_3620_[22])
);

INVX1 _13020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[23]),
    .Y(_3665_)
);

NAND2X1 _13021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [23]),
    .Y(_3666_)
);

OAI21X1 _13022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3665_),
    .B(vdd),
    .C(_3666_),
    .Y(_3620_[23])
);

INVX1 _13023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[24]),
    .Y(_3667_)
);

NAND2X1 _13024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [24]),
    .Y(_3668_)
);

OAI21X1 _13025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3667_),
    .B(vdd),
    .C(_3668_),
    .Y(_3620_[24])
);

INVX1 _13026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[25]),
    .Y(_3669_)
);

NAND2X1 _13027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [25]),
    .Y(_3670_)
);

OAI21X1 _13028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3669_),
    .B(vdd),
    .C(_3670_),
    .Y(_3620_[25])
);

INVX1 _13029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[26]),
    .Y(_3671_)
);

NAND2X1 _13030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [26]),
    .Y(_3672_)
);

OAI21X1 _13031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3671_),
    .B(vdd),
    .C(_3672_),
    .Y(_3620_[26])
);

INVX1 _13032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[27]),
    .Y(_3673_)
);

NAND2X1 _13033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [27]),
    .Y(_3674_)
);

OAI21X1 _13034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3673_),
    .B(vdd),
    .C(_3674_),
    .Y(_3620_[27])
);

INVX1 _13035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[28]),
    .Y(_3675_)
);

NAND2X1 _13036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [28]),
    .Y(_3676_)
);

OAI21X1 _13037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .B(vdd),
    .C(_3676_),
    .Y(_3620_[28])
);

INVX1 _13038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[29]),
    .Y(_3677_)
);

NAND2X1 _13039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [29]),
    .Y(_3678_)
);

OAI21X1 _13040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3677_),
    .B(vdd),
    .C(_3678_),
    .Y(_3620_[29])
);

INVX1 _13041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[30]),
    .Y(_3679_)
);

NAND2X1 _13042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [30]),
    .Y(_3680_)
);

OAI21X1 _13043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3679_),
    .B(vdd),
    .C(_3680_),
    .Y(_3620_[30])
);

INVX1 _13044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[31]),
    .Y(_3681_)
);

NAND2X1 _13045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(vdd),
    .B(\datapath_1.rd2 [31]),
    .Y(_3682_)
);

OAI21X1 _13046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3681_),
    .B(vdd),
    .C(_3682_),
    .Y(_3620_[31])
);

DFFSR _13047_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_3620_[0]),
    .Q(_2_[0]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _13048_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_3620_[1]),
    .Q(_2_[1]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _13049_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_3620_[2]),
    .Q(_2_[2]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _13050_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_3620_[3]),
    .Q(_2_[3]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _13051_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_3620_[4]),
    .Q(_2_[4]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _13052_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_3620_[5]),
    .Q(_2_[5]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _13053_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_3620_[6]),
    .Q(_2_[6]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _13054_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_3620_[7]),
    .Q(_2_[7]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _13055_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_3620_[8]),
    .Q(_2_[8]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _13056_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_3620_[9]),
    .Q(_2_[9]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _13057_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_3620_[10]),
    .Q(_2_[10]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _13058_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_3620_[11]),
    .Q(_2_[11]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _13059_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_3620_[12]),
    .Q(_2_[12]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _13060_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_3620_[13]),
    .Q(_2_[13]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _13061_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_3620_[14]),
    .Q(_2_[14]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _13062_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_3620_[15]),
    .Q(_2_[15]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _13063_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_3620_[16]),
    .Q(_2_[16]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _13064_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_3620_[17]),
    .Q(_2_[17]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _13065_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_3620_[18]),
    .Q(_2_[18]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _13066_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_3620_[19]),
    .Q(_2_[19]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _13067_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_3620_[20]),
    .Q(_2_[20]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _13068_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_3620_[21]),
    .Q(_2_[21]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _13069_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_3620_[22]),
    .Q(_2_[22]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _13070_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_3620_[23]),
    .Q(_2_[23]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _13071_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_3620_[24]),
    .Q(_2_[24]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _13072_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_3620_[25]),
    .Q(_2_[25]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _13073_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_3620_[26]),
    .Q(_2_[26]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _13074_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_3620_[27]),
    .Q(_2_[27]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _13075_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_3620_[28]),
    .Q(_2_[28]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _13076_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_3620_[29]),
    .Q(_2_[29]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _13077_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_3620_[30]),
    .Q(_2_[30]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _13078_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_3620_[31]),
    .Q(_2_[31]),
    .R(rst_bF$buf68),
    .S(vdd)
);

INVX1 _13079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [0]),
    .Y(_3748_)
);

NAND2X1 _13080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_pcsrc.dout [0]),
    .B(PCEn_bF$buf7),
    .Y(_3749_)
);

OAI21X1 _13081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3748_),
    .B(PCEn_bF$buf6),
    .C(_3749_),
    .Y(_3685_[0])
);

INVX1 _13082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [1]),
    .Y(_3686_)
);

NAND2X1 _13083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [1]),
    .Y(_3687_)
);

OAI21X1 _13084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3686_),
    .B(PCEn_bF$buf4),
    .C(_3687_),
    .Y(_3685_[1])
);

INVX1 _13085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [2]),
    .Y(_3688_)
);

NAND2X1 _13086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [2]),
    .Y(_3689_)
);

OAI21X1 _13087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3688_),
    .B(PCEn_bF$buf2),
    .C(_3689_),
    .Y(_3685_[2])
);

INVX1 _13088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [3]),
    .Y(_3690_)
);

NAND2X1 _13089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [3]),
    .Y(_3691_)
);

OAI21X1 _13090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3690_),
    .B(PCEn_bF$buf0),
    .C(_3691_),
    .Y(_3685_[3])
);

INVX1 _13091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [4]),
    .Y(_3692_)
);

NAND2X1 _13092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [4]),
    .Y(_3693_)
);

OAI21X1 _13093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3692_),
    .B(PCEn_bF$buf6),
    .C(_3693_),
    .Y(_3685_[4])
);

INVX1 _13094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [5]),
    .Y(_3694_)
);

NAND2X1 _13095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [5]),
    .Y(_3695_)
);

OAI21X1 _13096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3694_),
    .B(PCEn_bF$buf4),
    .C(_3695_),
    .Y(_3685_[5])
);

INVX1 _13097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [6]),
    .Y(_3696_)
);

NAND2X1 _13098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [6]),
    .Y(_3697_)
);

OAI21X1 _13099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3696_),
    .B(PCEn_bF$buf2),
    .C(_3697_),
    .Y(_3685_[6])
);

INVX1 _13100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [7]),
    .Y(_3698_)
);

NAND2X1 _13101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [7]),
    .Y(_3699_)
);

OAI21X1 _13102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3698_),
    .B(PCEn_bF$buf0),
    .C(_3699_),
    .Y(_3685_[7])
);

INVX1 _13103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [8]),
    .Y(_3700_)
);

NAND2X1 _13104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [8]),
    .Y(_3701_)
);

OAI21X1 _13105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3700_),
    .B(PCEn_bF$buf6),
    .C(_3701_),
    .Y(_3685_[8])
);

INVX1 _13106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [9]),
    .Y(_3702_)
);

NAND2X1 _13107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [9]),
    .Y(_3703_)
);

OAI21X1 _13108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3702_),
    .B(PCEn_bF$buf4),
    .C(_3703_),
    .Y(_3685_[9])
);

INVX1 _13109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [10]),
    .Y(_3704_)
);

NAND2X1 _13110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [10]),
    .Y(_3705_)
);

OAI21X1 _13111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3704_),
    .B(PCEn_bF$buf2),
    .C(_3705_),
    .Y(_3685_[10])
);

INVX1 _13112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [11]),
    .Y(_3706_)
);

NAND2X1 _13113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [11]),
    .Y(_3707_)
);

OAI21X1 _13114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3706_),
    .B(PCEn_bF$buf0),
    .C(_3707_),
    .Y(_3685_[11])
);

INVX1 _13115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [12]),
    .Y(_3708_)
);

NAND2X1 _13116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [12]),
    .Y(_3709_)
);

OAI21X1 _13117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3708_),
    .B(PCEn_bF$buf6),
    .C(_3709_),
    .Y(_3685_[12])
);

INVX1 _13118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [13]),
    .Y(_3710_)
);

NAND2X1 _13119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [13]),
    .Y(_3711_)
);

OAI21X1 _13120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3710_),
    .B(PCEn_bF$buf4),
    .C(_3711_),
    .Y(_3685_[13])
);

INVX1 _13121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [14]),
    .Y(_3712_)
);

NAND2X1 _13122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [14]),
    .Y(_3713_)
);

OAI21X1 _13123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3712_),
    .B(PCEn_bF$buf2),
    .C(_3713_),
    .Y(_3685_[14])
);

INVX1 _13124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [15]),
    .Y(_3714_)
);

NAND2X1 _13125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [15]),
    .Y(_3715_)
);

OAI21X1 _13126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3714_),
    .B(PCEn_bF$buf0),
    .C(_3715_),
    .Y(_3685_[15])
);

INVX1 _13127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [16]),
    .Y(_3716_)
);

NAND2X1 _13128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [16]),
    .Y(_3717_)
);

OAI21X1 _13129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3716_),
    .B(PCEn_bF$buf6),
    .C(_3717_),
    .Y(_3685_[16])
);

INVX1 _13130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [17]),
    .Y(_3718_)
);

NAND2X1 _13131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [17]),
    .Y(_3719_)
);

OAI21X1 _13132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3718_),
    .B(PCEn_bF$buf4),
    .C(_3719_),
    .Y(_3685_[17])
);

INVX1 _13133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [18]),
    .Y(_3720_)
);

NAND2X1 _13134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [18]),
    .Y(_3721_)
);

OAI21X1 _13135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3720_),
    .B(PCEn_bF$buf2),
    .C(_3721_),
    .Y(_3685_[18])
);

INVX1 _13136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [19]),
    .Y(_3722_)
);

NAND2X1 _13137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [19]),
    .Y(_3723_)
);

OAI21X1 _13138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3722_),
    .B(PCEn_bF$buf0),
    .C(_3723_),
    .Y(_3685_[19])
);

INVX1 _13139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [20]),
    .Y(_3724_)
);

NAND2X1 _13140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [20]),
    .Y(_3725_)
);

OAI21X1 _13141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3724_),
    .B(PCEn_bF$buf6),
    .C(_3725_),
    .Y(_3685_[20])
);

INVX1 _13142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [21]),
    .Y(_3726_)
);

NAND2X1 _13143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [21]),
    .Y(_3727_)
);

OAI21X1 _13144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3726_),
    .B(PCEn_bF$buf4),
    .C(_3727_),
    .Y(_3685_[21])
);

INVX1 _13145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [22]),
    .Y(_3728_)
);

NAND2X1 _13146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [22]),
    .Y(_3729_)
);

OAI21X1 _13147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3728_),
    .B(PCEn_bF$buf2),
    .C(_3729_),
    .Y(_3685_[22])
);

INVX1 _13148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [23]),
    .Y(_3730_)
);

NAND2X1 _13149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [23]),
    .Y(_3731_)
);

OAI21X1 _13150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3730_),
    .B(PCEn_bF$buf0),
    .C(_3731_),
    .Y(_3685_[23])
);

INVX1 _13151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [24]),
    .Y(_3732_)
);

NAND2X1 _13152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [24]),
    .Y(_3733_)
);

OAI21X1 _13153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3732_),
    .B(PCEn_bF$buf6),
    .C(_3733_),
    .Y(_3685_[24])
);

INVX1 _13154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [25]),
    .Y(_3734_)
);

NAND2X1 _13155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [25]),
    .Y(_3735_)
);

OAI21X1 _13156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3734_),
    .B(PCEn_bF$buf4),
    .C(_3735_),
    .Y(_3685_[25])
);

INVX1 _13157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [26]),
    .Y(_3736_)
);

NAND2X1 _13158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [26]),
    .Y(_3737_)
);

OAI21X1 _13159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3736_),
    .B(PCEn_bF$buf2),
    .C(_3737_),
    .Y(_3685_[26])
);

INVX1 _13160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_iord.din0 [27]),
    .Y(_3738_)
);

NAND2X1 _13161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [27]),
    .Y(_3739_)
);

OAI21X1 _13162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3738_),
    .B(PCEn_bF$buf0),
    .C(_3739_),
    .Y(_3685_[27])
);

INVX1 _13163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [28]),
    .Y(_3740_)
);

NAND2X1 _13164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf7),
    .B(\datapath_1.mux_pcsrc.dout [28]),
    .Y(_3741_)
);

OAI21X1 _13165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(PCEn_bF$buf6),
    .C(_3741_),
    .Y(_3685_[28])
);

INVX1 _13166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [29]),
    .Y(_3742_)
);

NAND2X1 _13167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf5),
    .B(\datapath_1.mux_pcsrc.dout [29]),
    .Y(_3743_)
);

OAI21X1 _13168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3742_),
    .B(PCEn_bF$buf4),
    .C(_3743_),
    .Y(_3685_[29])
);

INVX1 _13169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [30]),
    .Y(_3744_)
);

NAND2X1 _13170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf3),
    .B(\datapath_1.mux_pcsrc.dout [30]),
    .Y(_3745_)
);

OAI21X1 _13171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3744_),
    .B(PCEn_bF$buf2),
    .C(_3745_),
    .Y(_3685_[30])
);

INVX1 _13172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [31]),
    .Y(_3746_)
);

NAND2X1 _13173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PCEn_bF$buf1),
    .B(\datapath_1.mux_pcsrc.dout [31]),
    .Y(_3747_)
);

OAI21X1 _13174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3746_),
    .B(PCEn_bF$buf0),
    .C(_3747_),
    .Y(_3685_[31])
);

DFFSR _13175_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_3685_[0]),
    .Q(\datapath_1.mux_iord.din0 [0]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _13176_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_3685_[1]),
    .Q(\datapath_1.mux_iord.din0 [1]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _13177_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_3685_[2]),
    .Q(\datapath_1.mux_iord.din0 [2]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _13178_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_3685_[3]),
    .Q(\datapath_1.mux_iord.din0 [3]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _13179_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_3685_[4]),
    .Q(\datapath_1.mux_iord.din0 [4]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _13180_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_3685_[5]),
    .Q(\datapath_1.mux_iord.din0 [5]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _13181_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_3685_[6]),
    .Q(\datapath_1.mux_iord.din0 [6]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _13182_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_3685_[7]),
    .Q(\datapath_1.mux_iord.din0 [7]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _13183_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_3685_[8]),
    .Q(\datapath_1.mux_iord.din0 [8]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _13184_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_3685_[9]),
    .Q(\datapath_1.mux_iord.din0 [9]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _13185_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_3685_[10]),
    .Q(\datapath_1.mux_iord.din0 [10]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _13186_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_3685_[11]),
    .Q(\datapath_1.mux_iord.din0 [11]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _13187_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_3685_[12]),
    .Q(\datapath_1.mux_iord.din0 [12]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _13188_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_3685_[13]),
    .Q(\datapath_1.mux_iord.din0 [13]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _13189_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_3685_[14]),
    .Q(\datapath_1.mux_iord.din0 [14]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _13190_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_3685_[15]),
    .Q(\datapath_1.mux_iord.din0 [15]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _13191_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_3685_[16]),
    .Q(\datapath_1.mux_iord.din0 [16]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _13192_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_3685_[17]),
    .Q(\datapath_1.mux_iord.din0 [17]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _13193_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_3685_[18]),
    .Q(\datapath_1.mux_iord.din0 [18]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _13194_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_3685_[19]),
    .Q(\datapath_1.mux_iord.din0 [19]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _13195_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_3685_[20]),
    .Q(\datapath_1.mux_iord.din0 [20]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _13196_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_3685_[21]),
    .Q(\datapath_1.mux_iord.din0 [21]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _13197_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_3685_[22]),
    .Q(\datapath_1.mux_iord.din0 [22]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _13198_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_3685_[23]),
    .Q(\datapath_1.mux_iord.din0 [23]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _13199_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_3685_[24]),
    .Q(\datapath_1.mux_iord.din0 [24]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _13200_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_3685_[25]),
    .Q(\datapath_1.mux_iord.din0 [25]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _13201_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_3685_[26]),
    .Q(\datapath_1.mux_iord.din0 [26]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _13202_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_3685_[27]),
    .Q(\datapath_1.mux_iord.din0 [27]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _13203_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_3685_[28]),
    .Q(\datapath_1.PCJump [28]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _13204_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_3685_[29]),
    .Q(\datapath_1.PCJump [29]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _13205_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_3685_[30]),
    .Q(\datapath_1.PCJump [30]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _13206_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_3685_[31]),
    .Q(\datapath_1.PCJump [31]),
    .R(rst_bF$buf36),
    .S(vdd)
);

INVX4 _13207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .Y(_3750_)
);

INVX2 _13208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [0]),
    .Y(_3751_)
);

NOR2X1 _13209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .B(_3751_),
    .Y(_3752_)
);

NAND2X1 _13210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_3753_)
);

INVX2 _13211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3753_),
    .Y(_3754_)
);

AND2X2 _13212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3754_),
    .Y(_3755_)
);

INVX2 _13213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3755_),
    .Y(_3756_)
);

INVX1 _13214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .Y(_3757_)
);

NOR2X1 _13215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [2]),
    .B(_3757_),
    .Y(_3758_)
);

NAND2X1 _13216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_3759_)
);

INVX1 _13217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3759_),
    .Y(_3760_)
);

NAND2X1 _13218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3760_),
    .B(_3758_),
    .Y(_3761_)
);

AOI21X1 _13219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3761_),
    .B(_3756_),
    .C(_3750_),
    .Y(_3762_)
);

INVX2 _13220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .Y(_3763_)
);

NOR2X1 _13221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [0]),
    .B(_3763_),
    .Y(_3764_)
);

NOR2X1 _13222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3764_),
    .Y(_3765_)
);

NAND2X1 _13223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3758_),
    .Y(_3766_)
);

NAND2X1 _13224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3754_),
    .Y(_3767_)
);

OAI22X1 _13225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3767_),
    .C(_3765_),
    .D(_3766_),
    .Y(_3768_)
);

NOR2X1 _13226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3768_),
    .B(_3762_),
    .Y(_3769_)
);

NOR2X1 _13227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .Y(_3770_)
);

INVX1 _13228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [2]),
    .Y(_3771_)
);

NOR2X1 _13229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .B(_3771_),
    .Y(_3772_)
);

INVX2 _13230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3772_),
    .Y(_3773_)
);

NAND2X1 _13231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3770_),
    .B(_3758_),
    .Y(_3774_)
);

OAI21X1 _13232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3773_),
    .B(_3770_),
    .C(_3774_),
    .Y(_3775_)
);

INVX2 _13233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3770_),
    .Y(_3776_)
);

NOR2X1 _13234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .B(\datapath_1.a3 [2]),
    .Y(_3777_)
);

OAI21X1 _13235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .B(\datapath_1.a3 [0]),
    .C(_3777_),
    .Y(_3778_)
);

OAI21X1 _13236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3773_),
    .B(_3776_),
    .C(_3778_),
    .Y(_3779_)
);

OAI21X1 _13237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3775_),
    .B(_3779_),
    .C(\datapath_1.a3 [4]),
    .Y(_3780_)
);

NAND2X1 _13238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3780_),
    .B(_3769_),
    .Y(_3781_)
);

NOR2X1 _13239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3759_),
    .B(_3753_),
    .Y(_3782_)
);

NAND2X1 _13240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3777_),
    .Y(_3783_)
);

NOR2X1 _13241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3776_),
    .B(_3783_),
    .Y(_3784_)
);

AOI21X1 _13242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3750_),
    .B(_3782_),
    .C(_3784_),
    .Y(_3785_)
);

NAND2X1 _13243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3750_),
    .B(_3754_),
    .Y(_3786_)
);

OR2X2 _13244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3765_),
    .B(_3786_),
    .Y(_3787_)
);

AND2X2 _13245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3787_),
    .B(_3785_),
    .Y(_3788_)
);

NAND2X1 _13246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .B(_3771_),
    .Y(_3789_)
);

NOR2X1 _13247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3789_),
    .Y(_3790_)
);

INVX1 _13248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3790_),
    .Y(_3791_)
);

NOR2X1 _13249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3765_),
    .B(_3791_),
    .Y(_3792_)
);

NAND2X1 _13250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3770_),
    .B(_3754_),
    .Y(_3793_)
);

AOI21X1 _13251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3793_),
    .B(_3761_),
    .C(\datapath_1.a3 [4]),
    .Y(_3794_)
);

NOR2X1 _13252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3794_),
    .B(_3792_),
    .Y(_3795_)
);

NAND2X1 _13253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3788_),
    .B(_3795_),
    .Y(_3796_)
);

INVX4 _13254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite_bF$buf7),
    .Y(_3797_)
);

NAND2X1 _13255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(RegWrite_bF$buf6),
    .Y(_3798_)
);

INVX2 _13256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3777_),
    .Y(_3799_)
);

NAND2X1 _13257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3770_),
    .B(_3772_),
    .Y(_3800_)
);

OAI21X1 _13258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3759_),
    .B(_3799_),
    .C(_3800_),
    .Y(_3801_)
);

OAI21X1 _13259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3801_),
    .B(_3797_),
    .C(_3798_),
    .Y(_3802_)
);

NAND2X1 _13260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3750_),
    .B(_3775_),
    .Y(_3803_)
);

NOR2X1 _13261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3799_),
    .Y(_3804_)
);

NAND2X1 _13262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3751_),
    .B(_3804_),
    .Y(_3805_)
);

NAND3X1 _13263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3803_),
    .B(_3805_),
    .C(_3802_),
    .Y(_3806_)
);

OR2X2 _13264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3806_),
    .Y(_3807_)
);

NOR2X1 _13265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3807_),
    .Y(\datapath_1.regfile_1.regEn [1])
);

AOI22X1 _13266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_3804_),
    .C(_3775_),
    .D(_3750_),
    .Y(_3808_)
);

NAND2X1 _13267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .B(_3808_),
    .Y(_3809_)
);

OR2X2 _13268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3809_),
    .Y(_3810_)
);

NOR2X1 _13269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3810_),
    .Y(\datapath_1.regfile_1.regEn [2])
);

INVX1 _13270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3811_)
);

INVX2 _13271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3764_),
    .Y(_3812_)
);

NOR2X1 _13272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3799_),
    .B(_3812_),
    .Y(_3813_)
);

OAI21X1 _13273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3813_),
    .B(_3811_),
    .C(_3750_),
    .Y(_3814_)
);

NAND3X1 _13274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite_bF$buf5),
    .B(_3814_),
    .C(_3808_),
    .Y(_3815_)
);

OR2X2 _13275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3815_),
    .Y(_3816_)
);

NOR2X1 _13276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3816_),
    .Y(\datapath_1.regfile_1.regEn [3])
);

NOR2X1 _13277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3797_),
    .B(_3804_),
    .Y(_3817_)
);

NAND2X1 _13278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3817_),
    .B(_3803_),
    .Y(_3818_)
);

OR2X2 _13279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3818_),
    .Y(_3819_)
);

NOR2X1 _13280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3819_),
    .Y(\datapath_1.regfile_1.regEn [4])
);

OAI21X1 _13281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3773_),
    .B(_3759_),
    .C(_3774_),
    .Y(_3820_)
);

NAND2X1 _13282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3750_),
    .B(_3820_),
    .Y(_3821_)
);

NOR2X1 _13283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3812_),
    .B(_3773_),
    .Y(_3822_)
);

OAI21X1 _13284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3822_),
    .B(_3811_),
    .C(_3750_),
    .Y(_3823_)
);

NAND3X1 _13285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3821_),
    .B(_3817_),
    .C(_3823_),
    .Y(_3824_)
);

OR2X2 _13286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3824_),
    .Y(_3825_)
);

NOR2X1 _13287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3825_),
    .Y(\datapath_1.regfile_1.regEn [5])
);

NAND2X1 _13288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_3772_),
    .Y(_3826_)
);

OR2X2 _13289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3826_),
    .B(\datapath_1.a3 [4]),
    .Y(_3827_)
);

AND2X2 _13290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3827_),
    .B(_3817_),
    .Y(_3828_)
);

NAND2X1 _13291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3821_),
    .B(_3828_),
    .Y(_3829_)
);

OR2X2 _13292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3829_),
    .Y(_3830_)
);

NOR2X1 _13293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3830_),
    .Y(\datapath_1.regfile_1.regEn [6])
);

INVX1 _13294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3774_),
    .Y(_3831_)
);

OAI21X1 _13295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3822_),
    .B(_3831_),
    .C(_3750_),
    .Y(_3832_)
);

NAND2X1 _13296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3832_),
    .B(_3828_),
    .Y(_3833_)
);

NOR3X1 _13297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3833_),
    .C(_3781_),
    .Y(\datapath_1.regfile_1.regEn [7])
);

OAI21X1 _13298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3757_),
    .B(_3797_),
    .C(_3798_),
    .Y(_3834_)
);

INVX2 _13299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3834_),
    .Y(_3835_)
);

OR2X2 _13300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .B(_3835_),
    .Y(_3836_)
);

NOR2X1 _13301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3836_),
    .Y(\datapath_1.regfile_1.regEn [8])
);

OAI21X1 _13302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3764_),
    .C(_3754_),
    .Y(_3837_)
);

OAI21X1 _13303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3837_),
    .C(_3785_),
    .Y(_3838_)
);

NOR2X1 _13304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3794_),
    .B(_3838_),
    .Y(_3839_)
);

OAI21X1 _13305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [0]),
    .B(_3791_),
    .C(_3839_),
    .Y(_3840_)
);

NOR3X1 _13306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3835_),
    .C(_3840_),
    .Y(\datapath_1.regfile_1.regEn [9])
);

AOI21X1 _13307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_3790_),
    .C(_3835_),
    .Y(_3841_)
);

NAND2X1 _13308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3841_),
    .B(_3839_),
    .Y(_3842_)
);

NOR2X1 _13309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3842_),
    .Y(\datapath_1.regfile_1.regEn [10])
);

NOR2X1 _13310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3789_),
    .B(_3812_),
    .Y(_3843_)
);

INVX1 _13311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3793_),
    .Y(_3844_)
);

OAI21X1 _13312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3843_),
    .B(_3844_),
    .C(_3750_),
    .Y(_3845_)
);

NAND3X1 _13313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3841_),
    .B(_3845_),
    .C(_3788_),
    .Y(_3846_)
);

NOR2X1 _13314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3846_),
    .B(_3781_),
    .Y(\datapath_1.regfile_1.regEn [11])
);

NAND2X1 _13315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3834_),
    .B(_3785_),
    .Y(_3847_)
);

NOR2X1 _13316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3790_),
    .B(_3847_),
    .Y(_3848_)
);

OAI21X1 _13317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3837_),
    .C(_3848_),
    .Y(_3849_)
);

NOR2X1 _13318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3849_),
    .Y(\datapath_1.regfile_1.regEn [12])
);

OAI21X1 _13319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [0]),
    .B(_3786_),
    .C(_3848_),
    .Y(_3850_)
);

NOR2X1 _13320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3850_),
    .Y(\datapath_1.regfile_1.regEn [13])
);

NOR2X1 _13321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .B(_3753_),
    .Y(_3851_)
);

INVX1 _13322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3851_),
    .Y(_3852_)
);

OAI21X1 _13323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3852_),
    .C(_3848_),
    .Y(_3853_)
);

NOR2X1 _13324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3853_),
    .Y(\datapath_1.regfile_1.regEn [14])
);

NAND2X1 _13325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3750_),
    .B(_3782_),
    .Y(_3854_)
);

NOR2X1 _13326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3797_),
    .B(_3854_),
    .Y(\datapath_1.regfile_1.regEn [15])
);

AND2X2 _13327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3784_),
    .B(RegWrite_bF$buf4),
    .Y(\datapath_1.regfile_1.regEn [16])
);

NAND2X1 _13328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3777_),
    .B(_3752_),
    .Y(_3855_)
);

NOR2X1 _13329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3855_),
    .Y(\datapath_1.regfile_1.regEn [17])
);

INVX2 _13330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .Y(_3856_)
);

AND2X2 _13331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3813_),
    .B(_3856_),
    .Y(\datapath_1.regfile_1.regEn [18])
);

NAND2X1 _13332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3777_),
    .B(_3760_),
    .Y(_3857_)
);

NOR2X1 _13333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3857_),
    .Y(\datapath_1.regfile_1.regEn [19])
);

NOR2X1 _13334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3800_),
    .Y(\datapath_1.regfile_1.regEn [20])
);

INVX1 _13335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3769_),
    .Y(_3858_)
);

AOI21X1 _13336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3751_),
    .B(_3772_),
    .C(_3820_),
    .Y(_3859_)
);

NAND3X1 _13337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3799_),
    .B(_3856_),
    .C(_3859_),
    .Y(_3860_)
);

NOR2X1 _13338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3860_),
    .B(_3858_),
    .Y(\datapath_1.regfile_1.regEn [21])
);

NAND2X1 _13339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3822_),
    .Y(_3861_)
);

NOR2X1 _13340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3797_),
    .B(_3861_),
    .Y(\datapath_1.regfile_1.regEn [22])
);

OAI21X1 _13341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3776_),
    .B(_3789_),
    .C(_3856_),
    .Y(_3862_)
);

NAND3X1 _13342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_3826_),
    .C(_3861_),
    .Y(_3863_)
);

NOR2X1 _13343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3862_),
    .B(_3863_),
    .Y(_3864_)
);

AND2X2 _13344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3864_),
    .B(_3769_),
    .Y(\datapath_1.regfile_1.regEn [23])
);

NOR2X1 _13345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3774_),
    .Y(\datapath_1.regfile_1.regEn [24])
);

INVX1 _13346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3843_),
    .Y(_3865_)
);

AOI21X1 _13347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .B(_3865_),
    .C(_3750_),
    .Y(_3866_)
);

OR2X2 _13348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3866_),
    .B(_3762_),
    .Y(_3867_)
);

INVX1 _13349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3862_),
    .Y(_3868_)
);

OAI21X1 _13350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3767_),
    .C(_3868_),
    .Y(_3869_)
);

NOR2X1 _13351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3869_),
    .B(_3867_),
    .Y(\datapath_1.regfile_1.regEn [25])
);

NOR2X1 _13352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3865_),
    .Y(\datapath_1.regfile_1.regEn [26])
);

NAND3X1 _13353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [3]),
    .B(_3856_),
    .C(_3767_),
    .Y(_3870_)
);

OR2X2 _13354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3870_),
    .B(_3843_),
    .Y(_3871_)
);

OAI21X1 _13355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3766_),
    .B(\datapath_1.a3 [1]),
    .C(_3756_),
    .Y(_3872_)
);

NOR2X1 _13356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3872_),
    .B(_3871_),
    .Y(\datapath_1.regfile_1.regEn [27])
);

NAND2X1 _13357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [4]),
    .B(_3782_),
    .Y(_3873_)
);

NAND2X1 _13358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RegWrite_bF$buf3),
    .B(_3873_),
    .Y(_3874_)
);

INVX1 _13359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3767_),
    .Y(_3875_)
);

OAI21X1 _13360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3765_),
    .B(_3753_),
    .C(_3875_),
    .Y(_3876_)
);

NOR2X1 _13361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3874_),
    .B(_3876_),
    .Y(\datapath_1.regfile_1.regEn [28])
);

NOR2X1 _13362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3756_),
    .Y(\datapath_1.regfile_1.regEn [29])
);

NAND2X1 _13363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.a3 [1]),
    .B(_3875_),
    .Y(_3877_)
);

NOR2X1 _13364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3874_),
    .B(_3877_),
    .Y(\datapath_1.regfile_1.regEn [30])
);

NOR2X1 _13365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3797_),
    .B(_3873_),
    .Y(\datapath_1.regfile_1.regEn [31])
);

INVX1 _13366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [19]),
    .Y(_3878_)
);

AND2X2 _13367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3878_),
    .B(\datapath_1.PCJump [18]),
    .Y(_3879_)
);

AND2X2 _13368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3880_)
);

NAND3X1 _13369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3880_),
    .C(_3879_),
    .Y(_3881_)
);

INVX8 _13370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3881_),
    .Y(_3882_)
);

NOR2X1 _13371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [18]),
    .B(_3878_),
    .Y(_3883_)
);

NAND3X1 _13372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3880_),
    .C(_3883_),
    .Y(_3884_)
);

INVX8 _13373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf3),
    .Y(_3885_)
);

AOI22X1 _13374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [0]),
    .B(_3885_),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [0]),
    .Y(_3886_)
);

INVX1 _13375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [20]),
    .Y(_3887_)
);

NOR2X1 _13376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .B(_3887_),
    .Y(_3888_)
);

NOR3X1 _13377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(\datapath_1.PCJump [19]),
    .C(\datapath_1.PCJump [18]),
    .Y(_3889_)
);

NAND2X1 _13378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3889_),
    .B(_3888_),
    .Y(_3890_)
);

INVX8 _13379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3890_),
    .Y(_3891_)
);

NOR2X1 _13380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3892_)
);

NAND3X1 _13381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3892_),
    .C(_3880_),
    .Y(_3893_)
);

INVX8 _13382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893__bF$buf3),
    .Y(_3894_)
);

AOI22X1 _13383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .B(_3894_),
    .C(_3891__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_3895_)
);

INVX1 _13384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_3896_)
);

INVX1 _13385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_3897_)
);

INVX4 _13386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .Y(_3898_)
);

NAND2X1 _13387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3899_)
);

NAND2X1 _13388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3900_)
);

NOR2X1 _13389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3899_),
    .B(_3900_),
    .Y(_3901_)
);

NAND2X1 _13390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3901_),
    .Y(_3902_)
);

AND2X2 _13391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [19]),
    .B(\datapath_1.PCJump [18]),
    .Y(_3903_)
);

NOR2X1 _13392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .B(\datapath_1.PCJump [20]),
    .Y(_3904_)
);

NAND3X1 _13393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3904_),
    .C(_3903_),
    .Y(_3905_)
);

OAI22X1 _13394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905__bF$buf3),
    .B(_3896_),
    .C(_3902__bF$buf3),
    .D(_3897_),
    .Y(_3906_)
);

INVX1 _13395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_3907_)
);

INVX1 _13396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_3908_)
);

NAND3X1 _13397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3883_),
    .C(_3888_),
    .Y(_3909_)
);

NAND2X1 _13398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3880_),
    .B(_3889_),
    .Y(_3910_)
);

OAI22X1 _13399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3907_),
    .B(_3910_),
    .C(_3909_),
    .D(_3908_),
    .Y(_3911_)
);

NOR2X1 _13400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3906_),
    .B(_3911_),
    .Y(_3912_)
);

NAND3X1 _13401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3886_),
    .B(_3895_),
    .C(_3912_),
    .Y(_3913_)
);

INVX1 _13402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_3914_)
);

INVX1 _13403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_3915_)
);

NAND3X1 _13404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3903_),
    .C(_3888_),
    .Y(_3916_)
);

AND2X2 _13405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3892_),
    .B(\datapath_1.PCJump_22_bF$buf1 ),
    .Y(_3917_)
);

INVX1 _13406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [21]),
    .Y(_3918_)
);

NOR2X1 _13407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [20]),
    .B(_3918_),
    .Y(_3919_)
);

NAND2X1 _13408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3919_),
    .B(_3917_),
    .Y(_3920_)
);

OAI22X1 _13409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3915_),
    .B(_3916_),
    .C(_3920_),
    .D(_3914_),
    .Y(_3921_)
);

INVX1 _13410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [0]),
    .Y(_3922_)
);

INVX1 _13411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_3923_)
);

NAND2X1 _13412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3888_),
    .B(_3917_),
    .Y(_3924_)
);

NAND2X1 _13413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3901_),
    .Y(_3925_)
);

OAI22X1 _13414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3922_),
    .B(_3925_),
    .C(_3924__bF$buf3),
    .D(_3923_),
    .Y(_3926_)
);

NOR2X1 _13415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3926_),
    .B(_3921_),
    .Y(_3927_)
);

INVX1 _13416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_3928_)
);

INVX1 _13417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_3929_)
);

NAND2X1 _13418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3904_),
    .B(_3889_),
    .Y(_3930_)
);

NAND2X1 _13419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3889_),
    .B(_3919_),
    .Y(_3931_)
);

OAI22X1 _13420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3928_),
    .B(_3930__bF$buf3),
    .C(_3931__bF$buf3),
    .D(_3929_),
    .Y(_3932_)
);

INVX1 _13421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_3933_)
);

INVX1 _13422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_3934_)
);

NAND3X1 _13423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3883_),
    .C(_3919_),
    .Y(_3935_)
);

NAND3X1 _13424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3892_),
    .C(_3904_),
    .Y(_3936_)
);

OAI22X1 _13425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3933_),
    .B(_3936__bF$buf4),
    .C(_3935__bF$buf4),
    .D(_3934_),
    .Y(_3937_)
);

NOR2X1 _13426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3932_),
    .B(_3937_),
    .Y(_3938_)
);

NAND2X1 _13427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3938_),
    .B(_3927_),
    .Y(_3939_)
);

NOR2X1 _13428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3913_),
    .B(_3939_),
    .Y(_3940_)
);

NAND3X1 _13429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3904_),
    .C(_3903_),
    .Y(_3941_)
);

INVX8 _13430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3941_),
    .Y(_3942_)
);

INVX1 _13431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [0]),
    .Y(_3943_)
);

NAND3X1 _13432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3883_),
    .C(_3919_),
    .Y(_3944_)
);

NOR2X1 _13433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3943_),
    .B(_3944__bF$buf4),
    .Y(_3945_)
);

AOI21X1 _13434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .B(_3942__bF$buf3),
    .C(_3945_),
    .Y(_3946_)
);

NAND3X1 _13435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3903_),
    .C(_3888_),
    .Y(_3947_)
);

INVX8 _13436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf3),
    .Y(_3948_)
);

NAND3X1 _13437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3903_),
    .C(_3919_),
    .Y(_3949_)
);

INVX8 _13438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .Y(_3950_)
);

AOI22X1 _13439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [0]),
    .C(\datapath_1.regfile_1.regOut[11] [0]),
    .D(_3950__bF$buf3),
    .Y(_3951_)
);

INVX1 _13440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_3952_)
);

INVX1 _13441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_3953_)
);

NAND3X1 _13442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3888_),
    .C(_3879_),
    .Y(_3954_)
);

NAND3X1 _13443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3883_),
    .C(_3888_),
    .Y(_3955_)
);

OAI22X1 _13444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3952_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf4),
    .D(_3953_),
    .Y(_3956_)
);

INVX1 _13445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_3957_)
);

INVX1 _13446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_3958_)
);

NAND3X1 _13447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3904_),
    .C(_3879_),
    .Y(_3959_)
);

NAND3X1 _13448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3904_),
    .C(_3883_),
    .Y(_3960_)
);

OAI22X1 _13449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .B(_3960_),
    .C(_3959_),
    .D(_3957_),
    .Y(_3961_)
);

NOR2X1 _13450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .B(_3956_),
    .Y(_3962_)
);

NAND3X1 _13451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3946_),
    .B(_3951_),
    .C(_3962_),
    .Y(_3963_)
);

INVX1 _13452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [0]),
    .Y(_3964_)
);

INVX1 _13453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_3965_)
);

NAND3X1 _13454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf3 ),
    .B(_3919_),
    .C(_3879_),
    .Y(_3966_)
);

NAND3X1 _13455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf2 ),
    .B(_3903_),
    .C(_3919_),
    .Y(_3967_)
);

OAI22X1 _13456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf3),
    .B(_3964_),
    .C(_3966__bF$buf3),
    .D(_3965_),
    .Y(_3968_)
);

INVX1 _13457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_3969_)
);

INVX1 _13458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_3970_)
);

NAND3X1 _13459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3919_),
    .C(_3879_),
    .Y(_3971_)
);

NAND3X1 _13460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf1 ),
    .B(_3904_),
    .C(_3883_),
    .Y(_3972_)
);

OAI22X1 _13461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972__bF$buf3),
    .B(_3969_),
    .C(_3971__bF$buf4),
    .D(_3970_),
    .Y(_3973_)
);

NOR2X1 _13462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3968_),
    .B(_3973_),
    .Y(_3974_)
);

INVX1 _13463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_3975_)
);

INVX1 _13464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_3976_)
);

NAND3X1 _13465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3888_),
    .C(_3879_),
    .Y(_3977_)
);

NAND3X1 _13466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3880_),
    .C(_3879_),
    .Y(_3978_)
);

OAI22X1 _13467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_3975_),
    .C(_3977__bF$buf4),
    .D(_3976_),
    .Y(_3979_)
);

INVX1 _13468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_3980_)
);

INVX1 _13469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_3981_)
);

NAND3X1 _13470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3880_),
    .C(_3883_),
    .Y(_3982_)
);

NAND3X1 _13471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_22_bF$buf0 ),
    .B(_3904_),
    .C(_3879_),
    .Y(_3983_)
);

OAI22X1 _13472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3981_),
    .B(_3982__bF$buf3),
    .C(_3983__bF$buf4),
    .D(_3980_),
    .Y(_3984_)
);

NOR2X1 _13473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3984_),
    .B(_3979_),
    .Y(_3985_)
);

NAND2X1 _13474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .B(_3985_),
    .Y(_3986_)
);

NOR2X1 _13475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3986_),
    .B(_3963_),
    .Y(_3987_)
);

AOI21X1 _13476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3940_),
    .B(_3987_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [0])
);

INVX1 _13477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_3988_)
);

INVX1 _13478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_3989_)
);

OAI22X1 _13479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3989_),
    .B(_3949_),
    .C(_3983__bF$buf3),
    .D(_3988_),
    .Y(_3990_)
);

INVX1 _13480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_3991_)
);

INVX1 _13481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_3992_)
);

OAI22X1 _13482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3991_),
    .B(_3936__bF$buf3),
    .C(_3935__bF$buf3),
    .D(_3992_),
    .Y(_3993_)
);

NOR2X1 _13483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3993_),
    .B(_3990_),
    .Y(_3994_)
);

INVX8 _13484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3925_),
    .Y(_3995_)
);

AOI22X1 _13485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .B(_3995__bF$buf4),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_3996_)
);

INVX8 _13486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3959_),
    .Y(_3997_)
);

INVX8 _13487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3960_),
    .Y(_3998_)
);

AOI22X1 _13488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .B(_3998__bF$buf3),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_3999_)
);

NAND3X1 _13489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3996_),
    .B(_3999_),
    .C(_3994_),
    .Y(_4000_)
);

INVX8 _13490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3909_),
    .Y(_4001_)
);

INVX1 _13491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_4002_)
);

NOR2X1 _13492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4002_),
    .B(_3977__bF$buf3),
    .Y(_4003_)
);

AOI21X1 _13493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .B(_4001__bF$buf3),
    .C(_4003_),
    .Y(_4004_)
);

INVX8 _13494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3910_),
    .Y(_4005_)
);

AOI22X1 _13495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3942__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[3] [1]),
    .C(\datapath_1.regfile_1.regOut[12] [1]),
    .D(_4005__bF$buf3),
    .Y(_4006_)
);

INVX1 _13496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_4007_)
);

INVX1 _13497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_4008_)
);

OAI22X1 _13498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(_3930__bF$buf2),
    .C(_3967__bF$buf2),
    .D(_4008_),
    .Y(_4009_)
);

INVX1 _13499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_4010_)
);

INVX1 _13500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_4011_)
);

OAI22X1 _13501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4011_),
    .B(_3902__bF$buf2),
    .C(_3954__bF$buf3),
    .D(_4010_),
    .Y(_4012_)
);

NOR2X1 _13502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4009_),
    .B(_4012_),
    .Y(_4013_)
);

NAND3X1 _13503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4004_),
    .B(_4006_),
    .C(_4013_),
    .Y(_4014_)
);

NOR2X1 _13504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4014_),
    .B(_4000_),
    .Y(_4015_)
);

INVX1 _13505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_4016_)
);

INVX1 _13506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_4017_)
);

OAI22X1 _13507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4017_),
    .B(_3971__bF$buf3),
    .C(_3924__bF$buf2),
    .D(_4016_),
    .Y(_4018_)
);

INVX1 _13508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_4019_)
);

INVX1 _13509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_4020_)
);

OAI22X1 _13510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4020_),
    .B(_3972__bF$buf2),
    .C(_3920_),
    .D(_4019_),
    .Y(_4021_)
);

NOR2X1 _13511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4018_),
    .B(_4021_),
    .Y(_4022_)
);

INVX1 _13512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_4023_)
);

INVX1 _13513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_4024_)
);

OAI22X1 _13514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3890_),
    .B(_4024_),
    .C(_4023_),
    .D(_3931__bF$buf2),
    .Y(_4025_)
);

INVX1 _13515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_4026_)
);

INVX1 _13516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_4027_)
);

OAI22X1 _13517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4027_),
    .B(_3905__bF$buf2),
    .C(_3955__bF$buf3),
    .D(_4026_),
    .Y(_4028_)
);

NOR2X1 _13518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4025_),
    .B(_4028_),
    .Y(_4029_)
);

NAND2X1 _13519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4029_),
    .B(_4022_),
    .Y(_4030_)
);

INVX1 _13520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_4031_)
);

INVX1 _13521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_4032_)
);

OAI22X1 _13522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4031_),
    .B(_3982__bF$buf2),
    .C(_3978_),
    .D(_4032_),
    .Y(_4033_)
);

INVX1 _13523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [1]),
    .Y(_4034_)
);

INVX1 _13524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_4035_)
);

OAI22X1 _13525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf2),
    .B(_4035_),
    .C(_3944__bF$buf3),
    .D(_4034_),
    .Y(_4036_)
);

NOR2X1 _13526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4036_),
    .B(_4033_),
    .Y(_4037_)
);

INVX8 _13527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .Y(_4038_)
);

AOI22X1 _13528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .B(_3894_),
    .C(_4038__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_4039_)
);

INVX8 _13529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3966__bF$buf2),
    .Y(_4040_)
);

AOI22X1 _13530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .B(_3885_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_4041_)
);

NAND3X1 _13531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4039_),
    .B(_4041_),
    .C(_4037_),
    .Y(_4042_)
);

NOR2X1 _13532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4030_),
    .B(_4042_),
    .Y(_4043_)
);

AOI21X1 _13533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4043_),
    .B(_4015_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [1])
);

INVX1 _13534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_4044_)
);

INVX1 _13535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_4045_)
);

OAI22X1 _13536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4044_),
    .B(_3910_),
    .C(_3935__bF$buf2),
    .D(_4045_),
    .Y(_4046_)
);

INVX1 _13537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [2]),
    .Y(_4047_)
);

INVX1 _13538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_4048_)
);

OAI22X1 _13539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf1),
    .B(_4047_),
    .C(_4048_),
    .D(_3902__bF$buf1),
    .Y(_4049_)
);

NOR2X1 _13540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4049_),
    .B(_4046_),
    .Y(_4050_)
);

INVX8 _13541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .Y(_4051_)
);

AOI22X1 _13542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .B(_3891__bF$buf2),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_4052_)
);

AOI22X1 _13543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .B(_3942__bF$buf1),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_4053_)
);

NAND3X1 _13544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4052_),
    .B(_4053_),
    .C(_4050_),
    .Y(_4054_)
);

INVX1 _13545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_4055_)
);

INVX1 _13546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_4056_)
);

OAI22X1 _13547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf1),
    .B(_4055_),
    .C(_3971__bF$buf2),
    .D(_4056_),
    .Y(_4057_)
);

INVX1 _13548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_4058_)
);

INVX1 _13549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_4059_)
);

OAI22X1 _13550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4058_),
    .B(_3930__bF$buf1),
    .C(_3954__bF$buf2),
    .D(_4059_),
    .Y(_4060_)
);

NOR2X1 _13551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4057_),
    .B(_4060_),
    .Y(_4061_)
);

INVX1 _13552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [2]),
    .Y(_4062_)
);

INVX1 _13553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_4063_)
);

OAI22X1 _13554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3881_),
    .B(_4062_),
    .C(_3966__bF$buf1),
    .D(_4063_),
    .Y(_4064_)
);

INVX1 _13555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_4065_)
);

INVX1 _13556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_4066_)
);

OAI22X1 _13557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4065_),
    .B(_3955__bF$buf2),
    .C(_3924__bF$buf1),
    .D(_4066_),
    .Y(_4067_)
);

NOR2X1 _13558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4064_),
    .B(_4067_),
    .Y(_4068_)
);

NAND2X1 _13559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4061_),
    .B(_4068_),
    .Y(_4069_)
);

NOR2X1 _13560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4069_),
    .B(_4054_),
    .Y(_4070_)
);

INVX1 _13561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [2]),
    .Y(_4071_)
);

INVX1 _13562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_4072_)
);

OAI22X1 _13563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4071_),
    .B(_3893__bF$buf2),
    .C(_3972__bF$buf1),
    .D(_4072_),
    .Y(_4073_)
);

INVX1 _13564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_4074_)
);

INVX1 _13565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_4075_)
);

OAI22X1 _13566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4074_),
    .B(_3905__bF$buf1),
    .C(_3909_),
    .D(_4075_),
    .Y(_4076_)
);

NOR2X1 _13567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4073_),
    .B(_4076_),
    .Y(_4077_)
);

AOI22X1 _13568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .C(\datapath_1.regfile_1.regOut[31] [2]),
    .D(_3995__bF$buf3),
    .Y(_4078_)
);

INVX8 _13569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3920_),
    .Y(_4079_)
);

AOI22X1 _13570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .B(_4038__bF$buf2),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_4080_)
);

NAND3X1 _13571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4078_),
    .B(_4080_),
    .C(_4077_),
    .Y(_4081_)
);

INVX1 _13572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [2]),
    .Y(_4082_)
);

INVX1 _13573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_4083_)
);

OAI22X1 _13574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4083_),
    .B(_3936__bF$buf2),
    .C(_3944__bF$buf2),
    .D(_4082_),
    .Y(_4084_)
);

INVX1 _13575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_4085_)
);

INVX1 _13576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_4086_)
);

OAI22X1 _13577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf2),
    .B(_4085_),
    .C(_3977__bF$buf2),
    .D(_4086_),
    .Y(_4087_)
);

NOR2X1 _13578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4084_),
    .B(_4087_),
    .Y(_4088_)
);

AOI22X1 _13579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [2]),
    .C(\datapath_1.regfile_1.regOut[2] [2]),
    .D(_3998__bF$buf2),
    .Y(_4089_)
);

INVX8 _13580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931__bF$buf1),
    .Y(_4090_)
);

AOI22X1 _13581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .B(_4090_),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_4091_)
);

NAND3X1 _13582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4089_),
    .B(_4091_),
    .C(_4088_),
    .Y(_4092_)
);

NOR2X1 _13583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4092_),
    .Y(_4093_)
);

AOI21X1 _13584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4070_),
    .B(_4093_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [2])
);

INVX1 _13585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_4094_)
);

INVX1 _13586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_4095_)
);

OAI22X1 _13587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf1),
    .B(_4095_),
    .C(_3909_),
    .D(_4094_),
    .Y(_4096_)
);

INVX1 _13588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [3]),
    .Y(_4097_)
);

INVX1 _13589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_4098_)
);

OAI22X1 _13590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944__bF$buf1),
    .B(_4097_),
    .C(_4098_),
    .D(_3955__bF$buf1),
    .Y(_4099_)
);

NOR2X1 _13591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4096_),
    .B(_4099_),
    .Y(_4100_)
);

AOI22X1 _13592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[11] [3]),
    .C(\datapath_1.regfile_1.regOut[2] [3]),
    .D(_3998__bF$buf1),
    .Y(_4101_)
);

AND2X2 _13593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3889_),
    .B(_3904_),
    .Y(_4102_)
);

AOI22X1 _13594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .B(_4102_),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_4103_)
);

NAND3X1 _13595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4101_),
    .B(_4103_),
    .C(_4100_),
    .Y(_4104_)
);

INVX1 _13596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_4105_)
);

INVX1 _13597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_4106_)
);

OAI22X1 _13598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4106_),
    .B(_3936__bF$buf1),
    .C(_3966__bF$buf0),
    .D(_4105_),
    .Y(_4107_)
);

INVX1 _13599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_4108_)
);

INVX1 _13600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_4109_)
);

OAI22X1 _13601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4108_),
    .B(_3905__bF$buf0),
    .C(_3977__bF$buf1),
    .D(_4109_),
    .Y(_4110_)
);

NOR2X1 _13602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4110_),
    .B(_4107_),
    .Y(_4111_)
);

INVX1 _13603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_4112_)
);

NOR2X1 _13604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4112_),
    .B(_3935__bF$buf1),
    .Y(_4113_)
);

AOI21X1 _13605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .B(_3894_),
    .C(_4113_),
    .Y(_4114_)
);

INVX4 _13606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf0),
    .Y(_4115_)
);

INVX1 _13607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_4116_)
);

NOR2X1 _13608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .B(_3954__bF$buf1),
    .Y(_4117_)
);

AOI21X1 _13609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .B(_4115_),
    .C(_4117_),
    .Y(_4118_)
);

NAND3X1 _13610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4114_),
    .B(_4118_),
    .C(_4111_),
    .Y(_4119_)
);

NOR2X1 _13611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4104_),
    .B(_4119_),
    .Y(_4120_)
);

INVX1 _13612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_4121_)
);

INVX1 _13613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_4122_)
);

OAI22X1 _13614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4122_),
    .B(_3910_),
    .C(_3982__bF$buf0),
    .D(_4121_),
    .Y(_4123_)
);

INVX1 _13615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_4124_)
);

INVX1 _13616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_4125_)
);

OAI22X1 _13617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3890_),
    .B(_4125_),
    .C(_4124_),
    .D(_3931__bF$buf0),
    .Y(_4126_)
);

NOR2X1 _13618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4126_),
    .B(_4123_),
    .Y(_4127_)
);

AOI22X1 _13619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .B(_3942__bF$buf0),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_4128_)
);

INVX8 _13620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf0),
    .Y(_4129_)
);

AOI22X1 _13621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [3]),
    .B(_4129_),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_4130_)
);

NAND3X1 _13622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4128_),
    .B(_4130_),
    .C(_4127_),
    .Y(_4131_)
);

INVX1 _13623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_4132_)
);

NOR2X1 _13624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4132_),
    .B(_3983__bF$buf1),
    .Y(_4133_)
);

AOI21X1 _13625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [3]),
    .B(_4038__bF$buf1),
    .C(_4133_),
    .Y(_4134_)
);

INVX8 _13626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972__bF$buf0),
    .Y(_4135_)
);

AOI22X1 _13627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [3]),
    .C(\datapath_1.regfile_1.regOut[18] [3]),
    .D(_4135_),
    .Y(_4136_)
);

INVX1 _13628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [3]),
    .Y(_4137_)
);

INVX1 _13629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [3]),
    .Y(_4138_)
);

OAI22X1 _13630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4137_),
    .B(_3925_),
    .C(_3881_),
    .D(_4138_),
    .Y(_4139_)
);

INVX1 _13631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_4140_)
);

INVX1 _13632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_4141_)
);

OAI22X1 _13633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4141_),
    .B(_3971__bF$buf1),
    .C(_3924__bF$buf0),
    .D(_4140_),
    .Y(_4142_)
);

NOR2X1 _13634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4139_),
    .B(_4142_),
    .Y(_4143_)
);

NAND3X1 _13635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4134_),
    .B(_4136_),
    .C(_4143_),
    .Y(_4144_)
);

NOR2X1 _13636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4131_),
    .B(_4144_),
    .Y(_4145_)
);

AOI21X1 _13637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4120_),
    .B(_4145_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [3])
);

INVX1 _13638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_4146_)
);

INVX1 _13639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_4147_)
);

OAI22X1 _13640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4146_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf0),
    .D(_4147_),
    .Y(_4148_)
);

INVX1 _13641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_4149_)
);

INVX1 _13642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_4150_)
);

OAI22X1 _13643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4149_),
    .B(_3905__bF$buf3),
    .C(_3935__bF$buf0),
    .D(_4150_),
    .Y(_4151_)
);

NOR2X1 _13644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4151_),
    .B(_4148_),
    .Y(_4152_)
);

AOI22X1 _13645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .B(_3950__bF$buf0),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_4153_)
);

INVX8 _13646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf3),
    .Y(_4154_)
);

AOI22X1 _13647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .B(_4005__bF$buf2),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_4155_)
);

NAND3X1 _13648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4153_),
    .B(_4155_),
    .C(_4152_),
    .Y(_4156_)
);

INVX1 _13649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_4157_)
);

INVX1 _13650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_4158_)
);

OAI22X1 _13651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .B(_4157_),
    .C(_3971__bF$buf0),
    .D(_4158_),
    .Y(_4159_)
);

INVX1 _13652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_4160_)
);

INVX1 _13653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_4161_)
);

OAI22X1 _13654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4161_),
    .B(_3972__bF$buf3),
    .C(_3924__bF$buf3),
    .D(_4160_),
    .Y(_4162_)
);

NOR2X1 _13655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4159_),
    .B(_4162_),
    .Y(_4163_)
);

INVX1 _13656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_4164_)
);

INVX1 _13657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_4165_)
);

OAI22X1 _13658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4165_),
    .B(_3902__bF$buf3),
    .C(_3983__bF$buf0),
    .D(_4164_),
    .Y(_4166_)
);

INVX1 _13659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_4167_)
);

INVX1 _13660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_4168_)
);

OAI22X1 _13661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4167_),
    .B(_3936__bF$buf0),
    .C(_3978_),
    .D(_4168_),
    .Y(_4169_)
);

NOR2X1 _13662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4169_),
    .B(_4166_),
    .Y(_4170_)
);

NAND2X1 _13663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4170_),
    .B(_4163_),
    .Y(_4171_)
);

NOR2X1 _13664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4171_),
    .B(_4156_),
    .Y(_4172_)
);

AOI22X1 _13665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [4]),
    .C(\datapath_1.regfile_1.regOut[6] [4]),
    .D(_4001__bF$buf2),
    .Y(_4173_)
);

AOI22X1 _13666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [4]),
    .C(\datapath_1.regfile_1.regOut[31] [4]),
    .D(_3995__bF$buf2),
    .Y(_4174_)
);

INVX1 _13667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_4175_)
);

INVX1 _13668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_4176_)
);

OAI22X1 _13669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4176_),
    .B(_3941_),
    .C(_3960_),
    .D(_4175_),
    .Y(_4177_)
);

INVX1 _13670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [4]),
    .Y(_4178_)
);

INVX1 _13671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_4179_)
);

OAI22X1 _13672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4178_),
    .B(_3944__bF$buf0),
    .C(_3959_),
    .D(_4179_),
    .Y(_4180_)
);

NOR2X1 _13673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4177_),
    .B(_4180_),
    .Y(_4181_)
);

NAND3X1 _13674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4173_),
    .B(_4174_),
    .C(_4181_),
    .Y(_4182_)
);

INVX1 _13675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_4183_)
);

INVX1 _13676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_4184_)
);

OAI22X1 _13677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4183_),
    .B(_3931__bF$buf3),
    .C(_3977__bF$buf0),
    .D(_4184_),
    .Y(_4185_)
);

INVX1 _13678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .Y(_4186_)
);

INVX1 _13679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [4]),
    .Y(_4187_)
);

OAI22X1 _13680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4186_),
    .B(_3893__bF$buf1),
    .C(_3967__bF$buf3),
    .D(_4187_),
    .Y(_4188_)
);

NOR2X1 _13681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4188_),
    .B(_4185_),
    .Y(_4189_)
);

AOI22X1 _13682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[29] [4]),
    .C(\datapath_1.regfile_1.regOut[25] [4]),
    .D(_4040_),
    .Y(_4190_)
);

AOI22X1 _13683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .B(_4102_),
    .C(_3891__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_4191_)
);

NAND3X1 _13684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4190_),
    .B(_4191_),
    .C(_4189_),
    .Y(_4192_)
);

NOR2X1 _13685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4182_),
    .B(_4192_),
    .Y(_4193_)
);

AOI21X1 _13686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4172_),
    .B(_4193_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [4])
);

AOI22X1 _13687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [5]),
    .C(\datapath_1.regfile_1.regOut[31] [5]),
    .D(_3995__bF$buf1),
    .Y(_4194_)
);

INVX1 _13688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_4195_)
);

NOR2X1 _13689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4195_),
    .B(_3935__bF$buf4),
    .Y(_4196_)
);

AOI21X1 _13690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [5]),
    .B(_4001__bF$buf1),
    .C(_4196_),
    .Y(_4197_)
);

INVX1 _13691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_4198_)
);

INVX1 _13692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_4199_)
);

OAI22X1 _13693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4198_),
    .B(_3916_),
    .C(_3959_),
    .D(_4199_),
    .Y(_4200_)
);

INVX1 _13694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .Y(_4201_)
);

INVX1 _13695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_4202_)
);

OAI22X1 _13696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4201_),
    .B(_3893__bF$buf0),
    .C(_3966__bF$buf3),
    .D(_4202_),
    .Y(_4203_)
);

NOR2X1 _13697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4200_),
    .B(_4203_),
    .Y(_4204_)
);

NAND3X1 _13698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4194_),
    .B(_4197_),
    .C(_4204_),
    .Y(_4205_)
);

INVX1 _13699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [5]),
    .Y(_4206_)
);

INVX1 _13700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [5]),
    .Y(_4207_)
);

OAI22X1 _13701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf2),
    .B(_4207_),
    .C(_3944__bF$buf4),
    .D(_4206_),
    .Y(_4208_)
);

INVX1 _13702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [5]),
    .Y(_4209_)
);

INVX1 _13703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_4210_)
);

OAI22X1 _13704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf2),
    .B(_4209_),
    .C(_3955__bF$buf4),
    .D(_4210_),
    .Y(_4211_)
);

NOR2X1 _13705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4208_),
    .B(_4211_),
    .Y(_4212_)
);

INVX1 _13706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_4213_)
);

INVX1 _13707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_4214_)
);

OAI22X1 _13708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4214_),
    .B(_3902__bF$buf2),
    .C(_3954__bF$buf4),
    .D(_4213_),
    .Y(_4215_)
);

INVX1 _13709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_4216_)
);

INVX1 _13710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_4217_)
);

OAI22X1 _13711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4217_),
    .B(_3960_),
    .C(_3983__bF$buf4),
    .D(_4216_),
    .Y(_4218_)
);

NOR2X1 _13712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4218_),
    .B(_4215_),
    .Y(_4219_)
);

NAND2X1 _13713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4212_),
    .B(_4219_),
    .Y(_4220_)
);

NOR2X1 _13714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4220_),
    .B(_4205_),
    .Y(_4221_)
);

INVX1 _13715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_4222_)
);

NOR2X1 _13716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4222_),
    .B(_3971__bF$buf4),
    .Y(_4223_)
);

AOI21X1 _13717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .B(_4090_),
    .C(_4223_),
    .Y(_4224_)
);

AND2X2 _13718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .B(_3888_),
    .Y(_4225_)
);

AOI22X1 _13719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .B(_3942__bF$buf3),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_4226_)
);

INVX1 _13720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_4227_)
);

INVX1 _13721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_4228_)
);

OAI22X1 _13722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4227_),
    .B(_3910_),
    .C(_3978_),
    .D(_4228_),
    .Y(_4229_)
);

INVX1 _13723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [5]),
    .Y(_4230_)
);

INVX1 _13724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_4231_)
);

OAI22X1 _13725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4231_),
    .B(_3949_),
    .C(_3881_),
    .D(_4230_),
    .Y(_4232_)
);

NOR2X1 _13726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4229_),
    .B(_4232_),
    .Y(_4233_)
);

NAND3X1 _13727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4224_),
    .B(_4226_),
    .C(_4233_),
    .Y(_4234_)
);

INVX1 _13728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_4235_)
);

INVX1 _13729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_4236_)
);

OAI22X1 _13730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4235_),
    .B(_3905__bF$buf2),
    .C(_3977__bF$buf4),
    .D(_4236_),
    .Y(_4237_)
);

INVX1 _13731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_4238_)
);

INVX1 _13732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_4239_)
);

OAI22X1 _13733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4239_),
    .B(_3936__bF$buf4),
    .C(_3972__bF$buf2),
    .D(_4238_),
    .Y(_4240_)
);

NOR2X1 _13734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4240_),
    .B(_4237_),
    .Y(_4241_)
);

AOI22X1 _13735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .B(_3891__bF$buf0),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_4242_)
);

AOI22X1 _13736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .B(_4102_),
    .C(_4079__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_4243_)
);

NAND3X1 _13737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4242_),
    .B(_4243_),
    .C(_4241_),
    .Y(_4244_)
);

NOR2X1 _13738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4244_),
    .B(_4234_),
    .Y(_4245_)
);

AOI21X1 _13739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4221_),
    .B(_4245_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [5])
);

INVX8 _13740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905__bF$buf1),
    .Y(_4246_)
);

AOI22X1 _13741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4246_),
    .B(\datapath_1.regfile_1.regOut[19] [6]),
    .C(\datapath_1.regfile_1.regOut[12] [6]),
    .D(_4005__bF$buf1),
    .Y(_4247_)
);

AOI22X1 _13742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4154_),
    .B(\datapath_1.regfile_1.regOut[14] [6]),
    .C(\datapath_1.regfile_1.regOut[31] [6]),
    .D(_3995__bF$buf0),
    .Y(_4248_)
);

INVX1 _13743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [6]),
    .Y(_4249_)
);

INVX1 _13744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_4250_)
);

OAI22X1 _13745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3960_),
    .B(_4250_),
    .C(_3944__bF$buf3),
    .D(_4249_),
    .Y(_4251_)
);

INVX1 _13746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_4252_)
);

INVX1 _13747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_4253_)
);

OAI22X1 _13748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4253_),
    .B(_3902__bF$buf1),
    .C(_3966__bF$buf2),
    .D(_4252_),
    .Y(_4254_)
);

NOR2X1 _13749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4251_),
    .B(_4254_),
    .Y(_4255_)
);

NAND3X1 _13750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4247_),
    .B(_4248_),
    .C(_4255_),
    .Y(_4256_)
);

AOI22X1 _13751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .B(_4038__bF$buf0),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_4257_)
);

AOI22X1 _13752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .B(_3894_),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_4258_)
);

INVX1 _13753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_4259_)
);

INVX1 _13754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_4260_)
);

OAI22X1 _13755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4260_),
    .B(_3949_),
    .C(_3983__bF$buf3),
    .D(_4259_),
    .Y(_4261_)
);

INVX1 _13756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .Y(_4262_)
);

INVX1 _13757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_4263_)
);

OAI22X1 _13758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf1),
    .B(_4262_),
    .C(_3977__bF$buf3),
    .D(_4263_),
    .Y(_4264_)
);

NOR2X1 _13759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4261_),
    .B(_4264_),
    .Y(_4265_)
);

NAND3X1 _13760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4257_),
    .B(_4258_),
    .C(_4265_),
    .Y(_4266_)
);

NOR2X1 _13761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4256_),
    .B(_4266_),
    .Y(_4267_)
);

INVX1 _13762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_4268_)
);

NOR2X1 _13763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4268_),
    .B(_3959_),
    .Y(_4269_)
);

INVX1 _13764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_4270_)
);

NOR2X1 _13765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4270_),
    .B(_3931__bF$buf2),
    .Y(_4271_)
);

INVX1 _13766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_4272_)
);

INVX1 _13767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_4273_)
);

OAI22X1 _13768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3941_),
    .B(_4273_),
    .C(_3930__bF$buf0),
    .D(_4272_),
    .Y(_4274_)
);

NOR3X1 _13769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4271_),
    .B(_4274_),
    .C(_4269_),
    .Y(_4275_)
);

AOI22X1 _13770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [6]),
    .C(\datapath_1.regfile_1.regOut[6] [6]),
    .D(_4001__bF$buf0),
    .Y(_4276_)
);

AOI22X1 _13771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [6]),
    .C(\datapath_1.regfile_1.regOut[13] [6]),
    .D(_4051__bF$buf1),
    .Y(_4277_)
);

NAND3X1 _13772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4276_),
    .B(_4277_),
    .C(_4275_),
    .Y(_4278_)
);

INVX1 _13773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_4279_)
);

INVX1 _13774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_4280_)
);

OAI22X1 _13775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4279_),
    .B(_3936__bF$buf3),
    .C(_3971__bF$buf3),
    .D(_4280_),
    .Y(_4281_)
);

INVX1 _13776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_4282_)
);

INVX1 _13777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_4283_)
);

OAI22X1 _13778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4283_),
    .B(_3935__bF$buf3),
    .C(_3924__bF$buf2),
    .D(_4282_),
    .Y(_4284_)
);

NOR2X1 _13779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4281_),
    .B(_4284_),
    .Y(_4285_)
);

INVX1 _13780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_4286_)
);

INVX1 _13781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_4287_)
);

OAI22X1 _13782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4286_),
    .B(_3955__bF$buf3),
    .C(_3954__bF$buf3),
    .D(_4287_),
    .Y(_4288_)
);

INVX1 _13783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [6]),
    .Y(_4289_)
);

INVX1 _13784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_4290_)
);

OAI22X1 _13785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4290_),
    .B(_3890_),
    .C(_3967__bF$buf1),
    .D(_4289_),
    .Y(_4291_)
);

NOR2X1 _13786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4291_),
    .B(_4288_),
    .Y(_4292_)
);

NAND2X1 _13787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4292_),
    .B(_4285_),
    .Y(_4293_)
);

NOR2X1 _13788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4293_),
    .B(_4278_),
    .Y(_4294_)
);

AOI21X1 _13789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4267_),
    .B(_4294_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [6])
);

INVX1 _13790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .Y(_4295_)
);

NAND2X1 _13791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .B(_4102_),
    .Y(_4296_)
);

OAI21X1 _13792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4295_),
    .B(_3967__bF$buf0),
    .C(_4296_),
    .Y(_4297_)
);

INVX1 _13793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_4298_)
);

INVX1 _13794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_4299_)
);

OAI22X1 _13795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4299_),
    .B(_3972__bF$buf1),
    .C(_3920_),
    .D(_4298_),
    .Y(_4300_)
);

NOR2X1 _13796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4300_),
    .B(_4297_),
    .Y(_4301_)
);

INVX1 _13797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_4302_)
);

NOR2X1 _13798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4302_),
    .B(_3949_),
    .Y(_4303_)
);

INVX1 _13799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_4304_)
);

NOR2X1 _13800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4304_),
    .B(_3910_),
    .Y(_4305_)
);

INVX1 _13801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_4306_)
);

INVX1 _13802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_4307_)
);

OAI22X1 _13803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905__bF$buf0),
    .B(_4306_),
    .C(_3902__bF$buf0),
    .D(_4307_),
    .Y(_4308_)
);

NOR3X1 _13804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4303_),
    .B(_4305_),
    .C(_4308_),
    .Y(_4309_)
);

NAND2X1 _13805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4309_),
    .B(_4301_),
    .Y(_4310_)
);

AOI22X1 _13806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .B(_3894_),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_4311_)
);

AOI22X1 _13807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .B(_4038__bF$buf3),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_4312_)
);

INVX1 _13808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [7]),
    .Y(_4313_)
);

INVX1 _13809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_4314_)
);

OAI22X1 _13810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4313_),
    .B(_3944__bF$buf2),
    .C(_3959_),
    .D(_4314_),
    .Y(_4315_)
);

INVX1 _13811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_4316_)
);

INVX1 _13812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_4317_)
);

OAI22X1 _13813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_3936__bF$buf2),
    .C(_3935__bF$buf2),
    .D(_4317_),
    .Y(_4318_)
);

NOR2X1 _13814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4318_),
    .B(_4315_),
    .Y(_4319_)
);

NAND3X1 _13815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4311_),
    .B(_4312_),
    .C(_4319_),
    .Y(_4320_)
);

NOR2X1 _13816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4320_),
    .B(_4310_),
    .Y(_4321_)
);

AOI22X1 _13817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [7]),
    .C(\datapath_1.regfile_1.regOut[6] [7]),
    .D(_4001__bF$buf3),
    .Y(_4322_)
);

AOI22X1 _13818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [7]),
    .C(\datapath_1.regfile_1.regOut[8] [7]),
    .D(_4090_),
    .Y(_4323_)
);

INVX1 _13819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_4324_)
);

INVX1 _13820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_4325_)
);

OAI22X1 _13821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .B(_3941_),
    .C(_3960_),
    .D(_4324_),
    .Y(_4326_)
);

INVX1 _13822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_4327_)
);

INVX1 _13823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_4328_)
);

OAI22X1 _13824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4327_),
    .B(_3955__bF$buf2),
    .C(_3954__bF$buf2),
    .D(_4328_),
    .Y(_4329_)
);

NOR2X1 _13825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4326_),
    .B(_4329_),
    .Y(_4330_)
);

NAND3X1 _13826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4322_),
    .B(_4323_),
    .C(_4330_),
    .Y(_4331_)
);

AOI22X1 _13827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [7]),
    .C(\datapath_1.regfile_1.regOut[31] [7]),
    .D(_3995__bF$buf4),
    .Y(_4332_)
);

INVX1 _13828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_4333_)
);

NOR2X1 _13829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4333_),
    .B(_3971__bF$buf2),
    .Y(_4334_)
);

AOI21X1 _13830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .B(_4040_),
    .C(_4334_),
    .Y(_4335_)
);

INVX1 _13831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_4336_)
);

INVX1 _13832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_4337_)
);

OAI22X1 _13833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_4336_),
    .C(_3977__bF$buf2),
    .D(_4337_),
    .Y(_4338_)
);

INVX1 _13834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_4339_)
);

INVX1 _13835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_4340_)
);

OAI22X1 _13836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4340_),
    .B(_3982__bF$buf2),
    .C(_3983__bF$buf2),
    .D(_4339_),
    .Y(_4341_)
);

NOR2X1 _13837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(_4338_),
    .Y(_4342_)
);

NAND3X1 _13838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4332_),
    .B(_4335_),
    .C(_4342_),
    .Y(_4343_)
);

NOR2X1 _13839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4331_),
    .B(_4343_),
    .Y(_4344_)
);

AOI21X1 _13840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4321_),
    .B(_4344_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [7])
);

INVX1 _13841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_4345_)
);

INVX1 _13842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_4346_)
);

OAI22X1 _13843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4346_),
    .B(_3941_),
    .C(_3890_),
    .D(_4345_),
    .Y(_4347_)
);

INVX1 _13844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [8]),
    .Y(_4348_)
);

INVX1 _13845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_4349_)
);

OAI22X1 _13846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944__bF$buf1),
    .B(_4348_),
    .C(_4349_),
    .D(_3955__bF$buf1),
    .Y(_4350_)
);

NOR2X1 _13847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4347_),
    .B(_4350_),
    .Y(_4351_)
);

AOI22X1 _13848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .B(_4005__bF$buf0),
    .C(_4001__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_4352_)
);

INVX1 _13849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_4353_)
);

NOR2X1 _13850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4353_),
    .B(_3977__bF$buf1),
    .Y(_4354_)
);

AOI21X1 _13851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .B(_3894_),
    .C(_4354_),
    .Y(_4355_)
);

NAND3X1 _13852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4352_),
    .B(_4355_),
    .C(_4351_),
    .Y(_4356_)
);

AOI22X1 _13853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .B(_4115_),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_4357_)
);

AOI22X1 _13854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .B(_4246_),
    .C(_3998__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_4358_)
);

INVX1 _13855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_4359_)
);

INVX1 _13856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_4360_)
);

OAI22X1 _13857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4360_),
    .B(_3935__bF$buf1),
    .C(_3966__bF$buf1),
    .D(_4359_),
    .Y(_4361_)
);

INVX1 _13858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_4362_)
);

INVX1 _13859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_4363_)
);

OAI22X1 _13860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4363_),
    .B(_3936__bF$buf1),
    .C(_3954__bF$buf1),
    .D(_4362_),
    .Y(_4364_)
);

NOR2X1 _13861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4364_),
    .B(_4361_),
    .Y(_4365_)
);

NAND3X1 _13862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4357_),
    .B(_4358_),
    .C(_4365_),
    .Y(_4366_)
);

NOR2X1 _13863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4356_),
    .B(_4366_),
    .Y(_4367_)
);

AOI22X1 _13864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .B(_4154_),
    .C(_4051__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_4368_)
);

AOI22X1 _13865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .B(_4090_),
    .C(_3948_),
    .D(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_4369_)
);

INVX1 _13866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_4370_)
);

INVX1 _13867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_4371_)
);

OAI22X1 _13868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4371_),
    .B(_3949_),
    .C(_3983__bF$buf1),
    .D(_4370_),
    .Y(_4372_)
);

INVX1 _13869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [8]),
    .Y(_4373_)
);

INVX1 _13870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .Y(_4374_)
);

OAI22X1 _13871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf0),
    .B(_4373_),
    .C(_4374_),
    .D(_3967__bF$buf3),
    .Y(_4375_)
);

NOR2X1 _13872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4375_),
    .B(_4372_),
    .Y(_4376_)
);

NAND3X1 _13873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4368_),
    .B(_4369_),
    .C(_4376_),
    .Y(_4377_)
);

INVX1 _13874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_4378_)
);

INVX1 _13875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_4379_)
);

OAI22X1 _13876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_3972__bF$buf0),
    .C(_3920_),
    .D(_4378_),
    .Y(_4380_)
);

INVX1 _13877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [8]),
    .Y(_4381_)
);

INVX1 _13878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_4382_)
);

OAI22X1 _13879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4382_),
    .B(_3916_),
    .C(_3881_),
    .D(_4381_),
    .Y(_4383_)
);

NOR2X1 _13880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4383_),
    .B(_4380_),
    .Y(_4384_)
);

INVX1 _13881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_4385_)
);

NOR2X1 _13882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4385_),
    .B(_3971__bF$buf1),
    .Y(_4386_)
);

AOI21X1 _13883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .B(_4225_),
    .C(_4386_),
    .Y(_4387_)
);

AOI22X1 _13884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .B(_4102_),
    .C(_3995__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_4388_)
);

NAND3X1 _13885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4387_),
    .B(_4388_),
    .C(_4384_),
    .Y(_4389_)
);

NOR2X1 _13886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4377_),
    .B(_4389_),
    .Y(_4390_)
);

AOI21X1 _13887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4367_),
    .B(_4390_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [8])
);

INVX1 _13888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_4391_)
);

INVX1 _13889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_4392_)
);

OAI22X1 _13890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4392_),
    .B(_3983__bF$buf0),
    .C(_3920_),
    .D(_4391_),
    .Y(_4393_)
);

INVX1 _13891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .Y(_4394_)
);

INVX1 _13892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [9]),
    .Y(_4395_)
);

OAI22X1 _13893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4394_),
    .B(_3893__bF$buf3),
    .C(_3944__bF$buf0),
    .D(_4395_),
    .Y(_4396_)
);

NOR2X1 _13894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4396_),
    .B(_4393_),
    .Y(_4397_)
);

AOI22X1 _13895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .B(_4246_),
    .C(_4115_),
    .D(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_4398_)
);

AOI22X1 _13896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .B(_3942__bF$buf2),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_4399_)
);

NAND3X1 _13897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4398_),
    .B(_4399_),
    .C(_4397_),
    .Y(_4400_)
);

AOI22X1 _13898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .B(_4225_),
    .C(_3885_),
    .D(\datapath_1.regfile_1.regOut[30] [9]),
    .Y(_4401_)
);

AOI22X1 _13899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[23] [9]),
    .C(\datapath_1.regfile_1.regOut[18] [9]),
    .D(_4135_),
    .Y(_4402_)
);

INVX1 _13900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [9]),
    .Y(_4403_)
);

INVX1 _13901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_4404_)
);

OAI22X1 _13902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4404_),
    .B(_3931__bF$buf1),
    .C(_3966__bF$buf0),
    .D(_4403_),
    .Y(_4405_)
);

INVX1 _13903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_4406_)
);

INVX1 _13904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_4407_)
);

OAI22X1 _13905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4406_),
    .B(_3936__bF$buf0),
    .C(_3935__bF$buf0),
    .D(_4407_),
    .Y(_4408_)
);

NOR2X1 _13906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4408_),
    .B(_4405_),
    .Y(_4409_)
);

NAND3X1 _13907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4401_),
    .B(_4402_),
    .C(_4409_),
    .Y(_4410_)
);

NOR2X1 _13908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4410_),
    .B(_4400_),
    .Y(_4411_)
);

AOI22X1 _13909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .B(_4102_),
    .C(_4001__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_4412_)
);

AOI22X1 _13910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [9]),
    .B(_3891__bF$buf2),
    .C(_3998__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_4413_)
);

INVX1 _13911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_4414_)
);

INVX1 _13912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_4415_)
);

OAI22X1 _13913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4414_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf0),
    .D(_4415_),
    .Y(_4416_)
);

INVX1 _13914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_4417_)
);

INVX1 _13915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_4418_)
);

OAI22X1 _13916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf0),
    .B(_4417_),
    .C(_3977__bF$buf0),
    .D(_4418_),
    .Y(_4419_)
);

NOR2X1 _13917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4419_),
    .B(_4416_),
    .Y(_4420_)
);

NAND3X1 _13918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4412_),
    .B(_4413_),
    .C(_4420_),
    .Y(_4421_)
);

INVX1 _13919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [9]),
    .Y(_4422_)
);

INVX1 _13920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .Y(_4423_)
);

OAI22X1 _13921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4423_),
    .B(_3967__bF$buf2),
    .C(_3881_),
    .D(_4422_),
    .Y(_4424_)
);

INVX1 _13922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [9]),
    .Y(_4425_)
);

INVX1 _13923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_4426_)
);

OAI22X1 _13924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4425_),
    .B(_3925_),
    .C(_3971__bF$buf0),
    .D(_4426_),
    .Y(_4427_)
);

NOR2X1 _13925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4424_),
    .B(_4427_),
    .Y(_4428_)
);

AOI22X1 _13926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .B(_4154_),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_4429_)
);

AOI22X1 _13927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .B(_4005__bF$buf3),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_4430_)
);

NAND3X1 _13928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4429_),
    .B(_4430_),
    .C(_4428_),
    .Y(_4431_)
);

NOR2X1 _13929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4421_),
    .B(_4431_),
    .Y(_4432_)
);

AOI21X1 _13930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4432_),
    .B(_4411_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [9])
);

AOI22X1 _13931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .B(_3942__bF$buf1),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_4433_)
);

INVX1 _13932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [10]),
    .Y(_4434_)
);

NOR2X1 _13933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434_),
    .B(_3944__bF$buf4),
    .Y(_4435_)
);

AOI21X1 _13934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .B(_4102_),
    .C(_4435_),
    .Y(_4436_)
);

INVX1 _13935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_4437_)
);

INVX1 _13936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_4438_)
);

OAI22X1 _13937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf3),
    .B(_4438_),
    .C(_3954__bF$buf4),
    .D(_4437_),
    .Y(_4439_)
);

INVX1 _13938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_4440_)
);

INVX1 _13939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_4441_)
);

OAI22X1 _13940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4440_),
    .B(_3931__bF$buf0),
    .C(_3977__bF$buf4),
    .D(_4441_),
    .Y(_4442_)
);

NOR2X1 _13941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4442_),
    .B(_4439_),
    .Y(_4443_)
);

NAND3X1 _13942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4433_),
    .B(_4436_),
    .C(_4443_),
    .Y(_4444_)
);

INVX1 _13943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [10]),
    .Y(_4445_)
);

INVX1 _13944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_4446_)
);

OAI22X1 _13945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4446_),
    .B(_3909_),
    .C(_3881_),
    .D(_4445_),
    .Y(_4447_)
);

INVX1 _13946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_4448_)
);

INVX1 _13947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_4449_)
);

OAI22X1 _13948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4449_),
    .B(_3972__bF$buf3),
    .C(_3920_),
    .D(_4448_),
    .Y(_4450_)
);

NOR2X1 _13949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4447_),
    .B(_4450_),
    .Y(_4451_)
);

AOI22X1 _13950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .B(_4246_),
    .C(_4129_),
    .D(\datapath_1.regfile_1.regOut[27] [10]),
    .Y(_4452_)
);

AOI22X1 _13951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .B(_4225_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_4453_)
);

NAND3X1 _13952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4452_),
    .B(_4453_),
    .C(_4451_),
    .Y(_4454_)
);

NOR2X1 _13953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4444_),
    .B(_4454_),
    .Y(_4455_)
);

INVX1 _13954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_4456_)
);

INVX1 _13955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_4457_)
);

OAI22X1 _13956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4456_),
    .B(_3902__bF$buf3),
    .C(_3971__bF$buf4),
    .D(_4457_),
    .Y(_4458_)
);

INVX1 _13957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_4459_)
);

INVX1 _13958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_4460_)
);

OAI22X1 _13959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4459_),
    .B(_3936__bF$buf4),
    .C(_3935__bF$buf4),
    .D(_4460_),
    .Y(_4461_)
);

NOR2X1 _13960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4461_),
    .B(_4458_),
    .Y(_4462_)
);

AOI22X1 _13961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .B(_3891__bF$buf1),
    .C(_3998__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_4463_)
);

AOI22X1 _13962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .B(_4005__bF$buf2),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_4464_)
);

NAND3X1 _13963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4463_),
    .B(_4464_),
    .C(_4462_),
    .Y(_4465_)
);

INVX1 _13964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_4466_)
);

INVX1 _13965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_4467_)
);

OAI22X1 _13966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4466_),
    .B(_3916_),
    .C(_3983__bF$buf4),
    .D(_4467_),
    .Y(_4468_)
);

INVX1 _13967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .Y(_4469_)
);

INVX1 _13968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_4470_)
);

OAI22X1 _13969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf3),
    .B(_4469_),
    .C(_3955__bF$buf4),
    .D(_4470_),
    .Y(_4471_)
);

NOR2X1 _13970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4471_),
    .B(_4468_),
    .Y(_4472_)
);

AOI22X1 _13971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .B(_4154_),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_4473_)
);

AOI22X1 _13972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .B(_3894_),
    .C(_3995__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_4474_)
);

NAND3X1 _13973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4473_),
    .B(_4474_),
    .C(_4472_),
    .Y(_4475_)
);

NOR2X1 _13974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4475_),
    .B(_4465_),
    .Y(_4476_)
);

AOI21X1 _13975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4476_),
    .B(_4455_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [10])
);

AOI22X1 _13976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .B(_3891__bF$buf0),
    .C(_3998__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_4477_)
);

INVX1 _13977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_4478_)
);

NOR2X1 _13978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4478_),
    .B(_3935__bF$buf3),
    .Y(_4479_)
);

AOI21X1 _13979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .B(_4115_),
    .C(_4479_),
    .Y(_4480_)
);

INVX1 _13980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_4481_)
);

INVX1 _13981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_4482_)
);

OAI22X1 _13982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4481_),
    .B(_3930__bF$buf3),
    .C(_3977__bF$buf3),
    .D(_4482_),
    .Y(_4483_)
);

INVX1 _13983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [11]),
    .Y(_4484_)
);

INVX1 _13984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_4485_)
);

OAI22X1 _13985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4485_),
    .B(_3916_),
    .C(_3881_),
    .D(_4484_),
    .Y(_4486_)
);

NOR2X1 _13986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4486_),
    .B(_4483_),
    .Y(_4487_)
);

NAND3X1 _13987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4477_),
    .B(_4480_),
    .C(_4487_),
    .Y(_4488_)
);

AOI22X1 _13988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .B(_4005__bF$buf1),
    .C(_4001__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_4489_)
);

AOI22X1 _13989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .B(_3942__bF$buf0),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_4490_)
);

INVX1 _13990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_4491_)
);

INVX1 _13991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_4492_)
);

OAI22X1 _13992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4492_),
    .B(_3936__bF$buf3),
    .C(_3955__bF$buf3),
    .D(_4491_),
    .Y(_4493_)
);

INVX1 _13993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [11]),
    .Y(_4494_)
);

INVX1 _13994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [11]),
    .Y(_4495_)
);

OAI22X1 _13995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4494_),
    .B(_3893__bF$buf2),
    .C(_3944__bF$buf3),
    .D(_4495_),
    .Y(_4496_)
);

NOR2X1 _13996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4496_),
    .B(_4493_),
    .Y(_4497_)
);

NAND3X1 _13997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4489_),
    .B(_4490_),
    .C(_4497_),
    .Y(_4498_)
);

NOR2X1 _13998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4498_),
    .B(_4488_),
    .Y(_4499_)
);

INVX1 _13999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_4500_)
);

NOR2X1 _14000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4500_),
    .B(_3971__bF$buf3),
    .Y(_4501_)
);

AOI21X1 _14001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .B(_4225_),
    .C(_4501_),
    .Y(_4502_)
);

INVX1 _14002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_4503_)
);

NOR2X1 _14003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4503_),
    .B(_3983__bF$buf3),
    .Y(_4504_)
);

AOI21X1 _14004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [11]),
    .B(_4079__bF$buf2),
    .C(_4504_),
    .Y(_4505_)
);

INVX1 _14005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_4506_)
);

INVX1 _14006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_4507_)
);

OAI22X1 _14007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4506_),
    .B(_3931__bF$buf3),
    .C(_3947__bF$buf2),
    .D(_4507_),
    .Y(_4508_)
);

INVX1 _14008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_4509_)
);

INVX1 _14009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_4510_)
);

OAI22X1 _14010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4510_),
    .B(_3905__bF$buf3),
    .C(_3954__bF$buf3),
    .D(_4509_),
    .Y(_4511_)
);

NOR2X1 _14011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4508_),
    .B(_4511_),
    .Y(_4512_)
);

NAND3X1 _14012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4502_),
    .B(_4505_),
    .C(_4512_),
    .Y(_4513_)
);

INVX1 _14013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_4514_)
);

INVX1 _14014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_4515_)
);

OAI22X1 _14015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4515_),
    .B(_3949_),
    .C(_3978_),
    .D(_4514_),
    .Y(_4516_)
);

INVX1 _14016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [11]),
    .Y(_4517_)
);

INVX1 _14017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_4518_)
);

OAI22X1 _14018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf1),
    .B(_4518_),
    .C(_3966__bF$buf3),
    .D(_4517_),
    .Y(_4519_)
);

NOR2X1 _14019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4516_),
    .B(_4519_),
    .Y(_4520_)
);

AOI22X1 _14020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [11]),
    .C(\datapath_1.regfile_1.regOut[27] [11]),
    .D(_4129_),
    .Y(_4521_)
);

AOI22X1 _14021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4135_),
    .B(\datapath_1.regfile_1.regOut[18] [11]),
    .C(\datapath_1.regfile_1.regOut[31] [11]),
    .D(_3995__bF$buf1),
    .Y(_4522_)
);

NAND3X1 _14022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4521_),
    .B(_4522_),
    .C(_4520_),
    .Y(_4523_)
);

NOR2X1 _14023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4513_),
    .B(_4523_),
    .Y(_4524_)
);

AOI21X1 _14024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4524_),
    .B(_4499_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [11])
);

INVX1 _14025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [12]),
    .Y(_4525_)
);

INVX1 _14026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_4526_)
);

OAI22X1 _14027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4525_),
    .B(_3925_),
    .C(_3977__bF$buf2),
    .D(_4526_),
    .Y(_4527_)
);

INVX1 _14028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [12]),
    .Y(_4528_)
);

INVX1 _14029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_4529_)
);

OAI22X1 _14030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf0),
    .B(_4529_),
    .C(_3966__bF$buf2),
    .D(_4528_),
    .Y(_4530_)
);

NOR2X1 _14031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4530_),
    .B(_4527_),
    .Y(_4531_)
);

AOI22X1 _14032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .B(_4090_),
    .C(_3948_),
    .D(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_4532_)
);

INVX1 _14033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [12]),
    .Y(_4533_)
);

NOR2X1 _14034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4533_),
    .B(_3944__bF$buf2),
    .Y(_4534_)
);

AOI21X1 _14035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .B(_4079__bF$buf1),
    .C(_4534_),
    .Y(_4535_)
);

NAND3X1 _14036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4532_),
    .B(_4535_),
    .C(_4531_),
    .Y(_4536_)
);

AOI22X1 _14037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .B(_4005__bF$buf0),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_4537_)
);

AOI22X1 _14038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .B(_3885_),
    .C(_4051__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_4538_)
);

INVX1 _14039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_4539_)
);

NOR2X1 _14040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4539_),
    .B(_3960_),
    .Y(_4540_)
);

INVX1 _14041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_4541_)
);

NOR2X1 _14042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .B(_3890_),
    .Y(_4542_)
);

INVX1 _14043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_4543_)
);

INVX1 _14044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_4544_)
);

OAI22X1 _14045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3941_),
    .B(_4544_),
    .C(_3930__bF$buf2),
    .D(_4543_),
    .Y(_4545_)
);

NOR3X1 _14046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4542_),
    .B(_4545_),
    .C(_4540_),
    .Y(_4546_)
);

NAND3X1 _14047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4537_),
    .B(_4538_),
    .C(_4546_),
    .Y(_4547_)
);

NOR2X1 _14048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4547_),
    .B(_4536_),
    .Y(_4548_)
);

INVX1 _14049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_4549_)
);

INVX1 _14050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_4550_)
);

OAI22X1 _14051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4550_),
    .B(_3954__bF$buf2),
    .C(_3924__bF$buf1),
    .D(_4549_),
    .Y(_4551_)
);

INVX1 _14052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_4552_)
);

INVX1 _14053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_4553_)
);

OAI22X1 _14054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .B(_4552_),
    .C(_3935__bF$buf2),
    .D(_4553_),
    .Y(_4554_)
);

NOR2X1 _14055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4554_),
    .B(_4551_),
    .Y(_4555_)
);

INVX1 _14056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_4556_)
);

INVX1 _14057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_4557_)
);

OAI22X1 _14058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4557_),
    .B(_3905__bF$buf2),
    .C(_3972__bF$buf2),
    .D(_4556_),
    .Y(_4558_)
);

INVX1 _14059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_4559_)
);

INVX1 _14060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_4560_)
);

OAI22X1 _14061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4559_),
    .B(_3955__bF$buf2),
    .C(_3983__bF$buf2),
    .D(_4560_),
    .Y(_4561_)
);

NOR2X1 _14062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4558_),
    .B(_4561_),
    .Y(_4562_)
);

NAND2X1 _14063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4562_),
    .B(_4555_),
    .Y(_4563_)
);

AOI22X1 _14064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4129_),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .C(\datapath_1.regfile_1.regOut[6] [12]),
    .D(_4001__bF$buf3),
    .Y(_4564_)
);

AOI22X1 _14065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [12]),
    .B(_3950__bF$buf1),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [12]),
    .Y(_4565_)
);

INVX1 _14066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_4566_)
);

INVX1 _14067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_4567_)
);

OAI22X1 _14068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4566_),
    .B(_3936__bF$buf2),
    .C(_3902__bF$buf2),
    .D(_4567_),
    .Y(_4568_)
);

INVX1 _14069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .Y(_4569_)
);

INVX1 _14070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_4570_)
);

OAI22X1 _14071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4569_),
    .B(_3893__bF$buf1),
    .C(_3971__bF$buf2),
    .D(_4570_),
    .Y(_4571_)
);

NOR2X1 _14072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4568_),
    .B(_4571_),
    .Y(_4572_)
);

NAND3X1 _14073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4564_),
    .B(_4565_),
    .C(_4572_),
    .Y(_4573_)
);

NOR2X1 _14074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4563_),
    .B(_4573_),
    .Y(_4574_)
);

AOI21X1 _14075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4574_),
    .B(_4548_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [12])
);

AOI22X1 _14076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .B(_4005__bF$buf3),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_4575_)
);

AOI22X1 _14077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3998__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[2] [13]),
    .C(\datapath_1.regfile_1.regOut[27] [13]),
    .D(_4129_),
    .Y(_4576_)
);

INVX1 _14078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .Y(_4577_)
);

INVX1 _14079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_4578_)
);

OAI22X1 _14080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4577_),
    .B(_3893__bF$buf0),
    .C(_3977__bF$buf1),
    .D(_4578_),
    .Y(_4579_)
);

INVX1 _14081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [13]),
    .Y(_4580_)
);

INVX1 _14082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_4581_)
);

OAI22X1 _14083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4581_),
    .B(_3890_),
    .C(_3944__bF$buf1),
    .D(_4580_),
    .Y(_4582_)
);

NOR2X1 _14084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4582_),
    .B(_4579_),
    .Y(_4583_)
);

NAND3X1 _14085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4575_),
    .B(_4576_),
    .C(_4583_),
    .Y(_4584_)
);

INVX1 _14086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_4585_)
);

INVX1 _14087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_4586_)
);

OAI22X1 _14088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4586_),
    .B(_3941_),
    .C(_3916_),
    .D(_4585_),
    .Y(_4587_)
);

INVX1 _14089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [13]),
    .Y(_4588_)
);

INVX1 _14090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_4589_)
);

OAI22X1 _14091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4589_),
    .B(_3949_),
    .C(_3881_),
    .D(_4588_),
    .Y(_4590_)
);

NOR2X1 _14092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4587_),
    .B(_4590_),
    .Y(_4591_)
);

AOI22X1 _14093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .B(_4135_),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_4592_)
);

AOI22X1 _14094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .B(_3885_),
    .C(_4079__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_4593_)
);

NAND3X1 _14095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4592_),
    .B(_4593_),
    .C(_4591_),
    .Y(_4594_)
);

NOR2X1 _14096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4594_),
    .B(_4584_),
    .Y(_4595_)
);

AOI22X1 _14097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [13]),
    .C(\datapath_1.regfile_1.regOut[6] [13]),
    .D(_4001__bF$buf2),
    .Y(_4596_)
);

AOI22X1 _14098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[13] [13]),
    .C(\datapath_1.regfile_1.regOut[25] [13]),
    .D(_4040_),
    .Y(_4597_)
);

INVX1 _14099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_4598_)
);

INVX1 _14100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_4599_)
);

OAI22X1 _14101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4598_),
    .B(_3930__bF$buf1),
    .C(_3931__bF$buf2),
    .D(_4599_),
    .Y(_4600_)
);

INVX1 _14102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_4601_)
);

INVX1 _14103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_4602_)
);

OAI22X1 _14104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4602_),
    .B(_3936__bF$buf1),
    .C(_3905__bF$buf1),
    .D(_4601_),
    .Y(_4603_)
);

NOR2X1 _14105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4603_),
    .B(_4600_),
    .Y(_4604_)
);

NAND3X1 _14106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4604_),
    .B(_4596_),
    .C(_4597_),
    .Y(_4605_)
);

INVX1 _14107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_4606_)
);

NOR2X1 _14108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4606_),
    .B(_3971__bF$buf1),
    .Y(_4607_)
);

AOI21X1 _14109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .B(_4115_),
    .C(_4607_),
    .Y(_4608_)
);

INVX1 _14110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_4609_)
);

NOR2X1 _14111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4609_),
    .B(_3935__bF$buf1),
    .Y(_4610_)
);

AOI21X1 _14112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .B(_4225_),
    .C(_4610_),
    .Y(_4611_)
);

INVX1 _14113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_4612_)
);

INVX1 _14114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_4613_)
);

OAI22X1 _14115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4612_),
    .B(_3955__bF$buf1),
    .C(_3954__bF$buf1),
    .D(_4613_),
    .Y(_4614_)
);

INVX1 _14116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .Y(_4615_)
);

INVX1 _14117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_4616_)
);

OAI22X1 _14118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4615_),
    .B(_3925_),
    .C(_3983__bF$buf1),
    .D(_4616_),
    .Y(_4617_)
);

NOR2X1 _14119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4614_),
    .B(_4617_),
    .Y(_4618_)
);

NAND3X1 _14120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4608_),
    .B(_4611_),
    .C(_4618_),
    .Y(_4619_)
);

NOR2X1 _14121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4605_),
    .B(_4619_),
    .Y(_4620_)
);

AOI21X1 _14122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4620_),
    .B(_4595_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [13])
);

INVX1 _14123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [14]),
    .Y(_4621_)
);

INVX1 _14124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [14]),
    .Y(_4622_)
);

OAI22X1 _14125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4621_),
    .B(_3944__bF$buf0),
    .C(_3966__bF$buf1),
    .D(_4622_),
    .Y(_4623_)
);

INVX1 _14126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_4624_)
);

INVX1 _14127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_4625_)
);

OAI22X1 _14128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4625_),
    .B(_3972__bF$buf1),
    .C(_3920_),
    .D(_4624_),
    .Y(_4626_)
);

NOR2X1 _14129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4623_),
    .B(_4626_),
    .Y(_4627_)
);

AOI22X1 _14130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .B(_4005__bF$buf2),
    .C(_3950__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_4628_)
);

INVX2 _14131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936__bF$buf0),
    .Y(_4629_)
);

AOI22X1 _14132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_4630_)
);

NAND3X1 _14133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4628_),
    .B(_4630_),
    .C(_4627_),
    .Y(_4631_)
);

AOI22X1 _14134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .B(_4225_),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_4632_)
);

AOI22X1 _14135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[23] [14]),
    .C(\datapath_1.regfile_1.regOut[27] [14]),
    .D(_4129_),
    .Y(_4633_)
);

INVX1 _14136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_4634_)
);

INVX1 _14137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_4635_)
);

OAI22X1 _14138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4634_),
    .B(_3931__bF$buf1),
    .C(_3959_),
    .D(_4635_),
    .Y(_4636_)
);

INVX1 _14139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_4637_)
);

INVX1 _14140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_4638_)
);

OAI22X1 _14141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf1),
    .B(_4637_),
    .C(_4638_),
    .D(_3935__bF$buf0),
    .Y(_4639_)
);

NOR2X1 _14142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4639_),
    .B(_4636_),
    .Y(_4640_)
);

NAND3X1 _14143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4632_),
    .B(_4633_),
    .C(_4640_),
    .Y(_4641_)
);

NOR2X1 _14144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4641_),
    .B(_4631_),
    .Y(_4642_)
);

AOI22X1 _14145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [14]),
    .C(\datapath_1.regfile_1.regOut[6] [14]),
    .D(_4001__bF$buf1),
    .Y(_4643_)
);

AOI22X1 _14146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3894_),
    .B(\datapath_1.regfile_1.regOut[28] [14]),
    .C(\datapath_1.regfile_1.regOut[3] [14]),
    .D(_3942__bF$buf3),
    .Y(_4644_)
);

INVX1 _14147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_4645_)
);

INVX1 _14148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_4646_)
);

OAI22X1 _14149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4645_),
    .B(_3955__bF$buf0),
    .C(_3954__bF$buf0),
    .D(_4646_),
    .Y(_4647_)
);

INVX1 _14150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_4648_)
);

INVX1 _14151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_4649_)
);

OAI22X1 _14152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4648_),
    .B(_3890_),
    .C(_3960_),
    .D(_4649_),
    .Y(_4650_)
);

NOR2X1 _14153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4650_),
    .B(_4647_),
    .Y(_4651_)
);

NAND3X1 _14154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4643_),
    .B(_4644_),
    .C(_4651_),
    .Y(_4652_)
);

INVX1 _14155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [14]),
    .Y(_4653_)
);

INVX1 _14156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [14]),
    .Y(_4654_)
);

OAI22X1 _14157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf2),
    .B(_4653_),
    .C(_4654_),
    .D(_3925_),
    .Y(_4655_)
);

INVX1 _14158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_4656_)
);

INVX1 _14159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_4657_)
);

OAI22X1 _14160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4656_),
    .B(_3930__bF$buf0),
    .C(_3971__bF$buf0),
    .D(_4657_),
    .Y(_4658_)
);

NOR2X1 _14161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4655_),
    .B(_4658_),
    .Y(_4659_)
);

INVX1 _14162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_4660_)
);

INVX1 _14163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_4661_)
);

OAI22X1 _14164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_4660_),
    .C(_3977__bF$buf0),
    .D(_4661_),
    .Y(_4662_)
);

INVX1 _14165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_4663_)
);

INVX1 _14166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_4664_)
);

OAI22X1 _14167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4664_),
    .B(_3982__bF$buf3),
    .C(_3983__bF$buf0),
    .D(_4663_),
    .Y(_4665_)
);

NOR2X1 _14168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4665_),
    .B(_4662_),
    .Y(_4666_)
);

NAND2X1 _14169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4659_),
    .B(_4666_),
    .Y(_4667_)
);

NOR2X1 _14170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4667_),
    .B(_4652_),
    .Y(_4668_)
);

AOI21X1 _14171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4668_),
    .B(_4642_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [14])
);

INVX1 _14172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_4669_)
);

INVX1 _14173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [15]),
    .Y(_4670_)
);

OAI22X1 _14174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893__bF$buf3),
    .B(_4670_),
    .C(_3930__bF$buf3),
    .D(_4669_),
    .Y(_4671_)
);

INVX1 _14175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_4672_)
);

NOR2X1 _14176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .B(_3949_),
    .Y(_4673_)
);

INVX1 _14177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_4674_)
);

NOR2X1 _14178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4674_),
    .B(_3983__bF$buf4),
    .Y(_4675_)
);

NOR3X1 _14179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4673_),
    .B(_4671_),
    .C(_4675_),
    .Y(_4676_)
);

AOI22X1 _14180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .B(_3995__bF$buf0),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_4677_)
);

AOI22X1 _14181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .B(_4246_),
    .C(_4115_),
    .D(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_4678_)
);

NAND3X1 _14182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4677_),
    .B(_4678_),
    .C(_4676_),
    .Y(_4679_)
);

INVX1 _14183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_4680_)
);

NOR2X1 _14184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4680_),
    .B(_3977__bF$buf4),
    .Y(_4681_)
);

AOI21X1 _14185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [15]),
    .B(_4001__bF$buf0),
    .C(_4681_),
    .Y(_4682_)
);

AOI22X1 _14186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .B(_4005__bF$buf1),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_4683_)
);

INVX1 _14187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [15]),
    .Y(_4684_)
);

INVX1 _14188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_4685_)
);

OAI22X1 _14189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4684_),
    .B(_3944__bF$buf4),
    .C(_3959_),
    .D(_4685_),
    .Y(_4686_)
);

INVX1 _14190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_4687_)
);

INVX1 _14191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_4688_)
);

OAI22X1 _14192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4687_),
    .B(_3936__bF$buf4),
    .C(_3935__bF$buf4),
    .D(_4688_),
    .Y(_4689_)
);

NOR2X1 _14193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4689_),
    .B(_4686_),
    .Y(_4690_)
);

NAND3X1 _14194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4682_),
    .B(_4690_),
    .C(_4683_),
    .Y(_4691_)
);

NOR2X1 _14195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4691_),
    .B(_4679_),
    .Y(_4692_)
);

AOI22X1 _14196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [15]),
    .C(\datapath_1.regfile_1.regOut[8] [15]),
    .D(_4090_),
    .Y(_4693_)
);

AOI22X1 _14197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .B(_4135_),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_4694_)
);

INVX1 _14198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_4695_)
);

INVX1 _14199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_4696_)
);

OAI22X1 _14200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4696_),
    .B(_3941_),
    .C(_3960_),
    .D(_4695_),
    .Y(_4697_)
);

INVX1 _14201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_4698_)
);

INVX1 _14202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_4699_)
);

OAI22X1 _14203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4698_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf4),
    .D(_4699_),
    .Y(_4700_)
);

NOR2X1 _14204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4697_),
    .B(_4700_),
    .Y(_4701_)
);

NAND3X1 _14205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4693_),
    .B(_4694_),
    .C(_4701_),
    .Y(_4702_)
);

INVX1 _14206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_4703_)
);

INVX1 _14207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_4704_)
);

OAI22X1 _14208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4703_),
    .B(_3982__bF$buf2),
    .C(_3978_),
    .D(_4704_),
    .Y(_4705_)
);

INVX1 _14209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_4706_)
);

INVX1 _14210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_4707_)
);

OAI22X1 _14211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf1),
    .B(_4707_),
    .C(_3971__bF$buf4),
    .D(_4706_),
    .Y(_4708_)
);

NOR2X1 _14212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4705_),
    .B(_4708_),
    .Y(_4709_)
);

AOI22X1 _14213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[23] [15]),
    .C(\datapath_1.regfile_1.regOut[27] [15]),
    .D(_4129_),
    .Y(_4710_)
);

AOI22X1 _14214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .B(_3885_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_4711_)
);

NAND3X1 _14215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4710_),
    .B(_4711_),
    .C(_4709_),
    .Y(_4712_)
);

NOR2X1 _14216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4702_),
    .B(_4712_),
    .Y(_4713_)
);

AOI21X1 _14217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4713_),
    .B(_4692_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [15])
);

INVX1 _14218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_4714_)
);

INVX1 _14219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_4715_)
);

OAI22X1 _14220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4714_),
    .B(_3910_),
    .C(_3935__bF$buf3),
    .D(_4715_),
    .Y(_4716_)
);

INVX1 _14221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [16]),
    .Y(_4717_)
);

INVX1 _14222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_4718_)
);

OAI22X1 _14223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4718_),
    .B(_3936__bF$buf3),
    .C(_3967__bF$buf1),
    .D(_4717_),
    .Y(_4719_)
);

NOR2X1 _14224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4719_),
    .B(_4716_),
    .Y(_4720_)
);

AOI22X1 _14225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .B(_3891__bF$buf2),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_4721_)
);

AOI22X1 _14226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .B(_3942__bF$buf2),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_4722_)
);

NAND3X1 _14227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4721_),
    .B(_4722_),
    .C(_4720_),
    .Y(_4723_)
);

INVX1 _14228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_4724_)
);

INVX1 _14229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_4725_)
);

OAI22X1 _14230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf1),
    .B(_4724_),
    .C(_3971__bF$buf3),
    .D(_4725_),
    .Y(_4726_)
);

INVX1 _14231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_4727_)
);

INVX1 _14232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_4728_)
);

OAI22X1 _14233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3959_),
    .B(_4728_),
    .C(_3954__bF$buf3),
    .D(_4727_),
    .Y(_4729_)
);

NOR2X1 _14234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4726_),
    .B(_4729_),
    .Y(_4730_)
);

INVX1 _14235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_4731_)
);

INVX1 _14236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_4732_)
);

OAI22X1 _14237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4732_),
    .B(_3972__bF$buf0),
    .C(_3920_),
    .D(_4731_),
    .Y(_4733_)
);

INVX1 _14238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_4734_)
);

INVX1 _14239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_4735_)
);

OAI22X1 _14240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4734_),
    .B(_3955__bF$buf3),
    .C(_3924__bF$buf0),
    .D(_4735_),
    .Y(_4736_)
);

NOR2X1 _14241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4733_),
    .B(_4736_),
    .Y(_4737_)
);

NAND2X1 _14242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4730_),
    .B(_4737_),
    .Y(_4738_)
);

NOR2X1 _14243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4723_),
    .B(_4738_),
    .Y(_4739_)
);

INVX1 _14244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [16]),
    .Y(_4740_)
);

INVX1 _14245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [16]),
    .Y(_4741_)
);

OAI22X1 _14246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf1),
    .B(_4740_),
    .C(_3966__bF$buf0),
    .D(_4741_),
    .Y(_4742_)
);

INVX1 _14247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_4743_)
);

INVX1 _14248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_4744_)
);

OAI22X1 _14249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4743_),
    .B(_3905__bF$buf0),
    .C(_3909_),
    .D(_4744_),
    .Y(_4745_)
);

NOR2X1 _14250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4745_),
    .B(_4742_),
    .Y(_4746_)
);

AOI22X1 _14251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .B(_4038__bF$buf3),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [16]),
    .Y(_4747_)
);

AOI22X1 _14252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .B(_3894_),
    .C(_3995__bF$buf4),
    .D(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_4748_)
);

NAND3X1 _14253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4747_),
    .B(_4748_),
    .C(_4746_),
    .Y(_4749_)
);

INVX1 _14254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [16]),
    .Y(_4750_)
);

INVX1 _14255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_4751_)
);

OAI22X1 _14256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf0),
    .B(_4751_),
    .C(_4750_),
    .D(_3944__bF$buf3),
    .Y(_4752_)
);

INVX1 _14257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_4753_)
);

INVX1 _14258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_4754_)
);

OAI22X1 _14259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf3),
    .B(_4753_),
    .C(_3977__bF$buf3),
    .D(_4754_),
    .Y(_4755_)
);

NOR2X1 _14260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4752_),
    .B(_4755_),
    .Y(_4756_)
);

AOI22X1 _14261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [16]),
    .C(\datapath_1.regfile_1.regOut[2] [16]),
    .D(_3998__bF$buf3),
    .Y(_4757_)
);

AOI22X1 _14262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .B(_4102_),
    .C(_4090_),
    .D(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_4758_)
);

NAND3X1 _14263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4757_),
    .B(_4758_),
    .C(_4756_),
    .Y(_4759_)
);

NOR2X1 _14264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4749_),
    .B(_4759_),
    .Y(_4760_)
);

AOI21X1 _14265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4739_),
    .B(_4760_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [16])
);

INVX1 _14266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_4761_)
);

INVX1 _14267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_4762_)
);

OAI22X1 _14268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4761_),
    .B(_3910_),
    .C(_3935__bF$buf2),
    .D(_4762_),
    .Y(_4763_)
);

INVX1 _14269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .Y(_4764_)
);

INVX1 _14270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_4765_)
);

OAI22X1 _14271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4765_),
    .B(_3902__bF$buf3),
    .C(_3966__bF$buf3),
    .D(_4764_),
    .Y(_4766_)
);

NOR2X1 _14272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4763_),
    .B(_4766_),
    .Y(_4767_)
);

AOI22X1 _14273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .B(_3891__bF$buf1),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_4768_)
);

AOI22X1 _14274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .B(_3942__bF$buf1),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_4769_)
);

NAND3X1 _14275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4768_),
    .B(_4769_),
    .C(_4767_),
    .Y(_4770_)
);

INVX1 _14276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_4771_)
);

INVX1 _14277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_4772_)
);

OAI22X1 _14278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf0),
    .B(_4771_),
    .C(_3971__bF$buf2),
    .D(_4772_),
    .Y(_4773_)
);

INVX1 _14279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_4774_)
);

INVX1 _14280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_4775_)
);

OAI22X1 _14281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3959_),
    .B(_4775_),
    .C(_3954__bF$buf2),
    .D(_4774_),
    .Y(_4776_)
);

NOR2X1 _14282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4773_),
    .B(_4776_),
    .Y(_4777_)
);

AOI22X1 _14283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [17]),
    .B(_4135_),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_4778_)
);

INVX1 _14284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_4779_)
);

NOR2X1 _14285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4779_),
    .B(_3955__bF$buf2),
    .Y(_4780_)
);

AOI21X1 _14286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .B(_4225_),
    .C(_4780_),
    .Y(_4781_)
);

NAND3X1 _14287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4778_),
    .B(_4781_),
    .C(_4777_),
    .Y(_4782_)
);

NOR2X1 _14288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4770_),
    .B(_4782_),
    .Y(_4783_)
);

AOI22X1 _14289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .B(_4102_),
    .C(_3995__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [17]),
    .Y(_4784_)
);

AOI22X1 _14290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .B(_4246_),
    .C(_4001__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_4785_)
);

INVX1 _14291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [17]),
    .Y(_4786_)
);

INVX1 _14292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_4787_)
);

OAI22X1 _14293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4786_),
    .B(_3893__bF$buf2),
    .C(_3916_),
    .D(_4787_),
    .Y(_4788_)
);

INVX1 _14294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [17]),
    .Y(_4789_)
);

INVX1 _14295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [17]),
    .Y(_4790_)
);

OAI22X1 _14296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4789_),
    .B(_3884__bF$buf0),
    .C(_3881_),
    .D(_4790_),
    .Y(_4791_)
);

NOR2X1 _14297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4788_),
    .B(_4791_),
    .Y(_4792_)
);

NAND3X1 _14298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4784_),
    .B(_4785_),
    .C(_4792_),
    .Y(_4793_)
);

INVX1 _14299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .Y(_4794_)
);

INVX1 _14300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_4795_)
);

OAI22X1 _14301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4795_),
    .B(_3936__bF$buf2),
    .C(_3967__bF$buf0),
    .D(_4794_),
    .Y(_4796_)
);

INVX1 _14302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_4797_)
);

INVX1 _14303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_4798_)
);

OAI22X1 _14304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf2),
    .B(_4797_),
    .C(_3977__bF$buf2),
    .D(_4798_),
    .Y(_4799_)
);

NOR2X1 _14305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4796_),
    .B(_4799_),
    .Y(_4800_)
);

AOI22X1 _14306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [17]),
    .C(\datapath_1.regfile_1.regOut[2] [17]),
    .D(_3998__bF$buf2),
    .Y(_4801_)
);

INVX1 _14307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [17]),
    .Y(_4802_)
);

NOR2X1 _14308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4802_),
    .B(_3944__bF$buf2),
    .Y(_4803_)
);

AOI21X1 _14309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .B(_4090_),
    .C(_4803_),
    .Y(_4804_)
);

NAND3X1 _14310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4804_),
    .C(_4800_),
    .Y(_4805_)
);

NOR2X1 _14311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4793_),
    .B(_4805_),
    .Y(_4806_)
);

AOI21X1 _14312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4806_),
    .B(_4783_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [17])
);

AOI22X1 _14313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .B(_4154_),
    .C(_4051__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_4807_)
);

AOI22X1 _14314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [18]),
    .B(_4001__bF$buf2),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_4808_)
);

INVX1 _14315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_4809_)
);

INVX1 _14316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_4810_)
);

OAI22X1 _14317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4810_),
    .B(_3936__bF$buf1),
    .C(_3905__bF$buf3),
    .D(_4809_),
    .Y(_4811_)
);

INVX1 _14318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_4812_)
);

INVX1 _14319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_4813_)
);

OAI22X1 _14320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf0),
    .B(_4813_),
    .C(_3935__bF$buf1),
    .D(_4812_),
    .Y(_4814_)
);

NOR2X1 _14321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4811_),
    .B(_4814_),
    .Y(_4815_)
);

NAND3X1 _14322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4807_),
    .B(_4808_),
    .C(_4815_),
    .Y(_4816_)
);

AOI22X1 _14323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [18]),
    .B(_3950__bF$buf1),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_4817_)
);

AOI22X1 _14324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .B(_4005__bF$buf0),
    .C(_3995__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_4818_)
);

INVX1 _14325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_4819_)
);

INVX1 _14326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_4820_)
);

OAI22X1 _14327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .B(_4819_),
    .C(_3977__bF$buf1),
    .D(_4820_),
    .Y(_4821_)
);

INVX1 _14328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [18]),
    .Y(_4822_)
);

INVX1 _14329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_4823_)
);

OAI22X1 _14330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4822_),
    .B(_3884__bF$buf3),
    .C(_3920_),
    .D(_4823_),
    .Y(_4824_)
);

NOR2X1 _14331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4821_),
    .B(_4824_),
    .Y(_4825_)
);

NAND3X1 _14332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4817_),
    .B(_4818_),
    .C(_4825_),
    .Y(_4826_)
);

NOR2X1 _14333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4816_),
    .B(_4826_),
    .Y(_4827_)
);

INVX1 _14334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_4828_)
);

INVX1 _14335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_4829_)
);

OAI22X1 _14336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4828_),
    .B(_3955__bF$buf1),
    .C(_3924__bF$buf3),
    .D(_4829_),
    .Y(_4830_)
);

INVX1 _14337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_4831_)
);

INVX1 _14338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_4832_)
);

OAI22X1 _14339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf1),
    .B(_4831_),
    .C(_3971__bF$buf1),
    .D(_4832_),
    .Y(_4833_)
);

NOR2X1 _14340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4833_),
    .B(_4830_),
    .Y(_4834_)
);

INVX1 _14341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_4835_)
);

NOR2X1 _14342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4835_),
    .B(_3954__bF$buf1),
    .Y(_4836_)
);

AOI21X1 _14343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .B(_4115_),
    .C(_4836_),
    .Y(_4837_)
);

AOI22X1 _14344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .B(_4102_),
    .C(_3998__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_4838_)
);

NAND3X1 _14345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4837_),
    .B(_4838_),
    .C(_4834_),
    .Y(_4839_)
);

INVX1 _14346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [18]),
    .Y(_4840_)
);

INVX1 _14347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_4841_)
);

OAI22X1 _14348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4840_),
    .B(_3944__bF$buf1),
    .C(_3959_),
    .D(_4841_),
    .Y(_4842_)
);

INVX1 _14349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [18]),
    .Y(_4843_)
);

INVX1 _14350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_4844_)
);

OAI22X1 _14351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4844_),
    .B(_3941_),
    .C(_3967__bF$buf3),
    .D(_4843_),
    .Y(_4845_)
);

NOR2X1 _14352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4845_),
    .B(_4842_),
    .Y(_4846_)
);

AOI22X1 _14353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [18]),
    .C(\datapath_1.regfile_1.regOut[8] [18]),
    .D(_4090_),
    .Y(_4847_)
);

AOI22X1 _14354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .B(_3894_),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_4848_)
);

NAND3X1 _14355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4847_),
    .B(_4848_),
    .C(_4846_),
    .Y(_4849_)
);

NOR2X1 _14356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4849_),
    .B(_4839_),
    .Y(_4850_)
);

AOI21X1 _14357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4827_),
    .B(_4850_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [18])
);

AOI22X1 _14358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [19]),
    .B(_3995__bF$buf1),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_4851_)
);

AOI22X1 _14359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .B(_4102_),
    .C(_4129_),
    .D(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_4852_)
);

INVX1 _14360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_4853_)
);

INVX1 _14361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_4854_)
);

OAI22X1 _14362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4854_),
    .B(_3890_),
    .C(_3955__bF$buf0),
    .D(_4853_),
    .Y(_4855_)
);

INVX1 _14363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_4856_)
);

INVX1 _14364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_4857_)
);

OAI22X1 _14365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4856_),
    .B(_3931__bF$buf0),
    .C(_3960_),
    .D(_4857_),
    .Y(_4858_)
);

NOR2X1 _14366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4858_),
    .B(_4855_),
    .Y(_4859_)
);

NAND3X1 _14367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4851_),
    .B(_4852_),
    .C(_4859_),
    .Y(_4860_)
);

INVX1 _14368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_4861_)
);

INVX1 _14369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_4862_)
);

OAI22X1 _14370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4862_),
    .B(_3941_),
    .C(_3978_),
    .D(_4861_),
    .Y(_4863_)
);

INVX1 _14371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_4864_)
);

INVX1 _14372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_4865_)
);

OAI22X1 _14373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .B(_4864_),
    .C(_3977__bF$buf0),
    .D(_4865_),
    .Y(_4866_)
);

NOR2X1 _14374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4863_),
    .B(_4866_),
    .Y(_4867_)
);

AOI22X1 _14375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .B(_4246_),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_4868_)
);

INVX1 _14376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [19]),
    .Y(_4869_)
);

NOR2X1 _14377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4869_),
    .B(_3944__bF$buf0),
    .Y(_4870_)
);

AOI21X1 _14378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .B(_4225_),
    .C(_4870_),
    .Y(_4871_)
);

NAND3X1 _14379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4868_),
    .B(_4871_),
    .C(_4867_),
    .Y(_4872_)
);

NOR2X1 _14380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4860_),
    .B(_4872_),
    .Y(_4873_)
);

INVX1 _14381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_4874_)
);

INVX1 _14382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_4875_)
);

OAI22X1 _14383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4874_),
    .B(_3935__bF$buf0),
    .C(_3971__bF$buf0),
    .D(_4875_),
    .Y(_4876_)
);

INVX1 _14384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_4877_)
);

INVX1 _14385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_4878_)
);

OAI22X1 _14386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4877_),
    .B(_3936__bF$buf0),
    .C(_3902__bF$buf2),
    .D(_4878_),
    .Y(_4879_)
);

NOR2X1 _14387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4879_),
    .B(_4876_),
    .Y(_4880_)
);

AOI22X1 _14388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .B(_4135_),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_4881_)
);

AOI22X1 _14389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [19]),
    .B(_3894_),
    .C(_4038__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_4882_)
);

NAND3X1 _14390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4881_),
    .B(_4882_),
    .C(_4880_),
    .Y(_4883_)
);

INVX1 _14391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_4884_)
);

INVX1 _14392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_4885_)
);

OAI22X1 _14393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf3),
    .B(_4885_),
    .C(_3909_),
    .D(_4884_),
    .Y(_4886_)
);

INVX1 _14394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_4887_)
);

INVX1 _14395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_4888_)
);

OAI22X1 _14396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf0),
    .B(_4888_),
    .C(_3954__bF$buf0),
    .D(_4887_),
    .Y(_4889_)
);

NOR2X1 _14397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4886_),
    .B(_4889_),
    .Y(_4890_)
);

AOI22X1 _14398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .B(_3885_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_4891_)
);

AOI22X1 _14399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .B(_4005__bF$buf3),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_4892_)
);

NAND3X1 _14400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4891_),
    .B(_4892_),
    .C(_4890_),
    .Y(_4893_)
);

NOR2X1 _14401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4883_),
    .B(_4893_),
    .Y(_4894_)
);

AOI21X1 _14402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4873_),
    .B(_4894_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [19])
);

AOI22X1 _14403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .B(_4154_),
    .C(_4051__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_4895_)
);

AOI22X1 _14404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[31] [20]),
    .C(\datapath_1.regfile_1.regOut[6] [20]),
    .D(_4001__bF$buf1),
    .Y(_4896_)
);

INVX1 _14405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_4897_)
);

INVX1 _14406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_4898_)
);

OAI22X1 _14407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4898_),
    .B(_3936__bF$buf4),
    .C(_3905__bF$buf2),
    .D(_4897_),
    .Y(_4899_)
);

INVX1 _14408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_4900_)
);

INVX1 _14409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_4901_)
);

OAI22X1 _14410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf2),
    .B(_4901_),
    .C(_3935__bF$buf4),
    .D(_4900_),
    .Y(_4902_)
);

NOR2X1 _14411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4899_),
    .B(_4902_),
    .Y(_4903_)
);

NAND3X1 _14412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4895_),
    .B(_4896_),
    .C(_4903_),
    .Y(_4904_)
);

AOI22X1 _14413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [20]),
    .C(\datapath_1.regfile_1.regOut[27] [20]),
    .D(_4129_),
    .Y(_4905_)
);

AOI22X1 _14414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .B(_4005__bF$buf2),
    .C(_3885_),
    .D(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_4906_)
);

INVX1 _14415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_4907_)
);

INVX1 _14416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_4908_)
);

OAI22X1 _14417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .B(_4907_),
    .C(_3977__bF$buf4),
    .D(_4908_),
    .Y(_4909_)
);

INVX1 _14418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_4910_)
);

INVX1 _14419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_4911_)
);

OAI22X1 _14420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4910_),
    .B(_3930__bF$buf2),
    .C(_3920_),
    .D(_4911_),
    .Y(_4912_)
);

NOR2X1 _14421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4909_),
    .B(_4912_),
    .Y(_4913_)
);

NAND3X1 _14422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4905_),
    .B(_4906_),
    .C(_4913_),
    .Y(_4914_)
);

NOR2X1 _14423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4904_),
    .B(_4914_),
    .Y(_4915_)
);

INVX1 _14424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_4916_)
);

INVX1 _14425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_4917_)
);

OAI22X1 _14426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4916_),
    .B(_3955__bF$buf4),
    .C(_3924__bF$buf2),
    .D(_4917_),
    .Y(_4918_)
);

INVX1 _14427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_4919_)
);

INVX1 _14428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_4920_)
);

OAI22X1 _14429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf4),
    .B(_4919_),
    .C(_3971__bF$buf4),
    .D(_4920_),
    .Y(_4921_)
);

NOR2X1 _14430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4921_),
    .B(_4918_),
    .Y(_4922_)
);

INVX1 _14431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_4923_)
);

INVX1 _14432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_4924_)
);

OAI22X1 _14433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4924_),
    .B(_3902__bF$buf1),
    .C(_3954__bF$buf4),
    .D(_4923_),
    .Y(_4925_)
);

INVX1 _14434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [20]),
    .Y(_4926_)
);

INVX1 _14435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_4927_)
);

OAI22X1 _14436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3960_),
    .B(_4927_),
    .C(_3944__bF$buf4),
    .D(_4926_),
    .Y(_4928_)
);

NOR2X1 _14437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4928_),
    .B(_4925_),
    .Y(_4929_)
);

NAND2X1 _14438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4929_),
    .B(_4922_),
    .Y(_4930_)
);

INVX1 _14439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [20]),
    .Y(_4931_)
);

INVX1 _14440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_4932_)
);

OAI22X1 _14441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4931_),
    .B(_3893__bF$buf1),
    .C(_3959_),
    .D(_4932_),
    .Y(_4933_)
);

INVX1 _14442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [20]),
    .Y(_4934_)
);

INVX1 _14443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_4935_)
);

OAI22X1 _14444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4935_),
    .B(_3941_),
    .C(_3966__bF$buf2),
    .D(_4934_),
    .Y(_4936_)
);

NOR2X1 _14445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4933_),
    .B(_4936_),
    .Y(_4937_)
);

AOI22X1 _14446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[4] [20]),
    .C(\datapath_1.regfile_1.regOut[8] [20]),
    .D(_4090_),
    .Y(_4938_)
);

AOI22X1 _14447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .B(_4135_),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_4939_)
);

NAND3X1 _14448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4938_),
    .B(_4939_),
    .C(_4937_),
    .Y(_4940_)
);

NOR2X1 _14449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4930_),
    .B(_4940_),
    .Y(_4941_)
);

AOI21X1 _14450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4941_),
    .B(_4915_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [20])
);

INVX1 _14451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_4942_)
);

INVX1 _14452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_4943_)
);

OAI22X1 _14453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4942_),
    .B(_3982__bF$buf3),
    .C(_3978_),
    .D(_4943_),
    .Y(_4944_)
);

INVX1 _14454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [21]),
    .Y(_4945_)
);

INVX1 _14455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_4946_)
);

OAI22X1 _14456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4946_),
    .B(_3909_),
    .C(_3881_),
    .D(_4945_),
    .Y(_4947_)
);

NOR2X1 _14457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4944_),
    .B(_4947_),
    .Y(_4948_)
);

AOI22X1 _14458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .B(_4102_),
    .C(_3942__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_4949_)
);

AOI22X1 _14459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [21]),
    .C(\datapath_1.regfile_1.regOut[7] [21]),
    .D(_3948_),
    .Y(_4950_)
);

NAND3X1 _14460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4949_),
    .B(_4950_),
    .C(_4948_),
    .Y(_4951_)
);

INVX1 _14461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [21]),
    .Y(_4952_)
);

INVX1 _14462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_4953_)
);

OAI22X1 _14463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .B(_4953_),
    .C(_3966__bF$buf1),
    .D(_4952_),
    .Y(_4954_)
);

INVX1 _14464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [21]),
    .Y(_4955_)
);

INVX1 _14465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_4956_)
);

OAI22X1 _14466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4956_),
    .B(_3910_),
    .C(_3944__bF$buf3),
    .D(_4955_),
    .Y(_4957_)
);

NOR2X1 _14467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4957_),
    .B(_4954_),
    .Y(_4958_)
);

INVX1 _14468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_4959_)
);

NOR2X1 _14469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4959_),
    .B(_3977__bF$buf3),
    .Y(_4960_)
);

AOI21X1 _14470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .B(_4038__bF$buf1),
    .C(_4960_),
    .Y(_4961_)
);

AOI22X1 _14471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .B(_3894_),
    .C(_4079__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_4962_)
);

NAND3X1 _14472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4961_),
    .B(_4962_),
    .C(_4958_),
    .Y(_4963_)
);

NOR2X1 _14473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4963_),
    .B(_4951_),
    .Y(_4964_)
);

INVX1 _14474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_4965_)
);

INVX1 _14475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_4966_)
);

OAI22X1 _14476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4965_),
    .B(_3890_),
    .C(_3960_),
    .D(_4966_),
    .Y(_4967_)
);

INVX1 _14477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_4968_)
);

INVX1 _14478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_4969_)
);

OAI22X1 _14479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4969_),
    .B(_3931__bF$buf3),
    .C(_3983__bF$buf3),
    .D(_4968_),
    .Y(_4970_)
);

NOR2X1 _14480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4967_),
    .B(_4970_),
    .Y(_4971_)
);

AOI22X1 _14481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .B(_3995__bF$buf4),
    .C(_3997__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_4972_)
);

AOI22X1 _14482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_4973_)
);

NAND3X1 _14483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4972_),
    .B(_4973_),
    .C(_4971_),
    .Y(_4974_)
);

INVX1 _14484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_4975_)
);

INVX1 _14485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_4976_)
);

OAI22X1 _14486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4975_),
    .B(_3902__bF$buf0),
    .C(_3971__bF$buf3),
    .D(_4976_),
    .Y(_4977_)
);

INVX1 _14487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_4978_)
);

INVX1 _14488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_4979_)
);

OAI22X1 _14489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4979_),
    .B(_3935__bF$buf3),
    .C(_3924__bF$buf1),
    .D(_4978_),
    .Y(_4980_)
);

NOR2X1 _14490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4977_),
    .B(_4980_),
    .Y(_4981_)
);

INVX1 _14491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_4982_)
);

INVX1 _14492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_4983_)
);

OAI22X1 _14493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4982_),
    .B(_3955__bF$buf3),
    .C(_3954__bF$buf3),
    .D(_4983_),
    .Y(_4984_)
);

INVX1 _14494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .Y(_4985_)
);

INVX1 _14495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_4986_)
);

OAI22X1 _14496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf2),
    .B(_4985_),
    .C(_4986_),
    .D(_3972__bF$buf3),
    .Y(_4987_)
);

NOR2X1 _14497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4987_),
    .B(_4984_),
    .Y(_4988_)
);

NAND2X1 _14498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4988_),
    .B(_4981_),
    .Y(_4989_)
);

NOR2X1 _14499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4989_),
    .B(_4974_),
    .Y(_4990_)
);

AOI21X1 _14500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4990_),
    .B(_4964_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [21])
);

INVX1 _14501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_4991_)
);

INVX1 _14502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_4992_)
);

OAI22X1 _14503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf1),
    .B(_4992_),
    .C(_3909_),
    .D(_4991_),
    .Y(_4993_)
);

INVX1 _14504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [22]),
    .Y(_4994_)
);

INVX1 _14505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_4995_)
);

OAI22X1 _14506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf2),
    .B(_4994_),
    .C(_3955__bF$buf2),
    .D(_4995_),
    .Y(_4996_)
);

NOR2X1 _14507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4993_),
    .B(_4996_),
    .Y(_4997_)
);

INVX1 _14508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [22]),
    .Y(_4998_)
);

NOR2X1 _14509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4998_),
    .B(_3944__bF$buf2),
    .Y(_4999_)
);

AOI21X1 _14510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .B(_4079__bF$buf3),
    .C(_4999_),
    .Y(_5000_)
);

AOI22X1 _14511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .B(_4135_),
    .C(_3882__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_5001_)
);

NAND3X1 _14512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5000_),
    .B(_5001_),
    .C(_4997_),
    .Y(_5002_)
);

INVX1 _14513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_5003_)
);

INVX1 _14514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_5004_)
);

OAI22X1 _14515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5004_),
    .B(_3936__bF$buf3),
    .C(_3930__bF$buf1),
    .D(_5003_),
    .Y(_5005_)
);

INVX1 _14516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_5006_)
);

INVX1 _14517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_5007_)
);

OAI22X1 _14518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5006_),
    .B(_3905__bF$buf1),
    .C(_3977__bF$buf2),
    .D(_5007_),
    .Y(_5008_)
);

NOR2X1 _14519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5005_),
    .B(_5008_),
    .Y(_5009_)
);

INVX1 _14520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_5010_)
);

NOR2X1 _14521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5010_),
    .B(_3935__bF$buf2),
    .Y(_5011_)
);

AOI21X1 _14522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .B(_3995__bF$buf3),
    .C(_5011_),
    .Y(_5012_)
);

INVX1 _14523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_5013_)
);

NOR2X1 _14524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5013_),
    .B(_3954__bF$buf2),
    .Y(_5014_)
);

AOI21X1 _14525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .B(_4115_),
    .C(_5014_),
    .Y(_5015_)
);

NAND3X1 _14526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5012_),
    .B(_5015_),
    .C(_5009_),
    .Y(_5016_)
);

NOR2X1 _14527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5002_),
    .B(_5016_),
    .Y(_5017_)
);

AOI22X1 _14528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [22]),
    .B(_4129_),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_5018_)
);

AOI22X1 _14529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .B(_3894_),
    .C(_4090_),
    .D(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_5019_)
);

INVX1 _14530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_5020_)
);

INVX1 _14531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_5021_)
);

OAI22X1 _14532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5020_),
    .B(_3916_),
    .C(_3983__bF$buf2),
    .D(_5021_),
    .Y(_5022_)
);

INVX1 _14533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_5023_)
);

INVX1 _14534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_5024_)
);

OAI22X1 _14535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5024_),
    .B(_3941_),
    .C(_3949_),
    .D(_5023_),
    .Y(_5025_)
);

NOR2X1 _14536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5025_),
    .B(_5022_),
    .Y(_5026_)
);

NAND3X1 _14537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5018_),
    .B(_5019_),
    .C(_5026_),
    .Y(_5027_)
);

AOI22X1 _14538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .B(_3891__bF$buf2),
    .C(_3998__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_5028_)
);

AOI22X1 _14539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .B(_4005__bF$buf1),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_5029_)
);

INVX1 _14540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_5030_)
);

INVX1 _14541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_5031_)
);

OAI22X1 _14542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5030_),
    .B(_3982__bF$buf2),
    .C(_3978_),
    .D(_5031_),
    .Y(_5032_)
);

INVX1 _14543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_5033_)
);

INVX1 _14544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_5034_)
);

OAI22X1 _14545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5034_),
    .B(_3971__bF$buf2),
    .C(_3924__bF$buf0),
    .D(_5033_),
    .Y(_5035_)
);

NOR2X1 _14546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5032_),
    .B(_5035_),
    .Y(_5036_)
);

NAND3X1 _14547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5028_),
    .B(_5029_),
    .C(_5036_),
    .Y(_5037_)
);

NOR2X1 _14548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5027_),
    .B(_5037_),
    .Y(_5038_)
);

AOI21X1 _14549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5017_),
    .B(_5038_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [22])
);

INVX1 _14550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_5039_)
);

INVX1 _14551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_5040_)
);

OAI22X1 _14552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5040_),
    .B(_3972__bF$buf2),
    .C(_3920_),
    .D(_5039_),
    .Y(_5041_)
);

INVX1 _14553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [23]),
    .Y(_5042_)
);

INVX1 _14554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_5043_)
);

OAI22X1 _14555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5042_),
    .B(_3884__bF$buf1),
    .C(_3959_),
    .D(_5043_),
    .Y(_5044_)
);

NOR2X1 _14556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5044_),
    .B(_5041_),
    .Y(_5045_)
);

AOI22X1 _14557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .B(_4005__bF$buf0),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_5046_)
);

AOI22X1 _14558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_5047_)
);

NAND3X1 _14559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5046_),
    .B(_5047_),
    .C(_5045_),
    .Y(_5048_)
);

AOI22X1 _14560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .B(_4225_),
    .C(_4129_),
    .D(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_5049_)
);

AOI22X1 _14561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .B(_4038__bF$buf0),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_5050_)
);

INVX1 _14562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_5051_)
);

INVX1 _14563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_5052_)
);

OAI22X1 _14564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5051_),
    .B(_3930__bF$buf0),
    .C(_3931__bF$buf2),
    .D(_5052_),
    .Y(_5053_)
);

INVX1 _14565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_5054_)
);

INVX1 _14566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_5055_)
);

OAI22X1 _14567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf3),
    .B(_5054_),
    .C(_5055_),
    .D(_3935__bF$buf1),
    .Y(_5056_)
);

NOR2X1 _14568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5053_),
    .B(_5056_),
    .Y(_5057_)
);

NAND3X1 _14569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5049_),
    .B(_5050_),
    .C(_5057_),
    .Y(_5058_)
);

NOR2X1 _14570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5058_),
    .B(_5048_),
    .Y(_5059_)
);

AOI22X1 _14571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [23]),
    .C(\datapath_1.regfile_1.regOut[6] [23]),
    .D(_4001__bF$buf0),
    .Y(_5060_)
);

AOI22X1 _14572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .B(_3942__bF$buf3),
    .C(_3995__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_5061_)
);

INVX1 _14573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_5062_)
);

INVX1 _14574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_5063_)
);

OAI22X1 _14575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5062_),
    .B(_3955__bF$buf1),
    .C(_3954__bF$buf1),
    .D(_5063_),
    .Y(_5064_)
);

INVX1 _14576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_5065_)
);

INVX1 _14577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_5066_)
);

OAI22X1 _14578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5065_),
    .B(_3890_),
    .C(_3960_),
    .D(_5066_),
    .Y(_5067_)
);

NOR2X1 _14579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5067_),
    .B(_5064_),
    .Y(_5068_)
);

NAND3X1 _14580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5060_),
    .B(_5061_),
    .C(_5068_),
    .Y(_5069_)
);

INVX1 _14581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .Y(_5070_)
);

INVX1 _14582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [23]),
    .Y(_5071_)
);

OAI22X1 _14583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5070_),
    .B(_3893__bF$buf0),
    .C(_3944__bF$buf1),
    .D(_5071_),
    .Y(_5072_)
);

INVX1 _14584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [23]),
    .Y(_5073_)
);

INVX1 _14585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_5074_)
);

OAI22X1 _14586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3881_),
    .B(_5073_),
    .C(_3971__bF$buf1),
    .D(_5074_),
    .Y(_5075_)
);

NOR2X1 _14587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5072_),
    .B(_5075_),
    .Y(_5076_)
);

INVX1 _14588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_5077_)
);

INVX1 _14589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_5078_)
);

OAI22X1 _14590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_5077_),
    .C(_3977__bF$buf1),
    .D(_5078_),
    .Y(_5079_)
);

INVX1 _14591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_5080_)
);

INVX1 _14592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_5081_)
);

OAI22X1 _14593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5081_),
    .B(_3982__bF$buf1),
    .C(_3983__bF$buf1),
    .D(_5080_),
    .Y(_5082_)
);

NOR2X1 _14594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5082_),
    .B(_5079_),
    .Y(_5083_)
);

NAND2X1 _14595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5083_),
    .B(_5076_),
    .Y(_5084_)
);

NOR2X1 _14596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5084_),
    .B(_5069_),
    .Y(_5085_)
);

AOI21X1 _14597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5085_),
    .B(_5059_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [23])
);

INVX1 _14598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [24]),
    .Y(_5086_)
);

INVX1 _14599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [24]),
    .Y(_5087_)
);

OAI22X1 _14600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5086_),
    .B(_3884__bF$buf0),
    .C(_3881_),
    .D(_5087_),
    .Y(_5088_)
);

INVX1 _14601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_5089_)
);

INVX1 _14602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_5090_)
);

OAI22X1 _14603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5089_),
    .B(_3936__bF$buf2),
    .C(_3935__bF$buf0),
    .D(_5090_),
    .Y(_5091_)
);

NOR2X1 _14604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5091_),
    .B(_5088_),
    .Y(_5092_)
);

AOI22X1 _14605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .B(_4005__bF$buf3),
    .C(_3950__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_5093_)
);

AOI22X1 _14606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [24]),
    .B(_3998__bF$buf3),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_5094_)
);

NAND3X1 _14607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5093_),
    .B(_5094_),
    .C(_5092_),
    .Y(_5095_)
);

AOI22X1 _14608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .B(_4079__bF$buf2),
    .C(_4038__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_5096_)
);

AOI22X1 _14609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .B(_3942__bF$buf2),
    .C(_3995__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_5097_)
);

INVX1 _14610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_5098_)
);

INVX1 _14611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [24]),
    .Y(_5099_)
);

OAI22X1 _14612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3893__bF$buf3),
    .B(_5099_),
    .C(_3930__bF$buf3),
    .D(_5098_),
    .Y(_5100_)
);

INVX1 _14613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_5101_)
);

INVX1 _14614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_5102_)
);

OAI22X1 _14615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5102_),
    .B(_3902__bF$buf2),
    .C(_3954__bF$buf0),
    .D(_5101_),
    .Y(_5103_)
);

NOR2X1 _14616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5100_),
    .B(_5103_),
    .Y(_5104_)
);

NAND3X1 _14617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5096_),
    .B(_5097_),
    .C(_5104_),
    .Y(_5105_)
);

NOR2X1 _14618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5095_),
    .B(_5105_),
    .Y(_5106_)
);

INVX1 _14619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_5107_)
);

INVX1 _14620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_5108_)
);

OAI22X1 _14621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf0),
    .B(_5108_),
    .C(_3909_),
    .D(_5107_),
    .Y(_5109_)
);

INVX1 _14622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_5110_)
);

INVX1 _14623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_5111_)
);

OAI22X1 _14624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5111_),
    .B(_3971__bF$buf0),
    .C(_3924__bF$buf3),
    .D(_5110_),
    .Y(_5112_)
);

NOR2X1 _14625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5109_),
    .B(_5112_),
    .Y(_5113_)
);

AOI22X1 _14626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[4] [24]),
    .C(\datapath_1.regfile_1.regOut[8] [24]),
    .D(_4090_),
    .Y(_5114_)
);

INVX1 _14627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_5115_)
);

NOR2X1 _14628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5115_),
    .B(_3955__bF$buf0),
    .Y(_5116_)
);

AOI21X1 _14629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .B(_4246_),
    .C(_5116_),
    .Y(_5117_)
);

NAND3X1 _14630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5114_),
    .B(_5117_),
    .C(_5113_),
    .Y(_5118_)
);

INVX1 _14631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [24]),
    .Y(_5119_)
);

INVX1 _14632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [24]),
    .Y(_5120_)
);

OAI22X1 _14633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf1),
    .B(_5119_),
    .C(_3966__bF$buf0),
    .D(_5120_),
    .Y(_5121_)
);

INVX1 _14634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [24]),
    .Y(_5122_)
);

INVX1 _14635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_5123_)
);

OAI22X1 _14636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972__bF$buf1),
    .B(_5123_),
    .C(_3944__bF$buf0),
    .D(_5122_),
    .Y(_5124_)
);

NOR2X1 _14637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5124_),
    .B(_5121_),
    .Y(_5125_)
);

INVX1 _14638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_5126_)
);

INVX1 _14639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_5127_)
);

OAI22X1 _14640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_5126_),
    .C(_3977__bF$buf0),
    .D(_5127_),
    .Y(_5128_)
);

INVX1 _14641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_5129_)
);

INVX1 _14642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_5130_)
);

OAI22X1 _14643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5130_),
    .B(_3982__bF$buf0),
    .C(_3983__bF$buf0),
    .D(_5129_),
    .Y(_5131_)
);

NOR2X1 _14644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5131_),
    .B(_5128_),
    .Y(_5132_)
);

NAND2X1 _14645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5125_),
    .B(_5132_),
    .Y(_5133_)
);

NOR2X1 _14646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5133_),
    .B(_5118_),
    .Y(_5134_)
);

AOI21X1 _14647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5106_),
    .B(_5134_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd2 [24])
);

INVX1 _14648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_5135_)
);

INVX1 _14649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_5136_)
);

OAI22X1 _14650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5135_),
    .B(_3890_),
    .C(_3960_),
    .D(_5136_),
    .Y(_5137_)
);

INVX1 _14651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .Y(_5138_)
);

INVX1 _14652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [25]),
    .Y(_5139_)
);

OAI22X1 _14653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5138_),
    .B(_3893__bF$buf2),
    .C(_3944__bF$buf4),
    .D(_5139_),
    .Y(_5140_)
);

NOR2X1 _14654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5137_),
    .B(_5140_),
    .Y(_5141_)
);

AOI22X1 _14655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .B(_4629_),
    .C(_4246_),
    .D(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_5142_)
);

AOI22X1 _14656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .B(_4129_),
    .C(_4079__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_5143_)
);

NAND3X1 _14657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5142_),
    .B(_5143_),
    .C(_5141_),
    .Y(_5144_)
);

AOI22X1 _14658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .B(_4005__bF$buf2),
    .C(_4225_),
    .D(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_5145_)
);

AOI22X1 _14659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .B(_3942__bF$buf1),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_5146_)
);

INVX1 _14660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [25]),
    .Y(_5147_)
);

INVX1 _14661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_5148_)
);

OAI22X1 _14662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5148_),
    .B(_3931__bF$buf1),
    .C(_3966__bF$buf3),
    .D(_5147_),
    .Y(_5149_)
);

INVX1 _14663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_5150_)
);

INVX1 _14664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_5151_)
);

OAI22X1 _14665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf1),
    .B(_5150_),
    .C(_5151_),
    .D(_3935__bF$buf4),
    .Y(_5152_)
);

NOR2X1 _14666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5152_),
    .B(_5149_),
    .Y(_5153_)
);

NAND3X1 _14667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5145_),
    .B(_5146_),
    .C(_5153_),
    .Y(_5154_)
);

NOR2X1 _14668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5144_),
    .B(_5154_),
    .Y(_5155_)
);

AOI22X1 _14669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .B(_4102_),
    .C(_4001__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_5156_)
);

INVX1 _14670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_5157_)
);

NOR2X1 _14671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5157_),
    .B(_3983__bF$buf4),
    .Y(_5158_)
);

AOI21X1 _14672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .B(_4038__bF$buf2),
    .C(_5158_),
    .Y(_5159_)
);

INVX1 _14673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_5160_)
);

INVX1 _14674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_5161_)
);

OAI22X1 _14675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5160_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf4),
    .D(_5161_),
    .Y(_5162_)
);

INVX1 _14676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_5163_)
);

INVX1 _14677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_5164_)
);

OAI22X1 _14678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf3),
    .B(_5163_),
    .C(_3977__bF$buf4),
    .D(_5164_),
    .Y(_5165_)
);

NOR2X1 _14679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5165_),
    .B(_5162_),
    .Y(_5166_)
);

NAND3X1 _14680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5156_),
    .B(_5159_),
    .C(_5166_),
    .Y(_5167_)
);

INVX1 _14681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_5168_)
);

INVX1 _14682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_5169_)
);

OAI22X1 _14683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5169_),
    .B(_3949_),
    .C(_3978_),
    .D(_5168_),
    .Y(_5170_)
);

INVX1 _14684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_5171_)
);

INVX1 _14685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_5172_)
);

OAI22X1 _14686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3982__bF$buf3),
    .B(_5171_),
    .C(_3971__bF$buf4),
    .D(_5172_),
    .Y(_5173_)
);

NOR2X1 _14687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5170_),
    .B(_5173_),
    .Y(_5174_)
);

AOI22X1 _14688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .B(_3995__bF$buf0),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_5175_)
);

AOI22X1 _14689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [25]),
    .C(\datapath_1.regfile_1.regOut[18] [25]),
    .D(_4135_),
    .Y(_5176_)
);

NAND3X1 _14690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5175_),
    .B(_5176_),
    .C(_5174_),
    .Y(_5177_)
);

NOR2X1 _14691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5177_),
    .B(_5167_),
    .Y(_5178_)
);

AOI21X1 _14692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5155_),
    .B(_5178_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd2 [25])
);

AOI22X1 _14693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .B(_4154_),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_5179_)
);

AOI22X1 _14694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3995__bF$buf4),
    .B(\datapath_1.regfile_1.regOut[31] [26]),
    .C(\datapath_1.regfile_1.regOut[6] [26]),
    .D(_4001__bF$buf2),
    .Y(_5180_)
);

INVX1 _14695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_5181_)
);

INVX1 _14696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_5182_)
);

OAI22X1 _14697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5182_),
    .B(_3936__bF$buf1),
    .C(_3905__bF$buf0),
    .D(_5181_),
    .Y(_5183_)
);

INVX1 _14698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_5184_)
);

INVX1 _14699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_5185_)
);

OAI22X1 _14700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf2),
    .B(_5185_),
    .C(_3935__bF$buf3),
    .D(_5184_),
    .Y(_5186_)
);

NOR2X1 _14701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5183_),
    .B(_5186_),
    .Y(_5187_)
);

NAND3X1 _14702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5179_),
    .B(_5180_),
    .C(_5187_),
    .Y(_5188_)
);

INVX1 _14703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [26]),
    .Y(_5189_)
);

INVX1 _14704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_5190_)
);

OAI22X1 _14705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .B(_5190_),
    .C(_5189_),
    .D(_3967__bF$buf0),
    .Y(_5191_)
);

INVX1 _14706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [26]),
    .Y(_5192_)
);

INVX1 _14707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_5193_)
);

OAI22X1 _14708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5193_),
    .B(_3910_),
    .C(_3884__bF$buf3),
    .D(_5192_),
    .Y(_5194_)
);

NOR2X1 _14709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5194_),
    .B(_5191_),
    .Y(_5195_)
);

INVX1 _14710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_5196_)
);

NOR2X1 _14711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5196_),
    .B(_3977__bF$buf3),
    .Y(_5197_)
);

AOI21X1 _14712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .B(_4038__bF$buf1),
    .C(_5197_),
    .Y(_5198_)
);

AOI22X1 _14713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .B(_4102_),
    .C(_4079__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_5199_)
);

NAND3X1 _14714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5199_),
    .B(_5198_),
    .C(_5195_),
    .Y(_5200_)
);

NOR2X1 _14715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5200_),
    .B(_5188_),
    .Y(_5201_)
);

INVX1 _14716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_5202_)
);

INVX1 _14717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_5203_)
);

OAI22X1 _14718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5203_),
    .B(_3954__bF$buf3),
    .C(_3924__bF$buf2),
    .D(_5202_),
    .Y(_5204_)
);

INVX1 _14719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_5205_)
);

INVX1 _14720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_5206_)
);

OAI22X1 _14721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf3),
    .B(_5205_),
    .C(_3971__bF$buf3),
    .D(_5206_),
    .Y(_5207_)
);

NOR2X1 _14722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5207_),
    .B(_5204_),
    .Y(_5208_)
);

INVX1 _14723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_5209_)
);

INVX1 _14724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_5210_)
);

OAI22X1 _14725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf0),
    .B(_5210_),
    .C(_5209_),
    .D(_3955__bF$buf3),
    .Y(_5211_)
);

INVX1 _14726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_5212_)
);

INVX1 _14727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_5213_)
);

OAI22X1 _14728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5213_),
    .B(_3960_),
    .C(_3959_),
    .D(_5212_),
    .Y(_5214_)
);

NOR2X1 _14729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5211_),
    .B(_5214_),
    .Y(_5215_)
);

NAND2X1 _14730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5215_),
    .B(_5208_),
    .Y(_5216_)
);

INVX1 _14731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .Y(_5217_)
);

INVX1 _14732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [26]),
    .Y(_5218_)
);

OAI22X1 _14733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5217_),
    .B(_3893__bF$buf1),
    .C(_3944__bF$buf3),
    .D(_5218_),
    .Y(_5219_)
);

INVX1 _14734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [26]),
    .Y(_5220_)
);

INVX1 _14735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_5221_)
);

OAI22X1 _14736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5221_),
    .B(_3941_),
    .C(_3966__bF$buf2),
    .D(_5220_),
    .Y(_5222_)
);

NOR2X1 _14737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5219_),
    .B(_5222_),
    .Y(_5223_)
);

AOI22X1 _14738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[4] [26]),
    .C(\datapath_1.regfile_1.regOut[8] [26]),
    .D(_4090_),
    .Y(_5224_)
);

AOI22X1 _14739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .B(_4135_),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_5225_)
);

NAND3X1 _14740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5224_),
    .B(_5225_),
    .C(_5223_),
    .Y(_5226_)
);

NOR2X1 _14741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5216_),
    .B(_5226_),
    .Y(_5227_)
);

AOI21X1 _14742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5201_),
    .B(_5227_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd2 [26])
);

INVX1 _14743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_5228_)
);

NOR2X1 _14744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5228_),
    .B(_3977__bF$buf2),
    .Y(_5229_)
);

AOI21X1 _14745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [27]),
    .B(_3950__bF$buf1),
    .C(_5229_),
    .Y(_5230_)
);

AOI22X1 _14746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .B(_3894_),
    .C(_4051__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_5231_)
);

INVX1 _14747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_5232_)
);

INVX1 _14748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_5233_)
);

OAI22X1 _14749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5233_),
    .B(_3936__bF$buf0),
    .C(_3905__bF$buf3),
    .D(_5232_),
    .Y(_5234_)
);

INVX1 _14750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [27]),
    .Y(_5235_)
);

INVX1 _14751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_5236_)
);

OAI22X1 _14752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967__bF$buf3),
    .B(_5235_),
    .C(_3935__bF$buf2),
    .D(_5236_),
    .Y(_5237_)
);

NOR2X1 _14753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5234_),
    .B(_5237_),
    .Y(_5238_)
);

NAND3X1 _14754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5231_),
    .B(_5230_),
    .C(_5238_),
    .Y(_5239_)
);

INVX1 _14755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_5240_)
);

INVX1 _14756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_5241_)
);

OAI22X1 _14757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5240_),
    .B(_3916_),
    .C(_3983__bF$buf2),
    .D(_5241_),
    .Y(_5242_)
);

INVX1 _14758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_5243_)
);

INVX1 _14759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_5244_)
);

OAI22X1 _14760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5244_),
    .B(_3972__bF$buf0),
    .C(_3920_),
    .D(_5243_),
    .Y(_5245_)
);

NOR2X1 _14761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5242_),
    .B(_5245_),
    .Y(_5246_)
);

AOI22X1 _14762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .B(_3942__bF$buf0),
    .C(_4154_),
    .D(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_5247_)
);

AOI22X1 _14763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[29] [27]),
    .C(\datapath_1.regfile_1.regOut[1] [27]),
    .D(_3997__bF$buf1),
    .Y(_5248_)
);

NAND3X1 _14764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5247_),
    .B(_5248_),
    .C(_5246_),
    .Y(_5249_)
);

NOR2X1 _14765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5239_),
    .B(_5249_),
    .Y(_5250_)
);

INVX1 _14766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_5251_)
);

INVX1 _14767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_5252_)
);

OAI22X1 _14768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902__bF$buf3),
    .B(_5252_),
    .C(_5251_),
    .D(_3955__bF$buf2),
    .Y(_5253_)
);

INVX1 _14769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [27]),
    .Y(_5254_)
);

INVX1 _14770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_5255_)
);

OAI22X1 _14771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5254_),
    .B(_3884__bF$buf2),
    .C(_3924__bF$buf1),
    .D(_5255_),
    .Y(_5256_)
);

NOR2X1 _14772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5253_),
    .B(_5256_),
    .Y(_5257_)
);

AOI22X1 _14773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .B(_3891__bF$buf3),
    .C(_3998__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_5258_)
);

AOI22X1 _14774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .B(_4005__bF$buf1),
    .C(_3995__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_5259_)
);

NAND3X1 _14775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5258_),
    .B(_5259_),
    .C(_5257_),
    .Y(_5260_)
);

INVX1 _14776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_5261_)
);

INVX1 _14777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [27]),
    .Y(_5262_)
);

OAI22X1 _14778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5261_),
    .B(_3930__bF$buf2),
    .C(_3966__bF$buf1),
    .D(_5262_),
    .Y(_5263_)
);

INVX1 _14779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [27]),
    .Y(_5264_)
);

INVX1 _14780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_5265_)
);

OAI22X1 _14781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3909_),
    .B(_5265_),
    .C(_5264_),
    .D(_3944__bF$buf2),
    .Y(_5266_)
);

NOR2X1 _14782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5266_),
    .B(_5263_),
    .Y(_5267_)
);

AOI22X1 _14783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .B(_4090_),
    .C(_3948_),
    .D(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_5268_)
);

INVX1 _14784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_5269_)
);

NOR2X1 _14785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5269_),
    .B(_3971__bF$buf2),
    .Y(_5270_)
);

INVX1 _14786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_5271_)
);

NOR2X1 _14787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5271_),
    .B(_3954__bF$buf2),
    .Y(_5272_)
);

NOR2X1 _14788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5270_),
    .B(_5272_),
    .Y(_5273_)
);

NAND3X1 _14789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5268_),
    .B(_5273_),
    .C(_5267_),
    .Y(_5274_)
);

NOR2X1 _14790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5274_),
    .B(_5260_),
    .Y(_5275_)
);

AOI21X1 _14791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5250_),
    .B(_5275_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd2 [27])
);

AOI22X1 _14792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .B(_4005__bF$buf0),
    .C(_3998__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_5276_)
);

AOI22X1 _14793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4154_),
    .B(\datapath_1.regfile_1.regOut[14] [28]),
    .C(\datapath_1.regfile_1.regOut[31] [28]),
    .D(_3995__bF$buf2),
    .Y(_5277_)
);

INVX1 _14794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_5278_)
);

INVX1 _14795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_5279_)
);

OAI22X1 _14796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5279_),
    .B(_3936__bF$buf4),
    .C(_3905__bF$buf2),
    .D(_5278_),
    .Y(_5280_)
);

INVX1 _14797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [28]),
    .Y(_5281_)
);

INVX1 _14798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_5282_)
);

OAI22X1 _14799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935__bF$buf1),
    .B(_5282_),
    .C(_5281_),
    .D(_3944__bF$buf1),
    .Y(_5283_)
);

NOR2X1 _14800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5280_),
    .B(_5283_),
    .Y(_5284_)
);

NAND3X1 _14801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5276_),
    .B(_5277_),
    .C(_5284_),
    .Y(_5285_)
);

AOI22X1 _14802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .B(_4038__bF$buf0),
    .C(_4079__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_5286_)
);

AOI22X1 _14803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4129_),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .C(\datapath_1.regfile_1.regOut[18] [28]),
    .D(_4135_),
    .Y(_5287_)
);

INVX1 _14804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_5288_)
);

INVX1 _14805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_5289_)
);

OAI22X1 _14806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5289_),
    .B(_3949_),
    .C(_3983__bF$buf1),
    .D(_5288_),
    .Y(_5290_)
);

INVX1 _14807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [28]),
    .Y(_5291_)
);

INVX1 _14808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_5292_)
);

OAI22X1 _14809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf1),
    .B(_5291_),
    .C(_3977__bF$buf1),
    .D(_5292_),
    .Y(_5293_)
);

NOR2X1 _14810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5290_),
    .B(_5293_),
    .Y(_5294_)
);

NAND3X1 _14811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5286_),
    .B(_5287_),
    .C(_5294_),
    .Y(_5295_)
);

NOR2X1 _14812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5285_),
    .B(_5295_),
    .Y(_5296_)
);

INVX1 _14813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_5297_)
);

INVX1 _14814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_5298_)
);

OAI22X1 _14815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5298_),
    .B(_3902__bF$buf2),
    .C(_3954__bF$buf1),
    .D(_5297_),
    .Y(_5299_)
);

INVX1 _14816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_5300_)
);

INVX1 _14817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_5301_)
);

OAI22X1 _14818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5300_),
    .B(_3930__bF$buf1),
    .C(_3924__bF$buf0),
    .D(_5301_),
    .Y(_5302_)
);

NOR2X1 _14819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5299_),
    .B(_5302_),
    .Y(_5303_)
);

AOI22X1 _14820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3948_),
    .B(\datapath_1.regfile_1.regOut[7] [28]),
    .C(\datapath_1.regfile_1.regOut[6] [28]),
    .D(_4001__bF$buf1),
    .Y(_5304_)
);

AOI22X1 _14821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[29] [28]),
    .C(\datapath_1.regfile_1.regOut[13] [28]),
    .D(_4051__bF$buf1),
    .Y(_5305_)
);

NAND3X1 _14822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5304_),
    .B(_5305_),
    .C(_5303_),
    .Y(_5306_)
);

AOI22X1 _14823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [28]),
    .B(_3894_),
    .C(_3997__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_5307_)
);

AOI22X1 _14824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .B(_3942__bF$buf3),
    .C(_4040_),
    .D(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_5308_)
);

INVX1 _14825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_5309_)
);

INVX1 _14826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_5310_)
);

OAI22X1 _14827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3890_),
    .B(_5310_),
    .C(_5309_),
    .D(_3931__bF$buf0),
    .Y(_5311_)
);

INVX1 _14828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_5312_)
);

INVX1 _14829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_5313_)
);

OAI22X1 _14830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5312_),
    .B(_3955__bF$buf1),
    .C(_3971__bF$buf1),
    .D(_5313_),
    .Y(_5314_)
);

NOR2X1 _14831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5311_),
    .B(_5314_),
    .Y(_5315_)
);

NAND3X1 _14832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5307_),
    .B(_5308_),
    .C(_5315_),
    .Y(_5316_)
);

NOR2X1 _14833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5316_),
    .B(_5306_),
    .Y(_5317_)
);

AOI21X1 _14834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5296_),
    .B(_5317_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd2 [28])
);

AOI22X1 _14835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [29]),
    .B(_3942__bF$buf2),
    .C(_3891__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_5318_)
);

INVX1 _14836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_5319_)
);

NOR2X1 _14837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5319_),
    .B(_3935__bF$buf0),
    .Y(_5320_)
);

AOI21X1 _14838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .B(_4115_),
    .C(_5320_),
    .Y(_5321_)
);

INVX1 _14839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [29]),
    .Y(_5322_)
);

INVX1 _14840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_5323_)
);

OAI22X1 _14841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5322_),
    .B(_3944__bF$buf0),
    .C(_3954__bF$buf0),
    .D(_5323_),
    .Y(_5324_)
);

INVX1 _14842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [29]),
    .Y(_5325_)
);

INVX1 _14843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_5326_)
);

OAI22X1 _14844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5325_),
    .B(_3893__bF$buf0),
    .C(_3959_),
    .D(_5326_),
    .Y(_5327_)
);

NOR2X1 _14845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5327_),
    .B(_5324_),
    .Y(_5328_)
);

NAND3X1 _14846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5318_),
    .B(_5321_),
    .C(_5328_),
    .Y(_5329_)
);

AOI22X1 _14847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .B(_4090_),
    .C(_3998__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_5330_)
);

INVX1 _14848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_5331_)
);

NOR2X1 _14849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5331_),
    .B(_3971__bF$buf0),
    .Y(_5332_)
);

AOI21X1 _14850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .B(_4225_),
    .C(_5332_),
    .Y(_5333_)
);

INVX1 _14851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_5334_)
);

INVX1 _14852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_5335_)
);

OAI22X1 _14853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5335_),
    .B(_3936__bF$buf3),
    .C(_3955__bF$buf0),
    .D(_5334_),
    .Y(_5336_)
);

INVX1 _14854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_5337_)
);

INVX1 _14855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_5338_)
);

OAI22X1 _14856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3905__bF$buf1),
    .B(_5338_),
    .C(_3930__bF$buf0),
    .D(_5337_),
    .Y(_5339_)
);

NOR2X1 _14857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5339_),
    .B(_5336_),
    .Y(_5340_)
);

NAND3X1 _14858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5330_),
    .B(_5333_),
    .C(_5340_),
    .Y(_5341_)
);

NOR2X1 _14859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5341_),
    .B(_5329_),
    .Y(_5342_)
);

INVX1 _14860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_5343_)
);

INVX1 _14861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_5344_)
);

OAI22X1 _14862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5344_),
    .B(_3982__bF$buf2),
    .C(_3983__bF$buf0),
    .D(_5343_),
    .Y(_5345_)
);

INVX1 _14863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_5346_)
);

INVX1 _14864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_5347_)
);

OAI22X1 _14865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5346_),
    .B(_3910_),
    .C(_3977__bF$buf0),
    .D(_5347_),
    .Y(_5348_)
);

NOR2X1 _14866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5345_),
    .B(_5348_),
    .Y(_5349_)
);

AOI22X1 _14867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [29]),
    .B(_4038__bF$buf3),
    .C(_4079__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_5350_)
);

AOI22X1 _14868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(\datapath_1.regfile_1.regOut[30] [29]),
    .C(\datapath_1.regfile_1.regOut[18] [29]),
    .D(_4135_),
    .Y(_5351_)
);

NAND3X1 _14869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5350_),
    .B(_5351_),
    .C(_5349_),
    .Y(_5352_)
);

INVX1 _14870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [29]),
    .Y(_5353_)
);

INVX1 _14871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_5354_)
);

OAI22X1 _14872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf1),
    .B(_5354_),
    .C(_3966__bF$buf0),
    .D(_5353_),
    .Y(_5355_)
);

INVX1 _14873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [29]),
    .Y(_5356_)
);

INVX1 _14874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_5357_)
);

OAI22X1 _14875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5356_),
    .B(_3967__bF$buf2),
    .C(_3978_),
    .D(_5357_),
    .Y(_5358_)
);

NOR2X1 _14876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5358_),
    .B(_5355_),
    .Y(_5359_)
);

AOI22X1 _14877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[11] [29]),
    .C(\datapath_1.regfile_1.regOut[31] [29]),
    .D(_3995__bF$buf1),
    .Y(_5360_)
);

AOI22X1 _14878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .B(_4001__bF$buf0),
    .C(_3882__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_5361_)
);

NAND3X1 _14879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5360_),
    .B(_5361_),
    .C(_5359_),
    .Y(_5362_)
);

NOR2X1 _14880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5362_),
    .B(_5352_),
    .Y(_5363_)
);

AOI21X1 _14881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5342_),
    .B(_5363_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd2 [29])
);

INVX1 _14882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [30]),
    .Y(_5364_)
);

INVX1 _14883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [30]),
    .Y(_5365_)
);

OAI22X1 _14884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf0),
    .B(_5364_),
    .C(_5365_),
    .D(_3925_),
    .Y(_5366_)
);

INVX1 _14885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .Y(_5367_)
);

INVX1 _14886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_5368_)
);

OAI22X1 _14887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5367_),
    .B(_3967__bF$buf1),
    .C(_3920_),
    .D(_5368_),
    .Y(_5369_)
);

NOR2X1 _14888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5366_),
    .B(_5369_),
    .Y(_5370_)
);

AOI22X1 _14889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .B(_4246_),
    .C(_4115_),
    .D(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_5371_)
);

AOI22X1 _14890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .B(_3942__bF$buf1),
    .C(_3950__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_5372_)
);

NAND3X1 _14891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5371_),
    .B(_5372_),
    .C(_5370_),
    .Y(_5373_)
);

INVX1 _14892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [30]),
    .Y(_5374_)
);

INVX1 _14893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_5375_)
);

OAI22X1 _14894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5374_),
    .B(_3966__bF$buf3),
    .C(_3924__bF$buf3),
    .D(_5375_),
    .Y(_5376_)
);

INVX1 _14895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_5377_)
);

INVX1 _14896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_5378_)
);

OAI22X1 _14897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .B(_5377_),
    .C(_5378_),
    .D(_3972__bF$buf3),
    .Y(_5379_)
);

NOR2X1 _14898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5379_),
    .B(_5376_),
    .Y(_5380_)
);

INVX1 _14899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_5381_)
);

NAND2X1 _14900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .B(_4102_),
    .Y(_5382_)
);

OAI21X1 _14901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5381_),
    .B(_3931__bF$buf3),
    .C(_5382_),
    .Y(_5383_)
);

INVX1 _14902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_5384_)
);

INVX1 _14903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_5385_)
);

OAI22X1 _14904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5384_),
    .B(_3936__bF$buf2),
    .C(_3935__bF$buf4),
    .D(_5385_),
    .Y(_5386_)
);

NOR2X1 _14905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5386_),
    .B(_5383_),
    .Y(_5387_)
);

NAND2X1 _14906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5380_),
    .B(_5387_),
    .Y(_5388_)
);

NOR2X1 _14907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5388_),
    .B(_5373_),
    .Y(_5389_)
);

AOI22X1 _14908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [30]),
    .B(_4001__bF$buf3),
    .C(_3882__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_5390_)
);

AOI22X1 _14909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [30]),
    .B(_3891__bF$buf1),
    .C(_3998__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_5391_)
);

INVX1 _14910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_5392_)
);

INVX1 _14911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_5393_)
);

OAI22X1 _14912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5392_),
    .B(_3955__bF$buf4),
    .C(_3954__bF$buf4),
    .D(_5393_),
    .Y(_5394_)
);

INVX1 _14913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_5395_)
);

INVX1 _14914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_5396_)
);

OAI22X1 _14915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf0),
    .B(_5395_),
    .C(_3977__bF$buf4),
    .D(_5396_),
    .Y(_5397_)
);

NOR2X1 _14916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5397_),
    .B(_5394_),
    .Y(_5398_)
);

NAND3X1 _14917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5390_),
    .B(_5391_),
    .C(_5398_),
    .Y(_5399_)
);

INVX1 _14918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [30]),
    .Y(_5400_)
);

INVX1 _14919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [30]),
    .Y(_5401_)
);

OAI22X1 _14920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5400_),
    .B(_3893__bF$buf3),
    .C(_3944__bF$buf4),
    .D(_5401_),
    .Y(_5402_)
);

INVX1 _14921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_5403_)
);

INVX1 _14922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_5404_)
);

OAI22X1 _14923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3983__bF$buf4),
    .B(_5403_),
    .C(_3971__bF$buf4),
    .D(_5404_),
    .Y(_5405_)
);

NOR2X1 _14924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5402_),
    .B(_5405_),
    .Y(_5406_)
);

AOI22X1 _14925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .B(_4154_),
    .C(_4051__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_5407_)
);

AOI22X1 _14926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .B(_4005__bF$buf3),
    .C(_3997__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_5408_)
);

NAND3X1 _14927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5407_),
    .B(_5408_),
    .C(_5406_),
    .Y(_5409_)
);

NOR2X1 _14928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5399_),
    .B(_5409_),
    .Y(_5410_)
);

AOI21X1 _14929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5410_),
    .B(_5389_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd2 [30])
);

AOI22X1 _14930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .B(_4225_),
    .C(_4051__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_5411_)
);

AOI22X1 _14931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .B(_4005__bF$buf2),
    .C(_4135_),
    .D(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_5412_)
);

INVX1 _14932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[26] [31]),
    .Y(_5413_)
);

INVX1 _14933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_5414_)
);

OAI22X1 _14934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5414_),
    .B(_3936__bF$buf1),
    .C(_3944__bF$buf3),
    .D(_5413_),
    .Y(_5415_)
);

INVX1 _14935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_5416_)
);

INVX1 _14936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_5417_)
);

OAI22X1 _14937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5417_),
    .B(_3890_),
    .C(_3954__bF$buf3),
    .D(_5416_),
    .Y(_5418_)
);

NOR2X1 _14938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5415_),
    .B(_5418_),
    .Y(_5419_)
);

NAND3X1 _14939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5411_),
    .B(_5412_),
    .C(_5419_),
    .Y(_5420_)
);

INVX1 _14940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_5421_)
);

NOR2X1 _14941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5421_),
    .B(_3955__bF$buf3),
    .Y(_5422_)
);

AOI21X1 _14942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .B(_3894_),
    .C(_5422_),
    .Y(_5423_)
);

AOI22X1 _14943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [31]),
    .B(_3998__bF$buf2),
    .C(_3997__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_5424_)
);

INVX1 _14944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [31]),
    .Y(_5425_)
);

INVX1 _14945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_5426_)
);

OAI22X1 _14946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884__bF$buf3),
    .B(_5425_),
    .C(_5426_),
    .D(_3916_),
    .Y(_5427_)
);

INVX1 _14947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_5428_)
);

INVX1 _14948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_5429_)
);

OAI22X1 _14949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5428_),
    .B(_3930__bF$buf3),
    .C(_3971__bF$buf3),
    .D(_5429_),
    .Y(_5430_)
);

NOR2X1 _14950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5427_),
    .B(_5430_),
    .Y(_5431_)
);

NAND3X1 _14951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5423_),
    .B(_5424_),
    .C(_5431_),
    .Y(_5432_)
);

NOR2X1 _14952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .B(_5420_),
    .Y(_5433_)
);

INVX1 _14953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_5434_)
);

NOR2X1 _14954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .B(_3983__bF$buf3),
    .Y(_5435_)
);

AOI21X1 _14955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [31]),
    .B(_4154_),
    .C(_5435_),
    .Y(_5436_)
);

AOI22X1 _14956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4129_),
    .B(\datapath_1.regfile_1.regOut[27] [31]),
    .C(\datapath_1.regfile_1.regOut[31] [31]),
    .D(_3995__bF$buf0),
    .Y(_5437_)
);

INVX1 _14957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_5438_)
);

INVX1 _14958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_5439_)
);

OAI22X1 _14959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3947__bF$buf3),
    .B(_5439_),
    .C(_3909_),
    .D(_5438_),
    .Y(_5440_)
);

INVX1 _14960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_5441_)
);

INVX1 _14961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_5442_)
);

OAI22X1 _14962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5441_),
    .B(_3905__bF$buf0),
    .C(_3977__bF$buf3),
    .D(_5442_),
    .Y(_5443_)
);

NOR2X1 _14963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .B(_5443_),
    .Y(_5444_)
);

NAND3X1 _14964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .B(_5437_),
    .C(_5444_),
    .Y(_5445_)
);

AOI22X1 _14965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [31]),
    .B(_3950__bF$buf2),
    .C(_3882__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_5446_)
);

INVX1 _14966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_5447_)
);

NOR2X1 _14967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5447_),
    .B(_3935__bF$buf3),
    .Y(_5448_)
);

AOI21X1 _14968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [31]),
    .B(_4079__bF$buf1),
    .C(_5448_),
    .Y(_5449_)
);

INVX1 _14969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [31]),
    .Y(_5450_)
);

INVX1 _14970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_5451_)
);

OAI22X1 _14971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5451_),
    .B(_3931__bF$buf2),
    .C(_3966__bF$buf2),
    .D(_5450_),
    .Y(_5452_)
);

INVX1 _14972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_5453_)
);

INVX1 _14973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_5454_)
);

OAI22X1 _14974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3941_),
    .B(_5454_),
    .C(_3902__bF$buf1),
    .D(_5453_),
    .Y(_5455_)
);

NOR2X1 _14975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5455_),
    .B(_5452_),
    .Y(_5456_)
);

NAND3X1 _14976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .B(_5449_),
    .C(_5456_),
    .Y(_5457_)
);

NOR2X1 _14977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5457_),
    .B(_5445_),
    .Y(_5458_)
);

AOI21X1 _14978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458_),
    .B(_5433_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd2 [31])
);

INVX8 _14979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .Y(_5459_)
);

INVX2 _14980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [23]),
    .Y(_5460_)
);

NOR2X1 _14981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(_5460_),
    .Y(_5461_)
);

AND2X2 _14982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5462_)
);

NAND3X1 _14983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf3),
    .B(_5462_),
    .C(_5461_),
    .Y(_5463_)
);

INVX1 _14984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .Y(_5464_)
);

NOR2X1 _14985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [25]),
    .B(_5464_),
    .Y(_5465_)
);

NAND3X1 _14986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5461_),
    .C(_5465_),
    .Y(_5466_)
);

OAI22X1 _14987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf3),
    .B(_3975_),
    .C(_5466__bF$buf4),
    .D(_3965_),
    .Y(_5467_)
);

AND2X2 _14988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5468_)
);

NAND3X1 _14989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf2),
    .B(_5462_),
    .C(_5468_),
    .Y(_5469_)
);

INVX2 _14990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [25]),
    .Y(_5470_)
);

NOR2X1 _14991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .B(_5470_),
    .Y(_5471_)
);

NAND3X1 _14992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5461_),
    .C(_5471__bF$buf5),
    .Y(_5472_)
);

OAI22X1 _14993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3897_),
    .B(_5469__bF$buf3),
    .C(_5472__bF$buf3),
    .D(_3953_),
    .Y(_5473_)
);

NOR2X1 _14994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5473_),
    .B(_5467_),
    .Y(_5474_)
);

INVX2 _14995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .Y(_5475_)
);

NOR2X1 _14996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [23]),
    .B(_5475_),
    .Y(_5476_)
);

NOR2X1 _14997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5477_)
);

NAND3X1 _14998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf1),
    .B(_5477_),
    .C(_5476_),
    .Y(_5478_)
);

INVX4 _14999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .Y(_5479_)
);

NAND3X1 _15000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5462_),
    .C(_5476_),
    .Y(_5480_)
);

INVX4 _15001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .Y(_5481_)
);

AOI22X1 _15002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [0]),
    .C(\datapath_1.regfile_1.regOut[30] [0]),
    .D(_5481_),
    .Y(_5482_)
);

NAND3X1 _15003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(_5465_),
    .C(_5476_),
    .Y(_5483_)
);

INVX2 _15004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483__bF$buf4),
    .Y(_5484_)
);

NAND3X1 _15005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5462_),
    .C(_5461_),
    .Y(_5485_)
);

INVX4 _15006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf4),
    .Y(_5486_)
);

AOI22X1 _15007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .B(\datapath_1.regfile_1.regOut[29] [0]),
    .C(\datapath_1.regfile_1.regOut[26] [0]),
    .D(_5484_),
    .Y(_5487_)
);

NAND3X1 _15008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .B(_5487_),
    .C(_5474_),
    .Y(_5488_)
);

NAND3X1 _15009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf0),
    .B(_5468_),
    .C(_5471__bF$buf4),
    .Y(_5489_)
);

INVX8 _15010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf3),
    .Y(_5490_)
);

NAND2X1 _15011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .B(_5490_),
    .Y(_5491_)
);

NAND2X1 _15012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5492_)
);

OR2X2 _15013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .B(\datapath_1.PCJump [25]),
    .Y(_5493_)
);

NOR3X1 _15014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5492_),
    .C(_5493_),
    .Y(_5494_)
);

NAND3X1 _15015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf3),
    .B(_5468_),
    .C(_5465_),
    .Y(_5495_)
);

INVX8 _15016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495__bF$buf3),
    .Y(_5496_)
);

AOI22X1 _15017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_5497_)
);

INVX1 _15018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_5498_)
);

NAND3X1 _15019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf2),
    .B(_5477_),
    .C(_5461_),
    .Y(_5499_)
);

NOR3X1 _15020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(\datapath_1.PCJump [24]),
    .C(\datapath_1.PCJump [23]),
    .Y(_5500_)
);

NAND2X1 _15021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500__bF$buf3),
    .B(_5471__bF$buf3),
    .Y(_5501_)
);

OAI22X1 _15022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .B(_5501_),
    .C(_5499__bF$buf3),
    .D(_3957_),
    .Y(_5502_)
);

NAND2X1 _15023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .B(_5500__bF$buf2),
    .Y(_5503_)
);

NAND3X1 _15024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf1),
    .B(_5462_),
    .C(_5476_),
    .Y(_5504_)
);

OAI22X1 _15025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3907_),
    .B(_5503__bF$buf3),
    .C(_5504__bF$buf4),
    .D(_3981_),
    .Y(_5505_)
);

NOR2X1 _15026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .B(_5502_),
    .Y(_5506_)
);

NAND3X1 _15027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5491_),
    .B(_5497_),
    .C(_5506_),
    .Y(_5507_)
);

NOR2X1 _15028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5507_),
    .B(_5488_),
    .Y(_5508_)
);

NAND2X1 _15029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [25]),
    .B(_5464_),
    .Y(_5509_)
);

NAND2X1 _15030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(_5460_),
    .Y(_5510_)
);

AOI21X1 _15031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492_),
    .B(_5510_),
    .C(_5509_),
    .Y(_5511_)
);

NAND2X1 _15032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf0),
    .B(_5511_),
    .Y(_5512_)
);

NOR2X1 _15033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .Y(_5513_)
);

OAI21X1 _15034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5461_),
    .B(_5513_),
    .C(_5471__bF$buf2),
    .Y(_5514_)
);

OAI21X1 _15035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5514_),
    .C(_5512_),
    .Y(_5515_)
);

NOR2X1 _15036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(\datapath_1.PCJump [26]),
    .Y(_5516_)
);

OAI21X1 _15037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .B(_5493_),
    .C(_5516_),
    .Y(_5517_)
);

NAND3X1 _15038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf3),
    .B(_5477_),
    .C(_5468_),
    .Y(_5518_)
);

NAND3X1 _15039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5475_),
    .B(\datapath_1.PCJump [23]),
    .C(_5477_),
    .Y(_5519_)
);

OAI21X1 _15040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5519_),
    .B(\datapath_1.PCJump_27_bF$buf2 ),
    .C(_5518__bF$buf3),
    .Y(_5520_)
);

OR2X2 _15041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5520_),
    .B(_5517_),
    .Y(_5521_)
);

NOR3X1 _15042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf3),
    .B(_3928_),
    .C(_5521__bF$buf3),
    .Y(_5522_)
);

NAND3X1 _15043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf2),
    .B(_5471__bF$buf1),
    .C(_5476_),
    .Y(_5523_)
);

NAND3X1 _15044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf1),
    .B(_5461_),
    .C(_5471__bF$buf0),
    .Y(_5524_)
);

OAI22X1 _15045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5523_),
    .B(_3908_),
    .C(_3976_),
    .D(_5524__bF$buf3),
    .Y(_5525_)
);

NAND3X1 _15046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf0),
    .B(_5461_),
    .C(_5465_),
    .Y(_5526_)
);

NAND3X1 _15047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459__bF$buf3),
    .B(_5465_),
    .C(_5476_),
    .Y(_5527_)
);

OAI22X1 _15048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf4),
    .B(_3970_),
    .C(_3934_),
    .D(_5527__bF$buf4),
    .Y(_5528_)
);

NOR2X1 _15049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5525_),
    .B(_5528_),
    .Y(_5529_)
);

NAND3X1 _15050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5468_),
    .C(_5471__bF$buf5),
    .Y(_5530_)
);

NOR3X1 _15051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(\datapath_1.PCJump [23]),
    .C(_5459__bF$buf2),
    .Y(_5531_)
);

NAND2X1 _15052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5465_),
    .B(_5531__bF$buf4),
    .Y(_5532_)
);

OAI22X1 _15053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf3),
    .B(_3915_),
    .C(_5532__bF$buf3),
    .D(_3914_),
    .Y(_5533_)
);

NAND3X1 _15054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5477_),
    .C(_5461_),
    .Y(_5534_)
);

NAND3X1 _15055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5477_),
    .C(_5468_),
    .Y(_5535_)
);

OAI22X1 _15056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3896_),
    .B(_5535__bF$buf4),
    .C(_5534__bF$buf4),
    .D(_3980_),
    .Y(_5536_)
);

NOR2X1 _15057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5536_),
    .B(_5533_),
    .Y(_5537_)
);

NAND2X1 _15058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5537_),
    .B(_5529_),
    .Y(_5538_)
);

NAND3X1 _15059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(_5477_),
    .C(_5513_),
    .Y(_5539_)
);

NOR2X1 _15060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3933_),
    .B(_5539__bF$buf4),
    .Y(_5540_)
);

NAND3X1 _15061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .B(_5470_),
    .C(_5468_),
    .Y(_5541_)
);

NOR3X1 _15062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3964_),
    .B(_5459__bF$buf1),
    .C(_5541_),
    .Y(_5542_)
);

INVX1 _15063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [0]),
    .Y(_5543_)
);

NAND3X1 _15064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5513_),
    .C(_5462_),
    .Y(_5544_)
);

NAND3X1 _15065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5462_),
    .C(_5468_),
    .Y(_5545_)
);

OAI22X1 _15066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544__bF$buf3),
    .B(_5543_),
    .C(_5545__bF$buf3),
    .D(_3922_),
    .Y(_5546_)
);

NOR3X1 _15067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .B(_5540_),
    .C(_5542_),
    .Y(_5547_)
);

NAND2X1 _15068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500__bF$buf1),
    .B(_5465_),
    .Y(_5548_)
);

NAND3X1 _15069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf0 ),
    .B(_5477_),
    .C(_5476_),
    .Y(_5549_)
);

OAI22X1 _15070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3929_),
    .B(_5548__bF$buf4),
    .C(_5549__bF$buf4),
    .D(_3969_),
    .Y(_5550_)
);

NAND3X1 _15071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .B(_5471__bF$buf4),
    .C(_5531__bF$buf3),
    .Y(_5551_)
);

NAND3X1 _15072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf4 ),
    .B(_5471__bF$buf3),
    .C(_5476_),
    .Y(_5552_)
);

OAI21X1 _15073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552__bF$buf3),
    .B(_3952_),
    .C(_5551_),
    .Y(_5553_)
);

NOR2X1 _15074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5553_),
    .B(_5550_),
    .Y(_5554_)
);

NAND2X1 _15075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5547_),
    .B(_5554_),
    .Y(_5555_)
);

NOR3X1 _15076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5522_),
    .B(_5555_),
    .C(_5538_),
    .Y(_5556_)
);

AOI21X1 _15077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5508_),
    .B(_5556_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [0])
);

INVX1 _15078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf3),
    .Y(_5557_)
);

INVX1 _15079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf3),
    .Y(_5558_)
);

AOI22X1 _15080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5557_),
    .B(\datapath_1.regfile_1.regOut[17] [1]),
    .C(\datapath_1.regfile_1.regOut[18] [1]),
    .D(_5558_),
    .Y(_5559_)
);

INVX2 _15081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf3),
    .Y(_5560_)
);

NAND2X1 _15082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .B(_5560_),
    .Y(_5561_)
);

INVX2 _15083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .Y(_5562_)
);

NAND2X1 _15084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [1]),
    .B(_5562_),
    .Y(_5563_)
);

NAND3X1 _15085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5561_),
    .B(_5563_),
    .C(_5559_),
    .Y(_5564_)
);

INVX8 _15086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5523_),
    .Y(_5565_)
);

NAND2X1 _15087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .B(_5565__bF$buf3),
    .Y(_5566_)
);

INVX8 _15088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544__bF$buf2),
    .Y(_5567_)
);

NAND2X1 _15089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [1]),
    .B(_5567_),
    .Y(_5568_)
);

NAND3X1 _15090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf3 ),
    .B(_5468_),
    .C(_5465_),
    .Y(_5569_)
);

INVX8 _15091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .Y(_5570_)
);

INVX4 _15092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .Y(_5571_)
);

AOI22X1 _15093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [1]),
    .B(_5571_),
    .C(_5570__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[27] [1]),
    .Y(_5572_)
);

NAND3X1 _15094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5566_),
    .B(_5568_),
    .C(_5572_),
    .Y(_5573_)
);

OAI22X1 _15095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3991_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf2),
    .D(_4011_),
    .Y(_5574_)
);

AOI21X1 _15096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [1]),
    .B(_5494_),
    .C(_5574_),
    .Y(_5575_)
);

INVX8 _15097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf2),
    .Y(_5576_)
);

INVX4 _15098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503__bF$buf2),
    .Y(_5577_)
);

AOI22X1 _15099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [1]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_5578_)
);

INVX4 _15100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5548__bF$buf3),
    .Y(_5579_)
);

AOI22X1 _15101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .B(_5579_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_5580_)
);

NAND3X1 _15102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5575_),
    .B(_5580_),
    .C(_5578_),
    .Y(_5581_)
);

NOR3X1 _15103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .B(_5573_),
    .C(_5564_),
    .Y(_5582_)
);

NOR3X1 _15104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf2),
    .B(_4007_),
    .C(_5521__bF$buf2),
    .Y(_5583_)
);

INVX1 _15105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_5584_)
);

OAI22X1 _15106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf2),
    .B(_5584_),
    .C(_5532__bF$buf2),
    .D(_4019_),
    .Y(_5585_)
);

INVX1 _15107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_5586_)
);

OAI22X1 _15108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_5586_),
    .C(_5552__bF$buf2),
    .D(_4026_),
    .Y(_5587_)
);

NOR2X1 _15109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5587_),
    .B(_5585_),
    .Y(_5588_)
);

OAI22X1 _15110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_4010_),
    .C(_3992_),
    .D(_5527__bF$buf3),
    .Y(_5589_)
);

OAI22X1 _15111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf2),
    .B(_4035_),
    .C(_4031_),
    .D(_5504__bF$buf3),
    .Y(_5590_)
);

NOR2X1 _15112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5590_),
    .B(_5589_),
    .Y(_5591_)
);

NAND2X1 _15113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5588_),
    .B(_5591_),
    .Y(_5592_)
);

NAND3X1 _15114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf2),
    .Y(_5593_)
);

OAI21X1 _15115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf2),
    .B(_4002_),
    .C(_5593_),
    .Y(_5594_)
);

INVX1 _15116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [1]),
    .Y(_5595_)
);

INVX1 _15117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_5596_)
);

OAI22X1 _15118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_5595_),
    .C(_5596_),
    .D(_5499__bF$buf2),
    .Y(_5597_)
);

NOR2X1 _15119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5594_),
    .B(_5597_),
    .Y(_5598_)
);

NAND3X1 _15120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf2),
    .Y(_5599_)
);

OAI21X1 _15121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4027_),
    .B(_5535__bF$buf3),
    .C(_5599_),
    .Y(_5600_)
);

INVX1 _15122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [1]),
    .Y(_5601_)
);

OAI22X1 _15123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf3),
    .B(_5601_),
    .C(_5483__bF$buf3),
    .D(_4034_),
    .Y(_5602_)
);

NOR2X1 _15124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5600_),
    .B(_5602_),
    .Y(_5603_)
);

NAND2X1 _15125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5598_),
    .B(_5603_),
    .Y(_5604_)
);

NOR3X1 _15126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5604_),
    .B(_5583_),
    .C(_5592_),
    .Y(_5605_)
);

AOI21X1 _15127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5582_),
    .B(_5605_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [1])
);

INVX4 _15128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5469__bF$buf1),
    .Y(_5606_)
);

AOI22X1 _15129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .B(_5606_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_5607_)
);

AOI22X1 _15130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5481_),
    .B(\datapath_1.regfile_1.regOut[30] [2]),
    .C(\datapath_1.regfile_1.regOut[6] [2]),
    .D(_5565__bF$buf2),
    .Y(_5608_)
);

INVX1 _15131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_5609_)
);

OAI22X1 _15132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf1),
    .B(_5609_),
    .C(_5552__bF$buf1),
    .D(_4065_),
    .Y(_5610_)
);

INVX1 _15133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_5611_)
);

OAI22X1 _15134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4083_),
    .B(_5539__bF$buf2),
    .C(_5530__bF$buf1),
    .D(_5611_),
    .Y(_5612_)
);

NOR2X1 _15135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5612_),
    .B(_5610_),
    .Y(_5613_)
);

NAND3X1 _15136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5607_),
    .B(_5608_),
    .C(_5613_),
    .Y(_5614_)
);

NAND2X1 _15137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .B(_5494_),
    .Y(_5615_)
);

AOI22X1 _15138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_5616_)
);

OAI22X1 _15139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .B(_4047_),
    .C(_5483__bF$buf2),
    .D(_4082_),
    .Y(_5617_)
);

INVX1 _15140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_5618_)
);

OAI22X1 _15141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5618_),
    .B(_5548__bF$buf2),
    .C(_5504__bF$buf2),
    .D(_4055_),
    .Y(_5619_)
);

NOR2X1 _15142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5619_),
    .B(_5617_),
    .Y(_5620_)
);

NAND3X1 _15143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .B(_5616_),
    .C(_5620_),
    .Y(_5621_)
);

NOR2X1 _15144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5621_),
    .B(_5614_),
    .Y(_5622_)
);

NOR3X1 _15145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf1),
    .B(_4058_),
    .C(_5521__bF$buf1),
    .Y(_5623_)
);

NAND3X1 _15146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf0),
    .Y(_5624_)
);

OAI21X1 _15147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf1),
    .B(_4086_),
    .C(_5624_),
    .Y(_5625_)
);

INVX1 _15148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_5626_)
);

OAI22X1 _15149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4071_),
    .B(_5544__bF$buf1),
    .C(_5499__bF$buf1),
    .D(_5626_),
    .Y(_5627_)
);

NOR2X1 _15150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5625_),
    .B(_5627_),
    .Y(_5628_)
);

NAND3X1 _15151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf1),
    .Y(_5629_)
);

OAI21X1 _15152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4074_),
    .B(_5535__bF$buf2),
    .C(_5629_),
    .Y(_5630_)
);

INVX1 _15153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [2]),
    .Y(_5631_)
);

OAI22X1 _15154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5631_),
    .B(_5545__bF$buf1),
    .C(_5466__bF$buf2),
    .D(_4063_),
    .Y(_5632_)
);

NOR2X1 _15155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5630_),
    .B(_5632_),
    .Y(_5633_)
);

NAND2X1 _15156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5628_),
    .B(_5633_),
    .Y(_5634_)
);

OAI22X1 _15157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_4059_),
    .C(_4056_),
    .D(_5526__bF$buf2),
    .Y(_5635_)
);

INVX1 _15158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_5636_)
);

OAI22X1 _15159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527__bF$buf2),
    .B(_4045_),
    .C(_5636_),
    .D(_5532__bF$buf1),
    .Y(_5637_)
);

NOR2X1 _15160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5637_),
    .B(_5635_),
    .Y(_5638_)
);

INVX1 _15161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_5639_)
);

OAI22X1 _15162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495__bF$buf2),
    .B(_5639_),
    .C(_4085_),
    .D(_5534__bF$buf2),
    .Y(_5640_)
);

OAI22X1 _15163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf2),
    .B(_4062_),
    .C(_4072_),
    .D(_5549__bF$buf2),
    .Y(_5641_)
);

NOR2X1 _15164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5640_),
    .B(_5641_),
    .Y(_5642_)
);

NAND2X1 _15165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5642_),
    .B(_5638_),
    .Y(_5643_)
);

NOR3X1 _15166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5634_),
    .B(_5623_),
    .C(_5643_),
    .Y(_5644_)
);

AOI21X1 _15167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5622_),
    .B(_5644_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [2])
);

INVX1 _15168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_5645_)
);

OAI22X1 _15169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf1),
    .B(_4132_),
    .C(_5645_),
    .D(_5549__bF$buf1),
    .Y(_5646_)
);

OAI22X1 _15170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_4105_),
    .C(_4141_),
    .D(_5526__bF$buf1),
    .Y(_5647_)
);

NOR2X1 _15171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5646_),
    .B(_5647_),
    .Y(_5648_)
);

INVX8 _15172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf0),
    .Y(_5649_)
);

INVX8 _15173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552__bF$buf0),
    .Y(_5650_)
);

AOI22X1 _15174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5649_),
    .B(\datapath_1.regfile_1.regOut[23] [3]),
    .C(\datapath_1.regfile_1.regOut[22] [3]),
    .D(_5650_),
    .Y(_5651_)
);

AOI22X1 _15175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [3]),
    .B(_5567_),
    .C(_5565__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_5652_)
);

NAND3X1 _15176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5651_),
    .B(_5652_),
    .C(_5648_),
    .Y(_5653_)
);

NAND2X1 _15177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .B(_5494_),
    .Y(_5654_)
);

AOI22X1 _15178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .B(_5606_),
    .C(_5570__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[27] [3]),
    .Y(_5655_)
);

INVX1 _15179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_5656_)
);

OAI22X1 _15180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4122_),
    .B(_5503__bF$buf1),
    .C(_5463__bF$buf1),
    .D(_5656_),
    .Y(_5657_)
);

INVX1 _15181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_5658_)
);

OAI22X1 _15182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4124_),
    .B(_5548__bF$buf1),
    .C(_5495__bF$buf1),
    .D(_5658_),
    .Y(_5659_)
);

NOR2X1 _15183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5659_),
    .B(_5657_),
    .Y(_5660_)
);

NAND3X1 _15184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5654_),
    .B(_5655_),
    .C(_5660_),
    .Y(_5661_)
);

NOR2X1 _15185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5661_),
    .B(_5653_),
    .Y(_5662_)
);

INVX1 _15186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_5663_)
);

NOR3X1 _15187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf0),
    .B(_5663_),
    .C(_5521__bF$buf0),
    .Y(_5664_)
);

OAI22X1 _15188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4137_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf1),
    .D(_4138_),
    .Y(_5665_)
);

INVX1 _15189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [3]),
    .Y(_5666_)
);

INVX1 _15190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_5667_)
);

OAI22X1 _15191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf0),
    .B(_5667_),
    .C(_5666_),
    .D(_5480__bF$buf1),
    .Y(_5668_)
);

NOR2X1 _15192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5665_),
    .B(_5668_),
    .Y(_5669_)
);

OAI22X1 _15193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4106_),
    .B(_5539__bF$buf1),
    .C(_5527__bF$buf1),
    .D(_4112_),
    .Y(_5670_)
);

OAI22X1 _15194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf1),
    .B(_4095_),
    .C(_4121_),
    .D(_5504__bF$buf1),
    .Y(_5671_)
);

NOR2X1 _15195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5671_),
    .B(_5670_),
    .Y(_5672_)
);

NAND2X1 _15196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5669_),
    .B(_5672_),
    .Y(_5673_)
);

OAI22X1 _15197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4125_),
    .B(_5501_),
    .C(_5524__bF$buf0),
    .D(_4109_),
    .Y(_5674_)
);

INVX1 _15198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_5675_)
);

INVX1 _15199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_5676_)
);

OAI22X1 _15200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499__bF$buf0),
    .B(_5676_),
    .C(_5532__bF$buf0),
    .D(_5675_),
    .Y(_5677_)
);

NOR2X1 _15201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5674_),
    .B(_5677_),
    .Y(_5678_)
);

NAND3X1 _15202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .B(_5471__bF$buf4),
    .C(_5531__bF$buf0),
    .Y(_5679_)
);

OAI21X1 _15203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4108_),
    .B(_5535__bF$buf1),
    .C(_5679_),
    .Y(_5680_)
);

OAI22X1 _15204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_4116_),
    .C(_4097_),
    .D(_5483__bF$buf1),
    .Y(_5681_)
);

NOR2X1 _15205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5680_),
    .B(_5681_),
    .Y(_5682_)
);

NAND2X1 _15206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5678_),
    .B(_5682_),
    .Y(_5683_)
);

NOR3X1 _15207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5673_),
    .B(_5664_),
    .C(_5683_),
    .Y(_5684_)
);

AOI21X1 _15208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5662_),
    .B(_5684_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [3])
);

INVX4 _15209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .Y(_5685_)
);

AOI22X1 _15210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [4]),
    .C(\datapath_1.regfile_1.regOut[22] [4]),
    .D(_5650_),
    .Y(_5686_)
);

NOR2X1 _15211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4164_),
    .B(_5534__bF$buf0),
    .Y(_5687_)
);

NAND2X1 _15212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf2 ),
    .B(_5513_),
    .Y(_5688_)
);

NOR3X1 _15213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4160_),
    .B(_5509_),
    .C(_5688_),
    .Y(_5689_)
);

NOR2X1 _15214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4161_),
    .B(_5549__bF$buf0),
    .Y(_5690_)
);

NOR3X1 _15215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5687_),
    .B(_5689_),
    .C(_5690_),
    .Y(_5691_)
);

INVX4 _15216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5532__bF$buf3),
    .Y(_5692_)
);

INVX4 _15217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5535__bF$buf0),
    .Y(_5693_)
);

AOI22X1 _15218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .B(_5693_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_5694_)
);

NAND3X1 _15219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5686_),
    .B(_5694_),
    .C(_5691_),
    .Y(_5695_)
);

NAND2X1 _15220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [23]),
    .B(_5475_),
    .Y(_5696_)
);

NOR3X1 _15221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump_27_bF$buf1 ),
    .B(_5493_),
    .C(_5696_),
    .Y(_5697_)
);

INVX4 _15222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5501_),
    .Y(_5698_)
);

AOI22X1 _15223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_5699_)
);

INVX8 _15224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf3),
    .Y(_5700_)
);

AOI22X1 _15225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [4]),
    .C(\datapath_1.regfile_1.regOut[5] [4]),
    .D(_5700_),
    .Y(_5701_)
);

OAI22X1 _15226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf0),
    .B(_4158_),
    .C(_4150_),
    .D(_5527__bF$buf0),
    .Y(_5702_)
);

OAI22X1 _15227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4167_),
    .B(_5539__bF$buf0),
    .C(_5469__bF$buf0),
    .D(_4165_),
    .Y(_5703_)
);

NOR2X1 _15228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5703_),
    .B(_5702_),
    .Y(_5704_)
);

NAND3X1 _15229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5699_),
    .B(_5701_),
    .C(_5704_),
    .Y(_5705_)
);

NOR2X1 _15230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5705_),
    .B(_5695_),
    .Y(_5706_)
);

NAND2X1 _15231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .B(_5649_),
    .Y(_5707_)
);

INVX1 _15232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_5708_)
);

OAI22X1 _15233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_5708_),
    .C(_4178_),
    .D(_5483__bF$buf0),
    .Y(_5709_)
);

AOI21X1 _15234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [4]),
    .B(_5567_),
    .C(_5709_),
    .Y(_5710_)
);

INVX1 _15235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [4]),
    .Y(_5711_)
);

OAI22X1 _15236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_5711_),
    .C(_4187_),
    .D(_5569_),
    .Y(_5712_)
);

INVX1 _15237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [4]),
    .Y(_5713_)
);

INVX1 _15238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [4]),
    .Y(_5714_)
);

OAI22X1 _15239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5713_),
    .B(_5545__bF$buf3),
    .C(_5485__bF$buf0),
    .D(_5714_),
    .Y(_5715_)
);

NOR2X1 _15240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .B(_5712_),
    .Y(_5716_)
);

NAND3X1 _15241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5707_),
    .B(_5716_),
    .C(_5710_),
    .Y(_5717_)
);

NAND2X1 _15242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5475_),
    .B(_5460_),
    .Y(_5718_)
);

AOI21X1 _15243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5696_),
    .B(_5718_),
    .C(_5509_),
    .Y(_5719_)
);

OAI21X1 _15244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5719_),
    .B(_5511_),
    .C(_5459__bF$buf0),
    .Y(_5720_)
);

NOR3X1 _15245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .B(_5517_),
    .C(_5697_),
    .Y(_5721_)
);

NAND3X1 _15246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5722_)
);

OAI22X1 _15247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4176_),
    .B(_5518__bF$buf2),
    .C(_5478__bF$buf3),
    .D(_4175_),
    .Y(_5723_)
);

INVX1 _15248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_5724_)
);

OAI22X1 _15249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4183_),
    .B(_5548__bF$buf0),
    .C(_5489__bF$buf0),
    .D(_5724_),
    .Y(_5725_)
);

NOR2X1 _15250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5725_),
    .B(_5723_),
    .Y(_5726_)
);

INVX1 _15251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_5727_)
);

INVX1 _15252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_5728_)
);

OAI22X1 _15253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5727_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf0),
    .D(_5728_),
    .Y(_5729_)
);

INVX1 _15254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_5730_)
);

OAI22X1 _15255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf0),
    .B(_4168_),
    .C(_5730_),
    .D(_5504__bF$buf0),
    .Y(_5731_)
);

NOR2X1 _15256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5729_),
    .B(_5731_),
    .Y(_5732_)
);

NAND3X1 _15257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5726_),
    .B(_5732_),
    .C(_5722_),
    .Y(_5733_)
);

NOR2X1 _15258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5717_),
    .B(_5733_),
    .Y(_5734_)
);

AOI21X1 _15259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5734_),
    .B(_5706_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [4])
);

AOI22X1 _15260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_5735_)
);

AOI22X1 _15261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [5]),
    .B(_5567_),
    .C(_5565__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_5736_)
);

OAI22X1 _15262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_4217_),
    .C(_5552__bF$buf3),
    .D(_4210_),
    .Y(_5737_)
);

OAI22X1 _15263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4239_),
    .B(_5539__bF$buf4),
    .C(_5530__bF$buf3),
    .D(_4198_),
    .Y(_5738_)
);

NOR2X1 _15264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5738_),
    .B(_5737_),
    .Y(_5739_)
);

NAND3X1 _15265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5735_),
    .B(_5736_),
    .C(_5739_),
    .Y(_5740_)
);

NAND2X1 _15266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [5]),
    .B(_5490_),
    .Y(_5741_)
);

AOI22X1 _15267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_5742_)
);

INVX1 _15268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [5]),
    .Y(_5743_)
);

OAI22X1 _15269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5743_),
    .B(_5545__bF$buf2),
    .C(_5569_),
    .D(_4207_),
    .Y(_5744_)
);

INVX1 _15270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_5745_)
);

OAI22X1 _15271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4227_),
    .B(_5503__bF$buf3),
    .C(_5504__bF$buf4),
    .D(_5745_),
    .Y(_5746_)
);

NOR2X1 _15272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5744_),
    .B(_5746_),
    .Y(_5747_)
);

NAND3X1 _15273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5741_),
    .B(_5742_),
    .C(_5747_),
    .Y(_5748_)
);

NOR2X1 _15274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5748_),
    .B(_5740_),
    .Y(_5749_)
);

INVX1 _15275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_5750_)
);

NOR3X1 _15276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf3),
    .B(_5750_),
    .C(_5521__bF$buf3),
    .Y(_5751_)
);

NAND3X1 _15277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .B(_5500__bF$buf2),
    .C(_5471__bF$buf3),
    .Y(_5752_)
);

OAI21X1 _15278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf2),
    .B(_4236_),
    .C(_5752_),
    .Y(_5753_)
);

OAI22X1 _15279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_4209_),
    .C(_4199_),
    .D(_5499__bF$buf3),
    .Y(_5754_)
);

NOR2X1 _15280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5753_),
    .B(_5754_),
    .Y(_5755_)
);

NAND3X1 _15281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [5]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf4),
    .Y(_5756_)
);

OAI21X1 _15282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4235_),
    .B(_5535__bF$buf4),
    .C(_5756_),
    .Y(_5757_)
);

OAI22X1 _15283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf4),
    .B(_4230_),
    .C(_5483__bF$buf4),
    .D(_4206_),
    .Y(_5758_)
);

NOR2X1 _15284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5757_),
    .B(_5758_),
    .Y(_5759_)
);

NAND2X1 _15285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5755_),
    .B(_5759_),
    .Y(_5760_)
);

OAI22X1 _15286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_4213_),
    .C(_4222_),
    .D(_5526__bF$buf4),
    .Y(_5761_)
);

INVX1 _15287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_5762_)
);

OAI22X1 _15288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527__bF$buf4),
    .B(_4195_),
    .C(_5762_),
    .D(_5532__bF$buf2),
    .Y(_5763_)
);

NOR2X1 _15289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5763_),
    .B(_5761_),
    .Y(_5764_)
);

INVX1 _15290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_5765_)
);

OAI22X1 _15291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5765_),
    .B(_5548__bF$buf4),
    .C(_5534__bF$buf4),
    .D(_4216_),
    .Y(_5766_)
);

OAI22X1 _15292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf4),
    .B(_4238_),
    .C(_5466__bF$buf4),
    .D(_4202_),
    .Y(_5767_)
);

NOR2X1 _15293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5766_),
    .B(_5767_),
    .Y(_5768_)
);

NAND2X1 _15294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5768_),
    .B(_5764_),
    .Y(_5769_)
);

NOR3X1 _15295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .B(_5751_),
    .C(_5769_),
    .Y(_5770_)
);

AOI21X1 _15296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5749_),
    .B(_5770_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [5])
);

NAND2X1 _15297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [6]),
    .B(_5481_),
    .Y(_5771_)
);

AOI22X1 _15298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [6]),
    .B(_5571_),
    .C(_5486_),
    .D(\datapath_1.regfile_1.regOut[29] [6]),
    .Y(_5772_)
);

OAI22X1 _15299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_4252_),
    .C(_4249_),
    .D(_5483__bF$buf3),
    .Y(_5773_)
);

INVX1 _15300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [6]),
    .Y(_5774_)
);

OAI22X1 _15301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5774_),
    .B(_5544__bF$buf0),
    .C(_5569_),
    .D(_4289_),
    .Y(_5775_)
);

NOR2X1 _15302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5775_),
    .B(_5773_),
    .Y(_5776_)
);

NAND3X1 _15303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5771_),
    .B(_5772_),
    .C(_5776_),
    .Y(_5777_)
);

AOI22X1 _15304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_5778_)
);

AOI22X1 _15305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [6]),
    .C(\datapath_1.regfile_1.regOut[5] [6]),
    .D(_5700_),
    .Y(_5779_)
);

OAI22X1 _15306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf3),
    .B(_4280_),
    .C(_4283_),
    .D(_5527__bF$buf3),
    .Y(_5780_)
);

OAI22X1 _15307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4279_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf3),
    .D(_4253_),
    .Y(_5781_)
);

NOR2X1 _15308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5781_),
    .B(_5780_),
    .Y(_5782_)
);

NAND3X1 _15309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5778_),
    .B(_5779_),
    .C(_5782_),
    .Y(_5783_)
);

NOR2X1 _15310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5783_),
    .B(_5777_),
    .Y(_5784_)
);

NOR2X1 _15311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .B(_5688_),
    .Y(_5785_)
);

NAND2X1 _15312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .B(_5785_),
    .Y(_5786_)
);

NOR3X1 _15313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4259_),
    .B(_5459__bF$buf3),
    .C(_5519_),
    .Y(_5787_)
);

INVX1 _15314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_5788_)
);

NOR2X1 _15315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5788_),
    .B(_5549__bF$buf3),
    .Y(_5789_)
);

INVX1 _15316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_5790_)
);

NOR2X1 _15317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5790_),
    .B(_5535__bF$buf3),
    .Y(_5791_)
);

NOR3X1 _15318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5787_),
    .B(_5791_),
    .C(_5789_),
    .Y(_5792_)
);

INVX1 _15319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_5793_)
);

INVX1 _15320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_5794_)
);

OAI22X1 _15321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf2),
    .B(_5794_),
    .C(_5532__bF$buf1),
    .D(_5793_),
    .Y(_5795_)
);

OAI22X1 _15322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_4287_),
    .C(_4286_),
    .D(_5552__bF$buf2),
    .Y(_5796_)
);

NOR2X1 _15323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5795_),
    .B(_5796_),
    .Y(_5797_)
);

NAND3X1 _15324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5786_),
    .B(_5792_),
    .C(_5797_),
    .Y(_5798_)
);

NAND3X1 _15325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5799_)
);

OAI22X1 _15326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4273_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf1),
    .D(_4250_),
    .Y(_5800_)
);

INVX1 _15327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_5801_)
);

OAI22X1 _15328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4270_),
    .B(_5548__bF$buf3),
    .C(_5489__bF$buf3),
    .D(_5801_),
    .Y(_5802_)
);

NOR2X1 _15329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5802_),
    .B(_5800_),
    .Y(_5803_)
);

INVX1 _15330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_5804_)
);

OAI22X1 _15331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5804_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf3),
    .D(_4260_),
    .Y(_5805_)
);

INVX1 _15332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_5806_)
);

INVX1 _15333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_5807_)
);

OAI22X1 _15334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf3),
    .B(_5807_),
    .C(_5806_),
    .D(_5504__bF$buf3),
    .Y(_5808_)
);

NOR2X1 _15335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5805_),
    .B(_5808_),
    .Y(_5809_)
);

NAND3X1 _15336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5803_),
    .B(_5809_),
    .C(_5799_),
    .Y(_5810_)
);

NOR2X1 _15337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5798_),
    .B(_5810_),
    .Y(_5811_)
);

AOI21X1 _15338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5784_),
    .B(_5811_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [6])
);

NAND2X1 _15339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [7]),
    .B(_5785_),
    .Y(_5812_)
);

NOR2X1 _15340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4299_),
    .B(_5549__bF$buf2),
    .Y(_5813_)
);

NOR2X1 _15341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4339_),
    .B(_5534__bF$buf3),
    .Y(_5814_)
);

NOR2X1 _15342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4306_),
    .B(_5535__bF$buf2),
    .Y(_5815_)
);

NOR3X1 _15343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5813_),
    .B(_5815_),
    .C(_5814_),
    .Y(_5816_)
);

INVX1 _15344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_5817_)
);

OAI22X1 _15345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf1),
    .B(_5817_),
    .C(_5532__bF$buf0),
    .D(_4298_),
    .Y(_5818_)
);

OAI22X1 _15346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_4328_),
    .C(_4327_),
    .D(_5552__bF$buf1),
    .Y(_5819_)
);

NOR2X1 _15347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5818_),
    .B(_5819_),
    .Y(_5820_)
);

NAND3X1 _15348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5812_),
    .B(_5820_),
    .C(_5816_),
    .Y(_5821_)
);

AOI22X1 _15349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_5822_)
);

AOI22X1 _15350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [7]),
    .C(\datapath_1.regfile_1.regOut[5] [7]),
    .D(_5700_),
    .Y(_5823_)
);

OAI22X1 _15351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf2),
    .B(_4333_),
    .C(_4317_),
    .D(_5527__bF$buf2),
    .Y(_5824_)
);

OAI22X1 _15352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_5539__bF$buf2),
    .C(_5469__bF$buf2),
    .D(_4307_),
    .Y(_5825_)
);

NOR2X1 _15353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5825_),
    .B(_5824_),
    .Y(_5826_)
);

NAND3X1 _15354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5822_),
    .B(_5823_),
    .C(_5826_),
    .Y(_5827_)
);

NOR2X1 _15355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5827_),
    .B(_5821_),
    .Y(_5828_)
);

AOI22X1 _15356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [7]),
    .B(_5567_),
    .C(_5486_),
    .D(\datapath_1.regfile_1.regOut[29] [7]),
    .Y(_5829_)
);

AOI22X1 _15357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [7]),
    .B(_5571_),
    .C(_5481_),
    .D(\datapath_1.regfile_1.regOut[30] [7]),
    .Y(_5830_)
);

INVX1 _15358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_5831_)
);

OAI22X1 _15359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf2),
    .B(_5831_),
    .C(_4313_),
    .D(_5483__bF$buf2),
    .Y(_5832_)
);

AOI21X1 _15360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [7]),
    .B(_5570__bF$buf1),
    .C(_5832_),
    .Y(_5833_)
);

NAND3X1 _15361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5829_),
    .B(_5830_),
    .C(_5833_),
    .Y(_5834_)
);

NAND3X1 _15362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5835_)
);

OAI22X1 _15363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .B(_5518__bF$buf0),
    .C(_5478__bF$buf0),
    .D(_4324_),
    .Y(_5836_)
);

INVX1 _15364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_5837_)
);

INVX1 _15365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_5838_)
);

OAI22X1 _15366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5837_),
    .B(_5548__bF$buf2),
    .C(_5489__bF$buf2),
    .D(_5838_),
    .Y(_5839_)
);

NOR2X1 _15367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5839_),
    .B(_5836_),
    .Y(_5840_)
);

OAI22X1 _15368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4304_),
    .B(_5503__bF$buf1),
    .C(_5495__bF$buf2),
    .D(_4302_),
    .Y(_5841_)
);

OAI22X1 _15369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf2),
    .B(_4336_),
    .C(_4340_),
    .D(_5504__bF$buf2),
    .Y(_5842_)
);

NOR2X1 _15370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5841_),
    .B(_5842_),
    .Y(_5843_)
);

NAND3X1 _15371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5840_),
    .B(_5843_),
    .C(_5835_),
    .Y(_5844_)
);

NOR2X1 _15372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5834_),
    .B(_5844_),
    .Y(_5845_)
);

AOI21X1 _15373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5845_),
    .B(_5828_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [7])
);

AOI22X1 _15374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [8]),
    .C(\datapath_1.regfile_1.regOut[22] [8]),
    .D(_5650_),
    .Y(_5846_)
);

NOR2X1 _15375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_5549__bF$buf1),
    .Y(_5847_)
);

NOR2X1 _15376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4370_),
    .B(_5534__bF$buf2),
    .Y(_5848_)
);

INVX1 _15377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_5849_)
);

NOR2X1 _15378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5849_),
    .B(_5535__bF$buf1),
    .Y(_5850_)
);

NOR3X1 _15379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5847_),
    .B(_5850_),
    .C(_5848_),
    .Y(_5851_)
);

AOI22X1 _15380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .B(_5785_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_5852_)
);

NAND3X1 _15381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5846_),
    .B(_5852_),
    .C(_5851_),
    .Y(_5853_)
);

AOI22X1 _15382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [8]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_5854_)
);

AOI22X1 _15383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [8]),
    .C(\datapath_1.regfile_1.regOut[5] [8]),
    .D(_5700_),
    .Y(_5855_)
);

OAI22X1 _15384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf1),
    .B(_4385_),
    .C(_4360_),
    .D(_5527__bF$buf1),
    .Y(_5856_)
);

INVX1 _15385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_5857_)
);

OAI22X1 _15386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4363_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf1),
    .D(_5857_),
    .Y(_5858_)
);

NOR2X1 _15387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5858_),
    .B(_5856_),
    .Y(_5859_)
);

NAND3X1 _15388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5854_),
    .B(_5855_),
    .C(_5859_),
    .Y(_5860_)
);

NOR2X1 _15389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5860_),
    .B(_5853_),
    .Y(_5861_)
);

NAND2X1 _15390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .B(_5649_),
    .Y(_5862_)
);

INVX1 _15391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [8]),
    .Y(_5863_)
);

OAI22X1 _15392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5863_),
    .B(_5545__bF$buf1),
    .C(_5485__bF$buf3),
    .D(_4381_),
    .Y(_5864_)
);

INVX1 _15393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [8]),
    .Y(_5865_)
);

OAI22X1 _15394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5865_),
    .B(_5544__bF$buf3),
    .C(_5480__bF$buf2),
    .D(_4373_),
    .Y(_5866_)
);

NOR2X1 _15395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5864_),
    .B(_5866_),
    .Y(_5867_)
);

OAI22X1 _15396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_4359_),
    .C(_4348_),
    .D(_5483__bF$buf1),
    .Y(_5868_)
);

AOI21X1 _15397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [8]),
    .B(_5570__bF$buf0),
    .C(_5868_),
    .Y(_5869_)
);

NAND3X1 _15398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5862_),
    .B(_5867_),
    .C(_5869_),
    .Y(_5870_)
);

NAND3X1 _15399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5871_)
);

INVX1 _15400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_5872_)
);

OAI22X1 _15401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4346_),
    .B(_5518__bF$buf3),
    .C(_5478__bF$buf3),
    .D(_5872_),
    .Y(_5873_)
);

INVX1 _15402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_5874_)
);

INVX1 _15403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_5875_)
);

OAI22X1 _15404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5874_),
    .B(_5548__bF$buf1),
    .C(_5489__bF$buf1),
    .D(_5875_),
    .Y(_5876_)
);

NOR2X1 _15405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5876_),
    .B(_5873_),
    .Y(_5877_)
);

INVX1 _15406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_5878_)
);

OAI22X1 _15407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5878_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf1),
    .D(_4371_),
    .Y(_5879_)
);

INVX1 _15408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_5880_)
);

INVX1 _15409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_5881_)
);

OAI22X1 _15410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf1),
    .B(_5881_),
    .C(_5880_),
    .D(_5504__bF$buf1),
    .Y(_5882_)
);

NOR2X1 _15411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5879_),
    .B(_5882_),
    .Y(_5883_)
);

NAND3X1 _15412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5877_),
    .B(_5883_),
    .C(_5871_),
    .Y(_5884_)
);

NOR2X1 _15413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5870_),
    .B(_5884_),
    .Y(_5885_)
);

AOI21X1 _15414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5885_),
    .B(_5861_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [8])
);

NAND2X1 _15415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .B(_5693_),
    .Y(_5886_)
);

NOR2X1 _15416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4392_),
    .B(_5534__bF$buf1),
    .Y(_5887_)
);

INVX1 _15417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_5888_)
);

NOR3X1 _15418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_5509_),
    .C(_5688_),
    .Y(_5889_)
);

INVX1 _15419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_5890_)
);

NOR2X1 _15420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5890_),
    .B(_5549__bF$buf0),
    .Y(_5891_)
);

NOR3X1 _15421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5887_),
    .B(_5889_),
    .C(_5891_),
    .Y(_5892_)
);

INVX1 _15422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_5893_)
);

OAI22X1 _15423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf0),
    .B(_5893_),
    .C(_5532__bF$buf3),
    .D(_4391_),
    .Y(_5894_)
);

OAI22X1 _15424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_4415_),
    .C(_4414_),
    .D(_5552__bF$buf0),
    .Y(_5895_)
);

NOR2X1 _15425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .B(_5895_),
    .Y(_5896_)
);

NAND3X1 _15426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5886_),
    .B(_5896_),
    .C(_5892_),
    .Y(_5897_)
);

AOI22X1 _15427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [9]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_5898_)
);

AOI22X1 _15428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [9]),
    .C(\datapath_1.regfile_1.regOut[5] [9]),
    .D(_5700_),
    .Y(_5899_)
);

OAI22X1 _15429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf0),
    .B(_4426_),
    .C(_4407_),
    .D(_5527__bF$buf0),
    .Y(_5900_)
);

INVX1 _15430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_5901_)
);

OAI22X1 _15431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4406_),
    .B(_5539__bF$buf0),
    .C(_5469__bF$buf0),
    .D(_5901_),
    .Y(_5902_)
);

NOR2X1 _15432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5902_),
    .B(_5900_),
    .Y(_5903_)
);

NAND3X1 _15433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5898_),
    .B(_5899_),
    .C(_5903_),
    .Y(_5904_)
);

NOR2X1 _15434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5904_),
    .B(_5897_),
    .Y(_5905_)
);

NAND2X1 _15435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [9]),
    .B(_5570__bF$buf3),
    .Y(_5906_)
);

OAI22X1 _15436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_4403_),
    .C(_4395_),
    .D(_5483__bF$buf0),
    .Y(_5907_)
);

AOI21X1 _15437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [9]),
    .B(_5567_),
    .C(_5907_),
    .Y(_5908_)
);

OAI22X1 _15438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4425_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf2),
    .D(_4422_),
    .Y(_5909_)
);

AOI21X1 _15439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [9]),
    .B(_5481_),
    .C(_5909_),
    .Y(_5910_)
);

NAND3X1 _15440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5906_),
    .B(_5910_),
    .C(_5908_),
    .Y(_5911_)
);

NAND3X1 _15441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5912_)
);

INVX1 _15442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_5913_)
);

INVX1 _15443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_5914_)
);

OAI22X1 _15444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5914_),
    .B(_5518__bF$buf2),
    .C(_5478__bF$buf2),
    .D(_5913_),
    .Y(_5915_)
);

OAI22X1 _15445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4404_),
    .B(_5548__bF$buf0),
    .C(_5489__bF$buf0),
    .D(_4417_),
    .Y(_5916_)
);

NOR2X1 _15446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5916_),
    .B(_5915_),
    .Y(_5917_)
);

INVX1 _15447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_5918_)
);

INVX1 _15448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_5919_)
);

OAI22X1 _15449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5918_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf0),
    .D(_5919_),
    .Y(_5920_)
);

INVX1 _15450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_5921_)
);

INVX1 _15451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_5922_)
);

OAI22X1 _15452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf0),
    .B(_5922_),
    .C(_5921_),
    .D(_5504__bF$buf0),
    .Y(_5923_)
);

NOR2X1 _15453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5920_),
    .B(_5923_),
    .Y(_5924_)
);

NAND3X1 _15454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5917_),
    .B(_5924_),
    .C(_5912_),
    .Y(_5925_)
);

NOR2X1 _15455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5911_),
    .B(_5925_),
    .Y(_5926_)
);

AOI21X1 _15456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .B(_5905_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [9])
);

NAND2X1 _15457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .B(_5693_),
    .Y(_5927_)
);

NOR2X1 _15458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4467_),
    .B(_5534__bF$buf0),
    .Y(_5928_)
);

INVX1 _15459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_5929_)
);

NOR3X1 _15460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5929_),
    .B(_5509_),
    .C(_5688_),
    .Y(_5930_)
);

NOR2X1 _15461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4449_),
    .B(_5549__bF$buf4),
    .Y(_5931_)
);

NOR3X1 _15462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5928_),
    .B(_5930_),
    .C(_5931_),
    .Y(_5932_)
);

OAI22X1 _15463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf3),
    .B(_4466_),
    .C(_5532__bF$buf2),
    .D(_4448_),
    .Y(_5933_)
);

OAI22X1 _15464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_4437_),
    .C(_4470_),
    .D(_5552__bF$buf3),
    .Y(_5934_)
);

NOR2X1 _15465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5933_),
    .B(_5934_),
    .Y(_5935_)
);

NAND3X1 _15466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .B(_5935_),
    .C(_5932_),
    .Y(_5936_)
);

AOI22X1 _15467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [10]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_5937_)
);

AOI22X1 _15468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [10]),
    .C(\datapath_1.regfile_1.regOut[5] [10]),
    .D(_5700_),
    .Y(_5938_)
);

OAI22X1 _15469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf4),
    .B(_4457_),
    .C(_4460_),
    .D(_5527__bF$buf4),
    .Y(_5939_)
);

OAI22X1 _15470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4459_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf3),
    .D(_4456_),
    .Y(_5940_)
);

NOR2X1 _15471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5940_),
    .B(_5939_),
    .Y(_5941_)
);

NAND3X1 _15472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5937_),
    .B(_5938_),
    .C(_5941_),
    .Y(_5942_)
);

NOR2X1 _15473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5942_),
    .B(_5936_),
    .Y(_5943_)
);

NAND2X1 _15474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [10]),
    .B(_5570__bF$buf2),
    .Y(_5944_)
);

INVX1 _15475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [10]),
    .Y(_5945_)
);

OAI22X1 _15476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_5945_),
    .C(_4434_),
    .D(_5483__bF$buf4),
    .Y(_5946_)
);

AOI21X1 _15477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [10]),
    .B(_5567_),
    .C(_5946_),
    .Y(_5947_)
);

INVX1 _15478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [10]),
    .Y(_5948_)
);

OAI22X1 _15479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5948_),
    .B(_5545__bF$buf3),
    .C(_5485__bF$buf1),
    .D(_4445_),
    .Y(_5949_)
);

AOI21X1 _15480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [10]),
    .B(_5481_),
    .C(_5949_),
    .Y(_5950_)
);

NAND3X1 _15481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5944_),
    .B(_5950_),
    .C(_5947_),
    .Y(_5951_)
);

NAND3X1 _15482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .B(_5720_),
    .C(_5721_),
    .Y(_5952_)
);

INVX1 _15483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_5953_)
);

INVX1 _15484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_5954_)
);

OAI22X1 _15485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5954_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf1),
    .D(_5953_),
    .Y(_5955_)
);

OAI22X1 _15486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4440_),
    .B(_5548__bF$buf4),
    .C(_5489__bF$buf3),
    .D(_4438_),
    .Y(_5956_)
);

NOR2X1 _15487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5956_),
    .B(_5955_),
    .Y(_5957_)
);

INVX1 _15488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_5958_)
);

INVX1 _15489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_5959_)
);

OAI22X1 _15490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5958_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf3),
    .D(_5959_),
    .Y(_5960_)
);

INVX1 _15491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_5961_)
);

INVX1 _15492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_5962_)
);

OAI22X1 _15493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf3),
    .B(_5962_),
    .C(_5961_),
    .D(_5504__bF$buf4),
    .Y(_5963_)
);

NOR2X1 _15494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5960_),
    .B(_5963_),
    .Y(_5964_)
);

NAND3X1 _15495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5957_),
    .B(_5964_),
    .C(_5952_),
    .Y(_5965_)
);

NOR2X1 _15496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5951_),
    .B(_5965_),
    .Y(_5966_)
);

AOI21X1 _15497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5966_),
    .B(_5943_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [10])
);

OAI22X1 _15498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf2),
    .B(_4507_),
    .C(_5527__bF$buf3),
    .D(_4478_),
    .Y(_5967_)
);

OAI22X1 _15499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4492_),
    .B(_5539__bF$buf3),
    .C(_5552__bF$buf2),
    .D(_4491_),
    .Y(_5968_)
);

NOR2X1 _15500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5967_),
    .B(_5968_),
    .Y(_5969_)
);

AOI22X1 _15501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [11]),
    .C(\datapath_1.regfile_1.regOut[11] [11]),
    .D(_5496_),
    .Y(_5970_)
);

INVX4 _15502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504__bF$buf3),
    .Y(_5971_)
);

AOI22X1 _15503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .B(_5579_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_5972_)
);

NAND3X1 _15504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5970_),
    .B(_5972_),
    .C(_5969_),
    .Y(_5973_)
);

INVX1 _15505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_5974_)
);

OAI22X1 _15506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5974_),
    .B(_5469__bF$buf2),
    .C(_5472__bF$buf1),
    .D(_4509_),
    .Y(_5975_)
);

AOI21X1 _15507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .B(_5649_),
    .C(_5975_),
    .Y(_5976_)
);

AOI22X1 _15508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [11]),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_5977_)
);

AOI22X1 _15509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [11]),
    .B(_5571_),
    .C(_5570__bF$buf1),
    .D(\datapath_1.regfile_1.regOut[27] [11]),
    .Y(_5978_)
);

NAND3X1 _15510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5977_),
    .B(_5978_),
    .C(_5976_),
    .Y(_5979_)
);

NOR2X1 _15511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5979_),
    .B(_5973_),
    .Y(_5980_)
);

NOR3X1 _15512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf2),
    .B(_4481_),
    .C(_5521__bF$buf2),
    .Y(_5981_)
);

NAND3X1 _15513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf1),
    .Y(_5982_)
);

OAI21X1 _15514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf1),
    .B(_4482_),
    .C(_5982_),
    .Y(_5983_)
);

INVX1 _15515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [11]),
    .Y(_5984_)
);

INVX1 _15516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_5985_)
);

OAI22X1 _15517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_5984_),
    .C(_5985_),
    .D(_5499__bF$buf2),
    .Y(_5986_)
);

NOR2X1 _15518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5983_),
    .B(_5986_),
    .Y(_5987_)
);

NAND3X1 _15519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf3),
    .Y(_5988_)
);

OAI21X1 _15520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4510_),
    .B(_5535__bF$buf0),
    .C(_5988_),
    .Y(_5989_)
);

OAI22X1 _15521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf0),
    .B(_4484_),
    .C(_5483__bF$buf3),
    .D(_4495_),
    .Y(_5990_)
);

NOR2X1 _15522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5989_),
    .B(_5990_),
    .Y(_5991_)
);

NAND2X1 _15523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5987_),
    .B(_5991_),
    .Y(_5992_)
);

OAI22X1 _15524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_4517_),
    .C(_4500_),
    .D(_5526__bF$buf3),
    .Y(_5993_)
);

INVX1 _15525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_5994_)
);

INVX1 _15526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_5995_)
);

OAI22X1 _15527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518__bF$buf0),
    .B(_5995_),
    .C(_5503__bF$buf1),
    .D(_5994_),
    .Y(_5996_)
);

NOR2X1 _15528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5996_),
    .B(_5993_),
    .Y(_5997_)
);

INVX1 _15529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_5998_)
);

OAI22X1 _15530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf4),
    .B(_4503_),
    .C(_5998_),
    .D(_5549__bF$buf3),
    .Y(_5999_)
);

INVX1 _15531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_6000_)
);

OAI22X1 _15532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4494_),
    .B(_5544__bF$buf2),
    .C(_5523_),
    .D(_6000_),
    .Y(_6001_)
);

NOR2X1 _15533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5999_),
    .B(_6001_),
    .Y(_6002_)
);

NAND2X1 _15534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6002_),
    .B(_5997_),
    .Y(_6003_)
);

NOR3X1 _15535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5992_),
    .B(_5981_),
    .C(_6003_),
    .Y(_6004_)
);

AOI21X1 _15536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5980_),
    .B(_6004_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [11])
);

AOI22X1 _15537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [12]),
    .C(\datapath_1.regfile_1.regOut[9] [12]),
    .D(_5560_),
    .Y(_6005_)
);

AOI22X1 _15538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [12]),
    .C(\datapath_1.regfile_1.regOut[6] [12]),
    .D(_5565__bF$buf1),
    .Y(_6006_)
);

OAI22X1 _15539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf2),
    .B(_4552_),
    .C(_4560_),
    .D(_5534__bF$buf3),
    .Y(_6007_)
);

OAI22X1 _15540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf2),
    .B(_4556_),
    .C(_5466__bF$buf2),
    .D(_4528_),
    .Y(_6008_)
);

NOR2X1 _15541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6007_),
    .B(_6008_),
    .Y(_6009_)
);

NAND3X1 _15542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6005_),
    .B(_6006_),
    .C(_6009_),
    .Y(_6010_)
);

INVX1 _15543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_6011_)
);

OAI22X1 _15544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf1),
    .B(_6011_),
    .C(_5527__bF$buf2),
    .D(_4553_),
    .Y(_6012_)
);

AOI21X1 _15545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [12]),
    .B(_5486_),
    .C(_6012_),
    .Y(_6013_)
);

AOI22X1 _15546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .B(_5577_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_6014_)
);

AOI22X1 _15547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [12]),
    .B(_5567_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_6015_)
);

NAND3X1 _15548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6014_),
    .B(_6015_),
    .C(_6013_),
    .Y(_6016_)
);

NOR2X1 _15549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6016_),
    .B(_6010_),
    .Y(_6017_)
);

NOR3X1 _15550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf1),
    .B(_4543_),
    .C(_5521__bF$buf1),
    .Y(_6018_)
);

OAI22X1 _15551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .B(_5501_),
    .C(_5524__bF$buf0),
    .D(_4526_),
    .Y(_6019_)
);

INVX1 _15552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_6020_)
);

INVX1 _15553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_6021_)
);

OAI22X1 _15554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499__bF$buf1),
    .B(_6021_),
    .C(_5532__bF$buf1),
    .D(_6020_),
    .Y(_6022_)
);

NOR2X1 _15555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6019_),
    .B(_6022_),
    .Y(_6023_)
);

NAND3X1 _15556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf2),
    .Y(_6024_)
);

OAI21X1 _15557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4557_),
    .B(_5535__bF$buf4),
    .C(_6024_),
    .Y(_6025_)
);

OAI22X1 _15558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_4550_),
    .C(_4533_),
    .D(_5483__bF$buf2),
    .Y(_6026_)
);

NOR2X1 _15559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6025_),
    .B(_6026_),
    .Y(_6027_)
);

NAND2X1 _15560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6023_),
    .B(_6027_),
    .Y(_6028_)
);

INVX1 _15561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_6029_)
);

OAI22X1 _15562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4525_),
    .B(_5545__bF$buf2),
    .C(_5548__bF$buf3),
    .D(_6029_),
    .Y(_6030_)
);

OAI22X1 _15563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf0),
    .B(_4539_),
    .C(_5552__bF$buf1),
    .D(_4559_),
    .Y(_6031_)
);

NOR2X1 _15564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6030_),
    .B(_6031_),
    .Y(_6032_)
);

NOR2X1 _15565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4566_),
    .B(_5539__bF$buf2),
    .Y(_6033_)
);

INVX1 _15566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [12]),
    .Y(_6034_)
);

NAND3X1 _15567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [24]),
    .B(_5460_),
    .C(_5462_),
    .Y(_6035_)
);

NOR3X1 _15568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6034_),
    .B(_5459__bF$buf2),
    .C(_6035_),
    .Y(_6036_)
);

OAI22X1 _15569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518__bF$buf3),
    .B(_4544_),
    .C(_5469__bF$buf1),
    .D(_4567_),
    .Y(_6037_)
);

NOR3X1 _15570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6037_),
    .B(_6033_),
    .C(_6036_),
    .Y(_6038_)
);

NAND2X1 _15571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6038_),
    .B(_6032_),
    .Y(_6039_)
);

NOR3X1 _15572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6018_),
    .B(_6039_),
    .C(_6028_),
    .Y(_6040_)
);

AOI21X1 _15573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6017_),
    .B(_6040_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [12])
);

AOI22X1 _15574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_6041_)
);

AOI22X1 _15575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [13]),
    .B(_5567_),
    .C(_5565__bF$buf0),
    .D(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_6042_)
);

OAI22X1 _15576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_4613_),
    .C(_4612_),
    .D(_5552__bF$buf0),
    .Y(_6043_)
);

INVX1 _15577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_6044_)
);

OAI22X1 _15578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527__bF$buf1),
    .B(_4609_),
    .C(_6044_),
    .D(_5532__bF$buf0),
    .Y(_6045_)
);

NOR2X1 _15579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .B(_6043_),
    .Y(_6046_)
);

NAND3X1 _15580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .B(_6042_),
    .C(_6046_),
    .Y(_6047_)
);

OAI22X1 _15581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4586_),
    .B(_5518__bF$buf2),
    .C(_5548__bF$buf2),
    .D(_4599_),
    .Y(_6048_)
);

AOI21X1 _15582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [13]),
    .B(_5490_),
    .C(_6048_),
    .Y(_6049_)
);

AOI22X1 _15583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [13]),
    .B(_5571_),
    .C(_5570__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[27] [13]),
    .Y(_6050_)
);

AOI22X1 _15584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .B(_5577_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_6051_)
);

NAND3X1 _15585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6050_),
    .B(_6051_),
    .C(_6049_),
    .Y(_6052_)
);

NOR2X1 _15586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6052_),
    .B(_6047_),
    .Y(_6053_)
);

NOR3X1 _15587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf0),
    .B(_4598_),
    .C(_5521__bF$buf0),
    .Y(_6054_)
);

NAND3X1 _15588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf4),
    .Y(_6055_)
);

OAI21X1 _15589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf3),
    .B(_4578_),
    .C(_6055_),
    .Y(_6056_)
);

INVX1 _15590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [13]),
    .Y(_6057_)
);

INVX1 _15591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_6058_)
);

OAI22X1 _15592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_6057_),
    .C(_6058_),
    .D(_5499__bF$buf0),
    .Y(_6059_)
);

NOR2X1 _15593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6056_),
    .B(_6059_),
    .Y(_6060_)
);

NAND3X1 _15594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .B(_5471__bF$buf3),
    .C(_5531__bF$buf1),
    .Y(_6061_)
);

OAI21X1 _15595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4601_),
    .B(_5535__bF$buf3),
    .C(_6061_),
    .Y(_6062_)
);

OAI22X1 _15596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf4),
    .B(_4588_),
    .C(_5483__bF$buf1),
    .D(_4580_),
    .Y(_6063_)
);

NOR2X1 _15597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6062_),
    .B(_6063_),
    .Y(_6064_)
);

NAND2X1 _15598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6060_),
    .B(_6064_),
    .Y(_6065_)
);

OAI22X1 _15599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4602_),
    .B(_5539__bF$buf1),
    .C(_5526__bF$buf2),
    .D(_4606_),
    .Y(_6066_)
);

INVX1 _15600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_6067_)
);

OAI22X1 _15601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_6067_),
    .C(_4585_),
    .D(_5530__bF$buf1),
    .Y(_6068_)
);

NOR2X1 _15602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6068_),
    .B(_6066_),
    .Y(_6069_)
);

OAI22X1 _15603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495__bF$buf2),
    .B(_4589_),
    .C(_4616_),
    .D(_5534__bF$buf2),
    .Y(_6070_)
);

INVX1 _15604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [13]),
    .Y(_6071_)
);

INVX1 _15605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_6072_)
);

OAI22X1 _15606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf1),
    .B(_6072_),
    .C(_5466__bF$buf1),
    .D(_6071_),
    .Y(_6073_)
);

NOR2X1 _15607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6070_),
    .B(_6073_),
    .Y(_6074_)
);

NAND2X1 _15608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6069_),
    .B(_6074_),
    .Y(_6075_)
);

NOR3X1 _15609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6065_),
    .B(_6054_),
    .C(_6075_),
    .Y(_6076_)
);

AOI21X1 _15610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6053_),
    .B(_6076_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [13])
);

OAI22X1 _15611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504__bF$buf2),
    .B(_4664_),
    .C(_5527__bF$buf0),
    .D(_4638_),
    .Y(_6077_)
);

INVX1 _15612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [14]),
    .Y(_6078_)
);

INVX1 _15613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_6079_)
);

OAI22X1 _15614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .B(_6078_),
    .C(_5523_),
    .D(_6079_),
    .Y(_6080_)
);

NOR2X1 _15615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6077_),
    .B(_6080_),
    .Y(_6081_)
);

AOI22X1 _15616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [14]),
    .B(_5494_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_6082_)
);

AOI22X1 _15617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .B(_5577_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_6083_)
);

NAND3X1 _15618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6082_),
    .B(_6083_),
    .C(_6081_),
    .Y(_6084_)
);

NAND2X1 _15619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .B(_5606_),
    .Y(_6085_)
);

AOI22X1 _15620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [14]),
    .C(\datapath_1.regfile_1.regOut[22] [14]),
    .D(_5650_),
    .Y(_6086_)
);

INVX1 _15621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [14]),
    .Y(_6087_)
);

OAI22X1 _15622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544__bF$buf1),
    .B(_6087_),
    .C(_5545__bF$buf1),
    .D(_4654_),
    .Y(_6088_)
);

INVX1 _15623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_6089_)
);

NOR2X1 _15624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6089_),
    .B(_5539__bF$buf0),
    .Y(_6090_)
);

INVX1 _15625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_6091_)
);

NOR2X1 _15626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6091_),
    .B(_5530__bF$buf0),
    .Y(_6092_)
);

NOR3X1 _15627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6088_),
    .B(_6090_),
    .C(_6092_),
    .Y(_6093_)
);

NAND3X1 _15628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6085_),
    .B(_6086_),
    .C(_6093_),
    .Y(_6094_)
);

NOR2X1 _15629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6084_),
    .B(_6094_),
    .Y(_6095_)
);

NOR3X1 _15630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf3),
    .B(_4656_),
    .C(_5521__bF$buf3),
    .Y(_6096_)
);

NAND3X1 _15631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf2),
    .Y(_6097_)
);

OAI21X1 _15632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf2),
    .B(_4661_),
    .C(_6097_),
    .Y(_6098_)
);

OAI22X1 _15633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_4653_),
    .C(_4635_),
    .D(_5499__bF$buf3),
    .Y(_6099_)
);

NOR2X1 _15634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6098_),
    .B(_6099_),
    .Y(_6100_)
);

INVX1 _15635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_6101_)
);

NAND3X1 _15636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf0),
    .Y(_6102_)
);

OAI21X1 _15637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6101_),
    .B(_5535__bF$buf2),
    .C(_6102_),
    .Y(_6103_)
);

INVX1 _15638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [14]),
    .Y(_6104_)
);

OAI22X1 _15639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf3),
    .B(_6104_),
    .C(_5483__bF$buf0),
    .D(_4621_),
    .Y(_6105_)
);

NOR2X1 _15640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6103_),
    .B(_6105_),
    .Y(_6106_)
);

NAND2X1 _15641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6100_),
    .B(_6106_),
    .Y(_6107_)
);

OAI22X1 _15642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4634_),
    .B(_5548__bF$buf1),
    .C(_5526__bF$buf1),
    .D(_4657_),
    .Y(_6108_)
);

INVX1 _15643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_6109_)
);

OAI22X1 _15644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf2),
    .B(_4660_),
    .C(_6109_),
    .D(_5495__bF$buf1),
    .Y(_6110_)
);

NOR2X1 _15645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6110_),
    .B(_6108_),
    .Y(_6111_)
);

OAI22X1 _15646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_4649_),
    .C(_4663_),
    .D(_5534__bF$buf1),
    .Y(_6112_)
);

OAI22X1 _15647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf0),
    .B(_4625_),
    .C(_5466__bF$buf0),
    .D(_4622_),
    .Y(_6113_)
);

NOR2X1 _15648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6112_),
    .B(_6113_),
    .Y(_6114_)
);

NAND2X1 _15649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6111_),
    .B(_6114_),
    .Y(_6115_)
);

NOR3X1 _15650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .B(_6096_),
    .C(_6115_),
    .Y(_6116_)
);

AOI21X1 _15651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6095_),
    .B(_6116_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [14])
);

AOI22X1 _15652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [15]),
    .C(\datapath_1.regfile_1.regOut[22] [15]),
    .D(_5650_),
    .Y(_6117_)
);

INVX1 _15653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_6118_)
);

NOR2X1 _15654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6118_),
    .B(_5549__bF$buf4),
    .Y(_6119_)
);

INVX1 _15655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_6120_)
);

NOR3X1 _15656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6120_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6121_)
);

NOR2X1 _15657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4674_),
    .B(_5534__bF$buf0),
    .Y(_6122_)
);

NOR3X1 _15658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6119_),
    .B(_6121_),
    .C(_6122_),
    .Y(_6123_)
);

AOI22X1 _15659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .B(_5693_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_6124_)
);

NAND3X1 _15660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6117_),
    .B(_6124_),
    .C(_6123_),
    .Y(_6125_)
);

AOI22X1 _15661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_6126_)
);

AOI22X1 _15662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [15]),
    .C(\datapath_1.regfile_1.regOut[5] [15]),
    .D(_5700_),
    .Y(_6127_)
);

OAI22X1 _15663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf0),
    .B(_4706_),
    .C(_4688_),
    .D(_5527__bF$buf4),
    .Y(_6128_)
);

INVX1 _15664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_6129_)
);

OAI22X1 _15665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4687_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf0),
    .D(_6129_),
    .Y(_6130_)
);

NOR2X1 _15666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6130_),
    .B(_6128_),
    .Y(_6131_)
);

NAND3X1 _15667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6126_),
    .B(_6127_),
    .C(_6131_),
    .Y(_6132_)
);

NOR2X1 _15668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6132_),
    .B(_6125_),
    .Y(_6133_)
);

NAND2X1 _15669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [15]),
    .B(_5649_),
    .Y(_6134_)
);

INVX1 _15670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [15]),
    .Y(_6135_)
);

INVX1 _15671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [15]),
    .Y(_6136_)
);

OAI22X1 _15672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6135_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf2),
    .D(_6136_),
    .Y(_6137_)
);

INVX1 _15673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [15]),
    .Y(_6138_)
);

OAI22X1 _15674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4670_),
    .B(_5544__bF$buf0),
    .C(_5480__bF$buf2),
    .D(_6138_),
    .Y(_6139_)
);

NOR2X1 _15675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6139_),
    .B(_6137_),
    .Y(_6140_)
);

INVX1 _15676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [15]),
    .Y(_6141_)
);

OAI22X1 _15677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_6141_),
    .C(_4684_),
    .D(_5483__bF$buf4),
    .Y(_6142_)
);

AOI21X1 _15678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [15]),
    .B(_5570__bF$buf2),
    .C(_6142_),
    .Y(_6143_)
);

NAND3X1 _15679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6134_),
    .B(_6140_),
    .C(_6143_),
    .Y(_6144_)
);

NAND3X1 _15680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6145_)
);

OAI22X1 _15681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4696_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf1),
    .D(_4695_),
    .Y(_6146_)
);

INVX1 _15682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_6147_)
);

OAI22X1 _15683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6147_),
    .B(_5548__bF$buf0),
    .C(_5489__bF$buf0),
    .D(_4707_),
    .Y(_6148_)
);

NOR2X1 _15684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6148_),
    .B(_6146_),
    .Y(_6149_)
);

INVX1 _15685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_6150_)
);

OAI22X1 _15686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6150_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf0),
    .D(_4672_),
    .Y(_6151_)
);

OAI22X1 _15687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf1),
    .B(_4704_),
    .C(_4703_),
    .D(_5504__bF$buf1),
    .Y(_6152_)
);

NOR2X1 _15688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6151_),
    .B(_6152_),
    .Y(_6153_)
);

NAND3X1 _15689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6149_),
    .B(_6153_),
    .C(_6145_),
    .Y(_6154_)
);

NOR2X1 _15690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .B(_6154_),
    .Y(_6155_)
);

AOI21X1 _15691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6155_),
    .B(_6133_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [15])
);

OAI22X1 _15692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4743_),
    .B(_5535__bF$buf1),
    .C(_5569_),
    .D(_4717_),
    .Y(_6156_)
);

OAI22X1 _15693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf3),
    .B(_4732_),
    .C(_5532__bF$buf3),
    .D(_4731_),
    .Y(_6157_)
);

NOR2X1 _15694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6156_),
    .B(_6157_),
    .Y(_6158_)
);

AOI22X1 _15695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [16]),
    .C(\datapath_1.regfile_1.regOut[26] [16]),
    .D(_5484_),
    .Y(_6159_)
);

AOI22X1 _15696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5562_),
    .B(\datapath_1.regfile_1.regOut[25] [16]),
    .C(\datapath_1.regfile_1.regOut[22] [16]),
    .D(_5650_),
    .Y(_6160_)
);

NAND3X1 _15697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6159_),
    .B(_6160_),
    .C(_6158_),
    .Y(_6161_)
);

INVX1 _15698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [16]),
    .Y(_6162_)
);

NOR2X1 _15699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6162_),
    .B(_5544__bF$buf3),
    .Y(_6163_)
);

NOR2X1 _15700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4753_),
    .B(_5534__bF$buf4),
    .Y(_6164_)
);

NOR3X1 _15701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4735_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6165_)
);

NOR3X1 _15702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6163_),
    .B(_6165_),
    .C(_6164_),
    .Y(_6166_)
);

AOI22X1 _15703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .B(_5494_),
    .C(_5479_),
    .D(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_6167_)
);

AOI22X1 _15704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5481_),
    .B(\datapath_1.regfile_1.regOut[30] [16]),
    .C(\datapath_1.regfile_1.regOut[29] [16]),
    .D(_5486_),
    .Y(_6168_)
);

NAND3X1 _15705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6167_),
    .B(_6168_),
    .C(_6166_),
    .Y(_6169_)
);

NOR2X1 _15706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6161_),
    .B(_6169_),
    .Y(_6170_)
);

INVX1 _15707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_6171_)
);

NOR3X1 _15708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf2),
    .B(_6171_),
    .C(_5521__bF$buf2),
    .Y(_6172_)
);

INVX1 _15709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_6173_)
);

INVX1 _15710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_6174_)
);

OAI22X1 _15711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6173_),
    .B(_5548__bF$buf4),
    .C(_5489__bF$buf3),
    .D(_6174_),
    .Y(_6175_)
);

INVX1 _15712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_6176_)
);

OAI22X1 _15713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4714_),
    .B(_5503__bF$buf3),
    .C(_5495__bF$buf3),
    .D(_6176_),
    .Y(_6177_)
);

NOR2X1 _15714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6175_),
    .B(_6177_),
    .Y(_6178_)
);

NOR3X1 _15715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4728_),
    .B(\datapath_1.PCJump_27_bF$buf0 ),
    .C(_5519_),
    .Y(_6179_)
);

INVX1 _15716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_6180_)
);

NOR2X1 _15717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6180_),
    .B(_5501_),
    .Y(_6181_)
);

OAI22X1 _15718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4718_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf3),
    .D(_4751_),
    .Y(_6182_)
);

NOR3X1 _15719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6182_),
    .B(_6179_),
    .C(_6181_),
    .Y(_6183_)
);

NAND2X1 _15720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6183_),
    .B(_6178_),
    .Y(_6184_)
);

OAI22X1 _15721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504__bF$buf0),
    .B(_4724_),
    .C(_5527__bF$buf3),
    .D(_4715_),
    .Y(_6185_)
);

INVX1 _15722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [16]),
    .Y(_6186_)
);

INVX1 _15723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_6187_)
);

OAI22X1 _15724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6186_),
    .B(_5545__bF$buf3),
    .C(_5530__bF$buf3),
    .D(_6187_),
    .Y(_6188_)
);

NOR2X1 _15725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6188_),
    .B(_6185_),
    .Y(_6189_)
);

OAI22X1 _15726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5523_),
    .B(_4744_),
    .C(_4754_),
    .D(_5524__bF$buf1),
    .Y(_6190_)
);

INVX1 _15727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_6191_)
);

OAI22X1 _15728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf0),
    .B(_6191_),
    .C(_5526__bF$buf4),
    .D(_4725_),
    .Y(_6192_)
);

NOR2X1 _15729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6192_),
    .B(_6190_),
    .Y(_6193_)
);

NAND2X1 _15730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6189_),
    .B(_6193_),
    .Y(_6194_)
);

NOR3X1 _15731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6172_),
    .B(_6184_),
    .C(_6194_),
    .Y(_6195_)
);

AOI21X1 _15732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6170_),
    .B(_6195_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [16])
);

AOI22X1 _15733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5557_),
    .B(\datapath_1.regfile_1.regOut[17] [17]),
    .C(\datapath_1.regfile_1.regOut[18] [17]),
    .D(_5558_),
    .Y(_6196_)
);

NAND2X1 _15734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .B(_5560_),
    .Y(_6197_)
);

NAND2X1 _15735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [17]),
    .B(_5562_),
    .Y(_6198_)
);

NAND3X1 _15736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6197_),
    .B(_6198_),
    .C(_6196_),
    .Y(_6199_)
);

NAND2X1 _15737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [17]),
    .B(_5565__bF$buf2),
    .Y(_6200_)
);

NAND2X1 _15738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [17]),
    .B(_5570__bF$buf1),
    .Y(_6201_)
);

AOI22X1 _15739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5567_),
    .B(\datapath_1.regfile_1.regOut[28] [17]),
    .C(\datapath_1.regfile_1.regOut[31] [17]),
    .D(_5571_),
    .Y(_6202_)
);

NAND3X1 _15740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6202_),
    .B(_6201_),
    .C(_6200_),
    .Y(_6203_)
);

OAI22X1 _15741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4795_),
    .B(_5539__bF$buf2),
    .C(_5469__bF$buf2),
    .D(_4765_),
    .Y(_6204_)
);

AOI21X1 _15742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .B(_5494_),
    .C(_6204_),
    .Y(_6205_)
);

AOI22X1 _15743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_6206_)
);

AOI22X1 _15744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .B(_5579_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_6207_)
);

NAND3X1 _15745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6205_),
    .B(_6207_),
    .C(_6206_),
    .Y(_6208_)
);

NOR3X1 _15746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6208_),
    .B(_6203_),
    .C(_6199_),
    .Y(_6209_)
);

INVX1 _15747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_6210_)
);

NOR3X1 _15748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf1),
    .B(_6210_),
    .C(_5521__bF$buf1),
    .Y(_6211_)
);

INVX1 _15749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_6212_)
);

OAI22X1 _15750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf2),
    .B(_4787_),
    .C(_5532__bF$buf2),
    .D(_6212_),
    .Y(_6213_)
);

INVX1 _15751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_6214_)
);

OAI22X1 _15752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf0),
    .B(_6214_),
    .C(_5552__bF$buf3),
    .D(_4779_),
    .Y(_6215_)
);

NOR2X1 _15753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6215_),
    .B(_6213_),
    .Y(_6216_)
);

OAI22X1 _15754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_4774_),
    .C(_4762_),
    .D(_5527__bF$buf2),
    .Y(_6217_)
);

INVX1 _15755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_6218_)
);

OAI22X1 _15756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf2),
    .B(_6218_),
    .C(_4771_),
    .D(_5504__bF$buf4),
    .Y(_6219_)
);

NOR2X1 _15757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6219_),
    .B(_6217_),
    .Y(_6220_)
);

NAND2X1 _15758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6216_),
    .B(_6220_),
    .Y(_6221_)
);

NAND3X1 _15759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .B(_5500__bF$buf2),
    .C(_5471__bF$buf0),
    .Y(_6222_)
);

OAI21X1 _15760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf0),
    .B(_4798_),
    .C(_6222_),
    .Y(_6223_)
);

OAI22X1 _15761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_4789_),
    .C(_4775_),
    .D(_5499__bF$buf2),
    .Y(_6224_)
);

NOR2X1 _15762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6223_),
    .B(_6224_),
    .Y(_6225_)
);

INVX1 _15763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_6226_)
);

NAND3X1 _15764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf4),
    .Y(_6227_)
);

OAI21X1 _15765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6226_),
    .B(_5535__bF$buf0),
    .C(_6227_),
    .Y(_6228_)
);

OAI22X1 _15766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf1),
    .B(_4790_),
    .C(_5483__bF$buf3),
    .D(_4802_),
    .Y(_6229_)
);

NOR2X1 _15767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6228_),
    .B(_6229_),
    .Y(_6230_)
);

NAND2X1 _15768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6225_),
    .B(_6230_),
    .Y(_6231_)
);

NOR3X1 _15769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6231_),
    .B(_6211_),
    .C(_6221_),
    .Y(_6232_)
);

AOI21X1 _15770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6209_),
    .B(_6232_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [17])
);

AOI22X1 _15771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_6233_)
);

AOI22X1 _15772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5481_),
    .B(\datapath_1.regfile_1.regOut[30] [18]),
    .C(\datapath_1.regfile_1.regOut[6] [18]),
    .D(_5565__bF$buf1),
    .Y(_6234_)
);

INVX1 _15773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_6235_)
);

OAI22X1 _15774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_6235_),
    .C(_5527__bF$buf1),
    .D(_4812_),
    .Y(_6236_)
);

OAI22X1 _15775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4810_),
    .B(_5539__bF$buf1),
    .C(_5552__bF$buf2),
    .D(_4828_),
    .Y(_6237_)
);

NOR2X1 _15776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6236_),
    .B(_6237_),
    .Y(_6238_)
);

NAND3X1 _15777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6233_),
    .B(_6234_),
    .C(_6238_),
    .Y(_6239_)
);

NAND2X1 _15778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .B(_5490_),
    .Y(_6240_)
);

AOI22X1 _15779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_6241_)
);

OAI22X1 _15780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .B(_4843_),
    .C(_5483__bF$buf2),
    .D(_4840_),
    .Y(_6242_)
);

INVX1 _15781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_6243_)
);

INVX1 _15782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_6244_)
);

OAI22X1 _15783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6244_),
    .B(_5503__bF$buf2),
    .C(_5504__bF$buf3),
    .D(_6243_),
    .Y(_6245_)
);

NOR2X1 _15784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6245_),
    .B(_6242_),
    .Y(_6246_)
);

NAND3X1 _15785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6240_),
    .B(_6241_),
    .C(_6246_),
    .Y(_6247_)
);

NOR2X1 _15786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6247_),
    .B(_6239_),
    .Y(_6248_)
);

INVX1 _15787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_6249_)
);

NOR3X1 _15788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf0),
    .B(_6249_),
    .C(_5521__bF$buf0),
    .Y(_6250_)
);

NAND3X1 _15789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [18]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf4),
    .Y(_6251_)
);

OAI21X1 _15790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf3),
    .B(_4820_),
    .C(_6251_),
    .Y(_6252_)
);

INVX1 _15791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [18]),
    .Y(_6253_)
);

OAI22X1 _15792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6253_),
    .B(_5544__bF$buf2),
    .C(_5499__bF$buf1),
    .D(_4841_),
    .Y(_6254_)
);

NOR2X1 _15793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6252_),
    .B(_6254_),
    .Y(_6255_)
);

NAND3X1 _15794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .B(_5471__bF$buf3),
    .C(_5531__bF$buf3),
    .Y(_6256_)
);

OAI21X1 _15795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4809_),
    .B(_5535__bF$buf4),
    .C(_6256_),
    .Y(_6257_)
);

INVX1 _15796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [18]),
    .Y(_6258_)
);

INVX1 _15797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [18]),
    .Y(_6259_)
);

OAI22X1 _15798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6258_),
    .B(_5545__bF$buf2),
    .C(_5466__bF$buf3),
    .D(_6259_),
    .Y(_6260_)
);

NOR2X1 _15799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6257_),
    .B(_6260_),
    .Y(_6261_)
);

NAND2X1 _15800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6255_),
    .B(_6261_),
    .Y(_6262_)
);

OAI22X1 _15801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf1),
    .B(_4819_),
    .C(_5532__bF$buf1),
    .D(_4823_),
    .Y(_6263_)
);

OAI22X1 _15802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_4835_),
    .C(_4832_),
    .D(_5526__bF$buf3),
    .Y(_6264_)
);

NOR2X1 _15803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6263_),
    .B(_6264_),
    .Y(_6265_)
);

INVX1 _15804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_6266_)
);

OAI22X1 _15805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6266_),
    .B(_5548__bF$buf3),
    .C(_5534__bF$buf3),
    .D(_4831_),
    .Y(_6267_)
);

INVX1 _15806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [18]),
    .Y(_6268_)
);

INVX1 _15807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_6269_)
);

OAI22X1 _15808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf0),
    .B(_6268_),
    .C(_6269_),
    .D(_5549__bF$buf2),
    .Y(_6270_)
);

NOR2X1 _15809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6267_),
    .B(_6270_),
    .Y(_6271_)
);

NAND2X1 _15810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6271_),
    .B(_6265_),
    .Y(_6272_)
);

NOR3X1 _15811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6262_),
    .B(_6250_),
    .C(_6272_),
    .Y(_6273_)
);

AOI21X1 _15812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6248_),
    .B(_6273_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [18])
);

OAI22X1 _15813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf1),
    .B(_4885_),
    .C(_5527__bF$buf0),
    .D(_4874_),
    .Y(_6274_)
);

INVX1 _15814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [19]),
    .Y(_6275_)
);

OAI22X1 _15815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .B(_6275_),
    .C(_5523_),
    .D(_4884_),
    .Y(_6276_)
);

NOR2X1 _15816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6274_),
    .B(_6276_),
    .Y(_6277_)
);

AOI22X1 _15817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .B(_5494_),
    .C(_5479_),
    .D(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_6278_)
);

AOI22X1 _15818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .B(_5577_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_6279_)
);

NAND3X1 _15819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6278_),
    .B(_6279_),
    .C(_6277_),
    .Y(_6280_)
);

OAI22X1 _15820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4877_),
    .B(_5539__bF$buf0),
    .C(_5552__bF$buf1),
    .D(_4853_),
    .Y(_6281_)
);

AOI21X1 _15821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .B(_5606_),
    .C(_6281_),
    .Y(_6282_)
);

AOI22X1 _15822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5567_),
    .B(\datapath_1.regfile_1.regOut[28] [19]),
    .C(\datapath_1.regfile_1.regOut[31] [19]),
    .D(_5571_),
    .Y(_6283_)
);

AOI22X1 _15823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5649_),
    .B(\datapath_1.regfile_1.regOut[23] [19]),
    .C(\datapath_1.regfile_1.regOut[21] [19]),
    .D(_5685_),
    .Y(_6284_)
);

NAND3X1 _15824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6283_),
    .B(_6284_),
    .C(_6282_),
    .Y(_6285_)
);

NOR2X1 _15825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6285_),
    .B(_6280_),
    .Y(_6286_)
);

INVX1 _15826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_6287_)
);

NOR3X1 _15827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf3),
    .B(_6287_),
    .C(_5521__bF$buf3),
    .Y(_6288_)
);

NAND3X1 _15828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf2),
    .Y(_6289_)
);

OAI21X1 _15829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf2),
    .B(_4865_),
    .C(_6289_),
    .Y(_6290_)
);

INVX1 _15830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [19]),
    .Y(_6291_)
);

INVX1 _15831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_6292_)
);

OAI22X1 _15832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_6291_),
    .C(_6292_),
    .D(_5499__bF$buf0),
    .Y(_6293_)
);

NOR2X1 _15833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6290_),
    .B(_6293_),
    .Y(_6294_)
);

INVX1 _15834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_6295_)
);

NAND3X1 _15835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf2),
    .Y(_6296_)
);

OAI21X1 _15836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6295_),
    .B(_5535__bF$buf3),
    .C(_6296_),
    .Y(_6297_)
);

INVX1 _15837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [19]),
    .Y(_6298_)
);

OAI22X1 _15838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf4),
    .B(_6298_),
    .C(_5483__bF$buf1),
    .D(_4869_),
    .Y(_6299_)
);

NOR2X1 _15839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6297_),
    .B(_6299_),
    .Y(_6300_)
);

NAND2X1 _15840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6294_),
    .B(_6300_),
    .Y(_6301_)
);

OAI22X1 _15841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4856_),
    .B(_5548__bF$buf2),
    .C(_5526__bF$buf2),
    .D(_4875_),
    .Y(_6302_)
);

OAI22X1 _15842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf3),
    .B(_4861_),
    .C(_4864_),
    .D(_5495__bF$buf2),
    .Y(_6303_)
);

NOR2X1 _15843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6303_),
    .B(_6302_),
    .Y(_6304_)
);

INVX1 _15844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_6305_)
);

OAI22X1 _15845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf2),
    .B(_4888_),
    .C(_5532__bF$buf0),
    .D(_6305_),
    .Y(_6306_)
);

INVX1 _15846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [19]),
    .Y(_6307_)
);

INVX1 _15847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_6308_)
);

OAI22X1 _15848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf1),
    .B(_6308_),
    .C(_5466__bF$buf2),
    .D(_6307_),
    .Y(_6309_)
);

NOR2X1 _15849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6309_),
    .B(_6306_),
    .Y(_6310_)
);

NAND2X1 _15850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6304_),
    .B(_6310_),
    .Y(_6311_)
);

NOR3X1 _15851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6301_),
    .B(_6288_),
    .C(_6311_),
    .Y(_6312_)
);

AOI21X1 _15852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6286_),
    .B(_6312_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [19])
);

AOI22X1 _15853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [20]),
    .C(\datapath_1.regfile_1.regOut[22] [20]),
    .D(_5650_),
    .Y(_6313_)
);

INVX2 _15854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527__bF$buf4),
    .Y(_6314_)
);

AOI22X1 _15855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .B(\datapath_1.regfile_1.regOut[7] [20]),
    .C(\datapath_1.regfile_1.regOut[10] [20]),
    .D(_6314_),
    .Y(_6315_)
);

NAND2X1 _15856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6315_),
    .B(_6313_),
    .Y(_6316_)
);

AOI22X1 _15857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [20]),
    .C(\datapath_1.regfile_1.regOut[11] [20]),
    .D(_5496_),
    .Y(_6317_)
);

NAND2X1 _15858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [20]),
    .B(_5579_),
    .Y(_6318_)
);

NAND2X1 _15859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .B(_5971_),
    .Y(_6319_)
);

NAND3X1 _15860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6318_),
    .B(_6319_),
    .C(_6317_),
    .Y(_6320_)
);

OAI22X1 _15861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4898_),
    .B(_5539__bF$buf4),
    .C(_5469__bF$buf1),
    .D(_4924_),
    .Y(_6321_)
);

AOI21X1 _15862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .B(_5649_),
    .C(_6321_),
    .Y(_6322_)
);

AOI22X1 _15863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [20]),
    .C(\datapath_1.regfile_1.regOut[26] [20]),
    .D(_5484_),
    .Y(_6323_)
);

AOI22X1 _15864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [20]),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_6324_)
);

NAND3X1 _15865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6322_),
    .B(_6323_),
    .C(_6324_),
    .Y(_6325_)
);

NOR3X1 _15866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6320_),
    .B(_6316_),
    .C(_6325_),
    .Y(_6326_)
);

NOR3X1 _15867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf2),
    .B(_4910_),
    .C(_5521__bF$buf2),
    .Y(_6327_)
);

NAND3X1 _15868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [20]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf0),
    .Y(_6328_)
);

OAI21X1 _15869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf1),
    .B(_4908_),
    .C(_6328_),
    .Y(_6329_)
);

OAI22X1 _15870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4931_),
    .B(_5544__bF$buf1),
    .C(_5499__bF$buf3),
    .D(_4932_),
    .Y(_6330_)
);

NOR2X1 _15871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6329_),
    .B(_6330_),
    .Y(_6331_)
);

NAND3X1 _15872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf1),
    .Y(_6332_)
);

OAI21X1 _15873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4897_),
    .B(_5535__bF$buf2),
    .C(_6332_),
    .Y(_6333_)
);

INVX1 _15874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [20]),
    .Y(_6334_)
);

OAI22X1 _15875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6334_),
    .B(_5545__bF$buf1),
    .C(_5466__bF$buf1),
    .D(_4934_),
    .Y(_6335_)
);

NOR2X1 _15876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6333_),
    .B(_6335_),
    .Y(_6336_)
);

NAND2X1 _15877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6331_),
    .B(_6336_),
    .Y(_6337_)
);

INVX1 _15878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [20]),
    .Y(_6338_)
);

OAI22X1 _15879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf3),
    .B(_6338_),
    .C(_5526__bF$buf1),
    .D(_4920_),
    .Y(_6339_)
);

INVX1 _15880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_6340_)
);

OAI22X1 _15881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518__bF$buf0),
    .B(_4935_),
    .C(_5503__bF$buf1),
    .D(_6340_),
    .Y(_6341_)
);

NOR2X1 _15882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6341_),
    .B(_6339_),
    .Y(_6342_)
);

INVX1 _15883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_6343_)
);

OAI22X1 _15884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf1),
    .B(_4919_),
    .C(_6343_),
    .D(_5549__bF$buf0),
    .Y(_6344_)
);

INVX1 _15885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [20]),
    .Y(_6345_)
);

INVX1 _15886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_6346_)
);

OAI22X1 _15887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_6345_),
    .C(_5523_),
    .D(_6346_),
    .Y(_6347_)
);

NOR2X1 _15888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6344_),
    .B(_6347_),
    .Y(_6348_)
);

NAND2X1 _15889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6342_),
    .B(_6348_),
    .Y(_6349_)
);

NOR3X1 _15890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6337_),
    .B(_6327_),
    .C(_6349_),
    .Y(_6350_)
);

AOI21X1 _15891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6326_),
    .B(_6350_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [20])
);

NAND2X1 _15892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .B(_5693_),
    .Y(_6351_)
);

NOR2X1 _15893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4986_),
    .B(_5549__bF$buf4),
    .Y(_6352_)
);

NOR2X1 _15894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4968_),
    .B(_5534__bF$buf0),
    .Y(_6353_)
);

NOR3X1 _15895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4978_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6354_)
);

NOR3X1 _15896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6352_),
    .B(_6354_),
    .C(_6353_),
    .Y(_6355_)
);

INVX1 _15897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_6356_)
);

INVX1 _15898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_6357_)
);

OAI22X1 _15899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf0),
    .B(_6357_),
    .C(_5532__bF$buf3),
    .D(_6356_),
    .Y(_6358_)
);

OAI22X1 _15900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_4983_),
    .C(_4982_),
    .D(_5552__bF$buf0),
    .Y(_6359_)
);

NOR2X1 _15901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6358_),
    .B(_6359_),
    .Y(_6360_)
);

NAND3X1 _15902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6351_),
    .B(_6360_),
    .C(_6355_),
    .Y(_6361_)
);

AOI22X1 _15903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [21]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_6362_)
);

AOI22X1 _15904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[6] [21]),
    .C(\datapath_1.regfile_1.regOut[5] [21]),
    .D(_5700_),
    .Y(_6363_)
);

OAI22X1 _15905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf0),
    .B(_4976_),
    .C(_4979_),
    .D(_5527__bF$buf3),
    .Y(_6364_)
);

INVX1 _15906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_6365_)
);

OAI22X1 _15907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6365_),
    .B(_5539__bF$buf3),
    .C(_5469__bF$buf0),
    .D(_4975_),
    .Y(_6366_)
);

NOR2X1 _15908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6366_),
    .B(_6364_),
    .Y(_6367_)
);

NAND3X1 _15909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6362_),
    .B(_6363_),
    .C(_6367_),
    .Y(_6368_)
);

NOR2X1 _15910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6368_),
    .B(_6361_),
    .Y(_6369_)
);

NAND2X1 _15911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [21]),
    .B(_5570__bF$buf3),
    .Y(_6370_)
);

OAI22X1 _15912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_4952_),
    .C(_4955_),
    .D(_5483__bF$buf0),
    .Y(_6371_)
);

AOI21X1 _15913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [21]),
    .B(_5567_),
    .C(_6371_),
    .Y(_6372_)
);

INVX1 _15914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [21]),
    .Y(_6373_)
);

OAI22X1 _15915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6373_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf2),
    .D(_4945_),
    .Y(_6374_)
);

AOI21X1 _15916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [21]),
    .B(_5481_),
    .C(_6374_),
    .Y(_6375_)
);

NAND3X1 _15917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6370_),
    .B(_6375_),
    .C(_6372_),
    .Y(_6376_)
);

NAND3X1 _15918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6377_)
);

INVX1 _15919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_6378_)
);

OAI22X1 _15920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6378_),
    .B(_5518__bF$buf3),
    .C(_5478__bF$buf2),
    .D(_4966_),
    .Y(_6379_)
);

INVX1 _15921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_6380_)
);

OAI22X1 _15922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4969_),
    .B(_5548__bF$buf1),
    .C(_5489__bF$buf0),
    .D(_6380_),
    .Y(_6381_)
);

NOR2X1 _15923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6381_),
    .B(_6379_),
    .Y(_6382_)
);

OAI22X1 _15924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4956_),
    .B(_5503__bF$buf0),
    .C(_5495__bF$buf1),
    .D(_4953_),
    .Y(_6383_)
);

OAI22X1 _15925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf2),
    .B(_4943_),
    .C(_4942_),
    .D(_5504__bF$buf2),
    .Y(_6384_)
);

NOR2X1 _15926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6383_),
    .B(_6384_),
    .Y(_6385_)
);

NAND3X1 _15927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6382_),
    .B(_6385_),
    .C(_6377_),
    .Y(_6386_)
);

NOR2X1 _15928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6376_),
    .B(_6386_),
    .Y(_6387_)
);

AOI21X1 _15929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6387_),
    .B(_6369_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [21])
);

OAI22X1 _15930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504__bF$buf1),
    .B(_5030_),
    .C(_5527__bF$buf2),
    .D(_5010_),
    .Y(_6388_)
);

INVX1 _15931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [22]),
    .Y(_6389_)
);

OAI22X1 _15932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6389_),
    .B(_5544__bF$buf0),
    .C(_5523_),
    .D(_4991_),
    .Y(_6390_)
);

NOR2X1 _15933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6390_),
    .B(_6388_),
    .Y(_6391_)
);

AOI22X1 _15934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .B(_5494_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_6392_)
);

AOI22X1 _15935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .B(_5577_),
    .C(_5479_),
    .D(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_6393_)
);

NAND3X1 _15936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6392_),
    .B(_6393_),
    .C(_6391_),
    .Y(_6394_)
);

OAI22X1 _15937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_5013_),
    .C(_4995_),
    .D(_5552__bF$buf3),
    .Y(_6395_)
);

AOI21X1 _15938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .B(_5606_),
    .C(_6395_),
    .Y(_6396_)
);

AOI22X1 _15939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [22]),
    .B(_5571_),
    .C(_5570__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[27] [22]),
    .Y(_6397_)
);

NOR2X1 _15940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5004_),
    .B(_5539__bF$buf2),
    .Y(_6398_)
);

AOI21X1 _15941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .B(_5649_),
    .C(_6398_),
    .Y(_6399_)
);

NAND3X1 _15942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6399_),
    .C(_6396_),
    .Y(_6400_)
);

NOR2X1 _15943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6394_),
    .B(_6400_),
    .Y(_6401_)
);

NOR3X1 _15944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf1),
    .B(_5003_),
    .C(_5521__bF$buf1),
    .Y(_6402_)
);

NAND3X1 _15945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .B(_5500__bF$buf2),
    .C(_5471__bF$buf4),
    .Y(_6403_)
);

OAI21X1 _15946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf0),
    .B(_5007_),
    .C(_6403_),
    .Y(_6404_)
);

INVX1 _15947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_6405_)
);

OAI22X1 _15948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_4994_),
    .C(_6405_),
    .D(_5499__bF$buf2),
    .Y(_6406_)
);

NOR2X1 _15949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6404_),
    .B(_6406_),
    .Y(_6407_)
);

NAND3X1 _15950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .B(_5471__bF$buf3),
    .C(_5531__bF$buf0),
    .Y(_6408_)
);

OAI21X1 _15951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5006_),
    .B(_5535__bF$buf1),
    .C(_6408_),
    .Y(_6409_)
);

INVX1 _15952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [22]),
    .Y(_6410_)
);

OAI22X1 _15953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf1),
    .B(_6410_),
    .C(_5483__bF$buf4),
    .D(_4998_),
    .Y(_6411_)
);

NOR2X1 _15954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6409_),
    .B(_6411_),
    .Y(_6412_)
);

NAND2X1 _15955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6407_),
    .B(_6412_),
    .Y(_6413_)
);

OAI22X1 _15956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495__bF$buf0),
    .B(_5023_),
    .C(_5526__bF$buf4),
    .D(_5034_),
    .Y(_6414_)
);

INVX1 _15957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_6415_)
);

OAI22X1 _15958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6415_),
    .B(_5548__bF$buf0),
    .C(_5463__bF$buf1),
    .D(_5031_),
    .Y(_6416_)
);

NOR2X1 _15959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6416_),
    .B(_6414_),
    .Y(_6417_)
);

INVX1 _15960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_6418_)
);

OAI22X1 _15961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf4),
    .B(_5021_),
    .C(_5532__bF$buf2),
    .D(_6418_),
    .Y(_6419_)
);

INVX1 _15962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [22]),
    .Y(_6420_)
);

INVX1 _15963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_6421_)
);

OAI22X1 _15964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf3),
    .B(_6421_),
    .C(_5466__bF$buf4),
    .D(_6420_),
    .Y(_6422_)
);

NOR2X1 _15965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6422_),
    .B(_6419_),
    .Y(_6423_)
);

NAND2X1 _15966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6417_),
    .B(_6423_),
    .Y(_6424_)
);

NOR3X1 _15967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6413_),
    .B(_6402_),
    .C(_6424_),
    .Y(_6425_)
);

AOI21X1 _15968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6401_),
    .B(_6425_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [22])
);

AOI22X1 _15969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .B(_5606_),
    .C(_5490_),
    .D(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_6426_)
);

AOI22X1 _15970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [23]),
    .B(_5567_),
    .C(_5565__bF$buf3),
    .D(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_6427_)
);

INVX1 _15971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [23]),
    .Y(_6428_)
);

OAI22X1 _15972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6428_),
    .B(_5545__bF$buf3),
    .C(_5527__bF$buf1),
    .D(_5055_),
    .Y(_6429_)
);

INVX1 _15973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [23]),
    .Y(_6430_)
);

OAI22X1 _15974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_5042_),
    .C(_6430_),
    .D(_5569_),
    .Y(_6431_)
);

NOR2X1 _15975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6431_),
    .B(_6429_),
    .Y(_6432_)
);

NAND3X1 _15976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6426_),
    .B(_6427_),
    .C(_6432_),
    .Y(_6433_)
);

NAND2X1 _15977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .B(_5494_),
    .Y(_6434_)
);

AOI22X1 _15978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .B(_5577_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_6435_)
);

INVX1 _15979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_6436_)
);

OAI22X1 _15980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf3),
    .B(_6436_),
    .C(_5552__bF$buf2),
    .D(_5062_),
    .Y(_6437_)
);

OAI22X1 _15981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5052_),
    .B(_5548__bF$buf4),
    .C(_5504__bF$buf0),
    .D(_5081_),
    .Y(_6438_)
);

NOR2X1 _15982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6438_),
    .B(_6437_),
    .Y(_6439_)
);

NAND3X1 _15983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6434_),
    .B(_6435_),
    .C(_6439_),
    .Y(_6440_)
);

NOR2X1 _15984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6440_),
    .B(_6433_),
    .Y(_6441_)
);

NOR3X1 _15985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf0),
    .B(_5051_),
    .C(_5521__bF$buf0),
    .Y(_6442_)
);

OAI22X1 _15986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5065_),
    .B(_5501_),
    .C(_5524__bF$buf3),
    .D(_5078_),
    .Y(_6443_)
);

OAI22X1 _15987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5499__bF$buf1),
    .B(_5043_),
    .C(_5532__bF$buf1),
    .D(_5039_),
    .Y(_6444_)
);

NOR2X1 _15988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6443_),
    .B(_6444_),
    .Y(_6445_)
);

INVX1 _15989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_6446_)
);

NAND3X1 _15990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf4),
    .Y(_6447_)
);

OAI21X1 _15991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6446_),
    .B(_5535__bF$buf0),
    .C(_6447_),
    .Y(_6448_)
);

OAI22X1 _15992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_5063_),
    .C(_5071_),
    .D(_5483__bF$buf3),
    .Y(_6449_)
);

NOR2X1 _15993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6448_),
    .B(_6449_),
    .Y(_6450_)
);

NAND2X1 _15994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6445_),
    .B(_6450_),
    .Y(_6451_)
);

NAND3X1 _15995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .B(_5477_),
    .C(_5531__bF$buf3),
    .Y(_6452_)
);

OAI21X1 _15996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf3),
    .B(_5074_),
    .C(_6452_),
    .Y(_6453_)
);

OAI22X1 _15997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf1),
    .B(_5066_),
    .C(_5073_),
    .D(_5485__bF$buf0),
    .Y(_6454_)
);

NOR2X1 _15998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6453_),
    .B(_6454_),
    .Y(_6455_)
);

INVX1 _15999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_6456_)
);

OAI22X1 _16000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495__bF$buf3),
    .B(_6456_),
    .C(_5080_),
    .D(_5534__bF$buf3),
    .Y(_6457_)
);

INVX1 _16001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [23]),
    .Y(_6458_)
);

OAI22X1 _16002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf2),
    .B(_5040_),
    .C(_5466__bF$buf3),
    .D(_6458_),
    .Y(_6459_)
);

NOR2X1 _16003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6457_),
    .B(_6459_),
    .Y(_6460_)
);

NAND2X1 _16004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6455_),
    .B(_6460_),
    .Y(_6461_)
);

NOR3X1 _16005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6461_),
    .B(_6442_),
    .C(_6451_),
    .Y(_6462_)
);

AOI21X1 _16006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6441_),
    .B(_6462_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [23])
);

OAI22X1 _16007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5102_),
    .B(_5469__bF$buf3),
    .C(_5463__bF$buf0),
    .D(_5126_),
    .Y(_6463_)
);

OAI22X1 _16008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5099_),
    .B(_5544__bF$buf3),
    .C(_5523_),
    .D(_5107_),
    .Y(_6464_)
);

NOR2X1 _16009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6463_),
    .B(_6464_),
    .Y(_6465_)
);

AOI22X1 _16010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [24]),
    .C(\datapath_1.regfile_1.regOut[22] [24]),
    .D(_5650_),
    .Y(_6466_)
);

AOI22X1 _16011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [24]),
    .C(\datapath_1.regfile_1.regOut[10] [24]),
    .D(_6314_),
    .Y(_6467_)
);

NAND3X1 _16012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6466_),
    .B(_6467_),
    .C(_6465_),
    .Y(_6468_)
);

NAND2X1 _16013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .B(_5490_),
    .Y(_6469_)
);

AOI22X1 _16014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_6470_)
);

INVX1 _16015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [24]),
    .Y(_6471_)
);

OAI22X1 _16016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6471_),
    .B(_5545__bF$buf2),
    .C(_5569_),
    .D(_5119_),
    .Y(_6472_)
);

INVX1 _16017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_6473_)
);

OAI22X1 _16018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6473_),
    .B(_5503__bF$buf3),
    .C(_5504__bF$buf4),
    .D(_5130_),
    .Y(_6474_)
);

NOR2X1 _16019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6472_),
    .B(_6474_),
    .Y(_6475_)
);

NAND3X1 _16020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6469_),
    .B(_6470_),
    .C(_6475_),
    .Y(_6476_)
);

NOR2X1 _16021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6476_),
    .B(_6468_),
    .Y(_6477_)
);

NOR3X1 _16022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf3),
    .B(_5098_),
    .C(_5521__bF$buf3),
    .Y(_6478_)
);

INVX1 _16023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_6479_)
);

OAI22X1 _16024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6479_),
    .B(_5501_),
    .C(_5524__bF$buf2),
    .D(_5127_),
    .Y(_6480_)
);

INVX1 _16025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_6481_)
);

OAI22X1 _16026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_5086_),
    .C(_6481_),
    .D(_5499__bF$buf0),
    .Y(_6482_)
);

NOR2X1 _16027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6482_),
    .B(_6480_),
    .Y(_6483_)
);

INVX1 _16028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_6484_)
);

NAND3X1 _16029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .B(_5471__bF$buf1),
    .C(_5531__bF$buf2),
    .Y(_6485_)
);

OAI21X1 _16030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6484_),
    .B(_5535__bF$buf4),
    .C(_6485_),
    .Y(_6486_)
);

OAI22X1 _16031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf4),
    .B(_5087_),
    .C(_5483__bF$buf2),
    .D(_5122_),
    .Y(_6487_)
);

NOR2X1 _16032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6486_),
    .B(_6487_),
    .Y(_6488_)
);

NAND2X1 _16033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6488_),
    .B(_6483_),
    .Y(_6489_)
);

INVX1 _16034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_6490_)
);

NAND3X1 _16035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .B(_5465_),
    .C(_5531__bF$buf1),
    .Y(_6491_)
);

OAI21X1 _16036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf2),
    .B(_6490_),
    .C(_6491_),
    .Y(_6492_)
);

NAND3X1 _16037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .B(_5477_),
    .C(_5531__bF$buf0),
    .Y(_6493_)
);

OAI21X1 _16038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf2),
    .B(_5111_),
    .C(_6493_),
    .Y(_6494_)
);

NOR2X1 _16039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6492_),
    .B(_6494_),
    .Y(_6495_)
);

INVX1 _16040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_6496_)
);

OAI22X1 _16041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6496_),
    .B(_5548__bF$buf3),
    .C(_5534__bF$buf2),
    .D(_5129_),
    .Y(_6497_)
);

OAI22X1 _16042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf1),
    .B(_5123_),
    .C(_5466__bF$buf2),
    .D(_5120_),
    .Y(_6498_)
);

NOR2X1 _16043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6497_),
    .B(_6498_),
    .Y(_6499_)
);

NAND2X1 _16044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6495_),
    .B(_6499_),
    .Y(_6500_)
);

NOR3X1 _16045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6500_),
    .B(_6478_),
    .C(_6489_),
    .Y(_6501_)
);

AOI21X1 _16046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6477_),
    .B(_6501_),
    .C(RegWrite_bF$buf2),
    .Y(\datapath_1.rd1 [24])
);

NAND2X1 _16047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .B(_5693_),
    .Y(_6502_)
);

NOR2X1 _16048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5157_),
    .B(_5534__bF$buf1),
    .Y(_6503_)
);

INVX1 _16049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_6504_)
);

NOR3X1 _16050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6504_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6505_)
);

INVX1 _16051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_6506_)
);

NOR2X1 _16052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6506_),
    .B(_5549__bF$buf0),
    .Y(_6507_)
);

NOR3X1 _16053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6503_),
    .B(_6505_),
    .C(_6507_),
    .Y(_6508_)
);

INVX1 _16054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_6509_)
);

INVX1 _16055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_6510_)
);

OAI22X1 _16056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf1),
    .B(_6510_),
    .C(_5532__bF$buf0),
    .D(_6509_),
    .Y(_6511_)
);

OAI22X1 _16057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_5161_),
    .C(_5160_),
    .D(_5552__bF$buf1),
    .Y(_6512_)
);

NOR2X1 _16058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6511_),
    .B(_6512_),
    .Y(_6513_)
);

NAND3X1 _16059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6502_),
    .B(_6513_),
    .C(_6508_),
    .Y(_6514_)
);

AOI22X1 _16060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [25]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_6515_)
);

AOI22X1 _16061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf2),
    .B(\datapath_1.regfile_1.regOut[6] [25]),
    .C(\datapath_1.regfile_1.regOut[5] [25]),
    .D(_5700_),
    .Y(_6516_)
);

OAI22X1 _16062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf1),
    .B(_5172_),
    .C(_5151_),
    .D(_5527__bF$buf0),
    .Y(_6517_)
);

INVX1 _16063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_6518_)
);

OAI22X1 _16064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6518_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf2),
    .D(_5150_),
    .Y(_6519_)
);

NOR2X1 _16065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6519_),
    .B(_6517_),
    .Y(_6520_)
);

NAND3X1 _16066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6515_),
    .B(_6516_),
    .C(_6520_),
    .Y(_6521_)
);

NOR2X1 _16067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6521_),
    .B(_6514_),
    .Y(_6522_)
);

NAND2X1 _16068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [25]),
    .B(_5570__bF$buf1),
    .Y(_6523_)
);

OAI22X1 _16069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_5147_),
    .C(_5139_),
    .D(_5483__bF$buf1),
    .Y(_6524_)
);

AOI21X1 _16070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [25]),
    .B(_5567_),
    .C(_6524_),
    .Y(_6525_)
);

INVX1 _16071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [25]),
    .Y(_6526_)
);

INVX1 _16072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [25]),
    .Y(_6527_)
);

OAI22X1 _16073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6526_),
    .B(_5545__bF$buf1),
    .C(_5485__bF$buf3),
    .D(_6527_),
    .Y(_6528_)
);

AOI21X1 _16074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [25]),
    .B(_5481_),
    .C(_6528_),
    .Y(_6529_)
);

NAND3X1 _16075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6523_),
    .B(_6529_),
    .C(_6525_),
    .Y(_6530_)
);

NAND3X1 _16076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6531_)
);

INVX1 _16077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_6532_)
);

OAI22X1 _16078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6532_),
    .B(_5518__bF$buf2),
    .C(_5478__bF$buf0),
    .D(_5136_),
    .Y(_6533_)
);

OAI22X1 _16079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5148_),
    .B(_5548__bF$buf2),
    .C(_5489__bF$buf3),
    .D(_5163_),
    .Y(_6534_)
);

NOR2X1 _16080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6534_),
    .B(_6533_),
    .Y(_6535_)
);

INVX1 _16081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_6536_)
);

OAI22X1 _16082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6536_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf2),
    .D(_5169_),
    .Y(_6537_)
);

OAI22X1 _16083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf3),
    .B(_5168_),
    .C(_5171_),
    .D(_5504__bF$buf3),
    .Y(_6538_)
);

NOR2X1 _16084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6537_),
    .B(_6538_),
    .Y(_6539_)
);

NAND3X1 _16085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6535_),
    .B(_6539_),
    .C(_6531_),
    .Y(_6540_)
);

NOR2X1 _16086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6530_),
    .B(_6540_),
    .Y(_6541_)
);

AOI21X1 _16087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6541_),
    .B(_6522_),
    .C(RegWrite_bF$buf1),
    .Y(\datapath_1.rd1 [25])
);

AOI22X1 _16088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [26]),
    .C(\datapath_1.regfile_1.regOut[22] [26]),
    .D(_5650_),
    .Y(_6542_)
);

NOR2X1 _16089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5205_),
    .B(_5534__bF$buf0),
    .Y(_6543_)
);

NOR2X1 _16090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5181_),
    .B(_5535__bF$buf3),
    .Y(_6544_)
);

INVX1 _16091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_6545_)
);

NOR2X1 _16092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6545_),
    .B(_5549__bF$buf4),
    .Y(_6546_)
);

NOR3X1 _16093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6543_),
    .B(_6544_),
    .C(_6546_),
    .Y(_6547_)
);

AOI22X1 _16094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .B(_5785_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_6548_)
);

NAND3X1 _16095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6542_),
    .B(_6548_),
    .C(_6547_),
    .Y(_6549_)
);

AOI22X1 _16096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_6550_)
);

AOI22X1 _16097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf1),
    .B(\datapath_1.regfile_1.regOut[6] [26]),
    .C(\datapath_1.regfile_1.regOut[5] [26]),
    .D(_5700_),
    .Y(_6551_)
);

OAI22X1 _16098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf0),
    .B(_5206_),
    .C(_5184_),
    .D(_5527__bF$buf4),
    .Y(_6552_)
);

OAI22X1 _16099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5182_),
    .B(_5539__bF$buf0),
    .C(_5469__bF$buf1),
    .D(_5210_),
    .Y(_6553_)
);

NOR2X1 _16100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6553_),
    .B(_6552_),
    .Y(_6554_)
);

NAND3X1 _16101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6550_),
    .B(_6551_),
    .C(_6554_),
    .Y(_6555_)
);

NOR2X1 _16102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6555_),
    .B(_6549_),
    .Y(_6556_)
);

NAND2X1 _16103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .B(_5649_),
    .Y(_6557_)
);

OAI22X1 _16104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_5220_),
    .C(_5218_),
    .D(_5483__bF$buf0),
    .Y(_6558_)
);

AOI21X1 _16105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [26]),
    .B(_5567_),
    .C(_6558_),
    .Y(_6559_)
);

OAI22X1 _16106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_5192_),
    .C(_5189_),
    .D(_5569_),
    .Y(_6560_)
);

INVX1 _16107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [26]),
    .Y(_6561_)
);

INVX1 _16108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [26]),
    .Y(_6562_)
);

OAI22X1 _16109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6561_),
    .B(_5545__bF$buf0),
    .C(_5485__bF$buf2),
    .D(_6562_),
    .Y(_6563_)
);

NOR2X1 _16110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6563_),
    .B(_6560_),
    .Y(_6564_)
);

NAND3X1 _16111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6557_),
    .B(_6564_),
    .C(_6559_),
    .Y(_6565_)
);

NAND3X1 _16112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6566_)
);

OAI22X1 _16113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5221_),
    .B(_5518__bF$buf1),
    .C(_5478__bF$buf3),
    .D(_5213_),
    .Y(_6567_)
);

INVX1 _16114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_6568_)
);

OAI22X1 _16115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6568_),
    .B(_5548__bF$buf1),
    .C(_5489__bF$buf2),
    .D(_5185_),
    .Y(_6569_)
);

NOR2X1 _16116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6569_),
    .B(_6567_),
    .Y(_6570_)
);

OAI22X1 _16117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5193_),
    .B(_5503__bF$buf1),
    .C(_5495__bF$buf1),
    .D(_5190_),
    .Y(_6571_)
);

INVX1 _16118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_6572_)
);

INVX1 _16119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_6573_)
);

OAI22X1 _16120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf2),
    .B(_6573_),
    .C(_6572_),
    .D(_5504__bF$buf2),
    .Y(_6574_)
);

NOR2X1 _16121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6571_),
    .B(_6574_),
    .Y(_6575_)
);

NAND3X1 _16122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6570_),
    .B(_6575_),
    .C(_6566_),
    .Y(_6576_)
);

NOR2X1 _16123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6576_),
    .Y(_6577_)
);

AOI21X1 _16124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6577_),
    .B(_6556_),
    .C(RegWrite_bF$buf0),
    .Y(\datapath_1.rd1 [26])
);

INVX1 _16125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_6578_)
);

OAI22X1 _16126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5252_),
    .B(_5469__bF$buf0),
    .C(_5463__bF$buf1),
    .D(_6578_),
    .Y(_6579_)
);

OAI22X1 _16127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_5254_),
    .C(_5523_),
    .D(_5265_),
    .Y(_6580_)
);

NOR2X1 _16128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6579_),
    .B(_6580_),
    .Y(_6581_)
);

AOI22X1 _16129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [27]),
    .C(\datapath_1.regfile_1.regOut[22] [27]),
    .D(_5650_),
    .Y(_6582_)
);

AOI22X1 _16130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5649_),
    .B(\datapath_1.regfile_1.regOut[23] [27]),
    .C(\datapath_1.regfile_1.regOut[21] [27]),
    .D(_5685_),
    .Y(_6583_)
);

NAND3X1 _16131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582_),
    .B(_6583_),
    .C(_6581_),
    .Y(_6584_)
);

NAND2X1 _16132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [27]),
    .B(_5490_),
    .Y(_6585_)
);

AOI22X1 _16133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .B(_5494_),
    .C(_5496_),
    .D(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_6586_)
);

OAI22X1 _16134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .B(_5235_),
    .C(_5483__bF$buf4),
    .D(_5264_),
    .Y(_6587_)
);

INVX1 _16135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_6588_)
);

INVX1 _16136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_6589_)
);

OAI22X1 _16137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6589_),
    .B(_5503__bF$buf0),
    .C(_5504__bF$buf1),
    .D(_6588_),
    .Y(_6590_)
);

NOR2X1 _16138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6590_),
    .B(_6587_),
    .Y(_6591_)
);

NAND3X1 _16139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6585_),
    .B(_6586_),
    .C(_6591_),
    .Y(_6592_)
);

NOR2X1 _16140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6584_),
    .B(_6592_),
    .Y(_6593_)
);

NOR3X1 _16141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf2),
    .B(_5261_),
    .C(_5521__bF$buf2),
    .Y(_6594_)
);

NAND3X1 _16142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .B(_5500__bF$buf1),
    .C(_5471__bF$buf0),
    .Y(_6595_)
);

OAI21X1 _16143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf1),
    .B(_5228_),
    .C(_6595_),
    .Y(_6596_)
);

INVX1 _16144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [27]),
    .Y(_6597_)
);

INVX1 _16145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_6598_)
);

OAI22X1 _16146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6597_),
    .B(_5544__bF$buf2),
    .C(_5499__bF$buf3),
    .D(_6598_),
    .Y(_6599_)
);

NOR2X1 _16147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6596_),
    .B(_6599_),
    .Y(_6600_)
);

NAND3X1 _16148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .B(_5471__bF$buf5),
    .C(_5531__bF$buf4),
    .Y(_6601_)
);

OAI21X1 _16149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5232_),
    .B(_5535__bF$buf2),
    .C(_6601_),
    .Y(_6602_)
);

INVX1 _16150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [27]),
    .Y(_6603_)
);

OAI22X1 _16151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6603_),
    .B(_5545__bF$buf3),
    .C(_5466__bF$buf4),
    .D(_5262_),
    .Y(_6604_)
);

NOR2X1 _16152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6602_),
    .B(_6604_),
    .Y(_6605_)
);

NAND2X1 _16153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6600_),
    .B(_6605_),
    .Y(_6606_)
);

OAI22X1 _16154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5233_),
    .B(_5539__bF$buf4),
    .C(_5526__bF$buf4),
    .D(_5269_),
    .Y(_6607_)
);

OAI22X1 _16155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527__bF$buf3),
    .B(_5236_),
    .C(_5243_),
    .D(_5532__bF$buf3),
    .Y(_6608_)
);

NOR2X1 _16156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6607_),
    .B(_6608_),
    .Y(_6609_)
);

INVX1 _16157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_6610_)
);

OAI22X1 _16158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6610_),
    .B(_5548__bF$buf0),
    .C(_5534__bF$buf4),
    .D(_5241_),
    .Y(_6611_)
);

INVX1 _16159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [27]),
    .Y(_6612_)
);

OAI22X1 _16160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf1),
    .B(_6612_),
    .C(_5244_),
    .D(_5549__bF$buf3),
    .Y(_6613_)
);

NOR2X1 _16161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6611_),
    .B(_6613_),
    .Y(_6614_)
);

NAND2X1 _16162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6614_),
    .B(_6609_),
    .Y(_6615_)
);

NOR3X1 _16163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6606_),
    .B(_6594_),
    .C(_6615_),
    .Y(_6616_)
);

AOI21X1 _16164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6593_),
    .B(_6616_),
    .C(RegWrite_bF$buf7),
    .Y(\datapath_1.rd1 [27])
);

AOI22X1 _16165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .B(_5606_),
    .C(_5576_),
    .D(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_6617_)
);

AOI22X1 _16166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570__bF$buf0),
    .B(\datapath_1.regfile_1.regOut[27] [28]),
    .C(\datapath_1.regfile_1.regOut[6] [28]),
    .D(_5565__bF$buf0),
    .Y(_6618_)
);

INVX1 _16167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_6619_)
);

OAI22X1 _16168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_6619_),
    .C(_5552__bF$buf0),
    .D(_5312_),
    .Y(_6620_)
);

INVX1 _16169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_6621_)
);

OAI22X1 _16170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530__bF$buf0),
    .B(_6621_),
    .C(_5472__bF$buf0),
    .D(_5297_),
    .Y(_6622_)
);

NOR2X1 _16171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6620_),
    .B(_6622_),
    .Y(_6623_)
);

NAND3X1 _16172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6617_),
    .B(_6618_),
    .C(_6623_),
    .Y(_6624_)
);

INVX1 _16173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_6625_)
);

OAI22X1 _16174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6625_),
    .B(_5518__bF$buf0),
    .C(_5548__bF$buf4),
    .D(_5309_),
    .Y(_6626_)
);

AOI21X1 _16175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [28]),
    .B(_5490_),
    .C(_6626_),
    .Y(_6627_)
);

AOI22X1 _16176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5567_),
    .B(\datapath_1.regfile_1.regOut[28] [28]),
    .C(\datapath_1.regfile_1.regOut[31] [28]),
    .D(_5571_),
    .Y(_6628_)
);

AOI22X1 _16177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .B(_5577_),
    .C(_5971_),
    .D(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_6629_)
);

NAND3X1 _16178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6628_),
    .B(_6629_),
    .C(_6627_),
    .Y(_6630_)
);

NOR2X1 _16179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6630_),
    .B(_6624_),
    .Y(_6631_)
);

NOR3X1 _16180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf1),
    .B(_5300_),
    .C(_5521__bF$buf1),
    .Y(_6632_)
);

OAI22X1 _16181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5310_),
    .B(_5501_),
    .C(_5524__bF$buf0),
    .D(_5292_),
    .Y(_6633_)
);

INVX1 _16182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_6634_)
);

OAI22X1 _16183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_5291_),
    .C(_6634_),
    .D(_5499__bF$buf2),
    .Y(_6635_)
);

NOR2X1 _16184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6635_),
    .B(_6633_),
    .Y(_6636_)
);

NAND3X1 _16185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .B(_5471__bF$buf4),
    .C(_5531__bF$buf3),
    .Y(_6637_)
);

OAI21X1 _16186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5278_),
    .B(_5535__bF$buf1),
    .C(_6637_),
    .Y(_6638_)
);

INVX1 _16187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [28]),
    .Y(_6639_)
);

OAI22X1 _16188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf0),
    .B(_6639_),
    .C(_5483__bF$buf3),
    .D(_5281_),
    .Y(_6640_)
);

NOR2X1 _16189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6638_),
    .B(_6640_),
    .Y(_6641_)
);

NAND2X1 _16190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6641_),
    .B(_6636_),
    .Y(_6642_)
);

NAND3X1 _16191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .B(_5477_),
    .C(_5531__bF$buf2),
    .Y(_6643_)
);

OAI21X1 _16192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf3),
    .B(_5313_),
    .C(_6643_),
    .Y(_6644_)
);

NAND3X1 _16193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [28]),
    .B(_5465_),
    .C(_5531__bF$buf1),
    .Y(_6645_)
);

OAI21X1 _16194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527__bF$buf2),
    .B(_5282_),
    .C(_6645_),
    .Y(_6646_)
);

NOR2X1 _16195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6644_),
    .B(_6646_),
    .Y(_6647_)
);

OAI22X1 _16196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495__bF$buf0),
    .B(_5289_),
    .C(_5288_),
    .D(_5534__bF$buf3),
    .Y(_6648_)
);

INVX1 _16197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [28]),
    .Y(_6649_)
);

INVX1 _16198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_6650_)
);

OAI22X1 _16199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549__bF$buf2),
    .B(_6650_),
    .C(_5466__bF$buf3),
    .D(_6649_),
    .Y(_6651_)
);

NOR2X1 _16200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6648_),
    .B(_6651_),
    .Y(_6652_)
);

NAND2X1 _16201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6647_),
    .B(_6652_),
    .Y(_6653_)
);

NOR3X1 _16202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6653_),
    .B(_6632_),
    .C(_6642_),
    .Y(_6654_)
);

AOI21X1 _16203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6631_),
    .B(_6654_),
    .C(RegWrite_bF$buf6),
    .Y(\datapath_1.rd1 [28])
);

AOI22X1 _16204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .B(_5579_),
    .C(_5649_),
    .D(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_6655_)
);

AOI22X1 _16205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5576_),
    .B(\datapath_1.regfile_1.regOut[13] [29]),
    .C(\datapath_1.regfile_1.regOut[11] [29]),
    .D(_5496_),
    .Y(_6656_)
);

OAI22X1 _16206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5489__bF$buf1),
    .B(_5354_),
    .C(_5527__bF$buf1),
    .D(_5319_),
    .Y(_6657_)
);

INVX1 _16207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_6658_)
);

OAI22X1 _16208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6658_),
    .B(_5469__bF$buf3),
    .C(_5472__bF$buf3),
    .D(_5323_),
    .Y(_6659_)
);

NOR2X1 _16209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6659_),
    .B(_6657_),
    .Y(_6660_)
);

NAND3X1 _16210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6655_),
    .B(_6656_),
    .C(_6660_),
    .Y(_6661_)
);

NAND2X1 _16211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [29]),
    .B(_5479_),
    .Y(_6662_)
);

AOI22X1 _16212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5971_),
    .B(\datapath_1.regfile_1.regOut[14] [29]),
    .C(\datapath_1.regfile_1.regOut[22] [29]),
    .D(_5650_),
    .Y(_6663_)
);

OAI22X1 _16213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5335_),
    .B(_5539__bF$buf3),
    .C(_5503__bF$buf3),
    .D(_5346_),
    .Y(_6664_)
);

AND2X2 _16214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .B(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_6665_)
);

INVX1 _16215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_6666_)
);

NAND2X1 _16216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.PCJump [26]),
    .B(_5470_),
    .Y(_6667_)
);

NOR3X1 _16217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6666_),
    .B(_6667_),
    .C(_5688_),
    .Y(_6668_)
);

NOR3X1 _16218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6664_),
    .B(_6668_),
    .C(_6665_),
    .Y(_6669_)
);

NAND3X1 _16219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6662_),
    .B(_6663_),
    .C(_6669_),
    .Y(_6670_)
);

NOR2X1 _16220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6670_),
    .B(_6661_),
    .Y(_6671_)
);

NOR3X1 _16221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf0),
    .B(_5337_),
    .C(_5521__bF$buf0),
    .Y(_6672_)
);

INVX1 _16222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_6673_)
);

OAI22X1 _16223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf2),
    .B(_5343_),
    .C(_6673_),
    .D(_5549__bF$buf1),
    .Y(_6674_)
);

INVX1 _16224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [29]),
    .Y(_6675_)
);

OAI22X1 _16225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6675_),
    .B(_5545__bF$buf2),
    .C(_5569_),
    .D(_5356_),
    .Y(_6676_)
);

NOR2X1 _16226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6676_),
    .B(_6674_),
    .Y(_6677_)
);

INVX1 _16227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_6678_)
);

OAI22X1 _16228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5325_),
    .B(_5544__bF$buf1),
    .C(_5523_),
    .D(_6678_),
    .Y(_6679_)
);

OAI22X1 _16229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf2),
    .B(_5353_),
    .C(_5331_),
    .D(_5526__bF$buf2),
    .Y(_6680_)
);

NOR2X1 _16230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6679_),
    .B(_6680_),
    .Y(_6681_)
);

NAND2X1 _16231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6677_),
    .B(_6681_),
    .Y(_6682_)
);

NAND3X1 _16232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .B(_5500__bF$buf0),
    .C(_5471__bF$buf3),
    .Y(_6683_)
);

OAI21X1 _16233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf3),
    .B(_5347_),
    .C(_6683_),
    .Y(_6684_)
);

INVX1 _16234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[30] [29]),
    .Y(_6685_)
);

OAI22X1 _16235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_6685_),
    .C(_5326_),
    .D(_5499__bF$buf1),
    .Y(_6686_)
);

NOR2X1 _16236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6684_),
    .B(_6686_),
    .Y(_6687_)
);

NAND3X1 _16237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .B(_5471__bF$buf2),
    .C(_5531__bF$buf0),
    .Y(_6688_)
);

OAI21X1 _16238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5338_),
    .B(_5535__bF$buf0),
    .C(_6688_),
    .Y(_6689_)
);

INVX1 _16239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [29]),
    .Y(_6690_)
);

OAI22X1 _16240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf4),
    .B(_6690_),
    .C(_5483__bF$buf2),
    .D(_5322_),
    .Y(_6691_)
);

NOR2X1 _16241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6689_),
    .B(_6691_),
    .Y(_6692_)
);

NAND2X1 _16242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6687_),
    .B(_6692_),
    .Y(_6693_)
);

NOR3X1 _16243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6693_),
    .B(_6672_),
    .C(_6682_),
    .Y(_6694_)
);

AOI21X1 _16244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6671_),
    .B(_6694_),
    .C(RegWrite_bF$buf5),
    .Y(\datapath_1.rd1 [29])
);

NAND2X1 _16245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[27] [30]),
    .B(_5570__bF$buf3),
    .Y(_6695_)
);

INVX1 _16246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [30]),
    .Y(_6696_)
);

OAI22X1 _16247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5400_),
    .B(_5544__bF$buf0),
    .C(_5485__bF$buf3),
    .D(_6696_),
    .Y(_6697_)
);

OAI22X1 _16248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5365_),
    .B(_5545__bF$buf1),
    .C(_5480__bF$buf3),
    .D(_5364_),
    .Y(_6698_)
);

NOR2X1 _16249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6698_),
    .B(_6697_),
    .Y(_6699_)
);

AOI22X1 _16250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5562_),
    .B(\datapath_1.regfile_1.regOut[25] [30]),
    .C(\datapath_1.regfile_1.regOut[26] [30]),
    .D(_5484_),
    .Y(_6700_)
);

NAND3X1 _16251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6695_),
    .B(_6700_),
    .C(_6699_),
    .Y(_6701_)
);

AOI22X1 _16252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [30]),
    .B(_5697_),
    .C(_5698_),
    .D(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_6702_)
);

AOI22X1 _16253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565__bF$buf3),
    .B(\datapath_1.regfile_1.regOut[6] [30]),
    .C(\datapath_1.regfile_1.regOut[5] [30]),
    .D(_5700_),
    .Y(_6703_)
);

OAI22X1 _16254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5526__bF$buf1),
    .B(_5404_),
    .C(_5385_),
    .D(_5527__bF$buf0),
    .Y(_6704_)
);

INVX1 _16255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_6705_)
);

OAI22X1 _16256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5384_),
    .B(_5539__bF$buf2),
    .C(_5469__bF$buf2),
    .D(_6705_),
    .Y(_6706_)
);

NOR2X1 _16257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6706_),
    .B(_6704_),
    .Y(_6707_)
);

NAND3X1 _16258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6702_),
    .B(_6703_),
    .C(_6707_),
    .Y(_6708_)
);

NOR2X1 _16259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6701_),
    .B(_6708_),
    .Y(_6709_)
);

AOI22X1 _16260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .B(_5693_),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_6710_)
);

OAI22X1 _16261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_5393_),
    .C(_5392_),
    .D(_5552__bF$buf3),
    .Y(_6711_)
);

AOI21X1 _16262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .B(_5649_),
    .C(_6711_),
    .Y(_6712_)
);

NOR3X1 _16263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5403_),
    .B(_5459__bF$buf1),
    .C(_5519_),
    .Y(_6713_)
);

NOR2X1 _16264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5378_),
    .B(_5549__bF$buf0),
    .Y(_6714_)
);

NOR3X1 _16265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5375_),
    .B(_5509_),
    .C(_5688_),
    .Y(_6715_)
);

NOR3X1 _16266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6713_),
    .B(_6715_),
    .C(_6714_),
    .Y(_6716_)
);

NAND3X1 _16267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6710_),
    .B(_6716_),
    .C(_6712_),
    .Y(_6717_)
);

NAND3X1 _16268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .B(_5720_),
    .C(_5721_),
    .Y(_6718_)
);

INVX1 _16269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_6719_)
);

INVX1 _16270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_6720_)
);

OAI22X1 _16271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6720_),
    .B(_5518__bF$buf3),
    .C(_5478__bF$buf1),
    .D(_6719_),
    .Y(_6721_)
);

OAI22X1 _16272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5381_),
    .B(_5548__bF$buf3),
    .C(_5489__bF$buf0),
    .D(_5395_),
    .Y(_6722_)
);

NOR2X1 _16273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6722_),
    .B(_6721_),
    .Y(_6723_)
);

INVX1 _16274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_6724_)
);

INVX1 _16275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_6725_)
);

OAI22X1 _16276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6724_),
    .B(_5503__bF$buf2),
    .C(_5495__bF$buf3),
    .D(_6725_),
    .Y(_6726_)
);

INVX1 _16277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_6727_)
);

INVX1 _16278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_6728_)
);

OAI22X1 _16279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5463__bF$buf0),
    .B(_6728_),
    .C(_6727_),
    .D(_5504__bF$buf0),
    .Y(_6729_)
);

NOR2X1 _16280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6726_),
    .B(_6729_),
    .Y(_6730_)
);

NAND3X1 _16281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6723_),
    .B(_6730_),
    .C(_6718_),
    .Y(_6731_)
);

NOR2X1 _16282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6717_),
    .B(_6731_),
    .Y(_6732_)
);

AOI21X1 _16283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6709_),
    .B(_6732_),
    .C(RegWrite_bF$buf4),
    .Y(\datapath_1.rd1 [30])
);

AOI22X1 _16284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(\datapath_1.regfile_1.regOut[21] [31]),
    .C(\datapath_1.regfile_1.regOut[22] [31]),
    .D(_5650_),
    .Y(_6733_)
);

AOI22X1 _16285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .B(\datapath_1.regfile_1.regOut[7] [31]),
    .C(\datapath_1.regfile_1.regOut[10] [31]),
    .D(_6314_),
    .Y(_6734_)
);

NAND2X1 _16286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6734_),
    .B(_6733_),
    .Y(_6735_)
);

NAND2X1 _16287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .B(_5579_),
    .Y(_6736_)
);

NAND2X1 _16288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [31]),
    .B(_5576_),
    .Y(_6737_)
);

AOI22X1 _16289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .B(\datapath_1.regfile_1.regOut[11] [31]),
    .C(\datapath_1.regfile_1.regOut[14] [31]),
    .D(_5971_),
    .Y(_6738_)
);

NAND3X1 _16290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6736_),
    .B(_6737_),
    .C(_6738_),
    .Y(_6739_)
);

OAI22X1 _16291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5414_),
    .B(_5539__bF$buf1),
    .C(_5469__bF$buf1),
    .D(_5453_),
    .Y(_6740_)
);

AOI21X1 _16292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .B(_5649_),
    .C(_6740_),
    .Y(_6741_)
);

AOI22X1 _16293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(\datapath_1.regfile_1.regOut[2] [31]),
    .C(_5692_),
    .D(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_6742_)
);

AOI22X1 _16294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[31] [31]),
    .B(_5571_),
    .C(_5570__bF$buf2),
    .D(\datapath_1.regfile_1.regOut[27] [31]),
    .Y(_6743_)
);

NAND3X1 _16295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6741_),
    .B(_6743_),
    .C(_6742_),
    .Y(_6744_)
);

NOR3X1 _16296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6739_),
    .B(_6735_),
    .C(_6744_),
    .Y(_6745_)
);

NOR3X1 _16297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515__bF$buf3),
    .B(_5428_),
    .C(_5521__bF$buf3),
    .Y(_6746_)
);

NAND3X1 _16298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .B(_5500__bF$buf3),
    .C(_5471__bF$buf1),
    .Y(_6747_)
);

OAI21X1 _16299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524__bF$buf2),
    .B(_5442_),
    .C(_6747_),
    .Y(_6748_)
);

INVX1 _16300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_6749_)
);

OAI22X1 _16301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_5425_),
    .C(_6749_),
    .D(_5499__bF$buf0),
    .Y(_6750_)
);

NOR2X1 _16302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6748_),
    .B(_6750_),
    .Y(_6751_)
);

NAND3X1 _16303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .B(_5471__bF$buf0),
    .C(_5531__bF$buf4),
    .Y(_6752_)
);

OAI21X1 _16304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5441_),
    .B(_5535__bF$buf4),
    .C(_6752_),
    .Y(_6753_)
);

INVX1 _16305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[29] [31]),
    .Y(_6754_)
);

OAI22X1 _16306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485__bF$buf2),
    .B(_6754_),
    .C(_5483__bF$buf1),
    .D(_5413_),
    .Y(_6755_)
);

NOR2X1 _16307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6753_),
    .B(_6755_),
    .Y(_6756_)
);

NAND2X1 _16308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6751_),
    .B(_6756_),
    .Y(_6757_)
);

OAI22X1 _16309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_5450_),
    .C(_5429_),
    .D(_5526__bF$buf0),
    .Y(_6758_)
);

INVX1 _16310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_6759_)
);

OAI22X1 _16311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5518__bF$buf2),
    .B(_5454_),
    .C(_5503__bF$buf1),
    .D(_6759_),
    .Y(_6760_)
);

NOR2X1 _16312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6760_),
    .B(_6758_),
    .Y(_6761_)
);

INVX1 _16313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_6762_)
);

OAI22X1 _16314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5534__bF$buf1),
    .B(_5434_),
    .C(_6762_),
    .D(_5549__bF$buf4),
    .Y(_6763_)
);

INVX1 _16315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[28] [31]),
    .Y(_6764_)
);

OAI22X1 _16316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6764_),
    .B(_5544__bF$buf3),
    .C(_5523_),
    .D(_5438_),
    .Y(_6765_)
);

NOR2X1 _16317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6763_),
    .B(_6765_),
    .Y(_6766_)
);

NAND2X1 _16318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6766_),
    .B(_6761_),
    .Y(_6767_)
);

NOR3X1 _16319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6757_),
    .B(_6746_),
    .C(_6767_),
    .Y(_6768_)
);

AOI21X1 _16320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6745_),
    .B(_6768_),
    .C(RegWrite_bF$buf3),
    .Y(\datapath_1.rd1 [31])
);

INVX1 _16321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [0]),
    .Y(_6832_)
);

NAND2X1 _16322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6833_)
);

OAI21X1 _16323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6832_),
    .B(gnd),
    .C(_6833_),
    .Y(_6769_[0])
);

INVX1 _16324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [1]),
    .Y(_6770_)
);

NAND2X1 _16325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6771_)
);

OAI21X1 _16326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6770_),
    .B(gnd),
    .C(_6771_),
    .Y(_6769_[1])
);

INVX1 _16327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [2]),
    .Y(_6772_)
);

NAND2X1 _16328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6773_)
);

OAI21X1 _16329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6772_),
    .B(gnd),
    .C(_6773_),
    .Y(_6769_[2])
);

INVX1 _16330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [3]),
    .Y(_6774_)
);

NAND2X1 _16331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6775_)
);

OAI21X1 _16332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6774_),
    .B(gnd),
    .C(_6775_),
    .Y(_6769_[3])
);

INVX1 _16333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [4]),
    .Y(_6776_)
);

NAND2X1 _16334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6777_)
);

OAI21X1 _16335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6776_),
    .B(gnd),
    .C(_6777_),
    .Y(_6769_[4])
);

INVX1 _16336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [5]),
    .Y(_6778_)
);

NAND2X1 _16337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6779_)
);

OAI21X1 _16338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6778_),
    .B(gnd),
    .C(_6779_),
    .Y(_6769_[5])
);

INVX1 _16339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [6]),
    .Y(_6780_)
);

NAND2X1 _16340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6781_)
);

OAI21X1 _16341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6780_),
    .B(gnd),
    .C(_6781_),
    .Y(_6769_[6])
);

INVX1 _16342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [7]),
    .Y(_6782_)
);

NAND2X1 _16343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6783_)
);

OAI21X1 _16344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6782_),
    .B(gnd),
    .C(_6783_),
    .Y(_6769_[7])
);

INVX1 _16345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [8]),
    .Y(_6784_)
);

NAND2X1 _16346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6785_)
);

OAI21X1 _16347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6784_),
    .B(gnd),
    .C(_6785_),
    .Y(_6769_[8])
);

INVX1 _16348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [9]),
    .Y(_6786_)
);

NAND2X1 _16349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6787_)
);

OAI21X1 _16350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6786_),
    .B(gnd),
    .C(_6787_),
    .Y(_6769_[9])
);

INVX1 _16351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [10]),
    .Y(_6788_)
);

NAND2X1 _16352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6789_)
);

OAI21X1 _16353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6788_),
    .B(gnd),
    .C(_6789_),
    .Y(_6769_[10])
);

INVX1 _16354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [11]),
    .Y(_6790_)
);

NAND2X1 _16355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6791_)
);

OAI21X1 _16356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6790_),
    .B(gnd),
    .C(_6791_),
    .Y(_6769_[11])
);

INVX1 _16357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [12]),
    .Y(_6792_)
);

NAND2X1 _16358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6793_)
);

OAI21X1 _16359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6792_),
    .B(gnd),
    .C(_6793_),
    .Y(_6769_[12])
);

INVX1 _16360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [13]),
    .Y(_6794_)
);

NAND2X1 _16361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6795_)
);

OAI21X1 _16362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6794_),
    .B(gnd),
    .C(_6795_),
    .Y(_6769_[13])
);

INVX1 _16363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [14]),
    .Y(_6796_)
);

NAND2X1 _16364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6797_)
);

OAI21X1 _16365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6796_),
    .B(gnd),
    .C(_6797_),
    .Y(_6769_[14])
);

INVX1 _16366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [15]),
    .Y(_6798_)
);

NAND2X1 _16367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6799_)
);

OAI21X1 _16368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6798_),
    .B(gnd),
    .C(_6799_),
    .Y(_6769_[15])
);

INVX1 _16369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [16]),
    .Y(_6800_)
);

NAND2X1 _16370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6801_)
);

OAI21X1 _16371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6800_),
    .B(gnd),
    .C(_6801_),
    .Y(_6769_[16])
);

INVX1 _16372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [17]),
    .Y(_6802_)
);

NAND2X1 _16373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6803_)
);

OAI21X1 _16374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6802_),
    .B(gnd),
    .C(_6803_),
    .Y(_6769_[17])
);

INVX1 _16375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [18]),
    .Y(_6804_)
);

NAND2X1 _16376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6805_)
);

OAI21X1 _16377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6804_),
    .B(gnd),
    .C(_6805_),
    .Y(_6769_[18])
);

INVX1 _16378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [19]),
    .Y(_6806_)
);

NAND2X1 _16379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6807_)
);

OAI21X1 _16380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6806_),
    .B(gnd),
    .C(_6807_),
    .Y(_6769_[19])
);

INVX1 _16381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [20]),
    .Y(_6808_)
);

NAND2X1 _16382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6809_)
);

OAI21X1 _16383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6808_),
    .B(gnd),
    .C(_6809_),
    .Y(_6769_[20])
);

INVX1 _16384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [21]),
    .Y(_6810_)
);

NAND2X1 _16385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6811_)
);

OAI21X1 _16386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6810_),
    .B(gnd),
    .C(_6811_),
    .Y(_6769_[21])
);

INVX1 _16387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [22]),
    .Y(_6812_)
);

NAND2X1 _16388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6813_)
);

OAI21X1 _16389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6812_),
    .B(gnd),
    .C(_6813_),
    .Y(_6769_[22])
);

INVX1 _16390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [23]),
    .Y(_6814_)
);

NAND2X1 _16391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6815_)
);

OAI21X1 _16392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6814_),
    .B(gnd),
    .C(_6815_),
    .Y(_6769_[23])
);

INVX1 _16393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [24]),
    .Y(_6816_)
);

NAND2X1 _16394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6817_)
);

OAI21X1 _16395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6816_),
    .B(gnd),
    .C(_6817_),
    .Y(_6769_[24])
);

INVX1 _16396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [25]),
    .Y(_6818_)
);

NAND2X1 _16397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6819_)
);

OAI21X1 _16398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6818_),
    .B(gnd),
    .C(_6819_),
    .Y(_6769_[25])
);

INVX1 _16399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [26]),
    .Y(_6820_)
);

NAND2X1 _16400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6821_)
);

OAI21X1 _16401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6820_),
    .B(gnd),
    .C(_6821_),
    .Y(_6769_[26])
);

INVX1 _16402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [27]),
    .Y(_6822_)
);

NAND2X1 _16403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6823_)
);

OAI21X1 _16404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6822_),
    .B(gnd),
    .C(_6823_),
    .Y(_6769_[27])
);

INVX1 _16405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [28]),
    .Y(_6824_)
);

NAND2X1 _16406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6825_)
);

OAI21X1 _16407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6824_),
    .B(gnd),
    .C(_6825_),
    .Y(_6769_[28])
);

INVX1 _16408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [29]),
    .Y(_6826_)
);

NAND2X1 _16409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6827_)
);

OAI21X1 _16410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6826_),
    .B(gnd),
    .C(_6827_),
    .Y(_6769_[29])
);

INVX1 _16411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [30]),
    .Y(_6828_)
);

NAND2X1 _16412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6829_)
);

OAI21X1 _16413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6828_),
    .B(gnd),
    .C(_6829_),
    .Y(_6769_[30])
);

INVX1 _16414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[0] [31]),
    .Y(_6830_)
);

NAND2X1 _16415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(gnd),
    .Y(_6831_)
);

OAI21X1 _16416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6830_),
    .B(gnd),
    .C(_6831_),
    .Y(_6769_[31])
);

DFFSR _16417_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_6769_[0]),
    .Q(\datapath_1.regfile_1.regOut[0] [0]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _16418_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_6769_[1]),
    .Q(\datapath_1.regfile_1.regOut[0] [1]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _16419_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_6769_[2]),
    .Q(\datapath_1.regfile_1.regOut[0] [2]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _16420_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_6769_[3]),
    .Q(\datapath_1.regfile_1.regOut[0] [3]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _16421_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_6769_[4]),
    .Q(\datapath_1.regfile_1.regOut[0] [4]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _16422_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_6769_[5]),
    .Q(\datapath_1.regfile_1.regOut[0] [5]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _16423_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_6769_[6]),
    .Q(\datapath_1.regfile_1.regOut[0] [6]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _16424_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_6769_[7]),
    .Q(\datapath_1.regfile_1.regOut[0] [7]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _16425_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_6769_[8]),
    .Q(\datapath_1.regfile_1.regOut[0] [8]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _16426_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_6769_[9]),
    .Q(\datapath_1.regfile_1.regOut[0] [9]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _16427_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_6769_[10]),
    .Q(\datapath_1.regfile_1.regOut[0] [10]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _16428_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_6769_[11]),
    .Q(\datapath_1.regfile_1.regOut[0] [11]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _16429_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_6769_[12]),
    .Q(\datapath_1.regfile_1.regOut[0] [12]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _16430_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_6769_[13]),
    .Q(\datapath_1.regfile_1.regOut[0] [13]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _16431_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_6769_[14]),
    .Q(\datapath_1.regfile_1.regOut[0] [14]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _16432_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_6769_[15]),
    .Q(\datapath_1.regfile_1.regOut[0] [15]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _16433_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_6769_[16]),
    .Q(\datapath_1.regfile_1.regOut[0] [16]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _16434_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_6769_[17]),
    .Q(\datapath_1.regfile_1.regOut[0] [17]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _16435_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_6769_[18]),
    .Q(\datapath_1.regfile_1.regOut[0] [18]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _16436_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_6769_[19]),
    .Q(\datapath_1.regfile_1.regOut[0] [19]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _16437_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_6769_[20]),
    .Q(\datapath_1.regfile_1.regOut[0] [20]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _16438_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_6769_[21]),
    .Q(\datapath_1.regfile_1.regOut[0] [21]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _16439_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_6769_[22]),
    .Q(\datapath_1.regfile_1.regOut[0] [22]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _16440_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_6769_[23]),
    .Q(\datapath_1.regfile_1.regOut[0] [23]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _16441_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_6769_[24]),
    .Q(\datapath_1.regfile_1.regOut[0] [24]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _16442_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_6769_[25]),
    .Q(\datapath_1.regfile_1.regOut[0] [25]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _16443_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_6769_[26]),
    .Q(\datapath_1.regfile_1.regOut[0] [26]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _16444_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_6769_[27]),
    .Q(\datapath_1.regfile_1.regOut[0] [27]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _16445_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_6769_[28]),
    .Q(\datapath_1.regfile_1.regOut[0] [28]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _16446_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_6769_[29]),
    .Q(\datapath_1.regfile_1.regOut[0] [29]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _16447_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_6769_[30]),
    .Q(\datapath_1.regfile_1.regOut[0] [30]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _16448_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_6769_[31]),
    .Q(\datapath_1.regfile_1.regOut[0] [31]),
    .R(rst_bF$buf4),
    .S(vdd)
);

INVX1 _16449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BranchNe),
    .Y(_6834_)
);

AOI21X1 _16450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Branch),
    .B(ALUZero),
    .C(PCWrite),
    .Y(_6835_)
);

OAI21X1 _16451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6834_),
    .B(ALUZero),
    .C(_6835_),
    .Y(PCEn)
);

BUFX2 _6836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(MemRead)
);

BUFX2 _6837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .Y(MemWrite)
);

BUFX2 _6838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[0]),
    .Y(memoryAddress[0])
);

BUFX2 _6839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[1]),
    .Y(memoryAddress[1])
);

BUFX2 _6840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[2]),
    .Y(memoryAddress[2])
);

BUFX2 _6841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[3]),
    .Y(memoryAddress[3])
);

BUFX2 _6842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[4]),
    .Y(memoryAddress[4])
);

BUFX2 _6843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[5]),
    .Y(memoryAddress[5])
);

BUFX2 _6844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[6]),
    .Y(memoryAddress[6])
);

BUFX2 _6845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[7]),
    .Y(memoryAddress[7])
);

BUFX2 _6846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[8]),
    .Y(memoryAddress[8])
);

BUFX2 _6847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[9]),
    .Y(memoryAddress[9])
);

BUFX2 _6848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[10]),
    .Y(memoryAddress[10])
);

BUFX2 _6849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[11]),
    .Y(memoryAddress[11])
);

BUFX2 _6850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[12]),
    .Y(memoryAddress[12])
);

BUFX2 _6851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[13]),
    .Y(memoryAddress[13])
);

BUFX2 _6852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[14]),
    .Y(memoryAddress[14])
);

BUFX2 _6853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[15]),
    .Y(memoryAddress[15])
);

BUFX2 _6854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[16]),
    .Y(memoryAddress[16])
);

BUFX2 _6855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[17]),
    .Y(memoryAddress[17])
);

BUFX2 _6856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[18]),
    .Y(memoryAddress[18])
);

BUFX2 _6857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[19]),
    .Y(memoryAddress[19])
);

BUFX2 _6858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[20]),
    .Y(memoryAddress[20])
);

BUFX2 _6859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[21]),
    .Y(memoryAddress[21])
);

BUFX2 _6860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[22]),
    .Y(memoryAddress[22])
);

BUFX2 _6861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[23]),
    .Y(memoryAddress[23])
);

BUFX2 _6862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[24]),
    .Y(memoryAddress[24])
);

BUFX2 _6863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[25]),
    .Y(memoryAddress[25])
);

BUFX2 _6864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[26]),
    .Y(memoryAddress[26])
);

BUFX2 _6865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[27]),
    .Y(memoryAddress[27])
);

BUFX2 _6866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[28]),
    .Y(memoryAddress[28])
);

BUFX2 _6867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[29]),
    .Y(memoryAddress[29])
);

BUFX2 _6868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[30]),
    .Y(memoryAddress[30])
);

BUFX2 _6869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[31]),
    .Y(memoryAddress[31])
);

BUFX2 _6870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[0]),
    .Y(memoryWriteData[0])
);

BUFX2 _6871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[1]),
    .Y(memoryWriteData[1])
);

BUFX2 _6872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[2]),
    .Y(memoryWriteData[2])
);

BUFX2 _6873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[3]),
    .Y(memoryWriteData[3])
);

BUFX2 _6874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[4]),
    .Y(memoryWriteData[4])
);

BUFX2 _6875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[5]),
    .Y(memoryWriteData[5])
);

BUFX2 _6876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[6]),
    .Y(memoryWriteData[6])
);

BUFX2 _6877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[7]),
    .Y(memoryWriteData[7])
);

BUFX2 _6878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[8]),
    .Y(memoryWriteData[8])
);

BUFX2 _6879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[9]),
    .Y(memoryWriteData[9])
);

BUFX2 _6880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[10]),
    .Y(memoryWriteData[10])
);

BUFX2 _6881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[11]),
    .Y(memoryWriteData[11])
);

BUFX2 _6882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[12]),
    .Y(memoryWriteData[12])
);

BUFX2 _6883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[13]),
    .Y(memoryWriteData[13])
);

BUFX2 _6884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[14]),
    .Y(memoryWriteData[14])
);

BUFX2 _6885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[15]),
    .Y(memoryWriteData[15])
);

BUFX2 _6886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[16]),
    .Y(memoryWriteData[16])
);

BUFX2 _6887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[17]),
    .Y(memoryWriteData[17])
);

BUFX2 _6888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[18]),
    .Y(memoryWriteData[18])
);

BUFX2 _6889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[19]),
    .Y(memoryWriteData[19])
);

BUFX2 _6890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[20]),
    .Y(memoryWriteData[20])
);

BUFX2 _6891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[21]),
    .Y(memoryWriteData[21])
);

BUFX2 _6892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[22]),
    .Y(memoryWriteData[22])
);

BUFX2 _6893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[23]),
    .Y(memoryWriteData[23])
);

BUFX2 _6894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[24]),
    .Y(memoryWriteData[24])
);

BUFX2 _6895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[25]),
    .Y(memoryWriteData[25])
);

BUFX2 _6896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[26]),
    .Y(memoryWriteData[26])
);

BUFX2 _6897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[27]),
    .Y(memoryWriteData[27])
);

BUFX2 _6898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[28]),
    .Y(memoryWriteData[28])
);

BUFX2 _6899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[29]),
    .Y(memoryWriteData[29])
);

BUFX2 _6900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[30]),
    .Y(memoryWriteData[30])
);

BUFX2 _6901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_[31]),
    .Y(memoryWriteData[31])
);

INVX1 _6902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [0]),
    .Y(_66_)
);

NAND2X1 _6903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .Y(_67_)
);

OAI21X1 _6904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_67_),
    .Y(_3_[0])
);

INVX1 _6905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [1]),
    .Y(_4_)
);

NAND2X1 _6906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_5_)
);

OAI21X1 _6907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_5_),
    .Y(_3_[1])
);

INVX1 _6908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [2]),
    .Y(_6_)
);

NAND2X1 _6909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_7_)
);

OAI21X1 _6910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_7_),
    .Y(_3_[2])
);

INVX1 _6911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [3]),
    .Y(_8_)
);

NAND2X1 _6912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_9_)
);

OAI21X1 _6913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_9_),
    .Y(_3_[3])
);

INVX1 _6914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [4]),
    .Y(_10_)
);

NAND2X1 _6915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_11_)
);

OAI21X1 _6916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_11_),
    .Y(_3_[4])
);

INVX1 _6917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [5]),
    .Y(_12_)
);

NAND2X1 _6918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_13_)
);

OAI21X1 _6919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_13_),
    .Y(_3_[5])
);

INVX1 _6920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [6]),
    .Y(_14_)
);

NAND2X1 _6921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_15_)
);

OAI21X1 _6922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_14_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_15_),
    .Y(_3_[6])
);

INVX1 _6923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [7]),
    .Y(_16_)
);

NAND2X1 _6924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_17_)
);

OAI21X1 _6925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_16_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_17_),
    .Y(_3_[7])
);

INVX1 _6926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [8]),
    .Y(_18_)
);

NAND2X1 _6927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_19_)
);

OAI21X1 _6928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_19_),
    .Y(_3_[8])
);

INVX1 _6929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [9]),
    .Y(_20_)
);

NAND2X1 _6930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_21_)
);

OAI21X1 _6931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_20_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_21_),
    .Y(_3_[9])
);

INVX1 _6932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [10]),
    .Y(_22_)
);

NAND2X1 _6933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_23_)
);

OAI21X1 _6934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_22_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_23_),
    .Y(_3_[10])
);

INVX1 _6935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [11]),
    .Y(_24_)
);

NAND2X1 _6936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_25_)
);

OAI21X1 _6937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_25_),
    .Y(_3_[11])
);

INVX1 _6938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [12]),
    .Y(_26_)
);

NAND2X1 _6939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_27_)
);

OAI21X1 _6940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_27_),
    .Y(_3_[12])
);

INVX1 _6941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [13]),
    .Y(_28_)
);

NAND2X1 _6942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_29_)
);

OAI21X1 _6943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_28_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_29_),
    .Y(_3_[13])
);

INVX1 _6944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [14]),
    .Y(_30_)
);

NAND2X1 _6945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_31_)
);

OAI21X1 _6946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_31_),
    .Y(_3_[14])
);

INVX1 _6947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [15]),
    .Y(_32_)
);

NAND2X1 _6948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_33_)
);

OAI21X1 _6949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_33_),
    .Y(_3_[15])
);

INVX1 _6950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [16]),
    .Y(_34_)
);

NAND2X1 _6951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_35_)
);

OAI21X1 _6952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_35_),
    .Y(_3_[16])
);

INVX1 _6953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [17]),
    .Y(_36_)
);

NAND2X1 _6954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_37_)
);

OAI21X1 _6955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_37_),
    .Y(_3_[17])
);

INVX1 _6956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [18]),
    .Y(_38_)
);

NAND2X1 _6957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_39_)
);

OAI21X1 _6958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_39_),
    .Y(_3_[18])
);

INVX1 _6959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [19]),
    .Y(_40_)
);

NAND2X1 _6960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_41_)
);

OAI21X1 _6961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_41_),
    .Y(_3_[19])
);

INVX1 _6962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [20]),
    .Y(_42_)
);

NAND2X1 _6963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_43_)
);

OAI21X1 _6964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_43_),
    .Y(_3_[20])
);

INVX1 _6965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [21]),
    .Y(_44_)
);

NAND2X1 _6966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_45_)
);

OAI21X1 _6967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_45_),
    .Y(_3_[21])
);

INVX1 _6968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [22]),
    .Y(_46_)
);

NAND2X1 _6969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_47_)
);

OAI21X1 _6970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_46_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_47_),
    .Y(_3_[22])
);

INVX1 _6971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [23]),
    .Y(_48_)
);

NAND2X1 _6972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_49_)
);

OAI21X1 _6973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_48_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_49_),
    .Y(_3_[23])
);

INVX1 _6974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [24]),
    .Y(_50_)
);

NAND2X1 _6975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_51_)
);

OAI21X1 _6976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_51_),
    .Y(_3_[24])
);

INVX1 _6977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [25]),
    .Y(_52_)
);

NAND2X1 _6978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_53_)
);

OAI21X1 _6979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_52_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_53_),
    .Y(_3_[25])
);

INVX1 _6980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [26]),
    .Y(_54_)
);

NAND2X1 _6981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_55_)
);

OAI21X1 _6982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_55_),
    .Y(_3_[26])
);

INVX1 _6983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [27]),
    .Y(_56_)
);

NAND2X1 _6984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_57_)
);

OAI21X1 _6985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_57_),
    .Y(_3_[27])
);

INVX1 _6986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [28]),
    .Y(_58_)
);

NAND2X1 _6987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_59_)
);

OAI21X1 _6988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf6 ),
    .C(_59_),
    .Y(_3_[28])
);

INVX1 _6989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [29]),
    .Y(_60_)
);

NAND2X1 _6990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_61_)
);

OAI21X1 _6991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf4 ),
    .C(_61_),
    .Y(_3_[29])
);

INVX1 _6992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [30]),
    .Y(_62_)
);

NAND2X1 _6993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_63_)
);

OAI21X1 _6994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf2 ),
    .C(_63_),
    .Y(_3_[30])
);

INVX1 _6995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[1] [31]),
    .Y(_64_)
);

NAND2X1 _6996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_1_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_65_)
);

OAI21X1 _6997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_64_),
    .B(\datapath_1.regfile_1.regEn_1_bF$buf0 ),
    .C(_65_),
    .Y(_3_[31])
);

DFFSR _6998_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_3_[0]),
    .Q(\datapath_1.regfile_1.regOut[1] [0]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _6999_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_3_[1]),
    .Q(\datapath_1.regfile_1.regOut[1] [1]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _7000_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_3_[2]),
    .Q(\datapath_1.regfile_1.regOut[1] [2]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _7001_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_3_[3]),
    .Q(\datapath_1.regfile_1.regOut[1] [3]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _7002_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_3_[4]),
    .Q(\datapath_1.regfile_1.regOut[1] [4]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _7003_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_3_[5]),
    .Q(\datapath_1.regfile_1.regOut[1] [5]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _7004_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_3_[6]),
    .Q(\datapath_1.regfile_1.regOut[1] [6]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _7005_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_3_[7]),
    .Q(\datapath_1.regfile_1.regOut[1] [7]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _7006_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_3_[8]),
    .Q(\datapath_1.regfile_1.regOut[1] [8]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _7007_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_3_[9]),
    .Q(\datapath_1.regfile_1.regOut[1] [9]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _7008_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_3_[10]),
    .Q(\datapath_1.regfile_1.regOut[1] [10]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _7009_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_3_[11]),
    .Q(\datapath_1.regfile_1.regOut[1] [11]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _7010_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_3_[12]),
    .Q(\datapath_1.regfile_1.regOut[1] [12]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _7011_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_3_[13]),
    .Q(\datapath_1.regfile_1.regOut[1] [13]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _7012_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_3_[14]),
    .Q(\datapath_1.regfile_1.regOut[1] [14]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _7013_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_3_[15]),
    .Q(\datapath_1.regfile_1.regOut[1] [15]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _7014_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_3_[16]),
    .Q(\datapath_1.regfile_1.regOut[1] [16]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _7015_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_3_[17]),
    .Q(\datapath_1.regfile_1.regOut[1] [17]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _7016_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_3_[18]),
    .Q(\datapath_1.regfile_1.regOut[1] [18]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _7017_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_3_[19]),
    .Q(\datapath_1.regfile_1.regOut[1] [19]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _7018_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_3_[20]),
    .Q(\datapath_1.regfile_1.regOut[1] [20]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _7019_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_3_[21]),
    .Q(\datapath_1.regfile_1.regOut[1] [21]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _7020_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_3_[22]),
    .Q(\datapath_1.regfile_1.regOut[1] [22]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _7021_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_3_[23]),
    .Q(\datapath_1.regfile_1.regOut[1] [23]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _7022_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_3_[24]),
    .Q(\datapath_1.regfile_1.regOut[1] [24]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _7023_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_3_[25]),
    .Q(\datapath_1.regfile_1.regOut[1] [25]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _7024_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_3_[26]),
    .Q(\datapath_1.regfile_1.regOut[1] [26]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _7025_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_3_[27]),
    .Q(\datapath_1.regfile_1.regOut[1] [27]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _7026_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_3_[28]),
    .Q(\datapath_1.regfile_1.regOut[1] [28]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _7027_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_3_[29]),
    .Q(\datapath_1.regfile_1.regOut[1] [29]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _7028_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_3_[30]),
    .Q(\datapath_1.regfile_1.regOut[1] [30]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _7029_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_3_[31]),
    .Q(\datapath_1.regfile_1.regOut[1] [31]),
    .R(rst_bF$buf86),
    .S(vdd)
);

INVX1 _7030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [0]),
    .Y(_131_)
);

NAND2X1 _7031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .Y(_132_)
);

OAI21X1 _7032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_131_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_132_),
    .Y(_68_[0])
);

INVX1 _7033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [1]),
    .Y(_69_)
);

NAND2X1 _7034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_70_)
);

OAI21X1 _7035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_70_),
    .Y(_68_[1])
);

INVX1 _7036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [2]),
    .Y(_71_)
);

NAND2X1 _7037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_72_)
);

OAI21X1 _7038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_72_),
    .Y(_68_[2])
);

INVX1 _7039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [3]),
    .Y(_73_)
);

NAND2X1 _7040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_74_)
);

OAI21X1 _7041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_74_),
    .Y(_68_[3])
);

INVX1 _7042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [4]),
    .Y(_75_)
);

NAND2X1 _7043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_76_)
);

OAI21X1 _7044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_76_),
    .Y(_68_[4])
);

INVX1 _7045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [5]),
    .Y(_77_)
);

NAND2X1 _7046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_78_)
);

OAI21X1 _7047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_78_),
    .Y(_68_[5])
);

INVX1 _7048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [6]),
    .Y(_79_)
);

NAND2X1 _7049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_80_)
);

OAI21X1 _7050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_80_),
    .Y(_68_[6])
);

INVX1 _7051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [7]),
    .Y(_81_)
);

NAND2X1 _7052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_82_)
);

OAI21X1 _7053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_82_),
    .Y(_68_[7])
);

INVX1 _7054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [8]),
    .Y(_83_)
);

NAND2X1 _7055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_84_)
);

OAI21X1 _7056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_84_),
    .Y(_68_[8])
);

INVX1 _7057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [9]),
    .Y(_85_)
);

NAND2X1 _7058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_86_)
);

OAI21X1 _7059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_86_),
    .Y(_68_[9])
);

INVX1 _7060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [10]),
    .Y(_87_)
);

NAND2X1 _7061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_88_)
);

OAI21X1 _7062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_88_),
    .Y(_68_[10])
);

INVX1 _7063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [11]),
    .Y(_89_)
);

NAND2X1 _7064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_90_)
);

OAI21X1 _7065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_90_),
    .Y(_68_[11])
);

INVX1 _7066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [12]),
    .Y(_91_)
);

NAND2X1 _7067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_92_)
);

OAI21X1 _7068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_92_),
    .Y(_68_[12])
);

INVX1 _7069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [13]),
    .Y(_93_)
);

NAND2X1 _7070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_94_)
);

OAI21X1 _7071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_94_),
    .Y(_68_[13])
);

INVX1 _7072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [14]),
    .Y(_95_)
);

NAND2X1 _7073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_96_)
);

OAI21X1 _7074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_96_),
    .Y(_68_[14])
);

INVX1 _7075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [15]),
    .Y(_97_)
);

NAND2X1 _7076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_98_)
);

OAI21X1 _7077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_98_),
    .Y(_68_[15])
);

INVX1 _7078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [16]),
    .Y(_99_)
);

NAND2X1 _7079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_100_)
);

OAI21X1 _7080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_100_),
    .Y(_68_[16])
);

INVX1 _7081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [17]),
    .Y(_101_)
);

NAND2X1 _7082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_102_)
);

OAI21X1 _7083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_102_),
    .Y(_68_[17])
);

INVX1 _7084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [18]),
    .Y(_103_)
);

NAND2X1 _7085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_104_)
);

OAI21X1 _7086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_104_),
    .Y(_68_[18])
);

INVX1 _7087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [19]),
    .Y(_105_)
);

NAND2X1 _7088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_106_)
);

OAI21X1 _7089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_106_),
    .Y(_68_[19])
);

INVX1 _7090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [20]),
    .Y(_107_)
);

NAND2X1 _7091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_108_)
);

OAI21X1 _7092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_108_),
    .Y(_68_[20])
);

INVX1 _7093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [21]),
    .Y(_109_)
);

NAND2X1 _7094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_110_)
);

OAI21X1 _7095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_110_),
    .Y(_68_[21])
);

INVX1 _7096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [22]),
    .Y(_111_)
);

NAND2X1 _7097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_112_)
);

OAI21X1 _7098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_112_),
    .Y(_68_[22])
);

INVX1 _7099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [23]),
    .Y(_113_)
);

NAND2X1 _7100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_114_)
);

OAI21X1 _7101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_114_),
    .Y(_68_[23])
);

INVX1 _7102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [24]),
    .Y(_115_)
);

NAND2X1 _7103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_116_)
);

OAI21X1 _7104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_116_),
    .Y(_68_[24])
);

INVX1 _7105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [25]),
    .Y(_117_)
);

NAND2X1 _7106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_118_)
);

OAI21X1 _7107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_118_),
    .Y(_68_[25])
);

INVX1 _7108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [26]),
    .Y(_119_)
);

NAND2X1 _7109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_120_)
);

OAI21X1 _7110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_120_),
    .Y(_68_[26])
);

INVX1 _7111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [27]),
    .Y(_121_)
);

NAND2X1 _7112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_122_)
);

OAI21X1 _7113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_122_),
    .Y(_68_[27])
);

INVX1 _7114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [28]),
    .Y(_123_)
);

NAND2X1 _7115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_124_)
);

OAI21X1 _7116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf6 ),
    .C(_124_),
    .Y(_68_[28])
);

INVX1 _7117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [29]),
    .Y(_125_)
);

NAND2X1 _7118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_126_)
);

OAI21X1 _7119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf4 ),
    .C(_126_),
    .Y(_68_[29])
);

INVX1 _7120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [30]),
    .Y(_127_)
);

NAND2X1 _7121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_128_)
);

OAI21X1 _7122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf2 ),
    .C(_128_),
    .Y(_68_[30])
);

INVX1 _7123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[2] [31]),
    .Y(_129_)
);

NAND2X1 _7124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_2_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_130_)
);

OAI21X1 _7125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(\datapath_1.regfile_1.regEn_2_bF$buf0 ),
    .C(_130_),
    .Y(_68_[31])
);

DFFSR _7126_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_68_[0]),
    .Q(\datapath_1.regfile_1.regOut[2] [0]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _7127_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_68_[1]),
    .Q(\datapath_1.regfile_1.regOut[2] [1]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _7128_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_68_[2]),
    .Q(\datapath_1.regfile_1.regOut[2] [2]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _7129_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_68_[3]),
    .Q(\datapath_1.regfile_1.regOut[2] [3]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _7130_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_68_[4]),
    .Q(\datapath_1.regfile_1.regOut[2] [4]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _7131_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_68_[5]),
    .Q(\datapath_1.regfile_1.regOut[2] [5]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _7132_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_68_[6]),
    .Q(\datapath_1.regfile_1.regOut[2] [6]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _7133_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_68_[7]),
    .Q(\datapath_1.regfile_1.regOut[2] [7]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _7134_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_68_[8]),
    .Q(\datapath_1.regfile_1.regOut[2] [8]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _7135_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_68_[9]),
    .Q(\datapath_1.regfile_1.regOut[2] [9]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _7136_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_68_[10]),
    .Q(\datapath_1.regfile_1.regOut[2] [10]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _7137_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_68_[11]),
    .Q(\datapath_1.regfile_1.regOut[2] [11]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _7138_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_68_[12]),
    .Q(\datapath_1.regfile_1.regOut[2] [12]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _7139_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_68_[13]),
    .Q(\datapath_1.regfile_1.regOut[2] [13]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _7140_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_68_[14]),
    .Q(\datapath_1.regfile_1.regOut[2] [14]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _7141_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_68_[15]),
    .Q(\datapath_1.regfile_1.regOut[2] [15]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _7142_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_68_[16]),
    .Q(\datapath_1.regfile_1.regOut[2] [16]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _7143_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_68_[17]),
    .Q(\datapath_1.regfile_1.regOut[2] [17]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _7144_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_68_[18]),
    .Q(\datapath_1.regfile_1.regOut[2] [18]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _7145_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_68_[19]),
    .Q(\datapath_1.regfile_1.regOut[2] [19]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _7146_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_68_[20]),
    .Q(\datapath_1.regfile_1.regOut[2] [20]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _7147_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_68_[21]),
    .Q(\datapath_1.regfile_1.regOut[2] [21]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _7148_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_68_[22]),
    .Q(\datapath_1.regfile_1.regOut[2] [22]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _7149_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_68_[23]),
    .Q(\datapath_1.regfile_1.regOut[2] [23]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _7150_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_68_[24]),
    .Q(\datapath_1.regfile_1.regOut[2] [24]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _7151_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_68_[25]),
    .Q(\datapath_1.regfile_1.regOut[2] [25]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _7152_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_68_[26]),
    .Q(\datapath_1.regfile_1.regOut[2] [26]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _7153_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_68_[27]),
    .Q(\datapath_1.regfile_1.regOut[2] [27]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _7154_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_68_[28]),
    .Q(\datapath_1.regfile_1.regOut[2] [28]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _7155_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_68_[29]),
    .Q(\datapath_1.regfile_1.regOut[2] [29]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _7156_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_68_[30]),
    .Q(\datapath_1.regfile_1.regOut[2] [30]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _7157_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_68_[31]),
    .Q(\datapath_1.regfile_1.regOut[2] [31]),
    .R(rst_bF$buf54),
    .S(vdd)
);

INVX1 _7158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [0]),
    .Y(_196_)
);

NAND2X1 _7159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .Y(_197_)
);

OAI21X1 _7160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_197_),
    .Y(_133_[0])
);

INVX1 _7161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [1]),
    .Y(_134_)
);

NAND2X1 _7162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_135_)
);

OAI21X1 _7163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_135_),
    .Y(_133_[1])
);

INVX1 _7164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [2]),
    .Y(_136_)
);

NAND2X1 _7165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_137_)
);

OAI21X1 _7166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_137_),
    .Y(_133_[2])
);

INVX1 _7167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [3]),
    .Y(_138_)
);

NAND2X1 _7168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_139_)
);

OAI21X1 _7169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_139_),
    .Y(_133_[3])
);

INVX1 _7170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [4]),
    .Y(_140_)
);

NAND2X1 _7171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_141_)
);

OAI21X1 _7172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_141_),
    .Y(_133_[4])
);

INVX1 _7173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [5]),
    .Y(_142_)
);

NAND2X1 _7174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_143_)
);

OAI21X1 _7175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_143_),
    .Y(_133_[5])
);

INVX1 _7176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [6]),
    .Y(_144_)
);

NAND2X1 _7177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_145_)
);

OAI21X1 _7178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_145_),
    .Y(_133_[6])
);

INVX1 _7179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [7]),
    .Y(_146_)
);

NAND2X1 _7180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_147_)
);

OAI21X1 _7181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_147_),
    .Y(_133_[7])
);

INVX1 _7182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [8]),
    .Y(_148_)
);

NAND2X1 _7183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_149_)
);

OAI21X1 _7184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_149_),
    .Y(_133_[8])
);

INVX1 _7185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [9]),
    .Y(_150_)
);

NAND2X1 _7186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_151_)
);

OAI21X1 _7187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_151_),
    .Y(_133_[9])
);

INVX1 _7188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [10]),
    .Y(_152_)
);

NAND2X1 _7189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_153_)
);

OAI21X1 _7190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_153_),
    .Y(_133_[10])
);

INVX1 _7191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [11]),
    .Y(_154_)
);

NAND2X1 _7192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_155_)
);

OAI21X1 _7193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_155_),
    .Y(_133_[11])
);

INVX1 _7194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [12]),
    .Y(_156_)
);

NAND2X1 _7195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_157_)
);

OAI21X1 _7196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_157_),
    .Y(_133_[12])
);

INVX1 _7197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [13]),
    .Y(_158_)
);

NAND2X1 _7198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_159_)
);

OAI21X1 _7199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_159_),
    .Y(_133_[13])
);

INVX1 _7200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [14]),
    .Y(_160_)
);

NAND2X1 _7201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_161_)
);

OAI21X1 _7202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_161_),
    .Y(_133_[14])
);

INVX1 _7203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [15]),
    .Y(_162_)
);

NAND2X1 _7204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_163_)
);

OAI21X1 _7205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_163_),
    .Y(_133_[15])
);

INVX1 _7206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [16]),
    .Y(_164_)
);

NAND2X1 _7207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_165_)
);

OAI21X1 _7208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_165_),
    .Y(_133_[16])
);

INVX1 _7209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [17]),
    .Y(_166_)
);

NAND2X1 _7210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_167_)
);

OAI21X1 _7211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_167_),
    .Y(_133_[17])
);

INVX1 _7212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [18]),
    .Y(_168_)
);

NAND2X1 _7213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_169_)
);

OAI21X1 _7214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_169_),
    .Y(_133_[18])
);

INVX1 _7215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [19]),
    .Y(_170_)
);

NAND2X1 _7216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_171_)
);

OAI21X1 _7217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_171_),
    .Y(_133_[19])
);

INVX1 _7218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [20]),
    .Y(_172_)
);

NAND2X1 _7219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_173_)
);

OAI21X1 _7220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_173_),
    .Y(_133_[20])
);

INVX1 _7221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [21]),
    .Y(_174_)
);

NAND2X1 _7222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_175_)
);

OAI21X1 _7223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_174_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_175_),
    .Y(_133_[21])
);

INVX1 _7224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [22]),
    .Y(_176_)
);

NAND2X1 _7225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_177_)
);

OAI21X1 _7226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_177_),
    .Y(_133_[22])
);

INVX1 _7227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [23]),
    .Y(_178_)
);

NAND2X1 _7228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_179_)
);

OAI21X1 _7229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_179_),
    .Y(_133_[23])
);

INVX1 _7230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [24]),
    .Y(_180_)
);

NAND2X1 _7231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_181_)
);

OAI21X1 _7232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_181_),
    .Y(_133_[24])
);

INVX1 _7233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [25]),
    .Y(_182_)
);

NAND2X1 _7234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_183_)
);

OAI21X1 _7235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_183_),
    .Y(_133_[25])
);

INVX1 _7236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [26]),
    .Y(_184_)
);

NAND2X1 _7237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_185_)
);

OAI21X1 _7238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_185_),
    .Y(_133_[26])
);

INVX1 _7239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [27]),
    .Y(_186_)
);

NAND2X1 _7240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_187_)
);

OAI21X1 _7241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_187_),
    .Y(_133_[27])
);

INVX1 _7242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [28]),
    .Y(_188_)
);

NAND2X1 _7243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_189_)
);

OAI21X1 _7244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf6 ),
    .C(_189_),
    .Y(_133_[28])
);

INVX1 _7245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [29]),
    .Y(_190_)
);

NAND2X1 _7246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_191_)
);

OAI21X1 _7247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf4 ),
    .C(_191_),
    .Y(_133_[29])
);

INVX1 _7248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [30]),
    .Y(_192_)
);

NAND2X1 _7249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_193_)
);

OAI21X1 _7250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf2 ),
    .C(_193_),
    .Y(_133_[30])
);

INVX1 _7251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[3] [31]),
    .Y(_194_)
);

NAND2X1 _7252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_3_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_195_)
);

OAI21X1 _7253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(\datapath_1.regfile_1.regEn_3_bF$buf0 ),
    .C(_195_),
    .Y(_133_[31])
);

DFFSR _7254_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_133_[0]),
    .Q(\datapath_1.regfile_1.regOut[3] [0]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _7255_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_133_[1]),
    .Q(\datapath_1.regfile_1.regOut[3] [1]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _7256_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_133_[2]),
    .Q(\datapath_1.regfile_1.regOut[3] [2]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _7257_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_133_[3]),
    .Q(\datapath_1.regfile_1.regOut[3] [3]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _7258_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_133_[4]),
    .Q(\datapath_1.regfile_1.regOut[3] [4]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _7259_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_133_[5]),
    .Q(\datapath_1.regfile_1.regOut[3] [5]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _7260_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_133_[6]),
    .Q(\datapath_1.regfile_1.regOut[3] [6]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _7261_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_133_[7]),
    .Q(\datapath_1.regfile_1.regOut[3] [7]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _7262_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_133_[8]),
    .Q(\datapath_1.regfile_1.regOut[3] [8]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _7263_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_133_[9]),
    .Q(\datapath_1.regfile_1.regOut[3] [9]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _7264_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_133_[10]),
    .Q(\datapath_1.regfile_1.regOut[3] [10]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _7265_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_133_[11]),
    .Q(\datapath_1.regfile_1.regOut[3] [11]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _7266_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_133_[12]),
    .Q(\datapath_1.regfile_1.regOut[3] [12]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _7267_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_133_[13]),
    .Q(\datapath_1.regfile_1.regOut[3] [13]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _7268_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_133_[14]),
    .Q(\datapath_1.regfile_1.regOut[3] [14]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _7269_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_133_[15]),
    .Q(\datapath_1.regfile_1.regOut[3] [15]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _7270_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_133_[16]),
    .Q(\datapath_1.regfile_1.regOut[3] [16]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _7271_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_133_[17]),
    .Q(\datapath_1.regfile_1.regOut[3] [17]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _7272_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_133_[18]),
    .Q(\datapath_1.regfile_1.regOut[3] [18]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _7273_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_133_[19]),
    .Q(\datapath_1.regfile_1.regOut[3] [19]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _7274_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_133_[20]),
    .Q(\datapath_1.regfile_1.regOut[3] [20]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _7275_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_133_[21]),
    .Q(\datapath_1.regfile_1.regOut[3] [21]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _7276_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_133_[22]),
    .Q(\datapath_1.regfile_1.regOut[3] [22]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _7277_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_133_[23]),
    .Q(\datapath_1.regfile_1.regOut[3] [23]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _7278_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_133_[24]),
    .Q(\datapath_1.regfile_1.regOut[3] [24]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _7279_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_133_[25]),
    .Q(\datapath_1.regfile_1.regOut[3] [25]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _7280_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_133_[26]),
    .Q(\datapath_1.regfile_1.regOut[3] [26]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _7281_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_133_[27]),
    .Q(\datapath_1.regfile_1.regOut[3] [27]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _7282_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_133_[28]),
    .Q(\datapath_1.regfile_1.regOut[3] [28]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _7283_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_133_[29]),
    .Q(\datapath_1.regfile_1.regOut[3] [29]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _7284_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_133_[30]),
    .Q(\datapath_1.regfile_1.regOut[3] [30]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _7285_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_133_[31]),
    .Q(\datapath_1.regfile_1.regOut[3] [31]),
    .R(rst_bF$buf22),
    .S(vdd)
);

INVX1 _7286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [0]),
    .Y(_261_)
);

NAND2X1 _7287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .Y(_262_)
);

OAI21X1 _7288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_262_),
    .Y(_198_[0])
);

INVX1 _7289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [1]),
    .Y(_199_)
);

NAND2X1 _7290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_200_)
);

OAI21X1 _7291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_200_),
    .Y(_198_[1])
);

INVX1 _7292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [2]),
    .Y(_201_)
);

NAND2X1 _7293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_202_)
);

OAI21X1 _7294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_201_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_202_),
    .Y(_198_[2])
);

INVX1 _7295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [3]),
    .Y(_203_)
);

NAND2X1 _7296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_204_)
);

OAI21X1 _7297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_204_),
    .Y(_198_[3])
);

INVX1 _7298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [4]),
    .Y(_205_)
);

NAND2X1 _7299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_206_)
);

OAI21X1 _7300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_206_),
    .Y(_198_[4])
);

INVX1 _7301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [5]),
    .Y(_207_)
);

NAND2X1 _7302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_208_)
);

OAI21X1 _7303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_208_),
    .Y(_198_[5])
);

INVX1 _7304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [6]),
    .Y(_209_)
);

NAND2X1 _7305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_210_)
);

OAI21X1 _7306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_210_),
    .Y(_198_[6])
);

INVX1 _7307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [7]),
    .Y(_211_)
);

NAND2X1 _7308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_212_)
);

OAI21X1 _7309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_212_),
    .Y(_198_[7])
);

INVX1 _7310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [8]),
    .Y(_213_)
);

NAND2X1 _7311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_214_)
);

OAI21X1 _7312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_214_),
    .Y(_198_[8])
);

INVX1 _7313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [9]),
    .Y(_215_)
);

NAND2X1 _7314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_216_)
);

OAI21X1 _7315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_216_),
    .Y(_198_[9])
);

INVX1 _7316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [10]),
    .Y(_217_)
);

NAND2X1 _7317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_218_)
);

OAI21X1 _7318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_218_),
    .Y(_198_[10])
);

INVX1 _7319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [11]),
    .Y(_219_)
);

NAND2X1 _7320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_220_)
);

OAI21X1 _7321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_220_),
    .Y(_198_[11])
);

INVX1 _7322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [12]),
    .Y(_221_)
);

NAND2X1 _7323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_222_)
);

OAI21X1 _7324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_222_),
    .Y(_198_[12])
);

INVX1 _7325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [13]),
    .Y(_223_)
);

NAND2X1 _7326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_224_)
);

OAI21X1 _7327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_224_),
    .Y(_198_[13])
);

INVX1 _7328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [14]),
    .Y(_225_)
);

NAND2X1 _7329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_226_)
);

OAI21X1 _7330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_226_),
    .Y(_198_[14])
);

INVX1 _7331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [15]),
    .Y(_227_)
);

NAND2X1 _7332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_228_)
);

OAI21X1 _7333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_228_),
    .Y(_198_[15])
);

INVX1 _7334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [16]),
    .Y(_229_)
);

NAND2X1 _7335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_230_)
);

OAI21X1 _7336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_230_),
    .Y(_198_[16])
);

INVX1 _7337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [17]),
    .Y(_231_)
);

NAND2X1 _7338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_232_)
);

OAI21X1 _7339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_232_),
    .Y(_198_[17])
);

INVX1 _7340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [18]),
    .Y(_233_)
);

NAND2X1 _7341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_234_)
);

OAI21X1 _7342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_234_),
    .Y(_198_[18])
);

INVX1 _7343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [19]),
    .Y(_235_)
);

NAND2X1 _7344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_236_)
);

OAI21X1 _7345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_236_),
    .Y(_198_[19])
);

INVX1 _7346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [20]),
    .Y(_237_)
);

NAND2X1 _7347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_238_)
);

OAI21X1 _7348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_238_),
    .Y(_198_[20])
);

INVX1 _7349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [21]),
    .Y(_239_)
);

NAND2X1 _7350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_240_)
);

OAI21X1 _7351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_240_),
    .Y(_198_[21])
);

INVX1 _7352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [22]),
    .Y(_241_)
);

NAND2X1 _7353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_242_)
);

OAI21X1 _7354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_242_),
    .Y(_198_[22])
);

INVX1 _7355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [23]),
    .Y(_243_)
);

NAND2X1 _7356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_244_)
);

OAI21X1 _7357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_244_),
    .Y(_198_[23])
);

INVX1 _7358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [24]),
    .Y(_245_)
);

NAND2X1 _7359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_246_)
);

OAI21X1 _7360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_246_),
    .Y(_198_[24])
);

INVX1 _7361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [25]),
    .Y(_247_)
);

NAND2X1 _7362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_248_)
);

OAI21X1 _7363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_248_),
    .Y(_198_[25])
);

INVX1 _7364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [26]),
    .Y(_249_)
);

NAND2X1 _7365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_250_)
);

OAI21X1 _7366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_250_),
    .Y(_198_[26])
);

INVX1 _7367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [27]),
    .Y(_251_)
);

NAND2X1 _7368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_252_)
);

OAI21X1 _7369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_252_),
    .Y(_198_[27])
);

INVX1 _7370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [28]),
    .Y(_253_)
);

NAND2X1 _7371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_254_)
);

OAI21X1 _7372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_253_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf6 ),
    .C(_254_),
    .Y(_198_[28])
);

INVX1 _7373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [29]),
    .Y(_255_)
);

NAND2X1 _7374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_256_)
);

OAI21X1 _7375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf4 ),
    .C(_256_),
    .Y(_198_[29])
);

INVX1 _7376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [30]),
    .Y(_257_)
);

NAND2X1 _7377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_258_)
);

OAI21X1 _7378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf2 ),
    .C(_258_),
    .Y(_198_[30])
);

INVX1 _7379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[4] [31]),
    .Y(_259_)
);

NAND2X1 _7380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_4_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_260_)
);

OAI21X1 _7381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(\datapath_1.regfile_1.regEn_4_bF$buf0 ),
    .C(_260_),
    .Y(_198_[31])
);

DFFSR _7382_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_198_[0]),
    .Q(\datapath_1.regfile_1.regOut[4] [0]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _7383_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_198_[1]),
    .Q(\datapath_1.regfile_1.regOut[4] [1]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _7384_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_198_[2]),
    .Q(\datapath_1.regfile_1.regOut[4] [2]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _7385_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_198_[3]),
    .Q(\datapath_1.regfile_1.regOut[4] [3]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _7386_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_198_[4]),
    .Q(\datapath_1.regfile_1.regOut[4] [4]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _7387_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_198_[5]),
    .Q(\datapath_1.regfile_1.regOut[4] [5]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _7388_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_198_[6]),
    .Q(\datapath_1.regfile_1.regOut[4] [6]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _7389_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_198_[7]),
    .Q(\datapath_1.regfile_1.regOut[4] [7]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _7390_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_198_[8]),
    .Q(\datapath_1.regfile_1.regOut[4] [8]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _7391_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_198_[9]),
    .Q(\datapath_1.regfile_1.regOut[4] [9]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _7392_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_198_[10]),
    .Q(\datapath_1.regfile_1.regOut[4] [10]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _7393_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_198_[11]),
    .Q(\datapath_1.regfile_1.regOut[4] [11]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _7394_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_198_[12]),
    .Q(\datapath_1.regfile_1.regOut[4] [12]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _7395_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_198_[13]),
    .Q(\datapath_1.regfile_1.regOut[4] [13]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _7396_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_198_[14]),
    .Q(\datapath_1.regfile_1.regOut[4] [14]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _7397_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_198_[15]),
    .Q(\datapath_1.regfile_1.regOut[4] [15]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _7398_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_198_[16]),
    .Q(\datapath_1.regfile_1.regOut[4] [16]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _7399_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_198_[17]),
    .Q(\datapath_1.regfile_1.regOut[4] [17]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _7400_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_198_[18]),
    .Q(\datapath_1.regfile_1.regOut[4] [18]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _7401_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_198_[19]),
    .Q(\datapath_1.regfile_1.regOut[4] [19]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _7402_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_198_[20]),
    .Q(\datapath_1.regfile_1.regOut[4] [20]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _7403_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_198_[21]),
    .Q(\datapath_1.regfile_1.regOut[4] [21]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _7404_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_198_[22]),
    .Q(\datapath_1.regfile_1.regOut[4] [22]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _7405_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_198_[23]),
    .Q(\datapath_1.regfile_1.regOut[4] [23]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _7406_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_198_[24]),
    .Q(\datapath_1.regfile_1.regOut[4] [24]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _7407_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_198_[25]),
    .Q(\datapath_1.regfile_1.regOut[4] [25]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _7408_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_198_[26]),
    .Q(\datapath_1.regfile_1.regOut[4] [26]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _7409_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_198_[27]),
    .Q(\datapath_1.regfile_1.regOut[4] [27]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _7410_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_198_[28]),
    .Q(\datapath_1.regfile_1.regOut[4] [28]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _7411_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_198_[29]),
    .Q(\datapath_1.regfile_1.regOut[4] [29]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _7412_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_198_[30]),
    .Q(\datapath_1.regfile_1.regOut[4] [30]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _7413_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_198_[31]),
    .Q(\datapath_1.regfile_1.regOut[4] [31]),
    .R(rst_bF$buf104),
    .S(vdd)
);

INVX1 _7414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [0]),
    .Y(_326_)
);

NAND2X1 _7415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .Y(_327_)
);

OAI21X1 _7416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_327_),
    .Y(_263_[0])
);

INVX1 _7417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [1]),
    .Y(_264_)
);

NAND2X1 _7418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_265_)
);

OAI21X1 _7419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_265_),
    .Y(_263_[1])
);

INVX1 _7420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [2]),
    .Y(_266_)
);

NAND2X1 _7421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_267_)
);

OAI21X1 _7422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_267_),
    .Y(_263_[2])
);

INVX1 _7423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [3]),
    .Y(_268_)
);

NAND2X1 _7424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_269_)
);

OAI21X1 _7425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_269_),
    .Y(_263_[3])
);

INVX1 _7426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [4]),
    .Y(_270_)
);

NAND2X1 _7427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_271_)
);

OAI21X1 _7428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_271_),
    .Y(_263_[4])
);

INVX1 _7429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [5]),
    .Y(_272_)
);

NAND2X1 _7430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_273_)
);

OAI21X1 _7431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_273_),
    .Y(_263_[5])
);

INVX1 _7432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [6]),
    .Y(_274_)
);

NAND2X1 _7433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_275_)
);

OAI21X1 _7434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_275_),
    .Y(_263_[6])
);

INVX1 _7435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [7]),
    .Y(_276_)
);

NAND2X1 _7436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_277_)
);

OAI21X1 _7437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_277_),
    .Y(_263_[7])
);

INVX1 _7438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [8]),
    .Y(_278_)
);

NAND2X1 _7439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_279_)
);

OAI21X1 _7440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_279_),
    .Y(_263_[8])
);

INVX1 _7441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [9]),
    .Y(_280_)
);

NAND2X1 _7442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_281_)
);

OAI21X1 _7443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_281_),
    .Y(_263_[9])
);

INVX1 _7444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [10]),
    .Y(_282_)
);

NAND2X1 _7445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_283_)
);

OAI21X1 _7446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_283_),
    .Y(_263_[10])
);

INVX1 _7447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [11]),
    .Y(_284_)
);

NAND2X1 _7448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_285_)
);

OAI21X1 _7449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_285_),
    .Y(_263_[11])
);

INVX1 _7450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [12]),
    .Y(_286_)
);

NAND2X1 _7451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_287_)
);

OAI21X1 _7452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_287_),
    .Y(_263_[12])
);

INVX1 _7453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [13]),
    .Y(_288_)
);

NAND2X1 _7454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_289_)
);

OAI21X1 _7455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_289_),
    .Y(_263_[13])
);

INVX1 _7456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [14]),
    .Y(_290_)
);

NAND2X1 _7457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_291_)
);

OAI21X1 _7458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_291_),
    .Y(_263_[14])
);

INVX1 _7459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [15]),
    .Y(_292_)
);

NAND2X1 _7460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_293_)
);

OAI21X1 _7461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_293_),
    .Y(_263_[15])
);

INVX1 _7462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [16]),
    .Y(_294_)
);

NAND2X1 _7463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_295_)
);

OAI21X1 _7464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_295_),
    .Y(_263_[16])
);

INVX1 _7465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [17]),
    .Y(_296_)
);

NAND2X1 _7466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_297_)
);

OAI21X1 _7467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_297_),
    .Y(_263_[17])
);

INVX1 _7468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [18]),
    .Y(_298_)
);

NAND2X1 _7469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_299_)
);

OAI21X1 _7470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_299_),
    .Y(_263_[18])
);

INVX1 _7471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [19]),
    .Y(_300_)
);

NAND2X1 _7472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_301_)
);

OAI21X1 _7473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_301_),
    .Y(_263_[19])
);

INVX1 _7474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [20]),
    .Y(_302_)
);

NAND2X1 _7475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_303_)
);

OAI21X1 _7476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_303_),
    .Y(_263_[20])
);

INVX1 _7477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [21]),
    .Y(_304_)
);

NAND2X1 _7478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_305_)
);

OAI21X1 _7479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_305_),
    .Y(_263_[21])
);

INVX1 _7480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [22]),
    .Y(_306_)
);

NAND2X1 _7481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_307_)
);

OAI21X1 _7482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_307_),
    .Y(_263_[22])
);

INVX1 _7483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [23]),
    .Y(_308_)
);

NAND2X1 _7484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_309_)
);

OAI21X1 _7485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_309_),
    .Y(_263_[23])
);

INVX1 _7486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [24]),
    .Y(_310_)
);

NAND2X1 _7487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_311_)
);

OAI21X1 _7488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_311_),
    .Y(_263_[24])
);

INVX1 _7489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [25]),
    .Y(_312_)
);

NAND2X1 _7490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_313_)
);

OAI21X1 _7491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_313_),
    .Y(_263_[25])
);

INVX1 _7492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [26]),
    .Y(_314_)
);

NAND2X1 _7493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_315_)
);

OAI21X1 _7494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_315_),
    .Y(_263_[26])
);

INVX1 _7495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [27]),
    .Y(_316_)
);

NAND2X1 _7496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_317_)
);

OAI21X1 _7497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_317_),
    .Y(_263_[27])
);

INVX1 _7498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [28]),
    .Y(_318_)
);

NAND2X1 _7499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_319_)
);

OAI21X1 _7500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf6 ),
    .C(_319_),
    .Y(_263_[28])
);

INVX1 _7501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [29]),
    .Y(_320_)
);

NAND2X1 _7502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_321_)
);

OAI21X1 _7503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf4 ),
    .C(_321_),
    .Y(_263_[29])
);

INVX1 _7504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [30]),
    .Y(_322_)
);

NAND2X1 _7505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_323_)
);

OAI21X1 _7506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf2 ),
    .C(_323_),
    .Y(_263_[30])
);

INVX1 _7507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[5] [31]),
    .Y(_324_)
);

NAND2X1 _7508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_5_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_325_)
);

OAI21X1 _7509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(\datapath_1.regfile_1.regEn_5_bF$buf0 ),
    .C(_325_),
    .Y(_263_[31])
);

DFFSR _7510_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_263_[0]),
    .Q(\datapath_1.regfile_1.regOut[5] [0]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _7511_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_263_[1]),
    .Q(\datapath_1.regfile_1.regOut[5] [1]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _7512_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_263_[2]),
    .Q(\datapath_1.regfile_1.regOut[5] [2]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _7513_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_263_[3]),
    .Q(\datapath_1.regfile_1.regOut[5] [3]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _7514_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_263_[4]),
    .Q(\datapath_1.regfile_1.regOut[5] [4]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _7515_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_263_[5]),
    .Q(\datapath_1.regfile_1.regOut[5] [5]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _7516_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_263_[6]),
    .Q(\datapath_1.regfile_1.regOut[5] [6]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _7517_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_263_[7]),
    .Q(\datapath_1.regfile_1.regOut[5] [7]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _7518_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_263_[8]),
    .Q(\datapath_1.regfile_1.regOut[5] [8]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _7519_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_263_[9]),
    .Q(\datapath_1.regfile_1.regOut[5] [9]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _7520_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_263_[10]),
    .Q(\datapath_1.regfile_1.regOut[5] [10]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _7521_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_263_[11]),
    .Q(\datapath_1.regfile_1.regOut[5] [11]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _7522_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_263_[12]),
    .Q(\datapath_1.regfile_1.regOut[5] [12]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _7523_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_263_[13]),
    .Q(\datapath_1.regfile_1.regOut[5] [13]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _7524_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_263_[14]),
    .Q(\datapath_1.regfile_1.regOut[5] [14]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _7525_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_263_[15]),
    .Q(\datapath_1.regfile_1.regOut[5] [15]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _7526_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_263_[16]),
    .Q(\datapath_1.regfile_1.regOut[5] [16]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _7527_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_263_[17]),
    .Q(\datapath_1.regfile_1.regOut[5] [17]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _7528_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_263_[18]),
    .Q(\datapath_1.regfile_1.regOut[5] [18]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _7529_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_263_[19]),
    .Q(\datapath_1.regfile_1.regOut[5] [19]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _7530_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_263_[20]),
    .Q(\datapath_1.regfile_1.regOut[5] [20]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _7531_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_263_[21]),
    .Q(\datapath_1.regfile_1.regOut[5] [21]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _7532_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_263_[22]),
    .Q(\datapath_1.regfile_1.regOut[5] [22]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _7533_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_263_[23]),
    .Q(\datapath_1.regfile_1.regOut[5] [23]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _7534_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_263_[24]),
    .Q(\datapath_1.regfile_1.regOut[5] [24]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _7535_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_263_[25]),
    .Q(\datapath_1.regfile_1.regOut[5] [25]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _7536_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_263_[26]),
    .Q(\datapath_1.regfile_1.regOut[5] [26]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _7537_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_263_[27]),
    .Q(\datapath_1.regfile_1.regOut[5] [27]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _7538_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_263_[28]),
    .Q(\datapath_1.regfile_1.regOut[5] [28]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _7539_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_263_[29]),
    .Q(\datapath_1.regfile_1.regOut[5] [29]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _7540_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_263_[30]),
    .Q(\datapath_1.regfile_1.regOut[5] [30]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _7541_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_263_[31]),
    .Q(\datapath_1.regfile_1.regOut[5] [31]),
    .R(rst_bF$buf72),
    .S(vdd)
);

INVX1 _7542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [0]),
    .Y(_391_)
);

NAND2X1 _7543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .Y(_392_)
);

OAI21X1 _7544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_392_),
    .Y(_328_[0])
);

INVX1 _7545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [1]),
    .Y(_329_)
);

NAND2X1 _7546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_330_)
);

OAI21X1 _7547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_330_),
    .Y(_328_[1])
);

INVX1 _7548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [2]),
    .Y(_331_)
);

NAND2X1 _7549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_332_)
);

OAI21X1 _7550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_331_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_332_),
    .Y(_328_[2])
);

INVX1 _7551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [3]),
    .Y(_333_)
);

NAND2X1 _7552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_334_)
);

OAI21X1 _7553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_334_),
    .Y(_328_[3])
);

INVX1 _7554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [4]),
    .Y(_335_)
);

NAND2X1 _7555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_336_)
);

OAI21X1 _7556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_336_),
    .Y(_328_[4])
);

INVX1 _7557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [5]),
    .Y(_337_)
);

NAND2X1 _7558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_338_)
);

OAI21X1 _7559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_337_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_338_),
    .Y(_328_[5])
);

INVX1 _7560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [6]),
    .Y(_339_)
);

NAND2X1 _7561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_340_)
);

OAI21X1 _7562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_340_),
    .Y(_328_[6])
);

INVX1 _7563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [7]),
    .Y(_341_)
);

NAND2X1 _7564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_342_)
);

OAI21X1 _7565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_342_),
    .Y(_328_[7])
);

INVX1 _7566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [8]),
    .Y(_343_)
);

NAND2X1 _7567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_344_)
);

OAI21X1 _7568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_344_),
    .Y(_328_[8])
);

INVX1 _7569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [9]),
    .Y(_345_)
);

NAND2X1 _7570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_346_)
);

OAI21X1 _7571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_346_),
    .Y(_328_[9])
);

INVX1 _7572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [10]),
    .Y(_347_)
);

NAND2X1 _7573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_348_)
);

OAI21X1 _7574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_348_),
    .Y(_328_[10])
);

INVX1 _7575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [11]),
    .Y(_349_)
);

NAND2X1 _7576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_350_)
);

OAI21X1 _7577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_350_),
    .Y(_328_[11])
);

INVX1 _7578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [12]),
    .Y(_351_)
);

NAND2X1 _7579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_352_)
);

OAI21X1 _7580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_352_),
    .Y(_328_[12])
);

INVX1 _7581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [13]),
    .Y(_353_)
);

NAND2X1 _7582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_354_)
);

OAI21X1 _7583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_354_),
    .Y(_328_[13])
);

INVX1 _7584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [14]),
    .Y(_355_)
);

NAND2X1 _7585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_356_)
);

OAI21X1 _7586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_356_),
    .Y(_328_[14])
);

INVX1 _7587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [15]),
    .Y(_357_)
);

NAND2X1 _7588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_358_)
);

OAI21X1 _7589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_357_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_358_),
    .Y(_328_[15])
);

INVX1 _7590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [16]),
    .Y(_359_)
);

NAND2X1 _7591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_360_)
);

OAI21X1 _7592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_360_),
    .Y(_328_[16])
);

INVX1 _7593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [17]),
    .Y(_361_)
);

NAND2X1 _7594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_362_)
);

OAI21X1 _7595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_362_),
    .Y(_328_[17])
);

INVX1 _7596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [18]),
    .Y(_363_)
);

NAND2X1 _7597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_364_)
);

OAI21X1 _7598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_364_),
    .Y(_328_[18])
);

INVX1 _7599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [19]),
    .Y(_365_)
);

NAND2X1 _7600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_366_)
);

OAI21X1 _7601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_366_),
    .Y(_328_[19])
);

INVX1 _7602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [20]),
    .Y(_367_)
);

NAND2X1 _7603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_368_)
);

OAI21X1 _7604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_368_),
    .Y(_328_[20])
);

INVX1 _7605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [21]),
    .Y(_369_)
);

NAND2X1 _7606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_370_)
);

OAI21X1 _7607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_370_),
    .Y(_328_[21])
);

INVX1 _7608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [22]),
    .Y(_371_)
);

NAND2X1 _7609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_372_)
);

OAI21X1 _7610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_372_),
    .Y(_328_[22])
);

INVX1 _7611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [23]),
    .Y(_373_)
);

NAND2X1 _7612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_374_)
);

OAI21X1 _7613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_374_),
    .Y(_328_[23])
);

INVX1 _7614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [24]),
    .Y(_375_)
);

NAND2X1 _7615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_376_)
);

OAI21X1 _7616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_376_),
    .Y(_328_[24])
);

INVX1 _7617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [25]),
    .Y(_377_)
);

NAND2X1 _7618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_378_)
);

OAI21X1 _7619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_378_),
    .Y(_328_[25])
);

INVX1 _7620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [26]),
    .Y(_379_)
);

NAND2X1 _7621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_380_)
);

OAI21X1 _7622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_379_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_380_),
    .Y(_328_[26])
);

INVX1 _7623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [27]),
    .Y(_381_)
);

NAND2X1 _7624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_382_)
);

OAI21X1 _7625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_382_),
    .Y(_328_[27])
);

INVX1 _7626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [28]),
    .Y(_383_)
);

NAND2X1 _7627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_384_)
);

OAI21X1 _7628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf6 ),
    .C(_384_),
    .Y(_328_[28])
);

INVX1 _7629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [29]),
    .Y(_385_)
);

NAND2X1 _7630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_386_)
);

OAI21X1 _7631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf4 ),
    .C(_386_),
    .Y(_328_[29])
);

INVX1 _7632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [30]),
    .Y(_387_)
);

NAND2X1 _7633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_388_)
);

OAI21X1 _7634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_387_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf2 ),
    .C(_388_),
    .Y(_328_[30])
);

INVX1 _7635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[6] [31]),
    .Y(_389_)
);

NAND2X1 _7636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_6_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_390_)
);

OAI21X1 _7637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(\datapath_1.regfile_1.regEn_6_bF$buf0 ),
    .C(_390_),
    .Y(_328_[31])
);

DFFSR _7638_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_328_[0]),
    .Q(\datapath_1.regfile_1.regOut[6] [0]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _7639_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_328_[1]),
    .Q(\datapath_1.regfile_1.regOut[6] [1]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _7640_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_328_[2]),
    .Q(\datapath_1.regfile_1.regOut[6] [2]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _7641_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_328_[3]),
    .Q(\datapath_1.regfile_1.regOut[6] [3]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _7642_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_328_[4]),
    .Q(\datapath_1.regfile_1.regOut[6] [4]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _7643_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_328_[5]),
    .Q(\datapath_1.regfile_1.regOut[6] [5]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _7644_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_328_[6]),
    .Q(\datapath_1.regfile_1.regOut[6] [6]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _7645_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_328_[7]),
    .Q(\datapath_1.regfile_1.regOut[6] [7]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _7646_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_328_[8]),
    .Q(\datapath_1.regfile_1.regOut[6] [8]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _7647_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_328_[9]),
    .Q(\datapath_1.regfile_1.regOut[6] [9]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _7648_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_328_[10]),
    .Q(\datapath_1.regfile_1.regOut[6] [10]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _7649_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_328_[11]),
    .Q(\datapath_1.regfile_1.regOut[6] [11]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _7650_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_328_[12]),
    .Q(\datapath_1.regfile_1.regOut[6] [12]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _7651_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_328_[13]),
    .Q(\datapath_1.regfile_1.regOut[6] [13]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _7652_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_328_[14]),
    .Q(\datapath_1.regfile_1.regOut[6] [14]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _7653_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_328_[15]),
    .Q(\datapath_1.regfile_1.regOut[6] [15]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _7654_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_328_[16]),
    .Q(\datapath_1.regfile_1.regOut[6] [16]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _7655_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_328_[17]),
    .Q(\datapath_1.regfile_1.regOut[6] [17]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _7656_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_328_[18]),
    .Q(\datapath_1.regfile_1.regOut[6] [18]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _7657_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_328_[19]),
    .Q(\datapath_1.regfile_1.regOut[6] [19]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _7658_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_328_[20]),
    .Q(\datapath_1.regfile_1.regOut[6] [20]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _7659_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_328_[21]),
    .Q(\datapath_1.regfile_1.regOut[6] [21]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _7660_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_328_[22]),
    .Q(\datapath_1.regfile_1.regOut[6] [22]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _7661_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_328_[23]),
    .Q(\datapath_1.regfile_1.regOut[6] [23]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _7662_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_328_[24]),
    .Q(\datapath_1.regfile_1.regOut[6] [24]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _7663_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_328_[25]),
    .Q(\datapath_1.regfile_1.regOut[6] [25]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _7664_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_328_[26]),
    .Q(\datapath_1.regfile_1.regOut[6] [26]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _7665_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_328_[27]),
    .Q(\datapath_1.regfile_1.regOut[6] [27]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _7666_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_328_[28]),
    .Q(\datapath_1.regfile_1.regOut[6] [28]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _7667_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_328_[29]),
    .Q(\datapath_1.regfile_1.regOut[6] [29]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _7668_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_328_[30]),
    .Q(\datapath_1.regfile_1.regOut[6] [30]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _7669_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_328_[31]),
    .Q(\datapath_1.regfile_1.regOut[6] [31]),
    .R(rst_bF$buf40),
    .S(vdd)
);

INVX1 _7670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [0]),
    .Y(_456_)
);

NAND2X1 _7671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .Y(_457_)
);

OAI21X1 _7672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_457_),
    .Y(_393_[0])
);

INVX1 _7673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [1]),
    .Y(_394_)
);

NAND2X1 _7674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_395_)
);

OAI21X1 _7675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_395_),
    .Y(_393_[1])
);

INVX1 _7676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [2]),
    .Y(_396_)
);

NAND2X1 _7677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_397_)
);

OAI21X1 _7678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_397_),
    .Y(_393_[2])
);

INVX1 _7679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [3]),
    .Y(_398_)
);

NAND2X1 _7680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_399_)
);

OAI21X1 _7681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_399_),
    .Y(_393_[3])
);

INVX1 _7682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [4]),
    .Y(_400_)
);

NAND2X1 _7683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_401_)
);

OAI21X1 _7684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_401_),
    .Y(_393_[4])
);

INVX1 _7685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [5]),
    .Y(_402_)
);

NAND2X1 _7686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_403_)
);

OAI21X1 _7687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_403_),
    .Y(_393_[5])
);

INVX1 _7688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [6]),
    .Y(_404_)
);

NAND2X1 _7689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_405_)
);

OAI21X1 _7690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_405_),
    .Y(_393_[6])
);

INVX1 _7691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [7]),
    .Y(_406_)
);

NAND2X1 _7692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_407_)
);

OAI21X1 _7693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_407_),
    .Y(_393_[7])
);

INVX1 _7694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [8]),
    .Y(_408_)
);

NAND2X1 _7695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_409_)
);

OAI21X1 _7696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_409_),
    .Y(_393_[8])
);

INVX1 _7697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [9]),
    .Y(_410_)
);

NAND2X1 _7698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_411_)
);

OAI21X1 _7699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_411_),
    .Y(_393_[9])
);

INVX1 _7700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [10]),
    .Y(_412_)
);

NAND2X1 _7701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_413_)
);

OAI21X1 _7702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_412_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_413_),
    .Y(_393_[10])
);

INVX1 _7703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [11]),
    .Y(_414_)
);

NAND2X1 _7704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_415_)
);

OAI21X1 _7705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_415_),
    .Y(_393_[11])
);

INVX1 _7706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [12]),
    .Y(_416_)
);

NAND2X1 _7707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_417_)
);

OAI21X1 _7708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_417_),
    .Y(_393_[12])
);

INVX1 _7709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [13]),
    .Y(_418_)
);

NAND2X1 _7710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_419_)
);

OAI21X1 _7711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_418_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_419_),
    .Y(_393_[13])
);

INVX1 _7712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [14]),
    .Y(_420_)
);

NAND2X1 _7713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_421_)
);

OAI21X1 _7714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_421_),
    .Y(_393_[14])
);

INVX1 _7715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [15]),
    .Y(_422_)
);

NAND2X1 _7716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_423_)
);

OAI21X1 _7717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_423_),
    .Y(_393_[15])
);

INVX1 _7718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [16]),
    .Y(_424_)
);

NAND2X1 _7719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_425_)
);

OAI21X1 _7720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_425_),
    .Y(_393_[16])
);

INVX1 _7721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [17]),
    .Y(_426_)
);

NAND2X1 _7722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_427_)
);

OAI21X1 _7723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_427_),
    .Y(_393_[17])
);

INVX1 _7724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [18]),
    .Y(_428_)
);

NAND2X1 _7725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_429_)
);

OAI21X1 _7726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_429_),
    .Y(_393_[18])
);

INVX1 _7727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [19]),
    .Y(_430_)
);

NAND2X1 _7728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_431_)
);

OAI21X1 _7729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_431_),
    .Y(_393_[19])
);

INVX1 _7730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [20]),
    .Y(_432_)
);

NAND2X1 _7731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_433_)
);

OAI21X1 _7732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_433_),
    .Y(_393_[20])
);

INVX1 _7733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [21]),
    .Y(_434_)
);

NAND2X1 _7734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_435_)
);

OAI21X1 _7735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_435_),
    .Y(_393_[21])
);

INVX1 _7736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [22]),
    .Y(_436_)
);

NAND2X1 _7737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_437_)
);

OAI21X1 _7738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_436_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_437_),
    .Y(_393_[22])
);

INVX1 _7739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [23]),
    .Y(_438_)
);

NAND2X1 _7740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_439_)
);

OAI21X1 _7741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_439_),
    .Y(_393_[23])
);

INVX1 _7742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [24]),
    .Y(_440_)
);

NAND2X1 _7743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_441_)
);

OAI21X1 _7744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_441_),
    .Y(_393_[24])
);

INVX1 _7745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [25]),
    .Y(_442_)
);

NAND2X1 _7746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_443_)
);

OAI21X1 _7747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_443_),
    .Y(_393_[25])
);

INVX1 _7748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [26]),
    .Y(_444_)
);

NAND2X1 _7749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_445_)
);

OAI21X1 _7750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_445_),
    .Y(_393_[26])
);

INVX1 _7751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [27]),
    .Y(_446_)
);

NAND2X1 _7752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_447_)
);

OAI21X1 _7753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_447_),
    .Y(_393_[27])
);

INVX1 _7754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [28]),
    .Y(_448_)
);

NAND2X1 _7755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_449_)
);

OAI21X1 _7756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_448_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf6 ),
    .C(_449_),
    .Y(_393_[28])
);

INVX1 _7757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [29]),
    .Y(_450_)
);

NAND2X1 _7758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_451_)
);

OAI21X1 _7759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf4 ),
    .C(_451_),
    .Y(_393_[29])
);

INVX1 _7760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [30]),
    .Y(_452_)
);

NAND2X1 _7761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_453_)
);

OAI21X1 _7762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_452_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf2 ),
    .C(_453_),
    .Y(_393_[30])
);

INVX1 _7763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[7] [31]),
    .Y(_454_)
);

NAND2X1 _7764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_7_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_455_)
);

OAI21X1 _7765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(\datapath_1.regfile_1.regEn_7_bF$buf0 ),
    .C(_455_),
    .Y(_393_[31])
);

DFFSR _7766_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_393_[0]),
    .Q(\datapath_1.regfile_1.regOut[7] [0]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _7767_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_393_[1]),
    .Q(\datapath_1.regfile_1.regOut[7] [1]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _7768_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_393_[2]),
    .Q(\datapath_1.regfile_1.regOut[7] [2]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _7769_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_393_[3]),
    .Q(\datapath_1.regfile_1.regOut[7] [3]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _7770_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_393_[4]),
    .Q(\datapath_1.regfile_1.regOut[7] [4]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _7771_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_393_[5]),
    .Q(\datapath_1.regfile_1.regOut[7] [5]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _7772_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_393_[6]),
    .Q(\datapath_1.regfile_1.regOut[7] [6]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _7773_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_393_[7]),
    .Q(\datapath_1.regfile_1.regOut[7] [7]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _7774_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_393_[8]),
    .Q(\datapath_1.regfile_1.regOut[7] [8]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _7775_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_393_[9]),
    .Q(\datapath_1.regfile_1.regOut[7] [9]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _7776_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_393_[10]),
    .Q(\datapath_1.regfile_1.regOut[7] [10]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _7777_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_393_[11]),
    .Q(\datapath_1.regfile_1.regOut[7] [11]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _7778_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_393_[12]),
    .Q(\datapath_1.regfile_1.regOut[7] [12]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _7779_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_393_[13]),
    .Q(\datapath_1.regfile_1.regOut[7] [13]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _7780_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_393_[14]),
    .Q(\datapath_1.regfile_1.regOut[7] [14]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _7781_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_393_[15]),
    .Q(\datapath_1.regfile_1.regOut[7] [15]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _7782_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_393_[16]),
    .Q(\datapath_1.regfile_1.regOut[7] [16]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _7783_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_393_[17]),
    .Q(\datapath_1.regfile_1.regOut[7] [17]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _7784_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_393_[18]),
    .Q(\datapath_1.regfile_1.regOut[7] [18]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _7785_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_393_[19]),
    .Q(\datapath_1.regfile_1.regOut[7] [19]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _7786_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_393_[20]),
    .Q(\datapath_1.regfile_1.regOut[7] [20]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _7787_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_393_[21]),
    .Q(\datapath_1.regfile_1.regOut[7] [21]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _7788_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_393_[22]),
    .Q(\datapath_1.regfile_1.regOut[7] [22]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _7789_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_393_[23]),
    .Q(\datapath_1.regfile_1.regOut[7] [23]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _7790_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_393_[24]),
    .Q(\datapath_1.regfile_1.regOut[7] [24]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _7791_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_393_[25]),
    .Q(\datapath_1.regfile_1.regOut[7] [25]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _7792_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_393_[26]),
    .Q(\datapath_1.regfile_1.regOut[7] [26]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _7793_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_393_[27]),
    .Q(\datapath_1.regfile_1.regOut[7] [27]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _7794_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_393_[28]),
    .Q(\datapath_1.regfile_1.regOut[7] [28]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _7795_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_393_[29]),
    .Q(\datapath_1.regfile_1.regOut[7] [29]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _7796_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_393_[30]),
    .Q(\datapath_1.regfile_1.regOut[7] [30]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _7797_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_393_[31]),
    .Q(\datapath_1.regfile_1.regOut[7] [31]),
    .R(rst_bF$buf8),
    .S(vdd)
);

INVX1 _7798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [0]),
    .Y(_521_)
);

NAND2X1 _7799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .Y(_522_)
);

OAI21X1 _7800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_522_),
    .Y(_458_[0])
);

INVX1 _7801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [1]),
    .Y(_459_)
);

NAND2X1 _7802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_460_)
);

OAI21X1 _7803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_460_),
    .Y(_458_[1])
);

INVX1 _7804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [2]),
    .Y(_461_)
);

NAND2X1 _7805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_462_)
);

OAI21X1 _7806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_462_),
    .Y(_458_[2])
);

INVX1 _7807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [3]),
    .Y(_463_)
);

NAND2X1 _7808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_464_)
);

OAI21X1 _7809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_464_),
    .Y(_458_[3])
);

INVX1 _7810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [4]),
    .Y(_465_)
);

NAND2X1 _7811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_466_)
);

OAI21X1 _7812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_466_),
    .Y(_458_[4])
);

INVX1 _7813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [5]),
    .Y(_467_)
);

NAND2X1 _7814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_468_)
);

OAI21X1 _7815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_467_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_468_),
    .Y(_458_[5])
);

INVX1 _7816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [6]),
    .Y(_469_)
);

NAND2X1 _7817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_470_)
);

OAI21X1 _7818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_469_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_470_),
    .Y(_458_[6])
);

INVX1 _7819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [7]),
    .Y(_471_)
);

NAND2X1 _7820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_472_)
);

OAI21X1 _7821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_471_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_472_),
    .Y(_458_[7])
);

INVX1 _7822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [8]),
    .Y(_473_)
);

NAND2X1 _7823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_474_)
);

OAI21X1 _7824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_474_),
    .Y(_458_[8])
);

INVX1 _7825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [9]),
    .Y(_475_)
);

NAND2X1 _7826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_476_)
);

OAI21X1 _7827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_476_),
    .Y(_458_[9])
);

INVX1 _7828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [10]),
    .Y(_477_)
);

NAND2X1 _7829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_478_)
);

OAI21X1 _7830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_478_),
    .Y(_458_[10])
);

INVX1 _7831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [11]),
    .Y(_479_)
);

NAND2X1 _7832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_480_)
);

OAI21X1 _7833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_480_),
    .Y(_458_[11])
);

INVX1 _7834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [12]),
    .Y(_481_)
);

NAND2X1 _7835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_482_)
);

OAI21X1 _7836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_481_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_482_),
    .Y(_458_[12])
);

INVX1 _7837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [13]),
    .Y(_483_)
);

NAND2X1 _7838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_484_)
);

OAI21X1 _7839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_484_),
    .Y(_458_[13])
);

INVX1 _7840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [14]),
    .Y(_485_)
);

NAND2X1 _7841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_486_)
);

OAI21X1 _7842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_486_),
    .Y(_458_[14])
);

INVX1 _7843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [15]),
    .Y(_487_)
);

NAND2X1 _7844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_488_)
);

OAI21X1 _7845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_488_),
    .Y(_458_[15])
);

INVX1 _7846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [16]),
    .Y(_489_)
);

NAND2X1 _7847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_490_)
);

OAI21X1 _7848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_490_),
    .Y(_458_[16])
);

INVX1 _7849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [17]),
    .Y(_491_)
);

NAND2X1 _7850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_492_)
);

OAI21X1 _7851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_492_),
    .Y(_458_[17])
);

INVX1 _7852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [18]),
    .Y(_493_)
);

NAND2X1 _7853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_494_)
);

OAI21X1 _7854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_494_),
    .Y(_458_[18])
);

INVX1 _7855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [19]),
    .Y(_495_)
);

NAND2X1 _7856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_496_)
);

OAI21X1 _7857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_496_),
    .Y(_458_[19])
);

INVX1 _7858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [20]),
    .Y(_497_)
);

NAND2X1 _7859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_498_)
);

OAI21X1 _7860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_498_),
    .Y(_458_[20])
);

INVX1 _7861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [21]),
    .Y(_499_)
);

NAND2X1 _7862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_500_)
);

OAI21X1 _7863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_500_),
    .Y(_458_[21])
);

INVX1 _7864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [22]),
    .Y(_501_)
);

NAND2X1 _7865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_502_)
);

OAI21X1 _7866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_502_),
    .Y(_458_[22])
);

INVX1 _7867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [23]),
    .Y(_503_)
);

NAND2X1 _7868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_504_)
);

OAI21X1 _7869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_504_),
    .Y(_458_[23])
);

INVX1 _7870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [24]),
    .Y(_505_)
);

NAND2X1 _7871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_506_)
);

OAI21X1 _7872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_506_),
    .Y(_458_[24])
);

INVX1 _7873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [25]),
    .Y(_507_)
);

NAND2X1 _7874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_508_)
);

OAI21X1 _7875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_507_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_508_),
    .Y(_458_[25])
);

INVX1 _7876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [26]),
    .Y(_509_)
);

NAND2X1 _7877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_510_)
);

OAI21X1 _7878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_509_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_510_),
    .Y(_458_[26])
);

INVX1 _7879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [27]),
    .Y(_511_)
);

NAND2X1 _7880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_512_)
);

OAI21X1 _7881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_512_),
    .Y(_458_[27])
);

INVX1 _7882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [28]),
    .Y(_513_)
);

NAND2X1 _7883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_514_)
);

OAI21X1 _7884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_513_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf6 ),
    .C(_514_),
    .Y(_458_[28])
);

INVX1 _7885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [29]),
    .Y(_515_)
);

NAND2X1 _7886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_516_)
);

OAI21X1 _7887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf4 ),
    .C(_516_),
    .Y(_458_[29])
);

INVX1 _7888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [30]),
    .Y(_517_)
);

NAND2X1 _7889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_518_)
);

OAI21X1 _7890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_517_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf2 ),
    .C(_518_),
    .Y(_458_[30])
);

INVX1 _7891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[8] [31]),
    .Y(_519_)
);

NAND2X1 _7892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_8_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_520_)
);

OAI21X1 _7893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_519_),
    .B(\datapath_1.regfile_1.regEn_8_bF$buf0 ),
    .C(_520_),
    .Y(_458_[31])
);

DFFSR _7894_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_458_[0]),
    .Q(\datapath_1.regfile_1.regOut[8] [0]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _7895_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_458_[1]),
    .Q(\datapath_1.regfile_1.regOut[8] [1]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _7896_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_458_[2]),
    .Q(\datapath_1.regfile_1.regOut[8] [2]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _7897_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_458_[3]),
    .Q(\datapath_1.regfile_1.regOut[8] [3]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _7898_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_458_[4]),
    .Q(\datapath_1.regfile_1.regOut[8] [4]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _7899_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_458_[5]),
    .Q(\datapath_1.regfile_1.regOut[8] [5]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _7900_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_458_[6]),
    .Q(\datapath_1.regfile_1.regOut[8] [6]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _7901_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_458_[7]),
    .Q(\datapath_1.regfile_1.regOut[8] [7]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _7902_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_458_[8]),
    .Q(\datapath_1.regfile_1.regOut[8] [8]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _7903_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_458_[9]),
    .Q(\datapath_1.regfile_1.regOut[8] [9]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _7904_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_458_[10]),
    .Q(\datapath_1.regfile_1.regOut[8] [10]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _7905_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_458_[11]),
    .Q(\datapath_1.regfile_1.regOut[8] [11]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _7906_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_458_[12]),
    .Q(\datapath_1.regfile_1.regOut[8] [12]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _7907_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_458_[13]),
    .Q(\datapath_1.regfile_1.regOut[8] [13]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _7908_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_458_[14]),
    .Q(\datapath_1.regfile_1.regOut[8] [14]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _7909_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_458_[15]),
    .Q(\datapath_1.regfile_1.regOut[8] [15]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _7910_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_458_[16]),
    .Q(\datapath_1.regfile_1.regOut[8] [16]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _7911_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_458_[17]),
    .Q(\datapath_1.regfile_1.regOut[8] [17]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _7912_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_458_[18]),
    .Q(\datapath_1.regfile_1.regOut[8] [18]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _7913_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_458_[19]),
    .Q(\datapath_1.regfile_1.regOut[8] [19]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _7914_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_458_[20]),
    .Q(\datapath_1.regfile_1.regOut[8] [20]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _7915_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_458_[21]),
    .Q(\datapath_1.regfile_1.regOut[8] [21]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _7916_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_458_[22]),
    .Q(\datapath_1.regfile_1.regOut[8] [22]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _7917_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_458_[23]),
    .Q(\datapath_1.regfile_1.regOut[8] [23]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _7918_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_458_[24]),
    .Q(\datapath_1.regfile_1.regOut[8] [24]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _7919_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_458_[25]),
    .Q(\datapath_1.regfile_1.regOut[8] [25]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _7920_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_458_[26]),
    .Q(\datapath_1.regfile_1.regOut[8] [26]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _7921_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_458_[27]),
    .Q(\datapath_1.regfile_1.regOut[8] [27]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _7922_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_458_[28]),
    .Q(\datapath_1.regfile_1.regOut[8] [28]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _7923_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_458_[29]),
    .Q(\datapath_1.regfile_1.regOut[8] [29]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _7924_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_458_[30]),
    .Q(\datapath_1.regfile_1.regOut[8] [30]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _7925_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_458_[31]),
    .Q(\datapath_1.regfile_1.regOut[8] [31]),
    .R(rst_bF$buf90),
    .S(vdd)
);

INVX1 _7926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [0]),
    .Y(_586_)
);

NAND2X1 _7927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .Y(_587_)
);

OAI21X1 _7928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_587_),
    .Y(_523_[0])
);

INVX1 _7929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [1]),
    .Y(_524_)
);

NAND2X1 _7930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_525_)
);

OAI21X1 _7931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_525_),
    .Y(_523_[1])
);

INVX1 _7932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [2]),
    .Y(_526_)
);

NAND2X1 _7933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_527_)
);

OAI21X1 _7934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_527_),
    .Y(_523_[2])
);

INVX1 _7935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [3]),
    .Y(_528_)
);

NAND2X1 _7936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_529_)
);

OAI21X1 _7937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_529_),
    .Y(_523_[3])
);

INVX1 _7938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [4]),
    .Y(_530_)
);

NAND2X1 _7939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_531_)
);

OAI21X1 _7940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_531_),
    .Y(_523_[4])
);

INVX1 _7941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [5]),
    .Y(_532_)
);

NAND2X1 _7942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_533_)
);

OAI21X1 _7943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_532_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_533_),
    .Y(_523_[5])
);

INVX1 _7944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [6]),
    .Y(_534_)
);

NAND2X1 _7945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_535_)
);

OAI21X1 _7946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_535_),
    .Y(_523_[6])
);

INVX1 _7947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [7]),
    .Y(_536_)
);

NAND2X1 _7948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_537_)
);

OAI21X1 _7949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_537_),
    .Y(_523_[7])
);

INVX1 _7950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [8]),
    .Y(_538_)
);

NAND2X1 _7951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_539_)
);

OAI21X1 _7952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_538_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_539_),
    .Y(_523_[8])
);

INVX1 _7953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [9]),
    .Y(_540_)
);

NAND2X1 _7954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_541_)
);

OAI21X1 _7955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_540_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_541_),
    .Y(_523_[9])
);

INVX1 _7956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [10]),
    .Y(_542_)
);

NAND2X1 _7957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_543_)
);

OAI21X1 _7958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_543_),
    .Y(_523_[10])
);

INVX1 _7959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [11]),
    .Y(_544_)
);

NAND2X1 _7960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_545_)
);

OAI21X1 _7961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_544_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_545_),
    .Y(_523_[11])
);

INVX1 _7962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [12]),
    .Y(_546_)
);

NAND2X1 _7963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_547_)
);

OAI21X1 _7964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_547_),
    .Y(_523_[12])
);

INVX1 _7965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [13]),
    .Y(_548_)
);

NAND2X1 _7966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_549_)
);

OAI21X1 _7967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_549_),
    .Y(_523_[13])
);

INVX1 _7968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [14]),
    .Y(_550_)
);

NAND2X1 _7969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_551_)
);

OAI21X1 _7970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_551_),
    .Y(_523_[14])
);

INVX1 _7971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [15]),
    .Y(_552_)
);

NAND2X1 _7972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_553_)
);

OAI21X1 _7973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_553_),
    .Y(_523_[15])
);

INVX1 _7974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [16]),
    .Y(_554_)
);

NAND2X1 _7975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_555_)
);

OAI21X1 _7976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_555_),
    .Y(_523_[16])
);

INVX1 _7977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [17]),
    .Y(_556_)
);

NAND2X1 _7978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_557_)
);

OAI21X1 _7979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_557_),
    .Y(_523_[17])
);

INVX1 _7980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [18]),
    .Y(_558_)
);

NAND2X1 _7981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_559_)
);

OAI21X1 _7982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_558_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_559_),
    .Y(_523_[18])
);

INVX1 _7983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [19]),
    .Y(_560_)
);

NAND2X1 _7984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_561_)
);

OAI21X1 _7985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_561_),
    .Y(_523_[19])
);

INVX1 _7986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [20]),
    .Y(_562_)
);

NAND2X1 _7987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_563_)
);

OAI21X1 _7988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_563_),
    .Y(_523_[20])
);

INVX1 _7989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [21]),
    .Y(_564_)
);

NAND2X1 _7990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_565_)
);

OAI21X1 _7991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_564_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_565_),
    .Y(_523_[21])
);

INVX1 _7992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [22]),
    .Y(_566_)
);

NAND2X1 _7993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_567_)
);

OAI21X1 _7994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_567_),
    .Y(_523_[22])
);

INVX1 _7995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [23]),
    .Y(_568_)
);

NAND2X1 _7996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_569_)
);

OAI21X1 _7997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_568_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_569_),
    .Y(_523_[23])
);

INVX1 _7998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [24]),
    .Y(_570_)
);

NAND2X1 _7999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_571_)
);

OAI21X1 _8000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_570_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_571_),
    .Y(_523_[24])
);

INVX1 _8001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [25]),
    .Y(_572_)
);

NAND2X1 _8002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_573_)
);

OAI21X1 _8003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_573_),
    .Y(_523_[25])
);

INVX1 _8004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [26]),
    .Y(_574_)
);

NAND2X1 _8005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_575_)
);

OAI21X1 _8006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_575_),
    .Y(_523_[26])
);

INVX1 _8007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [27]),
    .Y(_576_)
);

NAND2X1 _8008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_577_)
);

OAI21X1 _8009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_577_),
    .Y(_523_[27])
);

INVX1 _8010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [28]),
    .Y(_578_)
);

NAND2X1 _8011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_579_)
);

OAI21X1 _8012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf6 ),
    .C(_579_),
    .Y(_523_[28])
);

INVX1 _8013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [29]),
    .Y(_580_)
);

NAND2X1 _8014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_581_)
);

OAI21X1 _8015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_580_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf4 ),
    .C(_581_),
    .Y(_523_[29])
);

INVX1 _8016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [30]),
    .Y(_582_)
);

NAND2X1 _8017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_583_)
);

OAI21X1 _8018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf2 ),
    .C(_583_),
    .Y(_523_[30])
);

INVX1 _8019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[9] [31]),
    .Y(_584_)
);

NAND2X1 _8020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_9_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_585_)
);

OAI21X1 _8021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .B(\datapath_1.regfile_1.regEn_9_bF$buf0 ),
    .C(_585_),
    .Y(_523_[31])
);

DFFSR _8022_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_523_[0]),
    .Q(\datapath_1.regfile_1.regOut[9] [0]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _8023_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_523_[1]),
    .Q(\datapath_1.regfile_1.regOut[9] [1]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _8024_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_523_[2]),
    .Q(\datapath_1.regfile_1.regOut[9] [2]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _8025_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_523_[3]),
    .Q(\datapath_1.regfile_1.regOut[9] [3]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _8026_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_523_[4]),
    .Q(\datapath_1.regfile_1.regOut[9] [4]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _8027_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_523_[5]),
    .Q(\datapath_1.regfile_1.regOut[9] [5]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _8028_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_523_[6]),
    .Q(\datapath_1.regfile_1.regOut[9] [6]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _8029_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_523_[7]),
    .Q(\datapath_1.regfile_1.regOut[9] [7]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _8030_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_523_[8]),
    .Q(\datapath_1.regfile_1.regOut[9] [8]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _8031_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_523_[9]),
    .Q(\datapath_1.regfile_1.regOut[9] [9]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _8032_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_523_[10]),
    .Q(\datapath_1.regfile_1.regOut[9] [10]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _8033_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_523_[11]),
    .Q(\datapath_1.regfile_1.regOut[9] [11]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _8034_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_523_[12]),
    .Q(\datapath_1.regfile_1.regOut[9] [12]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _8035_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_523_[13]),
    .Q(\datapath_1.regfile_1.regOut[9] [13]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _8036_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_523_[14]),
    .Q(\datapath_1.regfile_1.regOut[9] [14]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _8037_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_523_[15]),
    .Q(\datapath_1.regfile_1.regOut[9] [15]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _8038_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_523_[16]),
    .Q(\datapath_1.regfile_1.regOut[9] [16]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _8039_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_523_[17]),
    .Q(\datapath_1.regfile_1.regOut[9] [17]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _8040_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_523_[18]),
    .Q(\datapath_1.regfile_1.regOut[9] [18]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _8041_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_523_[19]),
    .Q(\datapath_1.regfile_1.regOut[9] [19]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _8042_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_523_[20]),
    .Q(\datapath_1.regfile_1.regOut[9] [20]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _8043_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_523_[21]),
    .Q(\datapath_1.regfile_1.regOut[9] [21]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _8044_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_523_[22]),
    .Q(\datapath_1.regfile_1.regOut[9] [22]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _8045_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_523_[23]),
    .Q(\datapath_1.regfile_1.regOut[9] [23]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _8046_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_523_[24]),
    .Q(\datapath_1.regfile_1.regOut[9] [24]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _8047_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_523_[25]),
    .Q(\datapath_1.regfile_1.regOut[9] [25]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _8048_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_523_[26]),
    .Q(\datapath_1.regfile_1.regOut[9] [26]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _8049_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_523_[27]),
    .Q(\datapath_1.regfile_1.regOut[9] [27]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _8050_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_523_[28]),
    .Q(\datapath_1.regfile_1.regOut[9] [28]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _8051_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_523_[29]),
    .Q(\datapath_1.regfile_1.regOut[9] [29]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _8052_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_523_[30]),
    .Q(\datapath_1.regfile_1.regOut[9] [30]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _8053_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_523_[31]),
    .Q(\datapath_1.regfile_1.regOut[9] [31]),
    .R(rst_bF$buf58),
    .S(vdd)
);

INVX1 _8054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [0]),
    .Y(_651_)
);

NAND2X1 _8055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .Y(_652_)
);

OAI21X1 _8056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_651_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_652_),
    .Y(_588_[0])
);

INVX1 _8057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [1]),
    .Y(_589_)
);

NAND2X1 _8058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_590_)
);

OAI21X1 _8059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_590_),
    .Y(_588_[1])
);

INVX1 _8060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [2]),
    .Y(_591_)
);

NAND2X1 _8061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_592_)
);

OAI21X1 _8062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_592_),
    .Y(_588_[2])
);

INVX1 _8063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [3]),
    .Y(_593_)
);

NAND2X1 _8064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_594_)
);

OAI21X1 _8065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_594_),
    .Y(_588_[3])
);

INVX1 _8066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [4]),
    .Y(_595_)
);

NAND2X1 _8067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_596_)
);

OAI21X1 _8068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_596_),
    .Y(_588_[4])
);

INVX1 _8069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [5]),
    .Y(_597_)
);

NAND2X1 _8070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_598_)
);

OAI21X1 _8071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_598_),
    .Y(_588_[5])
);

INVX1 _8072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [6]),
    .Y(_599_)
);

NAND2X1 _8073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_600_)
);

OAI21X1 _8074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_600_),
    .Y(_588_[6])
);

INVX1 _8075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [7]),
    .Y(_601_)
);

NAND2X1 _8076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_602_)
);

OAI21X1 _8077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_602_),
    .Y(_588_[7])
);

INVX1 _8078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [8]),
    .Y(_603_)
);

NAND2X1 _8079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_604_)
);

OAI21X1 _8080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_604_),
    .Y(_588_[8])
);

INVX1 _8081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [9]),
    .Y(_605_)
);

NAND2X1 _8082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_606_)
);

OAI21X1 _8083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_605_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_606_),
    .Y(_588_[9])
);

INVX1 _8084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [10]),
    .Y(_607_)
);

NAND2X1 _8085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_608_)
);

OAI21X1 _8086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_608_),
    .Y(_588_[10])
);

INVX1 _8087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [11]),
    .Y(_609_)
);

NAND2X1 _8088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_610_)
);

OAI21X1 _8089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_610_),
    .Y(_588_[11])
);

INVX1 _8090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [12]),
    .Y(_611_)
);

NAND2X1 _8091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_612_)
);

OAI21X1 _8092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_612_),
    .Y(_588_[12])
);

INVX1 _8093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [13]),
    .Y(_613_)
);

NAND2X1 _8094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_614_)
);

OAI21X1 _8095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_614_),
    .Y(_588_[13])
);

INVX1 _8096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [14]),
    .Y(_615_)
);

NAND2X1 _8097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_616_)
);

OAI21X1 _8098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_616_),
    .Y(_588_[14])
);

INVX1 _8099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [15]),
    .Y(_617_)
);

NAND2X1 _8100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_618_)
);

OAI21X1 _8101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_618_),
    .Y(_588_[15])
);

INVX1 _8102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [16]),
    .Y(_619_)
);

NAND2X1 _8103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_620_)
);

OAI21X1 _8104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_620_),
    .Y(_588_[16])
);

INVX1 _8105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [17]),
    .Y(_621_)
);

NAND2X1 _8106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_622_)
);

OAI21X1 _8107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_621_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_622_),
    .Y(_588_[17])
);

INVX1 _8108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [18]),
    .Y(_623_)
);

NAND2X1 _8109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_624_)
);

OAI21X1 _8110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_624_),
    .Y(_588_[18])
);

INVX1 _8111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [19]),
    .Y(_625_)
);

NAND2X1 _8112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_626_)
);

OAI21X1 _8113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_626_),
    .Y(_588_[19])
);

INVX1 _8114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [20]),
    .Y(_627_)
);

NAND2X1 _8115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_628_)
);

OAI21X1 _8116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_628_),
    .Y(_588_[20])
);

INVX1 _8117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [21]),
    .Y(_629_)
);

NAND2X1 _8118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_630_)
);

OAI21X1 _8119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_630_),
    .Y(_588_[21])
);

INVX1 _8120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [22]),
    .Y(_631_)
);

NAND2X1 _8121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_632_)
);

OAI21X1 _8122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_632_),
    .Y(_588_[22])
);

INVX1 _8123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [23]),
    .Y(_633_)
);

NAND2X1 _8124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_634_)
);

OAI21X1 _8125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_634_),
    .Y(_588_[23])
);

INVX1 _8126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [24]),
    .Y(_635_)
);

NAND2X1 _8127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_636_)
);

OAI21X1 _8128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_636_),
    .Y(_588_[24])
);

INVX1 _8129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [25]),
    .Y(_637_)
);

NAND2X1 _8130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_638_)
);

OAI21X1 _8131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_638_),
    .Y(_588_[25])
);

INVX1 _8132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [26]),
    .Y(_639_)
);

NAND2X1 _8133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_640_)
);

OAI21X1 _8134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_639_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_640_),
    .Y(_588_[26])
);

INVX1 _8135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [27]),
    .Y(_641_)
);

NAND2X1 _8136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_642_)
);

OAI21X1 _8137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_642_),
    .Y(_588_[27])
);

INVX1 _8138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [28]),
    .Y(_643_)
);

NAND2X1 _8139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_644_)
);

OAI21X1 _8140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf6 ),
    .C(_644_),
    .Y(_588_[28])
);

INVX1 _8141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [29]),
    .Y(_645_)
);

NAND2X1 _8142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_646_)
);

OAI21X1 _8143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf4 ),
    .C(_646_),
    .Y(_588_[29])
);

INVX1 _8144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [30]),
    .Y(_647_)
);

NAND2X1 _8145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_648_)
);

OAI21X1 _8146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_647_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf2 ),
    .C(_648_),
    .Y(_588_[30])
);

INVX1 _8147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[10] [31]),
    .Y(_649_)
);

NAND2X1 _8148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_10_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_650_)
);

OAI21X1 _8149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(\datapath_1.regfile_1.regEn_10_bF$buf0 ),
    .C(_650_),
    .Y(_588_[31])
);

DFFSR _8150_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_588_[0]),
    .Q(\datapath_1.regfile_1.regOut[10] [0]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _8151_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_588_[1]),
    .Q(\datapath_1.regfile_1.regOut[10] [1]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _8152_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_588_[2]),
    .Q(\datapath_1.regfile_1.regOut[10] [2]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _8153_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_588_[3]),
    .Q(\datapath_1.regfile_1.regOut[10] [3]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _8154_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_588_[4]),
    .Q(\datapath_1.regfile_1.regOut[10] [4]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _8155_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_588_[5]),
    .Q(\datapath_1.regfile_1.regOut[10] [5]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _8156_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_588_[6]),
    .Q(\datapath_1.regfile_1.regOut[10] [6]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _8157_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_588_[7]),
    .Q(\datapath_1.regfile_1.regOut[10] [7]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _8158_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_588_[8]),
    .Q(\datapath_1.regfile_1.regOut[10] [8]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _8159_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_588_[9]),
    .Q(\datapath_1.regfile_1.regOut[10] [9]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _8160_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_588_[10]),
    .Q(\datapath_1.regfile_1.regOut[10] [10]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _8161_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_588_[11]),
    .Q(\datapath_1.regfile_1.regOut[10] [11]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _8162_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_588_[12]),
    .Q(\datapath_1.regfile_1.regOut[10] [12]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _8163_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_588_[13]),
    .Q(\datapath_1.regfile_1.regOut[10] [13]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _8164_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_588_[14]),
    .Q(\datapath_1.regfile_1.regOut[10] [14]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _8165_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_588_[15]),
    .Q(\datapath_1.regfile_1.regOut[10] [15]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _8166_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_588_[16]),
    .Q(\datapath_1.regfile_1.regOut[10] [16]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _8167_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_588_[17]),
    .Q(\datapath_1.regfile_1.regOut[10] [17]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _8168_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_588_[18]),
    .Q(\datapath_1.regfile_1.regOut[10] [18]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _8169_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_588_[19]),
    .Q(\datapath_1.regfile_1.regOut[10] [19]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _8170_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_588_[20]),
    .Q(\datapath_1.regfile_1.regOut[10] [20]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _8171_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_588_[21]),
    .Q(\datapath_1.regfile_1.regOut[10] [21]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _8172_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_588_[22]),
    .Q(\datapath_1.regfile_1.regOut[10] [22]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _8173_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_588_[23]),
    .Q(\datapath_1.regfile_1.regOut[10] [23]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _8174_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_588_[24]),
    .Q(\datapath_1.regfile_1.regOut[10] [24]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _8175_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_588_[25]),
    .Q(\datapath_1.regfile_1.regOut[10] [25]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _8176_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_588_[26]),
    .Q(\datapath_1.regfile_1.regOut[10] [26]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _8177_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_588_[27]),
    .Q(\datapath_1.regfile_1.regOut[10] [27]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _8178_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_588_[28]),
    .Q(\datapath_1.regfile_1.regOut[10] [28]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _8179_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_588_[29]),
    .Q(\datapath_1.regfile_1.regOut[10] [29]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _8180_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_588_[30]),
    .Q(\datapath_1.regfile_1.regOut[10] [30]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _8181_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_588_[31]),
    .Q(\datapath_1.regfile_1.regOut[10] [31]),
    .R(rst_bF$buf26),
    .S(vdd)
);

INVX1 _8182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [0]),
    .Y(_716_)
);

NAND2X1 _8183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .Y(_717_)
);

OAI21X1 _8184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_717_),
    .Y(_653_[0])
);

INVX1 _8185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [1]),
    .Y(_654_)
);

NAND2X1 _8186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_655_)
);

OAI21X1 _8187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_655_),
    .Y(_653_[1])
);

INVX1 _8188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [2]),
    .Y(_656_)
);

NAND2X1 _8189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_657_)
);

OAI21X1 _8190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_656_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_657_),
    .Y(_653_[2])
);

INVX1 _8191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [3]),
    .Y(_658_)
);

NAND2X1 _8192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_659_)
);

OAI21X1 _8193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_659_),
    .Y(_653_[3])
);

INVX1 _8194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [4]),
    .Y(_660_)
);

NAND2X1 _8195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_661_)
);

OAI21X1 _8196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_661_),
    .Y(_653_[4])
);

INVX1 _8197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [5]),
    .Y(_662_)
);

NAND2X1 _8198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_663_)
);

OAI21X1 _8199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_663_),
    .Y(_653_[5])
);

INVX1 _8200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [6]),
    .Y(_664_)
);

NAND2X1 _8201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_665_)
);

OAI21X1 _8202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_665_),
    .Y(_653_[6])
);

INVX1 _8203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [7]),
    .Y(_666_)
);

NAND2X1 _8204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_667_)
);

OAI21X1 _8205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_667_),
    .Y(_653_[7])
);

INVX1 _8206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [8]),
    .Y(_668_)
);

NAND2X1 _8207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_669_)
);

OAI21X1 _8208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_669_),
    .Y(_653_[8])
);

INVX1 _8209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [9]),
    .Y(_670_)
);

NAND2X1 _8210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_671_)
);

OAI21X1 _8211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_671_),
    .Y(_653_[9])
);

INVX1 _8212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [10]),
    .Y(_672_)
);

NAND2X1 _8213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_673_)
);

OAI21X1 _8214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_672_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_673_),
    .Y(_653_[10])
);

INVX1 _8215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [11]),
    .Y(_674_)
);

NAND2X1 _8216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_675_)
);

OAI21X1 _8217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_675_),
    .Y(_653_[11])
);

INVX1 _8218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [12]),
    .Y(_676_)
);

NAND2X1 _8219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_677_)
);

OAI21X1 _8220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_677_),
    .Y(_653_[12])
);

INVX1 _8221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [13]),
    .Y(_678_)
);

NAND2X1 _8222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_679_)
);

OAI21X1 _8223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_679_),
    .Y(_653_[13])
);

INVX1 _8224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [14]),
    .Y(_680_)
);

NAND2X1 _8225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_681_)
);

OAI21X1 _8226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_680_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_681_),
    .Y(_653_[14])
);

INVX1 _8227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [15]),
    .Y(_682_)
);

NAND2X1 _8228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_683_)
);

OAI21X1 _8229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_683_),
    .Y(_653_[15])
);

INVX1 _8230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [16]),
    .Y(_684_)
);

NAND2X1 _8231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_685_)
);

OAI21X1 _8232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_685_),
    .Y(_653_[16])
);

INVX1 _8233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [17]),
    .Y(_686_)
);

NAND2X1 _8234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_687_)
);

OAI21X1 _8235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_687_),
    .Y(_653_[17])
);

INVX1 _8236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [18]),
    .Y(_688_)
);

NAND2X1 _8237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_689_)
);

OAI21X1 _8238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_689_),
    .Y(_653_[18])
);

INVX1 _8239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [19]),
    .Y(_690_)
);

NAND2X1 _8240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_691_)
);

OAI21X1 _8241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_690_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_691_),
    .Y(_653_[19])
);

INVX1 _8242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [20]),
    .Y(_692_)
);

NAND2X1 _8243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_693_)
);

OAI21X1 _8244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_693_),
    .Y(_653_[20])
);

INVX1 _8245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [21]),
    .Y(_694_)
);

NAND2X1 _8246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_695_)
);

OAI21X1 _8247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_694_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_695_),
    .Y(_653_[21])
);

INVX1 _8248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [22]),
    .Y(_696_)
);

NAND2X1 _8249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_697_)
);

OAI21X1 _8250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_697_),
    .Y(_653_[22])
);

INVX1 _8251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [23]),
    .Y(_698_)
);

NAND2X1 _8252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_699_)
);

OAI21X1 _8253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_699_),
    .Y(_653_[23])
);

INVX1 _8254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [24]),
    .Y(_700_)
);

NAND2X1 _8255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_701_)
);

OAI21X1 _8256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_701_),
    .Y(_653_[24])
);

INVX1 _8257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [25]),
    .Y(_702_)
);

NAND2X1 _8258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_703_)
);

OAI21X1 _8259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_703_),
    .Y(_653_[25])
);

INVX1 _8260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [26]),
    .Y(_704_)
);

NAND2X1 _8261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_705_)
);

OAI21X1 _8262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_704_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_705_),
    .Y(_653_[26])
);

INVX1 _8263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [27]),
    .Y(_706_)
);

NAND2X1 _8264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_707_)
);

OAI21X1 _8265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_706_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_707_),
    .Y(_653_[27])
);

INVX1 _8266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [28]),
    .Y(_708_)
);

NAND2X1 _8267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_709_)
);

OAI21X1 _8268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf6 ),
    .C(_709_),
    .Y(_653_[28])
);

INVX1 _8269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [29]),
    .Y(_710_)
);

NAND2X1 _8270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_711_)
);

OAI21X1 _8271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf4 ),
    .C(_711_),
    .Y(_653_[29])
);

INVX1 _8272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [30]),
    .Y(_712_)
);

NAND2X1 _8273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_713_)
);

OAI21X1 _8274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf2 ),
    .C(_713_),
    .Y(_653_[30])
);

INVX1 _8275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[11] [31]),
    .Y(_714_)
);

NAND2X1 _8276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_11_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_715_)
);

OAI21X1 _8277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(\datapath_1.regfile_1.regEn_11_bF$buf0 ),
    .C(_715_),
    .Y(_653_[31])
);

DFFSR _8278_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_653_[0]),
    .Q(\datapath_1.regfile_1.regOut[11] [0]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _8279_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_653_[1]),
    .Q(\datapath_1.regfile_1.regOut[11] [1]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _8280_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_653_[2]),
    .Q(\datapath_1.regfile_1.regOut[11] [2]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _8281_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_653_[3]),
    .Q(\datapath_1.regfile_1.regOut[11] [3]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _8282_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_653_[4]),
    .Q(\datapath_1.regfile_1.regOut[11] [4]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _8283_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_653_[5]),
    .Q(\datapath_1.regfile_1.regOut[11] [5]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _8284_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_653_[6]),
    .Q(\datapath_1.regfile_1.regOut[11] [6]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _8285_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_653_[7]),
    .Q(\datapath_1.regfile_1.regOut[11] [7]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _8286_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_653_[8]),
    .Q(\datapath_1.regfile_1.regOut[11] [8]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _8287_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_653_[9]),
    .Q(\datapath_1.regfile_1.regOut[11] [9]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _8288_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_653_[10]),
    .Q(\datapath_1.regfile_1.regOut[11] [10]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _8289_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_653_[11]),
    .Q(\datapath_1.regfile_1.regOut[11] [11]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _8290_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_653_[12]),
    .Q(\datapath_1.regfile_1.regOut[11] [12]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _8291_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_653_[13]),
    .Q(\datapath_1.regfile_1.regOut[11] [13]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _8292_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_653_[14]),
    .Q(\datapath_1.regfile_1.regOut[11] [14]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _8293_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_653_[15]),
    .Q(\datapath_1.regfile_1.regOut[11] [15]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _8294_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_653_[16]),
    .Q(\datapath_1.regfile_1.regOut[11] [16]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _8295_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_653_[17]),
    .Q(\datapath_1.regfile_1.regOut[11] [17]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _8296_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_653_[18]),
    .Q(\datapath_1.regfile_1.regOut[11] [18]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _8297_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_653_[19]),
    .Q(\datapath_1.regfile_1.regOut[11] [19]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _8298_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_653_[20]),
    .Q(\datapath_1.regfile_1.regOut[11] [20]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _8299_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_653_[21]),
    .Q(\datapath_1.regfile_1.regOut[11] [21]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _8300_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_653_[22]),
    .Q(\datapath_1.regfile_1.regOut[11] [22]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _8301_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_653_[23]),
    .Q(\datapath_1.regfile_1.regOut[11] [23]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _8302_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_653_[24]),
    .Q(\datapath_1.regfile_1.regOut[11] [24]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _8303_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_653_[25]),
    .Q(\datapath_1.regfile_1.regOut[11] [25]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _8304_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_653_[26]),
    .Q(\datapath_1.regfile_1.regOut[11] [26]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _8305_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_653_[27]),
    .Q(\datapath_1.regfile_1.regOut[11] [27]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _8306_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_653_[28]),
    .Q(\datapath_1.regfile_1.regOut[11] [28]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _8307_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_653_[29]),
    .Q(\datapath_1.regfile_1.regOut[11] [29]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _8308_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_653_[30]),
    .Q(\datapath_1.regfile_1.regOut[11] [30]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _8309_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_653_[31]),
    .Q(\datapath_1.regfile_1.regOut[11] [31]),
    .R(rst_bF$buf108),
    .S(vdd)
);

INVX1 _8310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [0]),
    .Y(_781_)
);

NAND2X1 _8311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .Y(_782_)
);

OAI21X1 _8312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_782_),
    .Y(_718_[0])
);

INVX1 _8313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [1]),
    .Y(_719_)
);

NAND2X1 _8314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_720_)
);

OAI21X1 _8315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_720_),
    .Y(_718_[1])
);

INVX1 _8316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [2]),
    .Y(_721_)
);

NAND2X1 _8317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_722_)
);

OAI21X1 _8318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_722_),
    .Y(_718_[2])
);

INVX1 _8319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [3]),
    .Y(_723_)
);

NAND2X1 _8320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_724_)
);

OAI21X1 _8321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_724_),
    .Y(_718_[3])
);

INVX1 _8322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [4]),
    .Y(_725_)
);

NAND2X1 _8323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_726_)
);

OAI21X1 _8324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_726_),
    .Y(_718_[4])
);

INVX1 _8325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [5]),
    .Y(_727_)
);

NAND2X1 _8326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_728_)
);

OAI21X1 _8327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_728_),
    .Y(_718_[5])
);

INVX1 _8328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [6]),
    .Y(_729_)
);

NAND2X1 _8329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_730_)
);

OAI21X1 _8330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_730_),
    .Y(_718_[6])
);

INVX1 _8331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [7]),
    .Y(_731_)
);

NAND2X1 _8332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_732_)
);

OAI21X1 _8333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_732_),
    .Y(_718_[7])
);

INVX1 _8334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [8]),
    .Y(_733_)
);

NAND2X1 _8335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_734_)
);

OAI21X1 _8336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_734_),
    .Y(_718_[8])
);

INVX1 _8337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [9]),
    .Y(_735_)
);

NAND2X1 _8338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_736_)
);

OAI21X1 _8339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_735_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_736_),
    .Y(_718_[9])
);

INVX1 _8340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [10]),
    .Y(_737_)
);

NAND2X1 _8341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_738_)
);

OAI21X1 _8342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_737_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_738_),
    .Y(_718_[10])
);

INVX1 _8343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [11]),
    .Y(_739_)
);

NAND2X1 _8344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_740_)
);

OAI21X1 _8345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_740_),
    .Y(_718_[11])
);

INVX1 _8346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [12]),
    .Y(_741_)
);

NAND2X1 _8347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_742_)
);

OAI21X1 _8348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_741_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_742_),
    .Y(_718_[12])
);

INVX1 _8349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [13]),
    .Y(_743_)
);

NAND2X1 _8350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_744_)
);

OAI21X1 _8351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_744_),
    .Y(_718_[13])
);

INVX1 _8352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [14]),
    .Y(_745_)
);

NAND2X1 _8353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_746_)
);

OAI21X1 _8354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_746_),
    .Y(_718_[14])
);

INVX1 _8355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [15]),
    .Y(_747_)
);

NAND2X1 _8356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_748_)
);

OAI21X1 _8357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_748_),
    .Y(_718_[15])
);

INVX1 _8358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [16]),
    .Y(_749_)
);

NAND2X1 _8359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_750_)
);

OAI21X1 _8360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_750_),
    .Y(_718_[16])
);

INVX1 _8361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [17]),
    .Y(_751_)
);

NAND2X1 _8362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_752_)
);

OAI21X1 _8363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_752_),
    .Y(_718_[17])
);

INVX1 _8364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [18]),
    .Y(_753_)
);

NAND2X1 _8365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_754_)
);

OAI21X1 _8366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_754_),
    .Y(_718_[18])
);

INVX1 _8367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [19]),
    .Y(_755_)
);

NAND2X1 _8368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_756_)
);

OAI21X1 _8369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_756_),
    .Y(_718_[19])
);

INVX1 _8370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [20]),
    .Y(_757_)
);

NAND2X1 _8371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_758_)
);

OAI21X1 _8372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_757_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_758_),
    .Y(_718_[20])
);

INVX1 _8373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [21]),
    .Y(_759_)
);

NAND2X1 _8374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_760_)
);

OAI21X1 _8375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_760_),
    .Y(_718_[21])
);

INVX1 _8376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [22]),
    .Y(_761_)
);

NAND2X1 _8377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_762_)
);

OAI21X1 _8378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_761_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_762_),
    .Y(_718_[22])
);

INVX1 _8379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [23]),
    .Y(_763_)
);

NAND2X1 _8380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_764_)
);

OAI21X1 _8381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_764_),
    .Y(_718_[23])
);

INVX1 _8382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [24]),
    .Y(_765_)
);

NAND2X1 _8383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_766_)
);

OAI21X1 _8384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_766_),
    .Y(_718_[24])
);

INVX1 _8385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [25]),
    .Y(_767_)
);

NAND2X1 _8386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_768_)
);

OAI21X1 _8387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_767_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_768_),
    .Y(_718_[25])
);

INVX1 _8388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [26]),
    .Y(_769_)
);

NAND2X1 _8389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_770_)
);

OAI21X1 _8390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_770_),
    .Y(_718_[26])
);

INVX1 _8391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [27]),
    .Y(_771_)
);

NAND2X1 _8392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_772_)
);

OAI21X1 _8393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_772_),
    .Y(_718_[27])
);

INVX1 _8394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [28]),
    .Y(_773_)
);

NAND2X1 _8395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_774_)
);

OAI21X1 _8396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf6 ),
    .C(_774_),
    .Y(_718_[28])
);

INVX1 _8397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [29]),
    .Y(_775_)
);

NAND2X1 _8398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_776_)
);

OAI21X1 _8399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf4 ),
    .C(_776_),
    .Y(_718_[29])
);

INVX1 _8400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [30]),
    .Y(_777_)
);

NAND2X1 _8401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_778_)
);

OAI21X1 _8402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf2 ),
    .C(_778_),
    .Y(_718_[30])
);

INVX1 _8403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[12] [31]),
    .Y(_779_)
);

NAND2X1 _8404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_12_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_780_)
);

OAI21X1 _8405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(\datapath_1.regfile_1.regEn_12_bF$buf0 ),
    .C(_780_),
    .Y(_718_[31])
);

DFFSR _8406_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_718_[0]),
    .Q(\datapath_1.regfile_1.regOut[12] [0]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _8407_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_718_[1]),
    .Q(\datapath_1.regfile_1.regOut[12] [1]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _8408_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_718_[2]),
    .Q(\datapath_1.regfile_1.regOut[12] [2]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _8409_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_718_[3]),
    .Q(\datapath_1.regfile_1.regOut[12] [3]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _8410_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_718_[4]),
    .Q(\datapath_1.regfile_1.regOut[12] [4]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _8411_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_718_[5]),
    .Q(\datapath_1.regfile_1.regOut[12] [5]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _8412_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_718_[6]),
    .Q(\datapath_1.regfile_1.regOut[12] [6]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _8413_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_718_[7]),
    .Q(\datapath_1.regfile_1.regOut[12] [7]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _8414_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_718_[8]),
    .Q(\datapath_1.regfile_1.regOut[12] [8]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _8415_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_718_[9]),
    .Q(\datapath_1.regfile_1.regOut[12] [9]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _8416_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_718_[10]),
    .Q(\datapath_1.regfile_1.regOut[12] [10]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _8417_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_718_[11]),
    .Q(\datapath_1.regfile_1.regOut[12] [11]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _8418_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_718_[12]),
    .Q(\datapath_1.regfile_1.regOut[12] [12]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _8419_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_718_[13]),
    .Q(\datapath_1.regfile_1.regOut[12] [13]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _8420_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_718_[14]),
    .Q(\datapath_1.regfile_1.regOut[12] [14]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _8421_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_718_[15]),
    .Q(\datapath_1.regfile_1.regOut[12] [15]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _8422_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_718_[16]),
    .Q(\datapath_1.regfile_1.regOut[12] [16]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _8423_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_718_[17]),
    .Q(\datapath_1.regfile_1.regOut[12] [17]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _8424_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_718_[18]),
    .Q(\datapath_1.regfile_1.regOut[12] [18]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _8425_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_718_[19]),
    .Q(\datapath_1.regfile_1.regOut[12] [19]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _8426_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_718_[20]),
    .Q(\datapath_1.regfile_1.regOut[12] [20]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _8427_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_718_[21]),
    .Q(\datapath_1.regfile_1.regOut[12] [21]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _8428_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_718_[22]),
    .Q(\datapath_1.regfile_1.regOut[12] [22]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _8429_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_718_[23]),
    .Q(\datapath_1.regfile_1.regOut[12] [23]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _8430_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_718_[24]),
    .Q(\datapath_1.regfile_1.regOut[12] [24]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _8431_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_718_[25]),
    .Q(\datapath_1.regfile_1.regOut[12] [25]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _8432_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_718_[26]),
    .Q(\datapath_1.regfile_1.regOut[12] [26]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _8433_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_718_[27]),
    .Q(\datapath_1.regfile_1.regOut[12] [27]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _8434_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_718_[28]),
    .Q(\datapath_1.regfile_1.regOut[12] [28]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _8435_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_718_[29]),
    .Q(\datapath_1.regfile_1.regOut[12] [29]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _8436_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_718_[30]),
    .Q(\datapath_1.regfile_1.regOut[12] [30]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _8437_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_718_[31]),
    .Q(\datapath_1.regfile_1.regOut[12] [31]),
    .R(rst_bF$buf76),
    .S(vdd)
);

INVX1 _8438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [0]),
    .Y(_846_)
);

NAND2X1 _8439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .Y(_847_)
);

OAI21X1 _8440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_847_),
    .Y(_783_[0])
);

INVX1 _8441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [1]),
    .Y(_784_)
);

NAND2X1 _8442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_785_)
);

OAI21X1 _8443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_785_),
    .Y(_783_[1])
);

INVX1 _8444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [2]),
    .Y(_786_)
);

NAND2X1 _8445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_787_)
);

OAI21X1 _8446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_787_),
    .Y(_783_[2])
);

INVX1 _8447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [3]),
    .Y(_788_)
);

NAND2X1 _8448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_789_)
);

OAI21X1 _8449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_789_),
    .Y(_783_[3])
);

INVX1 _8450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [4]),
    .Y(_790_)
);

NAND2X1 _8451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_791_)
);

OAI21X1 _8452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_791_),
    .Y(_783_[4])
);

INVX1 _8453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [5]),
    .Y(_792_)
);

NAND2X1 _8454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_793_)
);

OAI21X1 _8455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_793_),
    .Y(_783_[5])
);

INVX1 _8456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [6]),
    .Y(_794_)
);

NAND2X1 _8457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_795_)
);

OAI21X1 _8458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_794_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_795_),
    .Y(_783_[6])
);

INVX1 _8459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [7]),
    .Y(_796_)
);

NAND2X1 _8460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_797_)
);

OAI21X1 _8461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_797_),
    .Y(_783_[7])
);

INVX1 _8462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [8]),
    .Y(_798_)
);

NAND2X1 _8463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_799_)
);

OAI21X1 _8464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_799_),
    .Y(_783_[8])
);

INVX1 _8465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [9]),
    .Y(_800_)
);

NAND2X1 _8466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_801_)
);

OAI21X1 _8467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_801_),
    .Y(_783_[9])
);

INVX1 _8468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [10]),
    .Y(_802_)
);

NAND2X1 _8469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_803_)
);

OAI21X1 _8470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_803_),
    .Y(_783_[10])
);

INVX1 _8471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [11]),
    .Y(_804_)
);

NAND2X1 _8472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_805_)
);

OAI21X1 _8473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_804_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_805_),
    .Y(_783_[11])
);

INVX1 _8474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [12]),
    .Y(_806_)
);

NAND2X1 _8475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_807_)
);

OAI21X1 _8476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_807_),
    .Y(_783_[12])
);

INVX1 _8477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [13]),
    .Y(_808_)
);

NAND2X1 _8478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_809_)
);

OAI21X1 _8479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_808_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_809_),
    .Y(_783_[13])
);

INVX1 _8480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [14]),
    .Y(_810_)
);

NAND2X1 _8481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_811_)
);

OAI21X1 _8482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_810_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_811_),
    .Y(_783_[14])
);

INVX1 _8483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [15]),
    .Y(_812_)
);

NAND2X1 _8484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_813_)
);

OAI21X1 _8485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_812_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_813_),
    .Y(_783_[15])
);

INVX1 _8486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [16]),
    .Y(_814_)
);

NAND2X1 _8487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_815_)
);

OAI21X1 _8488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_815_),
    .Y(_783_[16])
);

INVX1 _8489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [17]),
    .Y(_816_)
);

NAND2X1 _8490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_817_)
);

OAI21X1 _8491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_817_),
    .Y(_783_[17])
);

INVX1 _8492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [18]),
    .Y(_818_)
);

NAND2X1 _8493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_819_)
);

OAI21X1 _8494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_819_),
    .Y(_783_[18])
);

INVX1 _8495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [19]),
    .Y(_820_)
);

NAND2X1 _8496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_821_)
);

OAI21X1 _8497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_821_),
    .Y(_783_[19])
);

INVX1 _8498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [20]),
    .Y(_822_)
);

NAND2X1 _8499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_823_)
);

OAI21X1 _8500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_822_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_823_),
    .Y(_783_[20])
);

INVX1 _8501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [21]),
    .Y(_824_)
);

NAND2X1 _8502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_825_)
);

OAI21X1 _8503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_824_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_825_),
    .Y(_783_[21])
);

INVX1 _8504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [22]),
    .Y(_826_)
);

NAND2X1 _8505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_827_)
);

OAI21X1 _8506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_826_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_827_),
    .Y(_783_[22])
);

INVX1 _8507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [23]),
    .Y(_828_)
);

NAND2X1 _8508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_829_)
);

OAI21X1 _8509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_829_),
    .Y(_783_[23])
);

INVX1 _8510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [24]),
    .Y(_830_)
);

NAND2X1 _8511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_831_)
);

OAI21X1 _8512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_831_),
    .Y(_783_[24])
);

INVX1 _8513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [25]),
    .Y(_832_)
);

NAND2X1 _8514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_833_)
);

OAI21X1 _8515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_833_),
    .Y(_783_[25])
);

INVX1 _8516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [26]),
    .Y(_834_)
);

NAND2X1 _8517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_835_)
);

OAI21X1 _8518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_834_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_835_),
    .Y(_783_[26])
);

INVX1 _8519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [27]),
    .Y(_836_)
);

NAND2X1 _8520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_837_)
);

OAI21X1 _8521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_837_),
    .Y(_783_[27])
);

INVX1 _8522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [28]),
    .Y(_838_)
);

NAND2X1 _8523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_839_)
);

OAI21X1 _8524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_838_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf6 ),
    .C(_839_),
    .Y(_783_[28])
);

INVX1 _8525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [29]),
    .Y(_840_)
);

NAND2X1 _8526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_841_)
);

OAI21X1 _8527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf4 ),
    .C(_841_),
    .Y(_783_[29])
);

INVX1 _8528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [30]),
    .Y(_842_)
);

NAND2X1 _8529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_843_)
);

OAI21X1 _8530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf2 ),
    .C(_843_),
    .Y(_783_[30])
);

INVX1 _8531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[13] [31]),
    .Y(_844_)
);

NAND2X1 _8532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_13_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_845_)
);

OAI21X1 _8533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(\datapath_1.regfile_1.regEn_13_bF$buf0 ),
    .C(_845_),
    .Y(_783_[31])
);

DFFSR _8534_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_783_[0]),
    .Q(\datapath_1.regfile_1.regOut[13] [0]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _8535_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_783_[1]),
    .Q(\datapath_1.regfile_1.regOut[13] [1]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _8536_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_783_[2]),
    .Q(\datapath_1.regfile_1.regOut[13] [2]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _8537_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_783_[3]),
    .Q(\datapath_1.regfile_1.regOut[13] [3]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _8538_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_783_[4]),
    .Q(\datapath_1.regfile_1.regOut[13] [4]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _8539_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_783_[5]),
    .Q(\datapath_1.regfile_1.regOut[13] [5]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _8540_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_783_[6]),
    .Q(\datapath_1.regfile_1.regOut[13] [6]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _8541_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_783_[7]),
    .Q(\datapath_1.regfile_1.regOut[13] [7]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _8542_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_783_[8]),
    .Q(\datapath_1.regfile_1.regOut[13] [8]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _8543_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_783_[9]),
    .Q(\datapath_1.regfile_1.regOut[13] [9]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _8544_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_783_[10]),
    .Q(\datapath_1.regfile_1.regOut[13] [10]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _8545_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_783_[11]),
    .Q(\datapath_1.regfile_1.regOut[13] [11]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _8546_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_783_[12]),
    .Q(\datapath_1.regfile_1.regOut[13] [12]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _8547_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_783_[13]),
    .Q(\datapath_1.regfile_1.regOut[13] [13]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _8548_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_783_[14]),
    .Q(\datapath_1.regfile_1.regOut[13] [14]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _8549_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_783_[15]),
    .Q(\datapath_1.regfile_1.regOut[13] [15]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _8550_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_783_[16]),
    .Q(\datapath_1.regfile_1.regOut[13] [16]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _8551_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_783_[17]),
    .Q(\datapath_1.regfile_1.regOut[13] [17]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _8552_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_783_[18]),
    .Q(\datapath_1.regfile_1.regOut[13] [18]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _8553_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_783_[19]),
    .Q(\datapath_1.regfile_1.regOut[13] [19]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _8554_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_783_[20]),
    .Q(\datapath_1.regfile_1.regOut[13] [20]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _8555_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_783_[21]),
    .Q(\datapath_1.regfile_1.regOut[13] [21]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _8556_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_783_[22]),
    .Q(\datapath_1.regfile_1.regOut[13] [22]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _8557_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_783_[23]),
    .Q(\datapath_1.regfile_1.regOut[13] [23]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _8558_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_783_[24]),
    .Q(\datapath_1.regfile_1.regOut[13] [24]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _8559_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_783_[25]),
    .Q(\datapath_1.regfile_1.regOut[13] [25]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _8560_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_783_[26]),
    .Q(\datapath_1.regfile_1.regOut[13] [26]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _8561_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_783_[27]),
    .Q(\datapath_1.regfile_1.regOut[13] [27]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _8562_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_783_[28]),
    .Q(\datapath_1.regfile_1.regOut[13] [28]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _8563_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_783_[29]),
    .Q(\datapath_1.regfile_1.regOut[13] [29]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _8564_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_783_[30]),
    .Q(\datapath_1.regfile_1.regOut[13] [30]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _8565_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_783_[31]),
    .Q(\datapath_1.regfile_1.regOut[13] [31]),
    .R(rst_bF$buf44),
    .S(vdd)
);

INVX1 _8566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [0]),
    .Y(_911_)
);

NAND2X1 _8567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .Y(_912_)
);

OAI21X1 _8568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_911_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_912_),
    .Y(_848_[0])
);

INVX1 _8569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [1]),
    .Y(_849_)
);

NAND2X1 _8570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_850_)
);

OAI21X1 _8571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_849_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_850_),
    .Y(_848_[1])
);

INVX1 _8572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [2]),
    .Y(_851_)
);

NAND2X1 _8573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_852_)
);

OAI21X1 _8574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_851_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_852_),
    .Y(_848_[2])
);

INVX1 _8575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [3]),
    .Y(_853_)
);

NAND2X1 _8576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_854_)
);

OAI21X1 _8577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_854_),
    .Y(_848_[3])
);

INVX1 _8578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [4]),
    .Y(_855_)
);

NAND2X1 _8579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_856_)
);

OAI21X1 _8580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_856_),
    .Y(_848_[4])
);

INVX1 _8581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [5]),
    .Y(_857_)
);

NAND2X1 _8582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_858_)
);

OAI21X1 _8583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_858_),
    .Y(_848_[5])
);

INVX1 _8584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [6]),
    .Y(_859_)
);

NAND2X1 _8585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_860_)
);

OAI21X1 _8586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_860_),
    .Y(_848_[6])
);

INVX1 _8587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [7]),
    .Y(_861_)
);

NAND2X1 _8588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_862_)
);

OAI21X1 _8589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_862_),
    .Y(_848_[7])
);

INVX1 _8590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [8]),
    .Y(_863_)
);

NAND2X1 _8591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_864_)
);

OAI21X1 _8592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_864_),
    .Y(_848_[8])
);

INVX1 _8593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [9]),
    .Y(_865_)
);

NAND2X1 _8594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_866_)
);

OAI21X1 _8595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_865_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_866_),
    .Y(_848_[9])
);

INVX1 _8596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [10]),
    .Y(_867_)
);

NAND2X1 _8597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_868_)
);

OAI21X1 _8598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_868_),
    .Y(_848_[10])
);

INVX1 _8599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [11]),
    .Y(_869_)
);

NAND2X1 _8600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_870_)
);

OAI21X1 _8601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_870_),
    .Y(_848_[11])
);

INVX1 _8602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [12]),
    .Y(_871_)
);

NAND2X1 _8603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_872_)
);

OAI21X1 _8604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_871_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_872_),
    .Y(_848_[12])
);

INVX1 _8605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [13]),
    .Y(_873_)
);

NAND2X1 _8606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_874_)
);

OAI21X1 _8607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_874_),
    .Y(_848_[13])
);

INVX1 _8608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [14]),
    .Y(_875_)
);

NAND2X1 _8609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_876_)
);

OAI21X1 _8610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_876_),
    .Y(_848_[14])
);

INVX1 _8611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [15]),
    .Y(_877_)
);

NAND2X1 _8612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_878_)
);

OAI21X1 _8613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_878_),
    .Y(_848_[15])
);

INVX1 _8614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [16]),
    .Y(_879_)
);

NAND2X1 _8615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_880_)
);

OAI21X1 _8616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_880_),
    .Y(_848_[16])
);

INVX1 _8617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [17]),
    .Y(_881_)
);

NAND2X1 _8618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_882_)
);

OAI21X1 _8619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_882_),
    .Y(_848_[17])
);

INVX1 _8620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [18]),
    .Y(_883_)
);

NAND2X1 _8621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_884_)
);

OAI21X1 _8622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_883_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_884_),
    .Y(_848_[18])
);

INVX1 _8623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [19]),
    .Y(_885_)
);

NAND2X1 _8624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_886_)
);

OAI21X1 _8625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_885_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_886_),
    .Y(_848_[19])
);

INVX1 _8626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [20]),
    .Y(_887_)
);

NAND2X1 _8627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_888_)
);

OAI21X1 _8628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_888_),
    .Y(_848_[20])
);

INVX1 _8629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [21]),
    .Y(_889_)
);

NAND2X1 _8630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_890_)
);

OAI21X1 _8631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_889_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_890_),
    .Y(_848_[21])
);

INVX1 _8632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [22]),
    .Y(_891_)
);

NAND2X1 _8633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_892_)
);

OAI21X1 _8634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_891_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_892_),
    .Y(_848_[22])
);

INVX1 _8635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [23]),
    .Y(_893_)
);

NAND2X1 _8636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_894_)
);

OAI21X1 _8637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_893_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_894_),
    .Y(_848_[23])
);

INVX1 _8638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [24]),
    .Y(_895_)
);

NAND2X1 _8639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_896_)
);

OAI21X1 _8640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_896_),
    .Y(_848_[24])
);

INVX1 _8641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [25]),
    .Y(_897_)
);

NAND2X1 _8642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_898_)
);

OAI21X1 _8643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_897_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_898_),
    .Y(_848_[25])
);

INVX1 _8644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [26]),
    .Y(_899_)
);

NAND2X1 _8645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_900_)
);

OAI21X1 _8646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_899_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_900_),
    .Y(_848_[26])
);

INVX1 _8647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [27]),
    .Y(_901_)
);

NAND2X1 _8648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_902_)
);

OAI21X1 _8649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_902_),
    .Y(_848_[27])
);

INVX1 _8650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [28]),
    .Y(_903_)
);

NAND2X1 _8651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_904_)
);

OAI21X1 _8652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_903_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf6 ),
    .C(_904_),
    .Y(_848_[28])
);

INVX1 _8653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [29]),
    .Y(_905_)
);

NAND2X1 _8654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_906_)
);

OAI21X1 _8655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf4 ),
    .C(_906_),
    .Y(_848_[29])
);

INVX1 _8656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [30]),
    .Y(_907_)
);

NAND2X1 _8657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_908_)
);

OAI21X1 _8658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf2 ),
    .C(_908_),
    .Y(_848_[30])
);

INVX1 _8659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[14] [31]),
    .Y(_909_)
);

NAND2X1 _8660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_14_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_910_)
);

OAI21X1 _8661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .B(\datapath_1.regfile_1.regEn_14_bF$buf0 ),
    .C(_910_),
    .Y(_848_[31])
);

DFFSR _8662_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_848_[0]),
    .Q(\datapath_1.regfile_1.regOut[14] [0]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _8663_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_848_[1]),
    .Q(\datapath_1.regfile_1.regOut[14] [1]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _8664_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_848_[2]),
    .Q(\datapath_1.regfile_1.regOut[14] [2]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _8665_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_848_[3]),
    .Q(\datapath_1.regfile_1.regOut[14] [3]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _8666_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_848_[4]),
    .Q(\datapath_1.regfile_1.regOut[14] [4]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _8667_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_848_[5]),
    .Q(\datapath_1.regfile_1.regOut[14] [5]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _8668_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_848_[6]),
    .Q(\datapath_1.regfile_1.regOut[14] [6]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _8669_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_848_[7]),
    .Q(\datapath_1.regfile_1.regOut[14] [7]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _8670_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_848_[8]),
    .Q(\datapath_1.regfile_1.regOut[14] [8]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _8671_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_848_[9]),
    .Q(\datapath_1.regfile_1.regOut[14] [9]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _8672_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_848_[10]),
    .Q(\datapath_1.regfile_1.regOut[14] [10]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _8673_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_848_[11]),
    .Q(\datapath_1.regfile_1.regOut[14] [11]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _8674_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_848_[12]),
    .Q(\datapath_1.regfile_1.regOut[14] [12]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _8675_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_848_[13]),
    .Q(\datapath_1.regfile_1.regOut[14] [13]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _8676_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_848_[14]),
    .Q(\datapath_1.regfile_1.regOut[14] [14]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _8677_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_848_[15]),
    .Q(\datapath_1.regfile_1.regOut[14] [15]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _8678_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_848_[16]),
    .Q(\datapath_1.regfile_1.regOut[14] [16]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _8679_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_848_[17]),
    .Q(\datapath_1.regfile_1.regOut[14] [17]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _8680_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_848_[18]),
    .Q(\datapath_1.regfile_1.regOut[14] [18]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _8681_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_848_[19]),
    .Q(\datapath_1.regfile_1.regOut[14] [19]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _8682_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_848_[20]),
    .Q(\datapath_1.regfile_1.regOut[14] [20]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _8683_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_848_[21]),
    .Q(\datapath_1.regfile_1.regOut[14] [21]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _8684_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_848_[22]),
    .Q(\datapath_1.regfile_1.regOut[14] [22]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _8685_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_848_[23]),
    .Q(\datapath_1.regfile_1.regOut[14] [23]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _8686_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_848_[24]),
    .Q(\datapath_1.regfile_1.regOut[14] [24]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _8687_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_848_[25]),
    .Q(\datapath_1.regfile_1.regOut[14] [25]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _8688_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_848_[26]),
    .Q(\datapath_1.regfile_1.regOut[14] [26]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _8689_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_848_[27]),
    .Q(\datapath_1.regfile_1.regOut[14] [27]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _8690_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_848_[28]),
    .Q(\datapath_1.regfile_1.regOut[14] [28]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _8691_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_848_[29]),
    .Q(\datapath_1.regfile_1.regOut[14] [29]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _8692_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_848_[30]),
    .Q(\datapath_1.regfile_1.regOut[14] [30]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _8693_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_848_[31]),
    .Q(\datapath_1.regfile_1.regOut[14] [31]),
    .R(rst_bF$buf12),
    .S(vdd)
);

INVX1 _8694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [0]),
    .Y(_976_)
);

NAND2X1 _8695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .Y(_977_)
);

OAI21X1 _8696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_977_),
    .Y(_913_[0])
);

INVX1 _8697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [1]),
    .Y(_914_)
);

NAND2X1 _8698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_915_)
);

OAI21X1 _8699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_915_),
    .Y(_913_[1])
);

INVX1 _8700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [2]),
    .Y(_916_)
);

NAND2X1 _8701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_917_)
);

OAI21X1 _8702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_917_),
    .Y(_913_[2])
);

INVX1 _8703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [3]),
    .Y(_918_)
);

NAND2X1 _8704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_919_)
);

OAI21X1 _8705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_919_),
    .Y(_913_[3])
);

INVX1 _8706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [4]),
    .Y(_920_)
);

NAND2X1 _8707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_921_)
);

OAI21X1 _8708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_921_),
    .Y(_913_[4])
);

INVX1 _8709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [5]),
    .Y(_922_)
);

NAND2X1 _8710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_923_)
);

OAI21X1 _8711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_922_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_923_),
    .Y(_913_[5])
);

INVX1 _8712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [6]),
    .Y(_924_)
);

NAND2X1 _8713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_925_)
);

OAI21X1 _8714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_924_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_925_),
    .Y(_913_[6])
);

INVX1 _8715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [7]),
    .Y(_926_)
);

NAND2X1 _8716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_927_)
);

OAI21X1 _8717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_927_),
    .Y(_913_[7])
);

INVX1 _8718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [8]),
    .Y(_928_)
);

NAND2X1 _8719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_929_)
);

OAI21X1 _8720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_928_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_929_),
    .Y(_913_[8])
);

INVX1 _8721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [9]),
    .Y(_930_)
);

NAND2X1 _8722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_931_)
);

OAI21X1 _8723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_930_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_931_),
    .Y(_913_[9])
);

INVX1 _8724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [10]),
    .Y(_932_)
);

NAND2X1 _8725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_933_)
);

OAI21X1 _8726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_933_),
    .Y(_913_[10])
);

INVX1 _8727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [11]),
    .Y(_934_)
);

NAND2X1 _8728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_935_)
);

OAI21X1 _8729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_935_),
    .Y(_913_[11])
);

INVX1 _8730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [12]),
    .Y(_936_)
);

NAND2X1 _8731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_937_)
);

OAI21X1 _8732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_936_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_937_),
    .Y(_913_[12])
);

INVX1 _8733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [13]),
    .Y(_938_)
);

NAND2X1 _8734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_939_)
);

OAI21X1 _8735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_938_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_939_),
    .Y(_913_[13])
);

INVX1 _8736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [14]),
    .Y(_940_)
);

NAND2X1 _8737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_941_)
);

OAI21X1 _8738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_940_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_941_),
    .Y(_913_[14])
);

INVX1 _8739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [15]),
    .Y(_942_)
);

NAND2X1 _8740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_943_)
);

OAI21X1 _8741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_943_),
    .Y(_913_[15])
);

INVX1 _8742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [16]),
    .Y(_944_)
);

NAND2X1 _8743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_945_)
);

OAI21X1 _8744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_944_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_945_),
    .Y(_913_[16])
);

INVX1 _8745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [17]),
    .Y(_946_)
);

NAND2X1 _8746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_947_)
);

OAI21X1 _8747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_946_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_947_),
    .Y(_913_[17])
);

INVX1 _8748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [18]),
    .Y(_948_)
);

NAND2X1 _8749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_949_)
);

OAI21X1 _8750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_948_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_949_),
    .Y(_913_[18])
);

INVX1 _8751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [19]),
    .Y(_950_)
);

NAND2X1 _8752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_951_)
);

OAI21X1 _8753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_951_),
    .Y(_913_[19])
);

INVX1 _8754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [20]),
    .Y(_952_)
);

NAND2X1 _8755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_953_)
);

OAI21X1 _8756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_952_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_953_),
    .Y(_913_[20])
);

INVX1 _8757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [21]),
    .Y(_954_)
);

NAND2X1 _8758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_955_)
);

OAI21X1 _8759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_954_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_955_),
    .Y(_913_[21])
);

INVX1 _8760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [22]),
    .Y(_956_)
);

NAND2X1 _8761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_957_)
);

OAI21X1 _8762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_957_),
    .Y(_913_[22])
);

INVX1 _8763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [23]),
    .Y(_958_)
);

NAND2X1 _8764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_959_)
);

OAI21X1 _8765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_958_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_959_),
    .Y(_913_[23])
);

INVX1 _8766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [24]),
    .Y(_960_)
);

NAND2X1 _8767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_961_)
);

OAI21X1 _8768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_960_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_961_),
    .Y(_913_[24])
);

INVX1 _8769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [25]),
    .Y(_962_)
);

NAND2X1 _8770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_963_)
);

OAI21X1 _8771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_963_),
    .Y(_913_[25])
);

INVX1 _8772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [26]),
    .Y(_964_)
);

NAND2X1 _8773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_965_)
);

OAI21X1 _8774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_965_),
    .Y(_913_[26])
);

INVX1 _8775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [27]),
    .Y(_966_)
);

NAND2X1 _8776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_967_)
);

OAI21X1 _8777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_966_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_967_),
    .Y(_913_[27])
);

INVX1 _8778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [28]),
    .Y(_968_)
);

NAND2X1 _8779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_969_)
);

OAI21X1 _8780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf6 ),
    .C(_969_),
    .Y(_913_[28])
);

INVX1 _8781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [29]),
    .Y(_970_)
);

NAND2X1 _8782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_971_)
);

OAI21X1 _8783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf4 ),
    .C(_971_),
    .Y(_913_[29])
);

INVX1 _8784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [30]),
    .Y(_972_)
);

NAND2X1 _8785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_973_)
);

OAI21X1 _8786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf2 ),
    .C(_973_),
    .Y(_913_[30])
);

INVX1 _8787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[15] [31]),
    .Y(_974_)
);

NAND2X1 _8788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_15_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_975_)
);

OAI21X1 _8789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(\datapath_1.regfile_1.regEn_15_bF$buf0 ),
    .C(_975_),
    .Y(_913_[31])
);

DFFSR _8790_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_913_[0]),
    .Q(\datapath_1.regfile_1.regOut[15] [0]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _8791_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_913_[1]),
    .Q(\datapath_1.regfile_1.regOut[15] [1]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _8792_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_913_[2]),
    .Q(\datapath_1.regfile_1.regOut[15] [2]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _8793_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_913_[3]),
    .Q(\datapath_1.regfile_1.regOut[15] [3]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _8794_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_913_[4]),
    .Q(\datapath_1.regfile_1.regOut[15] [4]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _8795_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_913_[5]),
    .Q(\datapath_1.regfile_1.regOut[15] [5]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _8796_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_913_[6]),
    .Q(\datapath_1.regfile_1.regOut[15] [6]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _8797_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_913_[7]),
    .Q(\datapath_1.regfile_1.regOut[15] [7]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _8798_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_913_[8]),
    .Q(\datapath_1.regfile_1.regOut[15] [8]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _8799_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_913_[9]),
    .Q(\datapath_1.regfile_1.regOut[15] [9]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _8800_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_913_[10]),
    .Q(\datapath_1.regfile_1.regOut[15] [10]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _8801_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_913_[11]),
    .Q(\datapath_1.regfile_1.regOut[15] [11]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _8802_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_913_[12]),
    .Q(\datapath_1.regfile_1.regOut[15] [12]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _8803_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_913_[13]),
    .Q(\datapath_1.regfile_1.regOut[15] [13]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _8804_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_913_[14]),
    .Q(\datapath_1.regfile_1.regOut[15] [14]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _8805_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_913_[15]),
    .Q(\datapath_1.regfile_1.regOut[15] [15]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _8806_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_913_[16]),
    .Q(\datapath_1.regfile_1.regOut[15] [16]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _8807_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_913_[17]),
    .Q(\datapath_1.regfile_1.regOut[15] [17]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _8808_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_913_[18]),
    .Q(\datapath_1.regfile_1.regOut[15] [18]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _8809_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_913_[19]),
    .Q(\datapath_1.regfile_1.regOut[15] [19]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _8810_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_913_[20]),
    .Q(\datapath_1.regfile_1.regOut[15] [20]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _8811_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_913_[21]),
    .Q(\datapath_1.regfile_1.regOut[15] [21]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _8812_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_913_[22]),
    .Q(\datapath_1.regfile_1.regOut[15] [22]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _8813_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_913_[23]),
    .Q(\datapath_1.regfile_1.regOut[15] [23]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _8814_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_913_[24]),
    .Q(\datapath_1.regfile_1.regOut[15] [24]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _8815_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_913_[25]),
    .Q(\datapath_1.regfile_1.regOut[15] [25]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _8816_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_913_[26]),
    .Q(\datapath_1.regfile_1.regOut[15] [26]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _8817_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_913_[27]),
    .Q(\datapath_1.regfile_1.regOut[15] [27]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _8818_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_913_[28]),
    .Q(\datapath_1.regfile_1.regOut[15] [28]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _8819_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_913_[29]),
    .Q(\datapath_1.regfile_1.regOut[15] [29]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _8820_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_913_[30]),
    .Q(\datapath_1.regfile_1.regOut[15] [30]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _8821_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_913_[31]),
    .Q(\datapath_1.regfile_1.regOut[15] [31]),
    .R(rst_bF$buf94),
    .S(vdd)
);

INVX1 _8822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [0]),
    .Y(_1041_)
);

NAND2X1 _8823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .Y(_1042_)
);

OAI21X1 _8824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1041_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1042_),
    .Y(_978_[0])
);

INVX1 _8825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [1]),
    .Y(_979_)
);

NAND2X1 _8826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_980_)
);

OAI21X1 _8827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_980_),
    .Y(_978_[1])
);

INVX1 _8828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [2]),
    .Y(_981_)
);

NAND2X1 _8829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_982_)
);

OAI21X1 _8830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_981_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_982_),
    .Y(_978_[2])
);

INVX1 _8831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [3]),
    .Y(_983_)
);

NAND2X1 _8832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_984_)
);

OAI21X1 _8833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_983_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_984_),
    .Y(_978_[3])
);

INVX1 _8834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [4]),
    .Y(_985_)
);

NAND2X1 _8835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_986_)
);

OAI21X1 _8836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_985_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_986_),
    .Y(_978_[4])
);

INVX1 _8837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [5]),
    .Y(_987_)
);

NAND2X1 _8838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_988_)
);

OAI21X1 _8839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_987_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_988_),
    .Y(_978_[5])
);

INVX1 _8840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [6]),
    .Y(_989_)
);

NAND2X1 _8841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_990_)
);

OAI21X1 _8842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_989_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_990_),
    .Y(_978_[6])
);

INVX1 _8843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [7]),
    .Y(_991_)
);

NAND2X1 _8844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_992_)
);

OAI21X1 _8845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_991_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_992_),
    .Y(_978_[7])
);

INVX1 _8846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [8]),
    .Y(_993_)
);

NAND2X1 _8847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_994_)
);

OAI21X1 _8848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_993_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_994_),
    .Y(_978_[8])
);

INVX1 _8849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [9]),
    .Y(_995_)
);

NAND2X1 _8850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_996_)
);

OAI21X1 _8851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_995_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_996_),
    .Y(_978_[9])
);

INVX1 _8852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [10]),
    .Y(_997_)
);

NAND2X1 _8853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_998_)
);

OAI21X1 _8854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_997_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_998_),
    .Y(_978_[10])
);

INVX1 _8855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [11]),
    .Y(_999_)
);

NAND2X1 _8856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1000_)
);

OAI21X1 _8857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_999_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1000_),
    .Y(_978_[11])
);

INVX1 _8858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [12]),
    .Y(_1001_)
);

NAND2X1 _8859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1002_)
);

OAI21X1 _8860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1001_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1002_),
    .Y(_978_[12])
);

INVX1 _8861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [13]),
    .Y(_1003_)
);

NAND2X1 _8862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1004_)
);

OAI21X1 _8863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1003_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1004_),
    .Y(_978_[13])
);

INVX1 _8864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [14]),
    .Y(_1005_)
);

NAND2X1 _8865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1006_)
);

OAI21X1 _8866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1005_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1006_),
    .Y(_978_[14])
);

INVX1 _8867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [15]),
    .Y(_1007_)
);

NAND2X1 _8868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1008_)
);

OAI21X1 _8869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1007_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1008_),
    .Y(_978_[15])
);

INVX1 _8870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [16]),
    .Y(_1009_)
);

NAND2X1 _8871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1010_)
);

OAI21X1 _8872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1009_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1010_),
    .Y(_978_[16])
);

INVX1 _8873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [17]),
    .Y(_1011_)
);

NAND2X1 _8874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1012_)
);

OAI21X1 _8875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1011_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1012_),
    .Y(_978_[17])
);

INVX1 _8876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [18]),
    .Y(_1013_)
);

NAND2X1 _8877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1014_)
);

OAI21X1 _8878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1013_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1014_),
    .Y(_978_[18])
);

INVX1 _8879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [19]),
    .Y(_1015_)
);

NAND2X1 _8880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1016_)
);

OAI21X1 _8881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1015_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1016_),
    .Y(_978_[19])
);

INVX1 _8882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [20]),
    .Y(_1017_)
);

NAND2X1 _8883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1018_)
);

OAI21X1 _8884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1017_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1018_),
    .Y(_978_[20])
);

INVX1 _8885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [21]),
    .Y(_1019_)
);

NAND2X1 _8886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1020_)
);

OAI21X1 _8887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1019_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1020_),
    .Y(_978_[21])
);

INVX1 _8888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [22]),
    .Y(_1021_)
);

NAND2X1 _8889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1022_)
);

OAI21X1 _8890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1021_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1022_),
    .Y(_978_[22])
);

INVX1 _8891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [23]),
    .Y(_1023_)
);

NAND2X1 _8892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1024_)
);

OAI21X1 _8893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1023_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1024_),
    .Y(_978_[23])
);

INVX1 _8894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [24]),
    .Y(_1025_)
);

NAND2X1 _8895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1026_)
);

OAI21X1 _8896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1025_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1026_),
    .Y(_978_[24])
);

INVX1 _8897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [25]),
    .Y(_1027_)
);

NAND2X1 _8898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1028_)
);

OAI21X1 _8899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1027_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1028_),
    .Y(_978_[25])
);

INVX1 _8900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [26]),
    .Y(_1029_)
);

NAND2X1 _8901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1030_)
);

OAI21X1 _8902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1029_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1030_),
    .Y(_978_[26])
);

INVX1 _8903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [27]),
    .Y(_1031_)
);

NAND2X1 _8904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1032_)
);

OAI21X1 _8905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1032_),
    .Y(_978_[27])
);

INVX1 _8906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [28]),
    .Y(_1033_)
);

NAND2X1 _8907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1034_)
);

OAI21X1 _8908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1033_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf6 ),
    .C(_1034_),
    .Y(_978_[28])
);

INVX1 _8909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [29]),
    .Y(_1035_)
);

NAND2X1 _8910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1036_)
);

OAI21X1 _8911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1035_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf4 ),
    .C(_1036_),
    .Y(_978_[29])
);

INVX1 _8912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [30]),
    .Y(_1037_)
);

NAND2X1 _8913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1038_)
);

OAI21X1 _8914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1037_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf2 ),
    .C(_1038_),
    .Y(_978_[30])
);

INVX1 _8915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[16] [31]),
    .Y(_1039_)
);

NAND2X1 _8916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_16_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1040_)
);

OAI21X1 _8917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1039_),
    .B(\datapath_1.regfile_1.regEn_16_bF$buf0 ),
    .C(_1040_),
    .Y(_978_[31])
);

DFFSR _8918_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_978_[0]),
    .Q(\datapath_1.regfile_1.regOut[16] [0]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _8919_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_978_[1]),
    .Q(\datapath_1.regfile_1.regOut[16] [1]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _8920_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_978_[2]),
    .Q(\datapath_1.regfile_1.regOut[16] [2]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _8921_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_978_[3]),
    .Q(\datapath_1.regfile_1.regOut[16] [3]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _8922_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_978_[4]),
    .Q(\datapath_1.regfile_1.regOut[16] [4]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _8923_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_978_[5]),
    .Q(\datapath_1.regfile_1.regOut[16] [5]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _8924_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_978_[6]),
    .Q(\datapath_1.regfile_1.regOut[16] [6]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _8925_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_978_[7]),
    .Q(\datapath_1.regfile_1.regOut[16] [7]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _8926_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_978_[8]),
    .Q(\datapath_1.regfile_1.regOut[16] [8]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _8927_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_978_[9]),
    .Q(\datapath_1.regfile_1.regOut[16] [9]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _8928_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_978_[10]),
    .Q(\datapath_1.regfile_1.regOut[16] [10]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _8929_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_978_[11]),
    .Q(\datapath_1.regfile_1.regOut[16] [11]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _8930_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_978_[12]),
    .Q(\datapath_1.regfile_1.regOut[16] [12]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _8931_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_978_[13]),
    .Q(\datapath_1.regfile_1.regOut[16] [13]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _8932_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_978_[14]),
    .Q(\datapath_1.regfile_1.regOut[16] [14]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _8933_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_978_[15]),
    .Q(\datapath_1.regfile_1.regOut[16] [15]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _8934_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_978_[16]),
    .Q(\datapath_1.regfile_1.regOut[16] [16]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _8935_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_978_[17]),
    .Q(\datapath_1.regfile_1.regOut[16] [17]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _8936_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_978_[18]),
    .Q(\datapath_1.regfile_1.regOut[16] [18]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _8937_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_978_[19]),
    .Q(\datapath_1.regfile_1.regOut[16] [19]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _8938_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_978_[20]),
    .Q(\datapath_1.regfile_1.regOut[16] [20]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _8939_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_978_[21]),
    .Q(\datapath_1.regfile_1.regOut[16] [21]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _8940_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_978_[22]),
    .Q(\datapath_1.regfile_1.regOut[16] [22]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _8941_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_978_[23]),
    .Q(\datapath_1.regfile_1.regOut[16] [23]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _8942_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_978_[24]),
    .Q(\datapath_1.regfile_1.regOut[16] [24]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _8943_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_978_[25]),
    .Q(\datapath_1.regfile_1.regOut[16] [25]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _8944_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_978_[26]),
    .Q(\datapath_1.regfile_1.regOut[16] [26]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _8945_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_978_[27]),
    .Q(\datapath_1.regfile_1.regOut[16] [27]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _8946_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_978_[28]),
    .Q(\datapath_1.regfile_1.regOut[16] [28]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _8947_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_978_[29]),
    .Q(\datapath_1.regfile_1.regOut[16] [29]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _8948_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_978_[30]),
    .Q(\datapath_1.regfile_1.regOut[16] [30]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _8949_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_978_[31]),
    .Q(\datapath_1.regfile_1.regOut[16] [31]),
    .R(rst_bF$buf62),
    .S(vdd)
);

INVX1 _8950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [0]),
    .Y(_1106_)
);

NAND2X1 _8951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .Y(_1107_)
);

OAI21X1 _8952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1106_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1107_),
    .Y(_1043_[0])
);

INVX1 _8953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [1]),
    .Y(_1044_)
);

NAND2X1 _8954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1045_)
);

OAI21X1 _8955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1044_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1045_),
    .Y(_1043_[1])
);

INVX1 _8956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [2]),
    .Y(_1046_)
);

NAND2X1 _8957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1047_)
);

OAI21X1 _8958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1046_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1047_),
    .Y(_1043_[2])
);

INVX1 _8959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [3]),
    .Y(_1048_)
);

NAND2X1 _8960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1049_)
);

OAI21X1 _8961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1049_),
    .Y(_1043_[3])
);

INVX1 _8962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [4]),
    .Y(_1050_)
);

NAND2X1 _8963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1051_)
);

OAI21X1 _8964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1050_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1051_),
    .Y(_1043_[4])
);

INVX1 _8965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [5]),
    .Y(_1052_)
);

NAND2X1 _8966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1053_)
);

OAI21X1 _8967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1053_),
    .Y(_1043_[5])
);

INVX1 _8968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [6]),
    .Y(_1054_)
);

NAND2X1 _8969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1055_)
);

OAI21X1 _8970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1055_),
    .Y(_1043_[6])
);

INVX1 _8971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [7]),
    .Y(_1056_)
);

NAND2X1 _8972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1057_)
);

OAI21X1 _8973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1057_),
    .Y(_1043_[7])
);

INVX1 _8974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [8]),
    .Y(_1058_)
);

NAND2X1 _8975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1059_)
);

OAI21X1 _8976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1059_),
    .Y(_1043_[8])
);

INVX1 _8977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [9]),
    .Y(_1060_)
);

NAND2X1 _8978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1061_)
);

OAI21X1 _8979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1060_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1061_),
    .Y(_1043_[9])
);

INVX1 _8980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [10]),
    .Y(_1062_)
);

NAND2X1 _8981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1063_)
);

OAI21X1 _8982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1062_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1063_),
    .Y(_1043_[10])
);

INVX1 _8983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [11]),
    .Y(_1064_)
);

NAND2X1 _8984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1065_)
);

OAI21X1 _8985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1065_),
    .Y(_1043_[11])
);

INVX1 _8986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [12]),
    .Y(_1066_)
);

NAND2X1 _8987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1067_)
);

OAI21X1 _8988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1067_),
    .Y(_1043_[12])
);

INVX1 _8989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [13]),
    .Y(_1068_)
);

NAND2X1 _8990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1069_)
);

OAI21X1 _8991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1068_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1069_),
    .Y(_1043_[13])
);

INVX1 _8992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [14]),
    .Y(_1070_)
);

NAND2X1 _8993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1071_)
);

OAI21X1 _8994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1070_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1071_),
    .Y(_1043_[14])
);

INVX1 _8995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [15]),
    .Y(_1072_)
);

NAND2X1 _8996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1073_)
);

OAI21X1 _8997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1072_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1073_),
    .Y(_1043_[15])
);

INVX1 _8998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [16]),
    .Y(_1074_)
);

NAND2X1 _8999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1075_)
);

OAI21X1 _9000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1074_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1075_),
    .Y(_1043_[16])
);

INVX1 _9001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [17]),
    .Y(_1076_)
);

NAND2X1 _9002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1077_)
);

OAI21X1 _9003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1076_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1077_),
    .Y(_1043_[17])
);

INVX1 _9004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [18]),
    .Y(_1078_)
);

NAND2X1 _9005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1079_)
);

OAI21X1 _9006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1078_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1079_),
    .Y(_1043_[18])
);

INVX1 _9007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [19]),
    .Y(_1080_)
);

NAND2X1 _9008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1081_)
);

OAI21X1 _9009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1080_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1081_),
    .Y(_1043_[19])
);

INVX1 _9010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [20]),
    .Y(_1082_)
);

NAND2X1 _9011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1083_)
);

OAI21X1 _9012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1083_),
    .Y(_1043_[20])
);

INVX1 _9013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [21]),
    .Y(_1084_)
);

NAND2X1 _9014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1085_)
);

OAI21X1 _9015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1084_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1085_),
    .Y(_1043_[21])
);

INVX1 _9016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [22]),
    .Y(_1086_)
);

NAND2X1 _9017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_1087_)
);

OAI21X1 _9018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1086_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1087_),
    .Y(_1043_[22])
);

INVX1 _9019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [23]),
    .Y(_1088_)
);

NAND2X1 _9020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1089_)
);

OAI21X1 _9021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1089_),
    .Y(_1043_[23])
);

INVX1 _9022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [24]),
    .Y(_1090_)
);

NAND2X1 _9023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1091_)
);

OAI21X1 _9024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1090_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1091_),
    .Y(_1043_[24])
);

INVX1 _9025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [25]),
    .Y(_1092_)
);

NAND2X1 _9026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1093_)
);

OAI21X1 _9027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1093_),
    .Y(_1043_[25])
);

INVX1 _9028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [26]),
    .Y(_1094_)
);

NAND2X1 _9029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1095_)
);

OAI21X1 _9030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1094_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1095_),
    .Y(_1043_[26])
);

INVX1 _9031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [27]),
    .Y(_1096_)
);

NAND2X1 _9032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1097_)
);

OAI21X1 _9033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1097_),
    .Y(_1043_[27])
);

INVX1 _9034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [28]),
    .Y(_1098_)
);

NAND2X1 _9035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1099_)
);

OAI21X1 _9036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1098_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf6 ),
    .C(_1099_),
    .Y(_1043_[28])
);

INVX1 _9037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [29]),
    .Y(_1100_)
);

NAND2X1 _9038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1101_)
);

OAI21X1 _9039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1100_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf4 ),
    .C(_1101_),
    .Y(_1043_[29])
);

INVX1 _9040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [30]),
    .Y(_1102_)
);

NAND2X1 _9041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1103_)
);

OAI21X1 _9042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf2 ),
    .C(_1103_),
    .Y(_1043_[30])
);

INVX1 _9043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[17] [31]),
    .Y(_1104_)
);

NAND2X1 _9044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_17_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1105_)
);

OAI21X1 _9045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1104_),
    .B(\datapath_1.regfile_1.regEn_17_bF$buf0 ),
    .C(_1105_),
    .Y(_1043_[31])
);

DFFSR _9046_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_1043_[0]),
    .Q(\datapath_1.regfile_1.regOut[17] [0]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _9047_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_1043_[1]),
    .Q(\datapath_1.regfile_1.regOut[17] [1]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _9048_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_1043_[2]),
    .Q(\datapath_1.regfile_1.regOut[17] [2]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _9049_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_1043_[3]),
    .Q(\datapath_1.regfile_1.regOut[17] [3]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _9050_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_1043_[4]),
    .Q(\datapath_1.regfile_1.regOut[17] [4]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _9051_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_1043_[5]),
    .Q(\datapath_1.regfile_1.regOut[17] [5]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _9052_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_1043_[6]),
    .Q(\datapath_1.regfile_1.regOut[17] [6]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _9053_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_1043_[7]),
    .Q(\datapath_1.regfile_1.regOut[17] [7]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _9054_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_1043_[8]),
    .Q(\datapath_1.regfile_1.regOut[17] [8]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _9055_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_1043_[9]),
    .Q(\datapath_1.regfile_1.regOut[17] [9]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _9056_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_1043_[10]),
    .Q(\datapath_1.regfile_1.regOut[17] [10]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _9057_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_1043_[11]),
    .Q(\datapath_1.regfile_1.regOut[17] [11]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _9058_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_1043_[12]),
    .Q(\datapath_1.regfile_1.regOut[17] [12]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _9059_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_1043_[13]),
    .Q(\datapath_1.regfile_1.regOut[17] [13]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _9060_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_1043_[14]),
    .Q(\datapath_1.regfile_1.regOut[17] [14]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _9061_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_1043_[15]),
    .Q(\datapath_1.regfile_1.regOut[17] [15]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _9062_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_1043_[16]),
    .Q(\datapath_1.regfile_1.regOut[17] [16]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _9063_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_1043_[17]),
    .Q(\datapath_1.regfile_1.regOut[17] [17]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _9064_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_1043_[18]),
    .Q(\datapath_1.regfile_1.regOut[17] [18]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _9065_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_1043_[19]),
    .Q(\datapath_1.regfile_1.regOut[17] [19]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _9066_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_1043_[20]),
    .Q(\datapath_1.regfile_1.regOut[17] [20]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _9067_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_1043_[21]),
    .Q(\datapath_1.regfile_1.regOut[17] [21]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _9068_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_1043_[22]),
    .Q(\datapath_1.regfile_1.regOut[17] [22]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _9069_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_1043_[23]),
    .Q(\datapath_1.regfile_1.regOut[17] [23]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _9070_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_1043_[24]),
    .Q(\datapath_1.regfile_1.regOut[17] [24]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _9071_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_1043_[25]),
    .Q(\datapath_1.regfile_1.regOut[17] [25]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _9072_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_1043_[26]),
    .Q(\datapath_1.regfile_1.regOut[17] [26]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _9073_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_1043_[27]),
    .Q(\datapath_1.regfile_1.regOut[17] [27]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _9074_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_1043_[28]),
    .Q(\datapath_1.regfile_1.regOut[17] [28]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _9075_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_1043_[29]),
    .Q(\datapath_1.regfile_1.regOut[17] [29]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _9076_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_1043_[30]),
    .Q(\datapath_1.regfile_1.regOut[17] [30]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _9077_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_1043_[31]),
    .Q(\datapath_1.regfile_1.regOut[17] [31]),
    .R(rst_bF$buf30),
    .S(vdd)
);

INVX1 _9078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [0]),
    .Y(_1171_)
);

NAND2X1 _9079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .Y(_1172_)
);

OAI21X1 _9080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1172_),
    .Y(_1108_[0])
);

INVX1 _9081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [1]),
    .Y(_1109_)
);

NAND2X1 _9082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1110_)
);

OAI21X1 _9083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1109_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1110_),
    .Y(_1108_[1])
);

INVX1 _9084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [2]),
    .Y(_1111_)
);

NAND2X1 _9085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1112_)
);

OAI21X1 _9086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1111_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1112_),
    .Y(_1108_[2])
);

INVX1 _9087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [3]),
    .Y(_1113_)
);

NAND2X1 _9088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1114_)
);

OAI21X1 _9089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1113_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1114_),
    .Y(_1108_[3])
);

INVX1 _9090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [4]),
    .Y(_1115_)
);

NAND2X1 _9091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1116_)
);

OAI21X1 _9092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1115_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1116_),
    .Y(_1108_[4])
);

INVX1 _9093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [5]),
    .Y(_1117_)
);

NAND2X1 _9094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1118_)
);

OAI21X1 _9095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1117_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1118_),
    .Y(_1108_[5])
);

INVX1 _9096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [6]),
    .Y(_1119_)
);

NAND2X1 _9097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1120_)
);

OAI21X1 _9098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1120_),
    .Y(_1108_[6])
);

INVX1 _9099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [7]),
    .Y(_1121_)
);

NAND2X1 _9100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1122_)
);

OAI21X1 _9101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1121_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1122_),
    .Y(_1108_[7])
);

INVX1 _9102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [8]),
    .Y(_1123_)
);

NAND2X1 _9103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1124_)
);

OAI21X1 _9104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1124_),
    .Y(_1108_[8])
);

INVX1 _9105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [9]),
    .Y(_1125_)
);

NAND2X1 _9106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1126_)
);

OAI21X1 _9107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1126_),
    .Y(_1108_[9])
);

INVX1 _9108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [10]),
    .Y(_1127_)
);

NAND2X1 _9109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1128_)
);

OAI21X1 _9110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1127_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1128_),
    .Y(_1108_[10])
);

INVX1 _9111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [11]),
    .Y(_1129_)
);

NAND2X1 _9112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1130_)
);

OAI21X1 _9113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1130_),
    .Y(_1108_[11])
);

INVX1 _9114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [12]),
    .Y(_1131_)
);

NAND2X1 _9115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1132_)
);

OAI21X1 _9116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1131_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1132_),
    .Y(_1108_[12])
);

INVX1 _9117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [13]),
    .Y(_1133_)
);

NAND2X1 _9118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1134_)
);

OAI21X1 _9119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1134_),
    .Y(_1108_[13])
);

INVX1 _9120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [14]),
    .Y(_1135_)
);

NAND2X1 _9121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1136_)
);

OAI21X1 _9122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1136_),
    .Y(_1108_[14])
);

INVX1 _9123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [15]),
    .Y(_1137_)
);

NAND2X1 _9124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1138_)
);

OAI21X1 _9125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1138_),
    .Y(_1108_[15])
);

INVX1 _9126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [16]),
    .Y(_1139_)
);

NAND2X1 _9127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1140_)
);

OAI21X1 _9128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1140_),
    .Y(_1108_[16])
);

INVX1 _9129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [17]),
    .Y(_1141_)
);

NAND2X1 _9130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1142_)
);

OAI21X1 _9131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1142_),
    .Y(_1108_[17])
);

INVX1 _9132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [18]),
    .Y(_1143_)
);

NAND2X1 _9133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1144_)
);

OAI21X1 _9134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1143_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1144_),
    .Y(_1108_[18])
);

INVX1 _9135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [19]),
    .Y(_1145_)
);

NAND2X1 _9136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1146_)
);

OAI21X1 _9137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1146_),
    .Y(_1108_[19])
);

INVX1 _9138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [20]),
    .Y(_1147_)
);

NAND2X1 _9139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1148_)
);

OAI21X1 _9140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1147_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1148_),
    .Y(_1108_[20])
);

INVX1 _9141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [21]),
    .Y(_1149_)
);

NAND2X1 _9142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1150_)
);

OAI21X1 _9143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1150_),
    .Y(_1108_[21])
);

INVX1 _9144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [22]),
    .Y(_1151_)
);

NAND2X1 _9145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1152_)
);

OAI21X1 _9146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1151_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1152_),
    .Y(_1108_[22])
);

INVX1 _9147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [23]),
    .Y(_1153_)
);

NAND2X1 _9148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1154_)
);

OAI21X1 _9149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1153_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1154_),
    .Y(_1108_[23])
);

INVX1 _9150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [24]),
    .Y(_1155_)
);

NAND2X1 _9151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1156_)
);

OAI21X1 _9152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1155_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1156_),
    .Y(_1108_[24])
);

INVX1 _9153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [25]),
    .Y(_1157_)
);

NAND2X1 _9154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1158_)
);

OAI21X1 _9155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1157_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1158_),
    .Y(_1108_[25])
);

INVX1 _9156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [26]),
    .Y(_1159_)
);

NAND2X1 _9157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1160_)
);

OAI21X1 _9158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1160_),
    .Y(_1108_[26])
);

INVX1 _9159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [27]),
    .Y(_1161_)
);

NAND2X1 _9160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1162_)
);

OAI21X1 _9161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1161_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1162_),
    .Y(_1108_[27])
);

INVX1 _9162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [28]),
    .Y(_1163_)
);

NAND2X1 _9163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1164_)
);

OAI21X1 _9164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1163_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf6 ),
    .C(_1164_),
    .Y(_1108_[28])
);

INVX1 _9165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [29]),
    .Y(_1165_)
);

NAND2X1 _9166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1166_)
);

OAI21X1 _9167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf4 ),
    .C(_1166_),
    .Y(_1108_[29])
);

INVX1 _9168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [30]),
    .Y(_1167_)
);

NAND2X1 _9169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1168_)
);

OAI21X1 _9170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1167_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf2 ),
    .C(_1168_),
    .Y(_1108_[30])
);

INVX1 _9171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[18] [31]),
    .Y(_1169_)
);

NAND2X1 _9172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_18_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1170_)
);

OAI21X1 _9173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1169_),
    .B(\datapath_1.regfile_1.regEn_18_bF$buf0 ),
    .C(_1170_),
    .Y(_1108_[31])
);

DFFSR _9174_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_1108_[0]),
    .Q(\datapath_1.regfile_1.regOut[18] [0]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _9175_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_1108_[1]),
    .Q(\datapath_1.regfile_1.regOut[18] [1]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _9176_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_1108_[2]),
    .Q(\datapath_1.regfile_1.regOut[18] [2]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _9177_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_1108_[3]),
    .Q(\datapath_1.regfile_1.regOut[18] [3]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _9178_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_1108_[4]),
    .Q(\datapath_1.regfile_1.regOut[18] [4]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _9179_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_1108_[5]),
    .Q(\datapath_1.regfile_1.regOut[18] [5]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _9180_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_1108_[6]),
    .Q(\datapath_1.regfile_1.regOut[18] [6]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _9181_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_1108_[7]),
    .Q(\datapath_1.regfile_1.regOut[18] [7]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _9182_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_1108_[8]),
    .Q(\datapath_1.regfile_1.regOut[18] [8]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _9183_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_1108_[9]),
    .Q(\datapath_1.regfile_1.regOut[18] [9]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _9184_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_1108_[10]),
    .Q(\datapath_1.regfile_1.regOut[18] [10]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _9185_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_1108_[11]),
    .Q(\datapath_1.regfile_1.regOut[18] [11]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _9186_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_1108_[12]),
    .Q(\datapath_1.regfile_1.regOut[18] [12]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _9187_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_1108_[13]),
    .Q(\datapath_1.regfile_1.regOut[18] [13]),
    .R(rst_bF$buf16),
    .S(vdd)
);

DFFSR _9188_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_1108_[14]),
    .Q(\datapath_1.regfile_1.regOut[18] [14]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _9189_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_1108_[15]),
    .Q(\datapath_1.regfile_1.regOut[18] [15]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _9190_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_1108_[16]),
    .Q(\datapath_1.regfile_1.regOut[18] [16]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _9191_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_1108_[17]),
    .Q(\datapath_1.regfile_1.regOut[18] [17]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _9192_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_1108_[18]),
    .Q(\datapath_1.regfile_1.regOut[18] [18]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _9193_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_1108_[19]),
    .Q(\datapath_1.regfile_1.regOut[18] [19]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _9194_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_1108_[20]),
    .Q(\datapath_1.regfile_1.regOut[18] [20]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _9195_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_1108_[21]),
    .Q(\datapath_1.regfile_1.regOut[18] [21]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _9196_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1108_[22]),
    .Q(\datapath_1.regfile_1.regOut[18] [22]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _9197_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1108_[23]),
    .Q(\datapath_1.regfile_1.regOut[18] [23]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _9198_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1108_[24]),
    .Q(\datapath_1.regfile_1.regOut[18] [24]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _9199_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1108_[25]),
    .Q(\datapath_1.regfile_1.regOut[18] [25]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _9200_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1108_[26]),
    .Q(\datapath_1.regfile_1.regOut[18] [26]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _9201_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1108_[27]),
    .Q(\datapath_1.regfile_1.regOut[18] [27]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _9202_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1108_[28]),
    .Q(\datapath_1.regfile_1.regOut[18] [28]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _9203_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1108_[29]),
    .Q(\datapath_1.regfile_1.regOut[18] [29]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _9204_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_1108_[30]),
    .Q(\datapath_1.regfile_1.regOut[18] [30]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _9205_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_1108_[31]),
    .Q(\datapath_1.regfile_1.regOut[18] [31]),
    .R(rst_bF$buf112),
    .S(vdd)
);

INVX1 _9206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [0]),
    .Y(_1236_)
);

NAND2X1 _9207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .Y(_1237_)
);

OAI21X1 _9208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1237_),
    .Y(_1173_[0])
);

INVX1 _9209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [1]),
    .Y(_1174_)
);

NAND2X1 _9210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1175_)
);

OAI21X1 _9211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1174_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1175_),
    .Y(_1173_[1])
);

INVX1 _9212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [2]),
    .Y(_1176_)
);

NAND2X1 _9213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1177_)
);

OAI21X1 _9214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1176_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1177_),
    .Y(_1173_[2])
);

INVX1 _9215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [3]),
    .Y(_1178_)
);

NAND2X1 _9216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1179_)
);

OAI21X1 _9217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1179_),
    .Y(_1173_[3])
);

INVX1 _9218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [4]),
    .Y(_1180_)
);

NAND2X1 _9219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1181_)
);

OAI21X1 _9220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1180_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1181_),
    .Y(_1173_[4])
);

INVX1 _9221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [5]),
    .Y(_1182_)
);

NAND2X1 _9222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1183_)
);

OAI21X1 _9223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1182_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1183_),
    .Y(_1173_[5])
);

INVX1 _9224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [6]),
    .Y(_1184_)
);

NAND2X1 _9225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1185_)
);

OAI21X1 _9226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1185_),
    .Y(_1173_[6])
);

INVX1 _9227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [7]),
    .Y(_1186_)
);

NAND2X1 _9228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1187_)
);

OAI21X1 _9229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1186_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1187_),
    .Y(_1173_[7])
);

INVX1 _9230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [8]),
    .Y(_1188_)
);

NAND2X1 _9231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1189_)
);

OAI21X1 _9232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1188_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1189_),
    .Y(_1173_[8])
);

INVX1 _9233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [9]),
    .Y(_1190_)
);

NAND2X1 _9234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1191_)
);

OAI21X1 _9235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1190_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1191_),
    .Y(_1173_[9])
);

INVX1 _9236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [10]),
    .Y(_1192_)
);

NAND2X1 _9237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1193_)
);

OAI21X1 _9238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1192_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1193_),
    .Y(_1173_[10])
);

INVX1 _9239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [11]),
    .Y(_1194_)
);

NAND2X1 _9240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1195_)
);

OAI21X1 _9241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1194_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1195_),
    .Y(_1173_[11])
);

INVX1 _9242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [12]),
    .Y(_1196_)
);

NAND2X1 _9243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1197_)
);

OAI21X1 _9244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1197_),
    .Y(_1173_[12])
);

INVX1 _9245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [13]),
    .Y(_1198_)
);

NAND2X1 _9246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1199_)
);

OAI21X1 _9247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1198_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1199_),
    .Y(_1173_[13])
);

INVX1 _9248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [14]),
    .Y(_1200_)
);

NAND2X1 _9249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1201_)
);

OAI21X1 _9250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1200_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1201_),
    .Y(_1173_[14])
);

INVX1 _9251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [15]),
    .Y(_1202_)
);

NAND2X1 _9252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1203_)
);

OAI21X1 _9253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1203_),
    .Y(_1173_[15])
);

INVX1 _9254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [16]),
    .Y(_1204_)
);

NAND2X1 _9255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1205_)
);

OAI21X1 _9256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1204_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1205_),
    .Y(_1173_[16])
);

INVX1 _9257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [17]),
    .Y(_1206_)
);

NAND2X1 _9258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1207_)
);

OAI21X1 _9259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1206_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1207_),
    .Y(_1173_[17])
);

INVX1 _9260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [18]),
    .Y(_1208_)
);

NAND2X1 _9261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1209_)
);

OAI21X1 _9262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1209_),
    .Y(_1173_[18])
);

INVX1 _9263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [19]),
    .Y(_1210_)
);

NAND2X1 _9264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1211_)
);

OAI21X1 _9265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1210_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1211_),
    .Y(_1173_[19])
);

INVX1 _9266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [20]),
    .Y(_1212_)
);

NAND2X1 _9267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1213_)
);

OAI21X1 _9268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1212_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1213_),
    .Y(_1173_[20])
);

INVX1 _9269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [21]),
    .Y(_1214_)
);

NAND2X1 _9270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1215_)
);

OAI21X1 _9271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1215_),
    .Y(_1173_[21])
);

INVX1 _9272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [22]),
    .Y(_1216_)
);

NAND2X1 _9273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1217_)
);

OAI21X1 _9274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1216_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1217_),
    .Y(_1173_[22])
);

INVX1 _9275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [23]),
    .Y(_1218_)
);

NAND2X1 _9276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1219_)
);

OAI21X1 _9277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1218_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1219_),
    .Y(_1173_[23])
);

INVX1 _9278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [24]),
    .Y(_1220_)
);

NAND2X1 _9279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1221_)
);

OAI21X1 _9280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1221_),
    .Y(_1173_[24])
);

INVX1 _9281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [25]),
    .Y(_1222_)
);

NAND2X1 _9282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1223_)
);

OAI21X1 _9283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1222_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1223_),
    .Y(_1173_[25])
);

INVX1 _9284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [26]),
    .Y(_1224_)
);

NAND2X1 _9285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1225_)
);

OAI21X1 _9286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1224_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1225_),
    .Y(_1173_[26])
);

INVX1 _9287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [27]),
    .Y(_1226_)
);

NAND2X1 _9288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1227_)
);

OAI21X1 _9289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1227_),
    .Y(_1173_[27])
);

INVX1 _9290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [28]),
    .Y(_1228_)
);

NAND2X1 _9291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1229_)
);

OAI21X1 _9292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1228_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf6 ),
    .C(_1229_),
    .Y(_1173_[28])
);

INVX1 _9293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [29]),
    .Y(_1230_)
);

NAND2X1 _9294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1231_)
);

OAI21X1 _9295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf4 ),
    .C(_1231_),
    .Y(_1173_[29])
);

INVX1 _9296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [30]),
    .Y(_1232_)
);

NAND2X1 _9297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1233_)
);

OAI21X1 _9298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1232_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf2 ),
    .C(_1233_),
    .Y(_1173_[30])
);

INVX1 _9299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[19] [31]),
    .Y(_1234_)
);

NAND2X1 _9300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_19_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1235_)
);

OAI21X1 _9301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1234_),
    .B(\datapath_1.regfile_1.regEn_19_bF$buf0 ),
    .C(_1235_),
    .Y(_1173_[31])
);

DFFSR _9302_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_1173_[0]),
    .Q(\datapath_1.regfile_1.regOut[19] [0]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _9303_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_1173_[1]),
    .Q(\datapath_1.regfile_1.regOut[19] [1]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _9304_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_1173_[2]),
    .Q(\datapath_1.regfile_1.regOut[19] [2]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _9305_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_1173_[3]),
    .Q(\datapath_1.regfile_1.regOut[19] [3]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _9306_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_1173_[4]),
    .Q(\datapath_1.regfile_1.regOut[19] [4]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _9307_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_1173_[5]),
    .Q(\datapath_1.regfile_1.regOut[19] [5]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _9308_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_1173_[6]),
    .Q(\datapath_1.regfile_1.regOut[19] [6]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _9309_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_1173_[7]),
    .Q(\datapath_1.regfile_1.regOut[19] [7]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _9310_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_1173_[8]),
    .Q(\datapath_1.regfile_1.regOut[19] [8]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _9311_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_1173_[9]),
    .Q(\datapath_1.regfile_1.regOut[19] [9]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _9312_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_1173_[10]),
    .Q(\datapath_1.regfile_1.regOut[19] [10]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _9313_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_1173_[11]),
    .Q(\datapath_1.regfile_1.regOut[19] [11]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _9314_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_1173_[12]),
    .Q(\datapath_1.regfile_1.regOut[19] [12]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _9315_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_1173_[13]),
    .Q(\datapath_1.regfile_1.regOut[19] [13]),
    .R(rst_bF$buf98),
    .S(vdd)
);

DFFSR _9316_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_1173_[14]),
    .Q(\datapath_1.regfile_1.regOut[19] [14]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _9317_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_1173_[15]),
    .Q(\datapath_1.regfile_1.regOut[19] [15]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _9318_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_1173_[16]),
    .Q(\datapath_1.regfile_1.regOut[19] [16]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _9319_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_1173_[17]),
    .Q(\datapath_1.regfile_1.regOut[19] [17]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _9320_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_1173_[18]),
    .Q(\datapath_1.regfile_1.regOut[19] [18]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _9321_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_1173_[19]),
    .Q(\datapath_1.regfile_1.regOut[19] [19]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _9322_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_1173_[20]),
    .Q(\datapath_1.regfile_1.regOut[19] [20]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _9323_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_1173_[21]),
    .Q(\datapath_1.regfile_1.regOut[19] [21]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _9324_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_1173_[22]),
    .Q(\datapath_1.regfile_1.regOut[19] [22]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _9325_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_1173_[23]),
    .Q(\datapath_1.regfile_1.regOut[19] [23]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _9326_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_1173_[24]),
    .Q(\datapath_1.regfile_1.regOut[19] [24]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _9327_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_1173_[25]),
    .Q(\datapath_1.regfile_1.regOut[19] [25]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _9328_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_1173_[26]),
    .Q(\datapath_1.regfile_1.regOut[19] [26]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _9329_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_1173_[27]),
    .Q(\datapath_1.regfile_1.regOut[19] [27]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _9330_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_1173_[28]),
    .Q(\datapath_1.regfile_1.regOut[19] [28]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _9331_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_1173_[29]),
    .Q(\datapath_1.regfile_1.regOut[19] [29]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _9332_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_1173_[30]),
    .Q(\datapath_1.regfile_1.regOut[19] [30]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _9333_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_1173_[31]),
    .Q(\datapath_1.regfile_1.regOut[19] [31]),
    .R(rst_bF$buf80),
    .S(vdd)
);

INVX1 _9334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [0]),
    .Y(_1301_)
);

NAND2X1 _9335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .Y(_1302_)
);

OAI21X1 _9336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1301_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1302_),
    .Y(_1238_[0])
);

INVX1 _9337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [1]),
    .Y(_1239_)
);

NAND2X1 _9338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1240_)
);

OAI21X1 _9339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1239_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1240_),
    .Y(_1238_[1])
);

INVX1 _9340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [2]),
    .Y(_1241_)
);

NAND2X1 _9341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1242_)
);

OAI21X1 _9342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1242_),
    .Y(_1238_[2])
);

INVX1 _9343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [3]),
    .Y(_1243_)
);

NAND2X1 _9344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1244_)
);

OAI21X1 _9345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1243_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1244_),
    .Y(_1238_[3])
);

INVX1 _9346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [4]),
    .Y(_1245_)
);

NAND2X1 _9347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1246_)
);

OAI21X1 _9348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1245_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1246_),
    .Y(_1238_[4])
);

INVX1 _9349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [5]),
    .Y(_1247_)
);

NAND2X1 _9350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1248_)
);

OAI21X1 _9351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1248_),
    .Y(_1238_[5])
);

INVX1 _9352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [6]),
    .Y(_1249_)
);

NAND2X1 _9353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1250_)
);

OAI21X1 _9354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1249_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1250_),
    .Y(_1238_[6])
);

INVX1 _9355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [7]),
    .Y(_1251_)
);

NAND2X1 _9356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1252_)
);

OAI21X1 _9357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1252_),
    .Y(_1238_[7])
);

INVX1 _9358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [8]),
    .Y(_1253_)
);

NAND2X1 _9359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1254_)
);

OAI21X1 _9360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1253_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1254_),
    .Y(_1238_[8])
);

INVX1 _9361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [9]),
    .Y(_1255_)
);

NAND2X1 _9362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf3 ),
    .Y(_1256_)
);

OAI21X1 _9363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1255_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1256_),
    .Y(_1238_[9])
);

INVX1 _9364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [10]),
    .Y(_1257_)
);

NAND2X1 _9365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf3 ),
    .Y(_1258_)
);

OAI21X1 _9366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1258_),
    .Y(_1238_[10])
);

INVX1 _9367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [11]),
    .Y(_1259_)
);

NAND2X1 _9368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf3 ),
    .Y(_1260_)
);

OAI21X1 _9369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1259_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1260_),
    .Y(_1238_[11])
);

INVX1 _9370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [12]),
    .Y(_1261_)
);

NAND2X1 _9371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf3 ),
    .Y(_1262_)
);

OAI21X1 _9372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1261_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1262_),
    .Y(_1238_[12])
);

INVX1 _9373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [13]),
    .Y(_1263_)
);

NAND2X1 _9374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf3 ),
    .Y(_1264_)
);

OAI21X1 _9375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1263_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1264_),
    .Y(_1238_[13])
);

INVX1 _9376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [14]),
    .Y(_1265_)
);

NAND2X1 _9377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf3 ),
    .Y(_1266_)
);

OAI21X1 _9378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1265_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1266_),
    .Y(_1238_[14])
);

INVX1 _9379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [15]),
    .Y(_1267_)
);

NAND2X1 _9380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf3 ),
    .Y(_1268_)
);

OAI21X1 _9381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1268_),
    .Y(_1238_[15])
);

INVX1 _9382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [16]),
    .Y(_1269_)
);

NAND2X1 _9383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf3 ),
    .Y(_1270_)
);

OAI21X1 _9384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1269_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1270_),
    .Y(_1238_[16])
);

INVX1 _9385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [17]),
    .Y(_1271_)
);

NAND2X1 _9386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf3 ),
    .Y(_1272_)
);

OAI21X1 _9387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1271_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1272_),
    .Y(_1238_[17])
);

INVX1 _9388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [18]),
    .Y(_1273_)
);

NAND2X1 _9389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf3 ),
    .Y(_1274_)
);

OAI21X1 _9390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1273_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1274_),
    .Y(_1238_[18])
);

INVX1 _9391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [19]),
    .Y(_1275_)
);

NAND2X1 _9392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf3 ),
    .Y(_1276_)
);

OAI21X1 _9393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1275_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1276_),
    .Y(_1238_[19])
);

INVX1 _9394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [20]),
    .Y(_1277_)
);

NAND2X1 _9395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf3 ),
    .Y(_1278_)
);

OAI21X1 _9396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1277_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1278_),
    .Y(_1238_[20])
);

INVX1 _9397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [21]),
    .Y(_1279_)
);

NAND2X1 _9398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf3 ),
    .Y(_1280_)
);

OAI21X1 _9399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1279_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1280_),
    .Y(_1238_[21])
);

INVX1 _9400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [22]),
    .Y(_1281_)
);

NAND2X1 _9401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf3 ),
    .Y(_1282_)
);

OAI21X1 _9402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1282_),
    .Y(_1238_[22])
);

INVX1 _9403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [23]),
    .Y(_1283_)
);

NAND2X1 _9404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf3 ),
    .Y(_1284_)
);

OAI21X1 _9405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1283_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1284_),
    .Y(_1238_[23])
);

INVX1 _9406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [24]),
    .Y(_1285_)
);

NAND2X1 _9407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf3 ),
    .Y(_1286_)
);

OAI21X1 _9408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1285_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1286_),
    .Y(_1238_[24])
);

INVX1 _9409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [25]),
    .Y(_1287_)
);

NAND2X1 _9410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf3 ),
    .Y(_1288_)
);

OAI21X1 _9411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1287_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1288_),
    .Y(_1238_[25])
);

INVX1 _9412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [26]),
    .Y(_1289_)
);

NAND2X1 _9413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf3 ),
    .Y(_1290_)
);

OAI21X1 _9414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1289_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1290_),
    .Y(_1238_[26])
);

INVX1 _9415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [27]),
    .Y(_1291_)
);

NAND2X1 _9416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf3 ),
    .Y(_1292_)
);

OAI21X1 _9417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1291_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1292_),
    .Y(_1238_[27])
);

INVX1 _9418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [28]),
    .Y(_1293_)
);

NAND2X1 _9419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf3 ),
    .Y(_1294_)
);

OAI21X1 _9420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf6 ),
    .C(_1294_),
    .Y(_1238_[28])
);

INVX1 _9421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [29]),
    .Y(_1295_)
);

NAND2X1 _9422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf3 ),
    .Y(_1296_)
);

OAI21X1 _9423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf4 ),
    .C(_1296_),
    .Y(_1238_[29])
);

INVX1 _9424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [30]),
    .Y(_1297_)
);

NAND2X1 _9425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf3 ),
    .Y(_1298_)
);

OAI21X1 _9426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf2 ),
    .C(_1298_),
    .Y(_1238_[30])
);

INVX1 _9427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[20] [31]),
    .Y(_1299_)
);

NAND2X1 _9428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_20_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf3 ),
    .Y(_1300_)
);

OAI21X1 _9429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1299_),
    .B(\datapath_1.regfile_1.regEn_20_bF$buf0 ),
    .C(_1300_),
    .Y(_1238_[31])
);

DFFSR _9430_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_1238_[0]),
    .Q(\datapath_1.regfile_1.regOut[20] [0]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _9431_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_1238_[1]),
    .Q(\datapath_1.regfile_1.regOut[20] [1]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _9432_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_1238_[2]),
    .Q(\datapath_1.regfile_1.regOut[20] [2]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _9433_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_1238_[3]),
    .Q(\datapath_1.regfile_1.regOut[20] [3]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _9434_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_1238_[4]),
    .Q(\datapath_1.regfile_1.regOut[20] [4]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _9435_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_1238_[5]),
    .Q(\datapath_1.regfile_1.regOut[20] [5]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _9436_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_1238_[6]),
    .Q(\datapath_1.regfile_1.regOut[20] [6]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _9437_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_1238_[7]),
    .Q(\datapath_1.regfile_1.regOut[20] [7]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _9438_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_1238_[8]),
    .Q(\datapath_1.regfile_1.regOut[20] [8]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _9439_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_1238_[9]),
    .Q(\datapath_1.regfile_1.regOut[20] [9]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _9440_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_1238_[10]),
    .Q(\datapath_1.regfile_1.regOut[20] [10]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _9441_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_1238_[11]),
    .Q(\datapath_1.regfile_1.regOut[20] [11]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _9442_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_1238_[12]),
    .Q(\datapath_1.regfile_1.regOut[20] [12]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _9443_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_1238_[13]),
    .Q(\datapath_1.regfile_1.regOut[20] [13]),
    .R(rst_bF$buf66),
    .S(vdd)
);

DFFSR _9444_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_1238_[14]),
    .Q(\datapath_1.regfile_1.regOut[20] [14]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _9445_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_1238_[15]),
    .Q(\datapath_1.regfile_1.regOut[20] [15]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _9446_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_1238_[16]),
    .Q(\datapath_1.regfile_1.regOut[20] [16]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _9447_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_1238_[17]),
    .Q(\datapath_1.regfile_1.regOut[20] [17]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _9448_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_1238_[18]),
    .Q(\datapath_1.regfile_1.regOut[20] [18]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _9449_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_1238_[19]),
    .Q(\datapath_1.regfile_1.regOut[20] [19]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _9450_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_1238_[20]),
    .Q(\datapath_1.regfile_1.regOut[20] [20]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _9451_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_1238_[21]),
    .Q(\datapath_1.regfile_1.regOut[20] [21]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _9452_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_1238_[22]),
    .Q(\datapath_1.regfile_1.regOut[20] [22]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _9453_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_1238_[23]),
    .Q(\datapath_1.regfile_1.regOut[20] [23]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _9454_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_1238_[24]),
    .Q(\datapath_1.regfile_1.regOut[20] [24]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _9455_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_1238_[25]),
    .Q(\datapath_1.regfile_1.regOut[20] [25]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _9456_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_1238_[26]),
    .Q(\datapath_1.regfile_1.regOut[20] [26]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _9457_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_1238_[27]),
    .Q(\datapath_1.regfile_1.regOut[20] [27]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _9458_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_1238_[28]),
    .Q(\datapath_1.regfile_1.regOut[20] [28]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _9459_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_1238_[29]),
    .Q(\datapath_1.regfile_1.regOut[20] [29]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _9460_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_1238_[30]),
    .Q(\datapath_1.regfile_1.regOut[20] [30]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _9461_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_1238_[31]),
    .Q(\datapath_1.regfile_1.regOut[20] [31]),
    .R(rst_bF$buf48),
    .S(vdd)
);

INVX1 _9462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [0]),
    .Y(_1366_)
);

NAND2X1 _9463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf3 ),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .Y(_1367_)
);

OAI21X1 _9464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1366_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1367_),
    .Y(_1303_[0])
);

INVX1 _9465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [1]),
    .Y(_1304_)
);

NAND2X1 _9466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf3 ),
    .Y(_1305_)
);

OAI21X1 _9467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1304_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1305_),
    .Y(_1303_[1])
);

INVX1 _9468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [2]),
    .Y(_1306_)
);

NAND2X1 _9469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf3 ),
    .Y(_1307_)
);

OAI21X1 _9470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1306_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1307_),
    .Y(_1303_[2])
);

INVX1 _9471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [3]),
    .Y(_1308_)
);

NAND2X1 _9472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf3 ),
    .Y(_1309_)
);

OAI21X1 _9473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1308_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1309_),
    .Y(_1303_[3])
);

INVX1 _9474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [4]),
    .Y(_1310_)
);

NAND2X1 _9475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf3 ),
    .Y(_1311_)
);

OAI21X1 _9476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1310_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1311_),
    .Y(_1303_[4])
);

INVX1 _9477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [5]),
    .Y(_1312_)
);

NAND2X1 _9478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf3 ),
    .Y(_1313_)
);

OAI21X1 _9479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1312_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1313_),
    .Y(_1303_[5])
);

INVX1 _9480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [6]),
    .Y(_1314_)
);

NAND2X1 _9481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf3 ),
    .Y(_1315_)
);

OAI21X1 _9482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1314_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1315_),
    .Y(_1303_[6])
);

INVX1 _9483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [7]),
    .Y(_1316_)
);

NAND2X1 _9484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf3 ),
    .Y(_1317_)
);

OAI21X1 _9485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1317_),
    .Y(_1303_[7])
);

INVX1 _9486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [8]),
    .Y(_1318_)
);

NAND2X1 _9487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf3 ),
    .Y(_1319_)
);

OAI21X1 _9488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1318_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1319_),
    .Y(_1303_[8])
);

INVX1 _9489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [9]),
    .Y(_1320_)
);

NAND2X1 _9490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf2 ),
    .Y(_1321_)
);

OAI21X1 _9491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1320_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1321_),
    .Y(_1303_[9])
);

INVX1 _9492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [10]),
    .Y(_1322_)
);

NAND2X1 _9493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf2 ),
    .Y(_1323_)
);

OAI21X1 _9494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1322_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1323_),
    .Y(_1303_[10])
);

INVX1 _9495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [11]),
    .Y(_1324_)
);

NAND2X1 _9496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf2 ),
    .Y(_1325_)
);

OAI21X1 _9497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1325_),
    .Y(_1303_[11])
);

INVX1 _9498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [12]),
    .Y(_1326_)
);

NAND2X1 _9499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf2 ),
    .Y(_1327_)
);

OAI21X1 _9500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1327_),
    .Y(_1303_[12])
);

INVX1 _9501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [13]),
    .Y(_1328_)
);

NAND2X1 _9502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf2 ),
    .Y(_1329_)
);

OAI21X1 _9503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1328_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1329_),
    .Y(_1303_[13])
);

INVX1 _9504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [14]),
    .Y(_1330_)
);

NAND2X1 _9505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf2 ),
    .Y(_1331_)
);

OAI21X1 _9506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1330_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1331_),
    .Y(_1303_[14])
);

INVX1 _9507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [15]),
    .Y(_1332_)
);

NAND2X1 _9508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf2 ),
    .Y(_1333_)
);

OAI21X1 _9509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1332_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1333_),
    .Y(_1303_[15])
);

INVX1 _9510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [16]),
    .Y(_1334_)
);

NAND2X1 _9511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf2 ),
    .Y(_1335_)
);

OAI21X1 _9512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1335_),
    .Y(_1303_[16])
);

INVX1 _9513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [17]),
    .Y(_1336_)
);

NAND2X1 _9514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf2 ),
    .Y(_1337_)
);

OAI21X1 _9515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1336_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1337_),
    .Y(_1303_[17])
);

INVX1 _9516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [18]),
    .Y(_1338_)
);

NAND2X1 _9517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf2 ),
    .Y(_1339_)
);

OAI21X1 _9518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1338_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1339_),
    .Y(_1303_[18])
);

INVX1 _9519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [19]),
    .Y(_1340_)
);

NAND2X1 _9520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf2 ),
    .Y(_1341_)
);

OAI21X1 _9521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1340_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1341_),
    .Y(_1303_[19])
);

INVX1 _9522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [20]),
    .Y(_1342_)
);

NAND2X1 _9523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf2 ),
    .Y(_1343_)
);

OAI21X1 _9524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1343_),
    .Y(_1303_[20])
);

INVX1 _9525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [21]),
    .Y(_1344_)
);

NAND2X1 _9526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf2 ),
    .Y(_1345_)
);

OAI21X1 _9527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1344_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1345_),
    .Y(_1303_[21])
);

INVX1 _9528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [22]),
    .Y(_1346_)
);

NAND2X1 _9529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf2 ),
    .Y(_1347_)
);

OAI21X1 _9530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1346_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1347_),
    .Y(_1303_[22])
);

INVX1 _9531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [23]),
    .Y(_1348_)
);

NAND2X1 _9532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf2 ),
    .Y(_1349_)
);

OAI21X1 _9533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1348_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1349_),
    .Y(_1303_[23])
);

INVX1 _9534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [24]),
    .Y(_1350_)
);

NAND2X1 _9535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf2 ),
    .Y(_1351_)
);

OAI21X1 _9536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1351_),
    .Y(_1303_[24])
);

INVX1 _9537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [25]),
    .Y(_1352_)
);

NAND2X1 _9538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf2 ),
    .Y(_1353_)
);

OAI21X1 _9539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1353_),
    .Y(_1303_[25])
);

INVX1 _9540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [26]),
    .Y(_1354_)
);

NAND2X1 _9541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf2 ),
    .Y(_1355_)
);

OAI21X1 _9542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1355_),
    .Y(_1303_[26])
);

INVX1 _9543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [27]),
    .Y(_1356_)
);

NAND2X1 _9544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf2 ),
    .Y(_1357_)
);

OAI21X1 _9545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1357_),
    .Y(_1303_[27])
);

INVX1 _9546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [28]),
    .Y(_1358_)
);

NAND2X1 _9547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf2 ),
    .Y(_1359_)
);

OAI21X1 _9548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf6 ),
    .C(_1359_),
    .Y(_1303_[28])
);

INVX1 _9549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [29]),
    .Y(_1360_)
);

NAND2X1 _9550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf2 ),
    .Y(_1361_)
);

OAI21X1 _9551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1360_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf4 ),
    .C(_1361_),
    .Y(_1303_[29])
);

INVX1 _9552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [30]),
    .Y(_1362_)
);

NAND2X1 _9553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf2 ),
    .Y(_1363_)
);

OAI21X1 _9554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf2 ),
    .C(_1363_),
    .Y(_1303_[30])
);

INVX1 _9555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[21] [31]),
    .Y(_1364_)
);

NAND2X1 _9556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_21_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf2 ),
    .Y(_1365_)
);

OAI21X1 _9557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1364_),
    .B(\datapath_1.regfile_1.regEn_21_bF$buf0 ),
    .C(_1365_),
    .Y(_1303_[31])
);

DFFSR _9558_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_1303_[0]),
    .Q(\datapath_1.regfile_1.regOut[21] [0]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _9559_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_1303_[1]),
    .Q(\datapath_1.regfile_1.regOut[21] [1]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _9560_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_1303_[2]),
    .Q(\datapath_1.regfile_1.regOut[21] [2]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _9561_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_1303_[3]),
    .Q(\datapath_1.regfile_1.regOut[21] [3]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _9562_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_1303_[4]),
    .Q(\datapath_1.regfile_1.regOut[21] [4]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _9563_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_1303_[5]),
    .Q(\datapath_1.regfile_1.regOut[21] [5]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _9564_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_1303_[6]),
    .Q(\datapath_1.regfile_1.regOut[21] [6]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _9565_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_1303_[7]),
    .Q(\datapath_1.regfile_1.regOut[21] [7]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _9566_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_1303_[8]),
    .Q(\datapath_1.regfile_1.regOut[21] [8]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _9567_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_1303_[9]),
    .Q(\datapath_1.regfile_1.regOut[21] [9]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _9568_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_1303_[10]),
    .Q(\datapath_1.regfile_1.regOut[21] [10]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _9569_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_1303_[11]),
    .Q(\datapath_1.regfile_1.regOut[21] [11]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _9570_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_1303_[12]),
    .Q(\datapath_1.regfile_1.regOut[21] [12]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _9571_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_1303_[13]),
    .Q(\datapath_1.regfile_1.regOut[21] [13]),
    .R(rst_bF$buf34),
    .S(vdd)
);

DFFSR _9572_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf33),
    .D(_1303_[14]),
    .Q(\datapath_1.regfile_1.regOut[21] [14]),
    .R(rst_bF$buf33),
    .S(vdd)
);

DFFSR _9573_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf32),
    .D(_1303_[15]),
    .Q(\datapath_1.regfile_1.regOut[21] [15]),
    .R(rst_bF$buf32),
    .S(vdd)
);

DFFSR _9574_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf31),
    .D(_1303_[16]),
    .Q(\datapath_1.regfile_1.regOut[21] [16]),
    .R(rst_bF$buf31),
    .S(vdd)
);

DFFSR _9575_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf30),
    .D(_1303_[17]),
    .Q(\datapath_1.regfile_1.regOut[21] [17]),
    .R(rst_bF$buf30),
    .S(vdd)
);

DFFSR _9576_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf29),
    .D(_1303_[18]),
    .Q(\datapath_1.regfile_1.regOut[21] [18]),
    .R(rst_bF$buf29),
    .S(vdd)
);

DFFSR _9577_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf28),
    .D(_1303_[19]),
    .Q(\datapath_1.regfile_1.regOut[21] [19]),
    .R(rst_bF$buf28),
    .S(vdd)
);

DFFSR _9578_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf27),
    .D(_1303_[20]),
    .Q(\datapath_1.regfile_1.regOut[21] [20]),
    .R(rst_bF$buf27),
    .S(vdd)
);

DFFSR _9579_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf26),
    .D(_1303_[21]),
    .Q(\datapath_1.regfile_1.regOut[21] [21]),
    .R(rst_bF$buf26),
    .S(vdd)
);

DFFSR _9580_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf25),
    .D(_1303_[22]),
    .Q(\datapath_1.regfile_1.regOut[21] [22]),
    .R(rst_bF$buf25),
    .S(vdd)
);

DFFSR _9581_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf24),
    .D(_1303_[23]),
    .Q(\datapath_1.regfile_1.regOut[21] [23]),
    .R(rst_bF$buf24),
    .S(vdd)
);

DFFSR _9582_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf23),
    .D(_1303_[24]),
    .Q(\datapath_1.regfile_1.regOut[21] [24]),
    .R(rst_bF$buf23),
    .S(vdd)
);

DFFSR _9583_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf22),
    .D(_1303_[25]),
    .Q(\datapath_1.regfile_1.regOut[21] [25]),
    .R(rst_bF$buf22),
    .S(vdd)
);

DFFSR _9584_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf21),
    .D(_1303_[26]),
    .Q(\datapath_1.regfile_1.regOut[21] [26]),
    .R(rst_bF$buf21),
    .S(vdd)
);

DFFSR _9585_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf20),
    .D(_1303_[27]),
    .Q(\datapath_1.regfile_1.regOut[21] [27]),
    .R(rst_bF$buf20),
    .S(vdd)
);

DFFSR _9586_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf19),
    .D(_1303_[28]),
    .Q(\datapath_1.regfile_1.regOut[21] [28]),
    .R(rst_bF$buf19),
    .S(vdd)
);

DFFSR _9587_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf18),
    .D(_1303_[29]),
    .Q(\datapath_1.regfile_1.regOut[21] [29]),
    .R(rst_bF$buf18),
    .S(vdd)
);

DFFSR _9588_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf17),
    .D(_1303_[30]),
    .Q(\datapath_1.regfile_1.regOut[21] [30]),
    .R(rst_bF$buf17),
    .S(vdd)
);

DFFSR _9589_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf16),
    .D(_1303_[31]),
    .Q(\datapath_1.regfile_1.regOut[21] [31]),
    .R(rst_bF$buf16),
    .S(vdd)
);

INVX1 _9590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [0]),
    .Y(_1431_)
);

NAND2X1 _9591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf2 ),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .Y(_1432_)
);

OAI21X1 _9592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1431_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1432_),
    .Y(_1368_[0])
);

INVX1 _9593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [1]),
    .Y(_1369_)
);

NAND2X1 _9594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf2 ),
    .Y(_1370_)
);

OAI21X1 _9595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1370_),
    .Y(_1368_[1])
);

INVX1 _9596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [2]),
    .Y(_1371_)
);

NAND2X1 _9597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf2 ),
    .Y(_1372_)
);

OAI21X1 _9598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1372_),
    .Y(_1368_[2])
);

INVX1 _9599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [3]),
    .Y(_1373_)
);

NAND2X1 _9600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf2 ),
    .Y(_1374_)
);

OAI21X1 _9601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1373_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1374_),
    .Y(_1368_[3])
);

INVX1 _9602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [4]),
    .Y(_1375_)
);

NAND2X1 _9603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf2 ),
    .Y(_1376_)
);

OAI21X1 _9604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1375_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1376_),
    .Y(_1368_[4])
);

INVX1 _9605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [5]),
    .Y(_1377_)
);

NAND2X1 _9606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf2 ),
    .Y(_1378_)
);

OAI21X1 _9607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1377_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1378_),
    .Y(_1368_[5])
);

INVX1 _9608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [6]),
    .Y(_1379_)
);

NAND2X1 _9609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf2 ),
    .Y(_1380_)
);

OAI21X1 _9610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1379_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1380_),
    .Y(_1368_[6])
);

INVX1 _9611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [7]),
    .Y(_1381_)
);

NAND2X1 _9612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf2 ),
    .Y(_1382_)
);

OAI21X1 _9613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1381_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1382_),
    .Y(_1368_[7])
);

INVX1 _9614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [8]),
    .Y(_1383_)
);

NAND2X1 _9615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf2 ),
    .Y(_1384_)
);

OAI21X1 _9616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1384_),
    .Y(_1368_[8])
);

INVX1 _9617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [9]),
    .Y(_1385_)
);

NAND2X1 _9618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf1 ),
    .Y(_1386_)
);

OAI21X1 _9619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1386_),
    .Y(_1368_[9])
);

INVX1 _9620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [10]),
    .Y(_1387_)
);

NAND2X1 _9621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf1 ),
    .Y(_1388_)
);

OAI21X1 _9622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1387_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1388_),
    .Y(_1368_[10])
);

INVX1 _9623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [11]),
    .Y(_1389_)
);

NAND2X1 _9624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf1 ),
    .Y(_1390_)
);

OAI21X1 _9625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1389_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1390_),
    .Y(_1368_[11])
);

INVX1 _9626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [12]),
    .Y(_1391_)
);

NAND2X1 _9627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf1 ),
    .Y(_1392_)
);

OAI21X1 _9628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1391_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1392_),
    .Y(_1368_[12])
);

INVX1 _9629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [13]),
    .Y(_1393_)
);

NAND2X1 _9630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf1 ),
    .Y(_1394_)
);

OAI21X1 _9631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1393_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1394_),
    .Y(_1368_[13])
);

INVX1 _9632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [14]),
    .Y(_1395_)
);

NAND2X1 _9633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf1 ),
    .Y(_1396_)
);

OAI21X1 _9634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1395_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1396_),
    .Y(_1368_[14])
);

INVX1 _9635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [15]),
    .Y(_1397_)
);

NAND2X1 _9636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf1 ),
    .Y(_1398_)
);

OAI21X1 _9637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1397_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1398_),
    .Y(_1368_[15])
);

INVX1 _9638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [16]),
    .Y(_1399_)
);

NAND2X1 _9639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf1 ),
    .Y(_1400_)
);

OAI21X1 _9640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1399_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1400_),
    .Y(_1368_[16])
);

INVX1 _9641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [17]),
    .Y(_1401_)
);

NAND2X1 _9642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf1 ),
    .Y(_1402_)
);

OAI21X1 _9643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1401_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1402_),
    .Y(_1368_[17])
);

INVX1 _9644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [18]),
    .Y(_1403_)
);

NAND2X1 _9645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf1 ),
    .Y(_1404_)
);

OAI21X1 _9646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1404_),
    .Y(_1368_[18])
);

INVX1 _9647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [19]),
    .Y(_1405_)
);

NAND2X1 _9648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf1 ),
    .Y(_1406_)
);

OAI21X1 _9649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1406_),
    .Y(_1368_[19])
);

INVX1 _9650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [20]),
    .Y(_1407_)
);

NAND2X1 _9651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf1 ),
    .Y(_1408_)
);

OAI21X1 _9652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1407_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1408_),
    .Y(_1368_[20])
);

INVX1 _9653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [21]),
    .Y(_1409_)
);

NAND2X1 _9654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf1 ),
    .Y(_1410_)
);

OAI21X1 _9655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1409_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1410_),
    .Y(_1368_[21])
);

INVX1 _9656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [22]),
    .Y(_1411_)
);

NAND2X1 _9657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf1 ),
    .Y(_1412_)
);

OAI21X1 _9658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1411_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1412_),
    .Y(_1368_[22])
);

INVX1 _9659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [23]),
    .Y(_1413_)
);

NAND2X1 _9660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf1 ),
    .Y(_1414_)
);

OAI21X1 _9661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1413_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1414_),
    .Y(_1368_[23])
);

INVX1 _9662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [24]),
    .Y(_1415_)
);

NAND2X1 _9663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf1 ),
    .Y(_1416_)
);

OAI21X1 _9664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1416_),
    .Y(_1368_[24])
);

INVX1 _9665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [25]),
    .Y(_1417_)
);

NAND2X1 _9666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf1 ),
    .Y(_1418_)
);

OAI21X1 _9667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1417_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1418_),
    .Y(_1368_[25])
);

INVX1 _9668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [26]),
    .Y(_1419_)
);

NAND2X1 _9669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf1 ),
    .Y(_1420_)
);

OAI21X1 _9670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1419_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1420_),
    .Y(_1368_[26])
);

INVX1 _9671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [27]),
    .Y(_1421_)
);

NAND2X1 _9672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf1 ),
    .Y(_1422_)
);

OAI21X1 _9673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1421_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1422_),
    .Y(_1368_[27])
);

INVX1 _9674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [28]),
    .Y(_1423_)
);

NAND2X1 _9675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf1 ),
    .Y(_1424_)
);

OAI21X1 _9676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1423_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf6 ),
    .C(_1424_),
    .Y(_1368_[28])
);

INVX1 _9677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [29]),
    .Y(_1425_)
);

NAND2X1 _9678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf1 ),
    .Y(_1426_)
);

OAI21X1 _9679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1425_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf4 ),
    .C(_1426_),
    .Y(_1368_[29])
);

INVX1 _9680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [30]),
    .Y(_1427_)
);

NAND2X1 _9681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf1 ),
    .Y(_1428_)
);

OAI21X1 _9682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1427_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf2 ),
    .C(_1428_),
    .Y(_1368_[30])
);

INVX1 _9683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[22] [31]),
    .Y(_1429_)
);

NAND2X1 _9684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_22_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf1 ),
    .Y(_1430_)
);

OAI21X1 _9685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1429_),
    .B(\datapath_1.regfile_1.regEn_22_bF$buf0 ),
    .C(_1430_),
    .Y(_1368_[31])
);

DFFSR _9686_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf15),
    .D(_1368_[0]),
    .Q(\datapath_1.regfile_1.regOut[22] [0]),
    .R(rst_bF$buf15),
    .S(vdd)
);

DFFSR _9687_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf14),
    .D(_1368_[1]),
    .Q(\datapath_1.regfile_1.regOut[22] [1]),
    .R(rst_bF$buf14),
    .S(vdd)
);

DFFSR _9688_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf13),
    .D(_1368_[2]),
    .Q(\datapath_1.regfile_1.regOut[22] [2]),
    .R(rst_bF$buf13),
    .S(vdd)
);

DFFSR _9689_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf12),
    .D(_1368_[3]),
    .Q(\datapath_1.regfile_1.regOut[22] [3]),
    .R(rst_bF$buf12),
    .S(vdd)
);

DFFSR _9690_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf11),
    .D(_1368_[4]),
    .Q(\datapath_1.regfile_1.regOut[22] [4]),
    .R(rst_bF$buf11),
    .S(vdd)
);

DFFSR _9691_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf10),
    .D(_1368_[5]),
    .Q(\datapath_1.regfile_1.regOut[22] [5]),
    .R(rst_bF$buf10),
    .S(vdd)
);

DFFSR _9692_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(_1368_[6]),
    .Q(\datapath_1.regfile_1.regOut[22] [6]),
    .R(rst_bF$buf9),
    .S(vdd)
);

DFFSR _9693_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_1368_[7]),
    .Q(\datapath_1.regfile_1.regOut[22] [7]),
    .R(rst_bF$buf8),
    .S(vdd)
);

DFFSR _9694_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1368_[8]),
    .Q(\datapath_1.regfile_1.regOut[22] [8]),
    .R(rst_bF$buf7),
    .S(vdd)
);

DFFSR _9695_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1368_[9]),
    .Q(\datapath_1.regfile_1.regOut[22] [9]),
    .R(rst_bF$buf6),
    .S(vdd)
);

DFFSR _9696_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1368_[10]),
    .Q(\datapath_1.regfile_1.regOut[22] [10]),
    .R(rst_bF$buf5),
    .S(vdd)
);

DFFSR _9697_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1368_[11]),
    .Q(\datapath_1.regfile_1.regOut[22] [11]),
    .R(rst_bF$buf4),
    .S(vdd)
);

DFFSR _9698_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1368_[12]),
    .Q(\datapath_1.regfile_1.regOut[22] [12]),
    .R(rst_bF$buf3),
    .S(vdd)
);

DFFSR _9699_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1368_[13]),
    .Q(\datapath_1.regfile_1.regOut[22] [13]),
    .R(rst_bF$buf2),
    .S(vdd)
);

DFFSR _9700_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1368_[14]),
    .Q(\datapath_1.regfile_1.regOut[22] [14]),
    .R(rst_bF$buf1),
    .S(vdd)
);

DFFSR _9701_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1368_[15]),
    .Q(\datapath_1.regfile_1.regOut[22] [15]),
    .R(rst_bF$buf0),
    .S(vdd)
);

DFFSR _9702_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf113),
    .D(_1368_[16]),
    .Q(\datapath_1.regfile_1.regOut[22] [16]),
    .R(rst_bF$buf113),
    .S(vdd)
);

DFFSR _9703_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf112),
    .D(_1368_[17]),
    .Q(\datapath_1.regfile_1.regOut[22] [17]),
    .R(rst_bF$buf112),
    .S(vdd)
);

DFFSR _9704_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf111),
    .D(_1368_[18]),
    .Q(\datapath_1.regfile_1.regOut[22] [18]),
    .R(rst_bF$buf111),
    .S(vdd)
);

DFFSR _9705_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf110),
    .D(_1368_[19]),
    .Q(\datapath_1.regfile_1.regOut[22] [19]),
    .R(rst_bF$buf110),
    .S(vdd)
);

DFFSR _9706_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf109),
    .D(_1368_[20]),
    .Q(\datapath_1.regfile_1.regOut[22] [20]),
    .R(rst_bF$buf109),
    .S(vdd)
);

DFFSR _9707_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf108),
    .D(_1368_[21]),
    .Q(\datapath_1.regfile_1.regOut[22] [21]),
    .R(rst_bF$buf108),
    .S(vdd)
);

DFFSR _9708_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf107),
    .D(_1368_[22]),
    .Q(\datapath_1.regfile_1.regOut[22] [22]),
    .R(rst_bF$buf107),
    .S(vdd)
);

DFFSR _9709_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf106),
    .D(_1368_[23]),
    .Q(\datapath_1.regfile_1.regOut[22] [23]),
    .R(rst_bF$buf106),
    .S(vdd)
);

DFFSR _9710_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf105),
    .D(_1368_[24]),
    .Q(\datapath_1.regfile_1.regOut[22] [24]),
    .R(rst_bF$buf105),
    .S(vdd)
);

DFFSR _9711_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf104),
    .D(_1368_[25]),
    .Q(\datapath_1.regfile_1.regOut[22] [25]),
    .R(rst_bF$buf104),
    .S(vdd)
);

DFFSR _9712_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf103),
    .D(_1368_[26]),
    .Q(\datapath_1.regfile_1.regOut[22] [26]),
    .R(rst_bF$buf103),
    .S(vdd)
);

DFFSR _9713_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf102),
    .D(_1368_[27]),
    .Q(\datapath_1.regfile_1.regOut[22] [27]),
    .R(rst_bF$buf102),
    .S(vdd)
);

DFFSR _9714_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf101),
    .D(_1368_[28]),
    .Q(\datapath_1.regfile_1.regOut[22] [28]),
    .R(rst_bF$buf101),
    .S(vdd)
);

DFFSR _9715_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf100),
    .D(_1368_[29]),
    .Q(\datapath_1.regfile_1.regOut[22] [29]),
    .R(rst_bF$buf100),
    .S(vdd)
);

DFFSR _9716_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf99),
    .D(_1368_[30]),
    .Q(\datapath_1.regfile_1.regOut[22] [30]),
    .R(rst_bF$buf99),
    .S(vdd)
);

DFFSR _9717_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf98),
    .D(_1368_[31]),
    .Q(\datapath_1.regfile_1.regOut[22] [31]),
    .R(rst_bF$buf98),
    .S(vdd)
);

INVX1 _9718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [0]),
    .Y(_1496_)
);

NAND2X1 _9719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf1 ),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .Y(_1497_)
);

OAI21X1 _9720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1497_),
    .Y(_1433_[0])
);

INVX1 _9721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [1]),
    .Y(_1434_)
);

NAND2X1 _9722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf1 ),
    .Y(_1435_)
);

OAI21X1 _9723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1434_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1435_),
    .Y(_1433_[1])
);

INVX1 _9724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [2]),
    .Y(_1436_)
);

NAND2X1 _9725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf1 ),
    .Y(_1437_)
);

OAI21X1 _9726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1436_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1437_),
    .Y(_1433_[2])
);

INVX1 _9727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [3]),
    .Y(_1438_)
);

NAND2X1 _9728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf1 ),
    .Y(_1439_)
);

OAI21X1 _9729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1438_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1439_),
    .Y(_1433_[3])
);

INVX1 _9730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [4]),
    .Y(_1440_)
);

NAND2X1 _9731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf1 ),
    .Y(_1441_)
);

OAI21X1 _9732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1441_),
    .Y(_1433_[4])
);

INVX1 _9733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [5]),
    .Y(_1442_)
);

NAND2X1 _9734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf1 ),
    .Y(_1443_)
);

OAI21X1 _9735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1442_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1443_),
    .Y(_1433_[5])
);

INVX1 _9736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [6]),
    .Y(_1444_)
);

NAND2X1 _9737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf1 ),
    .Y(_1445_)
);

OAI21X1 _9738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1444_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1445_),
    .Y(_1433_[6])
);

INVX1 _9739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [7]),
    .Y(_1446_)
);

NAND2X1 _9740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf1 ),
    .Y(_1447_)
);

OAI21X1 _9741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1446_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1447_),
    .Y(_1433_[7])
);

INVX1 _9742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [8]),
    .Y(_1448_)
);

NAND2X1 _9743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf1 ),
    .Y(_1449_)
);

OAI21X1 _9744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1449_),
    .Y(_1433_[8])
);

INVX1 _9745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [9]),
    .Y(_1450_)
);

NAND2X1 _9746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf0 ),
    .Y(_1451_)
);

OAI21X1 _9747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1450_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1451_),
    .Y(_1433_[9])
);

INVX1 _9748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [10]),
    .Y(_1452_)
);

NAND2X1 _9749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf0 ),
    .Y(_1453_)
);

OAI21X1 _9750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1452_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1453_),
    .Y(_1433_[10])
);

INVX1 _9751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [11]),
    .Y(_1454_)
);

NAND2X1 _9752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf0 ),
    .Y(_1455_)
);

OAI21X1 _9753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1454_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1455_),
    .Y(_1433_[11])
);

INVX1 _9754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [12]),
    .Y(_1456_)
);

NAND2X1 _9755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf0 ),
    .Y(_1457_)
);

OAI21X1 _9756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1456_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1457_),
    .Y(_1433_[12])
);

INVX1 _9757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [13]),
    .Y(_1458_)
);

NAND2X1 _9758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf0 ),
    .Y(_1459_)
);

OAI21X1 _9759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1458_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1459_),
    .Y(_1433_[13])
);

INVX1 _9760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [14]),
    .Y(_1460_)
);

NAND2X1 _9761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf0 ),
    .Y(_1461_)
);

OAI21X1 _9762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1461_),
    .Y(_1433_[14])
);

INVX1 _9763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [15]),
    .Y(_1462_)
);

NAND2X1 _9764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf0 ),
    .Y(_1463_)
);

OAI21X1 _9765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1462_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1463_),
    .Y(_1433_[15])
);

INVX1 _9766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [16]),
    .Y(_1464_)
);

NAND2X1 _9767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf0 ),
    .Y(_1465_)
);

OAI21X1 _9768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1464_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1465_),
    .Y(_1433_[16])
);

INVX1 _9769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [17]),
    .Y(_1466_)
);

NAND2X1 _9770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf0 ),
    .Y(_1467_)
);

OAI21X1 _9771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1466_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1467_),
    .Y(_1433_[17])
);

INVX1 _9772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [18]),
    .Y(_1468_)
);

NAND2X1 _9773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf0 ),
    .Y(_1469_)
);

OAI21X1 _9774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1468_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1469_),
    .Y(_1433_[18])
);

INVX1 _9775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [19]),
    .Y(_1470_)
);

NAND2X1 _9776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf0 ),
    .Y(_1471_)
);

OAI21X1 _9777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1470_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1471_),
    .Y(_1433_[19])
);

INVX1 _9778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [20]),
    .Y(_1472_)
);

NAND2X1 _9779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf0 ),
    .Y(_1473_)
);

OAI21X1 _9780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1472_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1473_),
    .Y(_1433_[20])
);

INVX1 _9781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [21]),
    .Y(_1474_)
);

NAND2X1 _9782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf0 ),
    .Y(_1475_)
);

OAI21X1 _9783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1474_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1475_),
    .Y(_1433_[21])
);

INVX1 _9784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [22]),
    .Y(_1476_)
);

NAND2X1 _9785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf0 ),
    .Y(_1477_)
);

OAI21X1 _9786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1477_),
    .Y(_1433_[22])
);

INVX1 _9787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [23]),
    .Y(_1478_)
);

NAND2X1 _9788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf0 ),
    .Y(_1479_)
);

OAI21X1 _9789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1478_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1479_),
    .Y(_1433_[23])
);

INVX1 _9790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [24]),
    .Y(_1480_)
);

NAND2X1 _9791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf0 ),
    .Y(_1481_)
);

OAI21X1 _9792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1480_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1481_),
    .Y(_1433_[24])
);

INVX1 _9793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [25]),
    .Y(_1482_)
);

NAND2X1 _9794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf0 ),
    .Y(_1483_)
);

OAI21X1 _9795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1482_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1483_),
    .Y(_1433_[25])
);

INVX1 _9796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [26]),
    .Y(_1484_)
);

NAND2X1 _9797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf0 ),
    .Y(_1485_)
);

OAI21X1 _9798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1484_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1485_),
    .Y(_1433_[26])
);

INVX1 _9799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [27]),
    .Y(_1486_)
);

NAND2X1 _9800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf0 ),
    .Y(_1487_)
);

OAI21X1 _9801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1486_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1487_),
    .Y(_1433_[27])
);

INVX1 _9802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [28]),
    .Y(_1488_)
);

NAND2X1 _9803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf0 ),
    .Y(_1489_)
);

OAI21X1 _9804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1488_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf6 ),
    .C(_1489_),
    .Y(_1433_[28])
);

INVX1 _9805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [29]),
    .Y(_1490_)
);

NAND2X1 _9806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf0 ),
    .Y(_1491_)
);

OAI21X1 _9807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf4 ),
    .C(_1491_),
    .Y(_1433_[29])
);

INVX1 _9808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [30]),
    .Y(_1492_)
);

NAND2X1 _9809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf0 ),
    .Y(_1493_)
);

OAI21X1 _9810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1492_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf2 ),
    .C(_1493_),
    .Y(_1433_[30])
);

INVX1 _9811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[23] [31]),
    .Y(_1494_)
);

NAND2X1 _9812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_23_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf0 ),
    .Y(_1495_)
);

OAI21X1 _9813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1494_),
    .B(\datapath_1.regfile_1.regEn_23_bF$buf0 ),
    .C(_1495_),
    .Y(_1433_[31])
);

DFFSR _9814_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf97),
    .D(_1433_[0]),
    .Q(\datapath_1.regfile_1.regOut[23] [0]),
    .R(rst_bF$buf97),
    .S(vdd)
);

DFFSR _9815_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf96),
    .D(_1433_[1]),
    .Q(\datapath_1.regfile_1.regOut[23] [1]),
    .R(rst_bF$buf96),
    .S(vdd)
);

DFFSR _9816_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf95),
    .D(_1433_[2]),
    .Q(\datapath_1.regfile_1.regOut[23] [2]),
    .R(rst_bF$buf95),
    .S(vdd)
);

DFFSR _9817_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf94),
    .D(_1433_[3]),
    .Q(\datapath_1.regfile_1.regOut[23] [3]),
    .R(rst_bF$buf94),
    .S(vdd)
);

DFFSR _9818_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf93),
    .D(_1433_[4]),
    .Q(\datapath_1.regfile_1.regOut[23] [4]),
    .R(rst_bF$buf93),
    .S(vdd)
);

DFFSR _9819_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf92),
    .D(_1433_[5]),
    .Q(\datapath_1.regfile_1.regOut[23] [5]),
    .R(rst_bF$buf92),
    .S(vdd)
);

DFFSR _9820_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf91),
    .D(_1433_[6]),
    .Q(\datapath_1.regfile_1.regOut[23] [6]),
    .R(rst_bF$buf91),
    .S(vdd)
);

DFFSR _9821_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf90),
    .D(_1433_[7]),
    .Q(\datapath_1.regfile_1.regOut[23] [7]),
    .R(rst_bF$buf90),
    .S(vdd)
);

DFFSR _9822_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf89),
    .D(_1433_[8]),
    .Q(\datapath_1.regfile_1.regOut[23] [8]),
    .R(rst_bF$buf89),
    .S(vdd)
);

DFFSR _9823_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf88),
    .D(_1433_[9]),
    .Q(\datapath_1.regfile_1.regOut[23] [9]),
    .R(rst_bF$buf88),
    .S(vdd)
);

DFFSR _9824_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf87),
    .D(_1433_[10]),
    .Q(\datapath_1.regfile_1.regOut[23] [10]),
    .R(rst_bF$buf87),
    .S(vdd)
);

DFFSR _9825_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf86),
    .D(_1433_[11]),
    .Q(\datapath_1.regfile_1.regOut[23] [11]),
    .R(rst_bF$buf86),
    .S(vdd)
);

DFFSR _9826_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf85),
    .D(_1433_[12]),
    .Q(\datapath_1.regfile_1.regOut[23] [12]),
    .R(rst_bF$buf85),
    .S(vdd)
);

DFFSR _9827_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf84),
    .D(_1433_[13]),
    .Q(\datapath_1.regfile_1.regOut[23] [13]),
    .R(rst_bF$buf84),
    .S(vdd)
);

DFFSR _9828_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf83),
    .D(_1433_[14]),
    .Q(\datapath_1.regfile_1.regOut[23] [14]),
    .R(rst_bF$buf83),
    .S(vdd)
);

DFFSR _9829_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf82),
    .D(_1433_[15]),
    .Q(\datapath_1.regfile_1.regOut[23] [15]),
    .R(rst_bF$buf82),
    .S(vdd)
);

DFFSR _9830_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf81),
    .D(_1433_[16]),
    .Q(\datapath_1.regfile_1.regOut[23] [16]),
    .R(rst_bF$buf81),
    .S(vdd)
);

DFFSR _9831_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf80),
    .D(_1433_[17]),
    .Q(\datapath_1.regfile_1.regOut[23] [17]),
    .R(rst_bF$buf80),
    .S(vdd)
);

DFFSR _9832_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf79),
    .D(_1433_[18]),
    .Q(\datapath_1.regfile_1.regOut[23] [18]),
    .R(rst_bF$buf79),
    .S(vdd)
);

DFFSR _9833_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf78),
    .D(_1433_[19]),
    .Q(\datapath_1.regfile_1.regOut[23] [19]),
    .R(rst_bF$buf78),
    .S(vdd)
);

DFFSR _9834_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf77),
    .D(_1433_[20]),
    .Q(\datapath_1.regfile_1.regOut[23] [20]),
    .R(rst_bF$buf77),
    .S(vdd)
);

DFFSR _9835_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf76),
    .D(_1433_[21]),
    .Q(\datapath_1.regfile_1.regOut[23] [21]),
    .R(rst_bF$buf76),
    .S(vdd)
);

DFFSR _9836_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf75),
    .D(_1433_[22]),
    .Q(\datapath_1.regfile_1.regOut[23] [22]),
    .R(rst_bF$buf75),
    .S(vdd)
);

DFFSR _9837_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf74),
    .D(_1433_[23]),
    .Q(\datapath_1.regfile_1.regOut[23] [23]),
    .R(rst_bF$buf74),
    .S(vdd)
);

DFFSR _9838_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf73),
    .D(_1433_[24]),
    .Q(\datapath_1.regfile_1.regOut[23] [24]),
    .R(rst_bF$buf73),
    .S(vdd)
);

DFFSR _9839_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf72),
    .D(_1433_[25]),
    .Q(\datapath_1.regfile_1.regOut[23] [25]),
    .R(rst_bF$buf72),
    .S(vdd)
);

DFFSR _9840_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf71),
    .D(_1433_[26]),
    .Q(\datapath_1.regfile_1.regOut[23] [26]),
    .R(rst_bF$buf71),
    .S(vdd)
);

DFFSR _9841_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf70),
    .D(_1433_[27]),
    .Q(\datapath_1.regfile_1.regOut[23] [27]),
    .R(rst_bF$buf70),
    .S(vdd)
);

DFFSR _9842_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf69),
    .D(_1433_[28]),
    .Q(\datapath_1.regfile_1.regOut[23] [28]),
    .R(rst_bF$buf69),
    .S(vdd)
);

DFFSR _9843_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf68),
    .D(_1433_[29]),
    .Q(\datapath_1.regfile_1.regOut[23] [29]),
    .R(rst_bF$buf68),
    .S(vdd)
);

DFFSR _9844_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf67),
    .D(_1433_[30]),
    .Q(\datapath_1.regfile_1.regOut[23] [30]),
    .R(rst_bF$buf67),
    .S(vdd)
);

DFFSR _9845_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf66),
    .D(_1433_[31]),
    .Q(\datapath_1.regfile_1.regOut[23] [31]),
    .R(rst_bF$buf66),
    .S(vdd)
);

INVX1 _9846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [0]),
    .Y(_1561_)
);

NAND2X1 _9847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf0 ),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .Y(_1562_)
);

OAI21X1 _9848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1561_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1562_),
    .Y(_1498_[0])
);

INVX1 _9849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [1]),
    .Y(_1499_)
);

NAND2X1 _9850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf0 ),
    .Y(_1500_)
);

OAI21X1 _9851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1499_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1500_),
    .Y(_1498_[1])
);

INVX1 _9852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [2]),
    .Y(_1501_)
);

NAND2X1 _9853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf0 ),
    .Y(_1502_)
);

OAI21X1 _9854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1502_),
    .Y(_1498_[2])
);

INVX1 _9855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [3]),
    .Y(_1503_)
);

NAND2X1 _9856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf0 ),
    .Y(_1504_)
);

OAI21X1 _9857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1503_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1504_),
    .Y(_1498_[3])
);

INVX1 _9858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [4]),
    .Y(_1505_)
);

NAND2X1 _9859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf0 ),
    .Y(_1506_)
);

OAI21X1 _9860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1505_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1506_),
    .Y(_1498_[4])
);

INVX1 _9861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [5]),
    .Y(_1507_)
);

NAND2X1 _9862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf0 ),
    .Y(_1508_)
);

OAI21X1 _9863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1507_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1508_),
    .Y(_1498_[5])
);

INVX1 _9864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [6]),
    .Y(_1509_)
);

NAND2X1 _9865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf0 ),
    .Y(_1510_)
);

OAI21X1 _9866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1509_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1510_),
    .Y(_1498_[6])
);

INVX1 _9867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [7]),
    .Y(_1511_)
);

NAND2X1 _9868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf0 ),
    .Y(_1512_)
);

OAI21X1 _9869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1512_),
    .Y(_1498_[7])
);

INVX1 _9870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [8]),
    .Y(_1513_)
);

NAND2X1 _9871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf0 ),
    .Y(_1514_)
);

OAI21X1 _9872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1514_),
    .Y(_1498_[8])
);

INVX1 _9873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [9]),
    .Y(_1515_)
);

NAND2X1 _9874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_9_bF$buf4 ),
    .Y(_1516_)
);

OAI21X1 _9875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1516_),
    .Y(_1498_[9])
);

INVX1 _9876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [10]),
    .Y(_1517_)
);

NAND2X1 _9877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_10_bF$buf4 ),
    .Y(_1518_)
);

OAI21X1 _9878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1517_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1518_),
    .Y(_1498_[10])
);

INVX1 _9879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [11]),
    .Y(_1519_)
);

NAND2X1 _9880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_11_bF$buf4 ),
    .Y(_1520_)
);

OAI21X1 _9881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1519_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1520_),
    .Y(_1498_[11])
);

INVX1 _9882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [12]),
    .Y(_1521_)
);

NAND2X1 _9883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_12_bF$buf4 ),
    .Y(_1522_)
);

OAI21X1 _9884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1521_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1522_),
    .Y(_1498_[12])
);

INVX1 _9885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [13]),
    .Y(_1523_)
);

NAND2X1 _9886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_13_bF$buf4 ),
    .Y(_1524_)
);

OAI21X1 _9887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1523_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1524_),
    .Y(_1498_[13])
);

INVX1 _9888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [14]),
    .Y(_1525_)
);

NAND2X1 _9889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_14_bF$buf4 ),
    .Y(_1526_)
);

OAI21X1 _9890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1526_),
    .Y(_1498_[14])
);

INVX1 _9891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [15]),
    .Y(_1527_)
);

NAND2X1 _9892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_15_bF$buf4 ),
    .Y(_1528_)
);

OAI21X1 _9893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1528_),
    .Y(_1498_[15])
);

INVX1 _9894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [16]),
    .Y(_1529_)
);

NAND2X1 _9895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_16_bF$buf4 ),
    .Y(_1530_)
);

OAI21X1 _9896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1530_),
    .Y(_1498_[16])
);

INVX1 _9897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [17]),
    .Y(_1531_)
);

NAND2X1 _9898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_17_bF$buf4 ),
    .Y(_1532_)
);

OAI21X1 _9899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1531_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1532_),
    .Y(_1498_[17])
);

INVX1 _9900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [18]),
    .Y(_1533_)
);

NAND2X1 _9901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_18_bF$buf4 ),
    .Y(_1534_)
);

OAI21X1 _9902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1533_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1534_),
    .Y(_1498_[18])
);

INVX1 _9903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [19]),
    .Y(_1535_)
);

NAND2X1 _9904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_19_bF$buf4 ),
    .Y(_1536_)
);

OAI21X1 _9905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1535_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1536_),
    .Y(_1498_[19])
);

INVX1 _9906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [20]),
    .Y(_1537_)
);

NAND2X1 _9907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_20_bF$buf4 ),
    .Y(_1538_)
);

OAI21X1 _9908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1538_),
    .Y(_1498_[20])
);

INVX1 _9909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [21]),
    .Y(_1539_)
);

NAND2X1 _9910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_21_bF$buf4 ),
    .Y(_1540_)
);

OAI21X1 _9911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1540_),
    .Y(_1498_[21])
);

INVX1 _9912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [22]),
    .Y(_1541_)
);

NAND2X1 _9913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_22_bF$buf4 ),
    .Y(_1542_)
);

OAI21X1 _9914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1541_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1542_),
    .Y(_1498_[22])
);

INVX1 _9915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [23]),
    .Y(_1543_)
);

NAND2X1 _9916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_23_bF$buf4 ),
    .Y(_1544_)
);

OAI21X1 _9917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1543_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1544_),
    .Y(_1498_[23])
);

INVX1 _9918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [24]),
    .Y(_1545_)
);

NAND2X1 _9919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_24_bF$buf4 ),
    .Y(_1546_)
);

OAI21X1 _9920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1545_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1546_),
    .Y(_1498_[24])
);

INVX1 _9921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [25]),
    .Y(_1547_)
);

NAND2X1 _9922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_25_bF$buf4 ),
    .Y(_1548_)
);

OAI21X1 _9923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1548_),
    .Y(_1498_[25])
);

INVX1 _9924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [26]),
    .Y(_1549_)
);

NAND2X1 _9925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_26_bF$buf4 ),
    .Y(_1550_)
);

OAI21X1 _9926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1550_),
    .Y(_1498_[26])
);

INVX1 _9927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [27]),
    .Y(_1551_)
);

NAND2X1 _9928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_27_bF$buf4 ),
    .Y(_1552_)
);

OAI21X1 _9929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1551_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1552_),
    .Y(_1498_[27])
);

INVX1 _9930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [28]),
    .Y(_1553_)
);

NAND2X1 _9931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf7 ),
    .B(\datapath_1.mux_wd3.dout_28_bF$buf4 ),
    .Y(_1554_)
);

OAI21X1 _9932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf6 ),
    .C(_1554_),
    .Y(_1498_[28])
);

INVX1 _9933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [29]),
    .Y(_1555_)
);

NAND2X1 _9934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf5 ),
    .B(\datapath_1.mux_wd3.dout_29_bF$buf4 ),
    .Y(_1556_)
);

OAI21X1 _9935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf4 ),
    .C(_1556_),
    .Y(_1498_[29])
);

INVX1 _9936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [30]),
    .Y(_1557_)
);

NAND2X1 _9937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf3 ),
    .B(\datapath_1.mux_wd3.dout_30_bF$buf4 ),
    .Y(_1558_)
);

OAI21X1 _9938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf2 ),
    .C(_1558_),
    .Y(_1498_[30])
);

INVX1 _9939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[24] [31]),
    .Y(_1559_)
);

NAND2X1 _9940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_24_bF$buf1 ),
    .B(\datapath_1.mux_wd3.dout_31_bF$buf4 ),
    .Y(_1560_)
);

OAI21X1 _9941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1559_),
    .B(\datapath_1.regfile_1.regEn_24_bF$buf0 ),
    .C(_1560_),
    .Y(_1498_[31])
);

DFFSR _9942_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf65),
    .D(_1498_[0]),
    .Q(\datapath_1.regfile_1.regOut[24] [0]),
    .R(rst_bF$buf65),
    .S(vdd)
);

DFFSR _9943_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf64),
    .D(_1498_[1]),
    .Q(\datapath_1.regfile_1.regOut[24] [1]),
    .R(rst_bF$buf64),
    .S(vdd)
);

DFFSR _9944_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf63),
    .D(_1498_[2]),
    .Q(\datapath_1.regfile_1.regOut[24] [2]),
    .R(rst_bF$buf63),
    .S(vdd)
);

DFFSR _9945_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf62),
    .D(_1498_[3]),
    .Q(\datapath_1.regfile_1.regOut[24] [3]),
    .R(rst_bF$buf62),
    .S(vdd)
);

DFFSR _9946_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf61),
    .D(_1498_[4]),
    .Q(\datapath_1.regfile_1.regOut[24] [4]),
    .R(rst_bF$buf61),
    .S(vdd)
);

DFFSR _9947_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf60),
    .D(_1498_[5]),
    .Q(\datapath_1.regfile_1.regOut[24] [5]),
    .R(rst_bF$buf60),
    .S(vdd)
);

DFFSR _9948_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf59),
    .D(_1498_[6]),
    .Q(\datapath_1.regfile_1.regOut[24] [6]),
    .R(rst_bF$buf59),
    .S(vdd)
);

DFFSR _9949_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf58),
    .D(_1498_[7]),
    .Q(\datapath_1.regfile_1.regOut[24] [7]),
    .R(rst_bF$buf58),
    .S(vdd)
);

DFFSR _9950_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf57),
    .D(_1498_[8]),
    .Q(\datapath_1.regfile_1.regOut[24] [8]),
    .R(rst_bF$buf57),
    .S(vdd)
);

DFFSR _9951_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf56),
    .D(_1498_[9]),
    .Q(\datapath_1.regfile_1.regOut[24] [9]),
    .R(rst_bF$buf56),
    .S(vdd)
);

DFFSR _9952_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf55),
    .D(_1498_[10]),
    .Q(\datapath_1.regfile_1.regOut[24] [10]),
    .R(rst_bF$buf55),
    .S(vdd)
);

DFFSR _9953_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf54),
    .D(_1498_[11]),
    .Q(\datapath_1.regfile_1.regOut[24] [11]),
    .R(rst_bF$buf54),
    .S(vdd)
);

DFFSR _9954_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf53),
    .D(_1498_[12]),
    .Q(\datapath_1.regfile_1.regOut[24] [12]),
    .R(rst_bF$buf53),
    .S(vdd)
);

DFFSR _9955_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf52),
    .D(_1498_[13]),
    .Q(\datapath_1.regfile_1.regOut[24] [13]),
    .R(rst_bF$buf52),
    .S(vdd)
);

DFFSR _9956_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf51),
    .D(_1498_[14]),
    .Q(\datapath_1.regfile_1.regOut[24] [14]),
    .R(rst_bF$buf51),
    .S(vdd)
);

DFFSR _9957_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf50),
    .D(_1498_[15]),
    .Q(\datapath_1.regfile_1.regOut[24] [15]),
    .R(rst_bF$buf50),
    .S(vdd)
);

DFFSR _9958_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf49),
    .D(_1498_[16]),
    .Q(\datapath_1.regfile_1.regOut[24] [16]),
    .R(rst_bF$buf49),
    .S(vdd)
);

DFFSR _9959_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf48),
    .D(_1498_[17]),
    .Q(\datapath_1.regfile_1.regOut[24] [17]),
    .R(rst_bF$buf48),
    .S(vdd)
);

DFFSR _9960_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf47),
    .D(_1498_[18]),
    .Q(\datapath_1.regfile_1.regOut[24] [18]),
    .R(rst_bF$buf47),
    .S(vdd)
);

DFFSR _9961_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf46),
    .D(_1498_[19]),
    .Q(\datapath_1.regfile_1.regOut[24] [19]),
    .R(rst_bF$buf46),
    .S(vdd)
);

DFFSR _9962_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf45),
    .D(_1498_[20]),
    .Q(\datapath_1.regfile_1.regOut[24] [20]),
    .R(rst_bF$buf45),
    .S(vdd)
);

DFFSR _9963_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf44),
    .D(_1498_[21]),
    .Q(\datapath_1.regfile_1.regOut[24] [21]),
    .R(rst_bF$buf44),
    .S(vdd)
);

DFFSR _9964_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf43),
    .D(_1498_[22]),
    .Q(\datapath_1.regfile_1.regOut[24] [22]),
    .R(rst_bF$buf43),
    .S(vdd)
);

DFFSR _9965_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf42),
    .D(_1498_[23]),
    .Q(\datapath_1.regfile_1.regOut[24] [23]),
    .R(rst_bF$buf42),
    .S(vdd)
);

DFFSR _9966_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf41),
    .D(_1498_[24]),
    .Q(\datapath_1.regfile_1.regOut[24] [24]),
    .R(rst_bF$buf41),
    .S(vdd)
);

DFFSR _9967_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf40),
    .D(_1498_[25]),
    .Q(\datapath_1.regfile_1.regOut[24] [25]),
    .R(rst_bF$buf40),
    .S(vdd)
);

DFFSR _9968_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf39),
    .D(_1498_[26]),
    .Q(\datapath_1.regfile_1.regOut[24] [26]),
    .R(rst_bF$buf39),
    .S(vdd)
);

DFFSR _9969_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf38),
    .D(_1498_[27]),
    .Q(\datapath_1.regfile_1.regOut[24] [27]),
    .R(rst_bF$buf38),
    .S(vdd)
);

DFFSR _9970_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf37),
    .D(_1498_[28]),
    .Q(\datapath_1.regfile_1.regOut[24] [28]),
    .R(rst_bF$buf37),
    .S(vdd)
);

DFFSR _9971_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf36),
    .D(_1498_[29]),
    .Q(\datapath_1.regfile_1.regOut[24] [29]),
    .R(rst_bF$buf36),
    .S(vdd)
);

DFFSR _9972_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf35),
    .D(_1498_[30]),
    .Q(\datapath_1.regfile_1.regOut[24] [30]),
    .R(rst_bF$buf35),
    .S(vdd)
);

DFFSR _9973_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf34),
    .D(_1498_[31]),
    .Q(\datapath_1.regfile_1.regOut[24] [31]),
    .R(rst_bF$buf34),
    .S(vdd)
);

INVX1 _9974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [0]),
    .Y(_1626_)
);

NAND2X1 _9975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.mux_wd3.dout_0_bF$buf4 ),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .Y(_1627_)
);

OAI21X1 _9976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1626_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1627_),
    .Y(_1563_[0])
);

INVX1 _9977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [1]),
    .Y(_1564_)
);

NAND2X1 _9978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_1_bF$buf4 ),
    .Y(_1565_)
);

OAI21X1 _9979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1565_),
    .Y(_1563_[1])
);

INVX1 _9980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [2]),
    .Y(_1566_)
);

NAND2X1 _9981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_2_bF$buf4 ),
    .Y(_1567_)
);

OAI21X1 _9982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1567_),
    .Y(_1563_[2])
);

INVX1 _9983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [3]),
    .Y(_1568_)
);

NAND2X1 _9984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_3_bF$buf4 ),
    .Y(_1569_)
);

OAI21X1 _9985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1568_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1569_),
    .Y(_1563_[3])
);

INVX1 _9986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [4]),
    .Y(_1570_)
);

NAND2X1 _9987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_4_bF$buf4 ),
    .Y(_1571_)
);

OAI21X1 _9988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1570_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf7 ),
    .C(_1571_),
    .Y(_1563_[4])
);

INVX1 _9989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [5]),
    .Y(_1572_)
);

NAND2X1 _9990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf6 ),
    .B(\datapath_1.mux_wd3.dout_5_bF$buf4 ),
    .Y(_1573_)
);

OAI21X1 _9991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1572_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf5 ),
    .C(_1573_),
    .Y(_1563_[5])
);

INVX1 _9992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [6]),
    .Y(_1574_)
);

NAND2X1 _9993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf4 ),
    .B(\datapath_1.mux_wd3.dout_6_bF$buf4 ),
    .Y(_1575_)
);

OAI21X1 _9994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf3 ),
    .C(_1575_),
    .Y(_1563_[6])
);

INVX1 _9995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [7]),
    .Y(_1576_)
);

NAND2X1 _9996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf2 ),
    .B(\datapath_1.mux_wd3.dout_7_bF$buf4 ),
    .Y(_1577_)
);

OAI21X1 _9997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .B(\datapath_1.regfile_1.regEn_25_bF$buf1 ),
    .C(_1577_),
    .Y(_1563_[7])
);

INVX1 _9998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regOut[25] [8]),
    .Y(_1578_)
);

NAND2X1 _9999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath_1.regfile_1.regEn_25_bF$buf0 ),
    .B(\datapath_1.mux_wd3.dout_8_bF$buf4 ),
    .Y(_1579_)
);

endmodule
